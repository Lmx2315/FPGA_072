// (C) 2001-2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
tAcKgjPoRJlwf9j2xe/wEUmb9cWsV0LeOgWNh0LC6oa+e3STLvugxEqzkg0v9PS3hhSTPMZHUcDC
cKQ+uxD2Y/NpnI/sORh+2qPQVzzXN9LbPniHMelGQTj2W/SjhepKHbpFOSW0oYbSmrRMTUZKI7Vf
SZpxjAIQO2WFoyEwruR2OEg6HvWnW97yGAs/rLdD79qOhKSrxoE9Q82X6x7C+2uPUkomgWVE3vPV
rkZMaLBikThX9p9o/0k82jIzELNBeqY5rjRl0kSeMoawNxbbN1UvM7PQ7gM6iuX+DL0i1ed3iJCU
n+1I74hsmTiTNs1f/Mpdh1AIEvKCon0sUk4d9Q==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 9008)
neUYXXEOKrzDDXyxF2IX/2bZqwHn84/gpV5jDz1zg7KviH1NfYzRaWiWLxrTBIYPm8fHONUIzORy
uuuaNsP1fIgtZSwkVq7OBbXidCgKWXf5r+FvhiGuK2fARvR1ntiS3scVT/lVBNyEFqPoY3wAWLMO
Gq2X/SfoP8NIGccDfxmPf6fRAN3JbjmGgrz8ykJDjspRdXTWZxdzm6EnN2tiI4+ojg7zalpBR+CG
zogimUaHFeYFCdquJGZwkSDc5xs8m01d0gkS6LulI+kgOI3gLWf/8X0XjrY/mTHcCgKmoEpjeN/+
69vDDLIUnvglA9G/KWt6tzH9E2hz4SqxJtMpWv+LMTaQvp8REhlGmGONPlpi98eS8ZNAhlimejwj
ajGMkJnXh3HkbJc7R9iiJFhl2o5e1T33O3G4i7H3pFnMJhQ0uMmDJ9roxLILDMcnaCJrA0WMuG1X
iEvjHkf1qhFNuf1BFJ19u1xdlM9P8bn2lWbgJ9tE4H4BzRDcgphDVbEuoV1ggqPeVAp/U3umT8O+
z1hSCcm0oOHk/buhbmiAa2feSCnWzMKuCmS9d79gb+f15T60pfTpZLhRMWlLsOgr60ddYIRFqajp
qxUS8+BIc0WH2OouvzGYPUYJ00PCuCD6p4TXqLno3k9B4U0CcgsrEZ3iH67SsrRm6VVIqgvuRr/9
qaf+3iQrosfslResroiW+MHBXgesdrxtl+HBS8BWQkRpJJbcMrcNB70MBFo/w8YlyK4kYFSbJrAg
Y00qDMYCZnwk1URtrzObyZKvwjB0mx+qv11CwjHwzHB/n99FdZbdCPLmLa/RhXCSNAWJ5O1erBmR
Rx7puBH9B/28jcBkvvsF6zpZuURKcgT77pR0BFSkQu46ADDpCqHbRm5QI1RarnllhHFJAtROY9/N
SiqXi32hgBOn+0F07mrzZxIT4r6+7liO7RTMXdwdkH7I8DbhZjwbzojcpy3zynHd2bRQfnzOY2I3
mfPiowoOQmieKPek8XbHiroStkAD4z5v4/n1mK0T/7y8bvYok058lVb52HLUBAzbz9/aHaP8cKhJ
41x1J+va1I7wA/7OKt3xYvQ6M1sVVrFb3p1fzp5v85Z88VTNFQ/SLBbLgvHDoIA/KbdMUMFooJXk
COU6XRVEAf81RbTcTp/F5a3NdGPdqOxbrVQsaQlsGVVDvXrXh6+xzXLK4oxTASEolrh+H6QPXXhF
YsfBNygy4RJ+M6HApsOAXQCydgMkvfoNEoO7PcYmkkcDlOt81i8NFO2qTJJsjim7ZgzYbz0YhIvM
Gs1UGamhjjMgIQ7y4U6kxcfPMGLmWnhypkBBXnrvMZUrgo13EVF/qIg/mmBwyV0Y6dnyJcmOOVAg
H7DBNo3bRXyyHzSQ9QCwX0m1zfUI5YcCDxi+KsJDCxV2ufYFE0bXfdfWVF3NYmoLgzybfu69MgOg
LbBZsAM/mxoKXnyswNOohswFX573yHubg51ltvgax6R8MY87NivV/oFVmJwON3SCQlfELkohAvY8
aVwPrNek1u6/KpP1GZSPG/7RRGUh3SvaCLMQs5e5na5wCXl4zSXJCTPsJyy//F3OgmwlINJfZWqh
GnOlCm7mVQQJsbOwh1L8KJCguAznXZIFtEajKtgYR9g+pJ1mw/LxF5ukhiRupAJFA2ZyJrM04pgC
NPtO5aGZzpeJd8o7lQaRWR+deL7fKuLN8BIZ0Z6oYJEnfqDBpr070yC3Vv/RdhmrM6juhGutTZBp
yAWX7aH66eJcGVk+y2lKy0rHkb7tHKs6QvgOhhTu/bjQdwQF+zQtO5qfHzGxUFvB0vwU6WtcV2EY
7v22J4BOujig0bqcwZNjrxAUEMWV3W+K8lflCbf5XfuNZkYXB52C65iLi214ukfyn5ot0IQnW8IX
smWLrfEYwHQV1Hg94LRMOhAOcRNrKlPrsrMNPmFMzMSuHy+zEndXYCwxff3J3JGbNdz+l3mJJoIk
u/dcazFYwner9Rd8TbCZMqNEYmCDQrte5Y3Cl8SXe+gz9ySHFUsUZZOZQmC5itPXboUS97uuuWmx
yxXUEG6Rzr20VzuOp3nlLwzfsVOVZj25aZccON927kfOy8lH7T8gu0eRLgSIkyufMsuSIJ8fAN8U
LoI0uHyyf+ZbfZ2PUdh38+U6voZZ+bBnhjLRpKBhMXmJomsSV3byqvooswzAlPlVp+/dxFHf0GUN
3di1BeDghgSkqVeueuMdcXqo6gKXdTA63pwVta7Yh3FeaxlANbUOP1Hqfv6ODhmH4Gfl598EanUt
WMv/dMJ2hfLCC73lpbHei4AeYMQLPT9gOMdnAMKYoz4jNTGKHvttPcXJyM91efxlFZ6NsMUIjo8+
wIhJz4vK/efY6YgL30EuP1hu+AMu3xobp9P641hPsxVGJrQNelm4L4fNiJNg48CflWxBXQO8jsCD
teypLMyzrKiJCH9TwAWBvSWY8Kz3utR6ZRvbQoS4KIP94dybbdJ+yhKAqgKzW3cVQ7sDpLY5/jHB
0bUX75RrJC35tZNyCBXO3dQW91Rp3a0OL4sh9O5dmvAoEhW3bSDDyWQZS6QTe4fepSlZmhes/1sW
z0JxN3NAvoIBVF88lj0ARohB08W4W5lORnv0n0xJ8FMXFMyE7XzGQQn4pARJexmxxHdiDofzNTe5
CIJUtlVfScVrwlKN82bNyEA4AieKMJPvIlU0Mw2rBZq05q0GmFXJCr4T+qEKTSdg1pk9XDWIDMkM
pGZ5XKhpMOafBm5spYlPTOOT6T4vztF10NT7T2VDoTT4GcBZM8QwIRkB0M08GP12SCsHO4tw2BwJ
rMvS2IEjjgMjn+X/Z/GLpsPyjevY74zCfYVI0Q3FVaKLJGjoIK+dzyr0lKXjuj8977eIpSkMaWk7
Qwg3IQWl4mmDL8nHwtzJuDVMhSL2GtfKGvPO9siF9c8IICjzXKGK2EvJ7egjRee+BR62D33u5svo
zUl/UQaUv9si1jmCqfAkfPrj9sIr1j4IxvHUDeHa8JQBGpyU1XVKJZUfzWDXt9N+DMNUcHyS2PMZ
7ZlMGm7XfmFzJIDlmZBjWPSA7eTOG+FXoGJ11FrDp/x0vhOu5ZVbscchpjUEK2mCQBVXuepfOKee
HmTuZT+Xp9Y6chH7NTf1C1Mus3k6pslvx9A7YRd+sfRK3NBDjhnIkzxtBnpdAzzbSL9mr2aLKdEM
wSnGHCu0Agdm69uSwGmAxOXSb9OsUn/YxaTvh2/bD8OeDiugjq8jTEUvnz1zuIQCTU6dK8cHKKcE
pPhpp2idfgBZlzi/qLna5XEfDxK2dolG9i8RGhWUECxZGHZtJnFVgeOIwpLkFN4GKcQE8f63PfeK
0maOj6HFPTWyU1UNX3lX9b1wYP/SSyZ31cJP499dBg9I2YmyN80UKrlw/khxcMCqP876T9syP0kN
nN0Ih19MKk1cnl4gW57h9Ztzx/5zk2oW3naWICzW5oFXO4X8OH20vQWw8gytcMMpotMbFM9uX+SI
d65TUlvIiCit6lYKiQTUqGdGYXYievVIFN9V7CmmSlpbJWfEor6s00J3FE6ePWsoOhIk9S8ss8Z3
EXIAVxzQBs32sx9Upm2Z2z1+5awUL2nLSpfHs5ryt79iokPOhb8D2M8pjvEyTruvBCG8IdFTwJxS
7UgutuAzLpi5SJxCSEjjneJvUPjzSf/GfK0sW8sAVW4SKQM660XCJFc13Ysya3d4fByw3HA78X8/
A9vX/0goxq7UV8S6QycJKITwLMpPy1hbOGeojnTxvivoN1kmSjypMX3R4MSJXFWv7gLIbrVk6ERE
dUIyJDWe29VnN9VTnljE+sCDJFX9k3hue/1hZ+A4WwHte2IBnJ+OemXczpmvtgxCZH/6tdb0K06Y
QTKxsK/Ohi6PmJrj8tGGMyhAF0CcTCt2MFQOyBsU3OZoo7vXPmeWrtNAN/4pSrW1iA5mNKi2m91/
IjSuBDDcxlQG+lfdhE5ATYPGOCrlYDEyT3jn4ZrL3B/R+DEitf9DGLPXXZYGFF+0058kzEniYIed
DCqhN5Fccpx2etf3p/6KjjVwaARWuYjlYBaFCbIK/RFJaNgjO6kpL/72dhQ3O8FYw0cQUzy8V4Ec
d/C9yEMVGVnJF/f7sm3Ms5N4EHHC3PVDAM8cyW3xXQR7i5yzHyd8+zqwoLvw303wrCRysHTLB1fp
bFl3vUzh14XdpN0cl3W95Lc3ZlE/KCnxCxmOyJFja9GXg4nX8ouWMn7qy2iASGBAIpCEIsbq6/l1
N6BjsSOUlFFaeKYZjGffqJTva/DatyM7LSl4OMg2teRLN5ebhaFgCZXO/7Le4d2vQ7eGP8MmyLcT
Oc2rPEBEIvtXhtF+CXTC7c+J+wOXmW0Ss/lqzKcNWcVHJ1eACfNTmJftJUoJDRF9ShN7qbbzGpyL
RrG4OgSa5/5xLcrePjHIpsMGBISmrPXcV/pL9MPSUc+s9BfXoTBevqwKWKnetkeEvli+DuAqVqB7
MwdV8P+05UWbzu25s7Osgg0/lo26IT/IsOsO8VJXt07ZJfKNw9x6bC5wM0hyat1QkLeRgwIu33in
QrlqcIeM3BWe+HPir5DrR6Ar2IY8zIq1GBp6tenK+9Pi1ArZn/DunoX4ZTKNsdikW+c41z114jp2
xvDcCE6pDIpTr5p7IK51qKBaihIXBDu9ex/Yl0SYs9h4xDuNCgCiimW6NUrkONA+tRh5wo949dIH
EQ8mJTtJ5GkXgdekCCPuOVOn5lXG/VrWw0E5tlECEWO9xXfYpZwXIvgyEENxRFlKgTr5B8Z9gbPf
n5y2eK2apYjf17p4/uURwvz3Q21pWpZwQjY7pPVcVm/wPB3HljbeSqsbanfmmdQ2dD2F+AKDgNF7
L54fRaFMPKFyYYFnukc4w4x11xMsqAvo5aZSQP9V1ZA3DchvbGnKHcWyqh+tB6TdkH2UzzehsA/7
GGxQmqEy6w5abgUpmdUUmM0gzgAtND2GGeL/02pkaw7GU/Twz1FvmzGKwS9EAxCgDS30sqtUokB9
mTznDtxARReIzQzTQTvCjRmV5ceGgeigdgnYJYmtpEnYoq3EBUDcSYX2RjK1dlytz5wdxC4C1WxR
fBnafILEpuaiZqZ4RpLiPXTBcvL/LtnxK3FaUSzqknc9tZm/KJwfIlCEL+YvG9O49gW6tSFNh0eB
+6Ht8ZmwOfof3HRhtDTfSdkPCpkKs8EAJPc3n/Bk/hqixSemmzALTvL/MKsIEhSQNclyOlm3b0LD
iieUtWgFxvklDmW+bSV1mvm1n452m/SkMiogB1BtWpQ5biKRhK/0RoiIAWCTP6Gyhnb+nULo2zBz
dBuz+HF606gtmsUQvgD5GCPgWEqNHaIx6hRN2jOBRf+znmQQGRdKPNsqX2IP8h7EUNPEx2jEYuJP
og+xlGU1v/bkHQj147VT/zslcPjETNRXZFFQON8jY6h11/70puuknFm0gnjat6WrQXZ1Hq+F/kjS
ogbjUsjPZQb1qcQhkAQHnWy/6bzAcDcdDDFgPR9xaSXIQHi/jpf1+kGxJyjNwycGGlZnGqhM1BaX
5KK6XI1+HUQrI4RYQbNmixd/kZHejfy66cDNURm3aIEtghDjhs6CzbeHO2ahJZLcyVUWMQR+W/5W
FfRgK22fRfnCC6UR+NHnqwq3bwGWO1H205kIiMRaFrOLJUgU0+nGle2KmKY3K5cA+FOdixJor+iY
z8Jw+GcMopWJCu+akgHn5P9UmMoV07kN3lPORudioSfzs2Cx3zC14+nP8wPttI0hH90ahES7v9vG
Ak/BlKHBtwuhk4kXrDwO05ULb8Jyimo+LFCV9swpieRZBVjOFbKXas7tTyP9DC3eZXfdSDQqfG7r
C22cIjPIi+Szev9jO8jrkUFQqc7NoOAFsLpQUUInLvlLcZXnP45rR39H0pwmZIAIrQMqPh5cjnAe
E14Au28WZ3UC8NyFuZgwrOGOM26vADiRmSEWEBGAJQZQ+g0HV+TdXHgwwZ8e69/4+4IiuwayIti2
1ebt30G2uaA9LkEKfrJA64brvS+NuEmNb8eRquMIrt9RsH4idOSFqqkkRQ3WV2HFOzia1m3y0+lF
3IwWFBJvp1U8lAVJkGpBUiyF4fSJGRGjzrwOanSl8xjpl9MGDtb56k4EFmnuNEBAwTSacW4o2f8D
9SUfvhCkIPgwIcx19Ipv0BE6/p8o66y8PU42rNVBwOOwjwgHAfPkbr4ibHCeqc7JJrYTk8bxsXfN
5286Z0WOhW+zaoajwmFBGms6lL7lFoI0dju452IvwrrA35aL9PGvpCS3OWZzqbAba4akVGhWSy6G
GIf9bLFQPQCeZ+/Ul4nVbIVOuBfOlRyVLnI5HloIkPZAnQxEbvaradlcpIO24VnWlGK+kvV/YyuZ
FRurZpOZ7aNdlybrGzxYCmkSxOt1V7jdW3r5wAolFzIsyRJgt2Q4sOKFUU6NVVMCxPqxS838yqZq
YFLUObVozXcTJ5yqcHydYm/+uOYFDm8CxSwQ5OmH9GdAoRWecx2eW+ONUJTdYbP3zaOmtROnCkcK
2hVgSSAFbHzmLYhTIWZ+5Ntt4TndNdldiKyUuR2GlakID2x295PSqX4BdYLxLFuCcVvZPcPO3XHS
qQFwGS6FJYWplqv09/uuBlte7TY3U7aSkmRlb0Q689UPIUAmHY63wf55b42l8use3nphuUv0FyoN
0dUMloIzU44i+Hsccrs6FJRbtJc22ukYP6LfDPcEeiisiHK9VpNqOns1BI7k90bTFy+AjlxP0gJT
4WF1Y1aEfVdd+myZXddUr1Fuy8ewOHcTp3M0lF3EQudXeCbkzYCGpZVIRhkagPPmMQEROfrA6X4z
wl/qBl5I8W0ffmwklVCCBcpgkWZU7Np6HuVk9mBUe8ibATeGUbIJEgPs8k4VNsnMtpxwOehLIVX1
GXbpYGnMVRQTKp5b8nBWdrNgsLFqzU7VdsobsLSroYDfQDfNk3TjV31FX8CZbVRocJziZKeFCPwi
VNwsD3gC1dXcSco+in0obV/0rU1juTodugKqybR2y3mTXfwa7eH9RsoOk9Dt1bVFEQD5V+pk1+mI
RQgXMPIw0wJ8kSIZHSGdW042CMl+GF+PMQwSUqRJYKhZFp2HvpLuq2Y6n/efyGWHQJdFeRJjRjk7
w0OpBRBvYh9gyq4HZoCt0V5ATRnAJsR/EAEfSb+vpwEi8ox3ebyFwe7nTCyeQsMbVxyrgocu5Seh
3O61WkhysgGBOMgTi06TXZhgfWQTzTDtXVhrjAOb+CDJAW1xyPNEnfFsFSxVPaBm4xhP+HY4N+Sv
saj+j7DtQEqqqgmHr1uqVSRvRD4E5wncBSFNlz949AYHAOjrQdHVU8oBB6DJnSTsdY+e60rk8thG
kkUV+G9d7FF1NPfD6VpFrptO0VabWP/06tHJDqLCyWk7Pjg0WL5EHM6wgT/34Z4jpzXyPN6Q2Qu1
jrbHy/Iu02j9CtZdjscyoAe82oCdn/m8AMTAvXn1fwp9n2GthgBF52YiD1jWhOKCvabJxN4FC37B
lE/M03VHlbZx1XrS1O3knygGdAL8XcMNz+ooaY4kGUMipru08rgY7WPSS52eld5yPKv5Ua1a9+bo
3sMWFDOpGAPoj82R/n85o142R5xPzZFLxRCC7vpo3+EgBqI3pR2G8RDNmdzYgHkSW97MmrRHlVYE
kdu4Wg1KFpQSTDoFJI/57JFu/kQkhus+bNpV2/Xj+roBvfKt7RCb+l2iEtcrPkOeQXReTJBfZHR/
yMIaapgFCIffb+Rc4FF7lehbV1wCqQP3FiBb5gR58tc4xnA8Xfnhcndbl//Gd2Fs6rAfczK7nNke
60V8lydAy4AtSV/pwnAzlE0U3YC0D/vskIBTKSkWArHhcDNWcflOCsWzKb89s0ZQERhzid6Az6yA
+r4lmibECcMxp+JTqPO1frKRZN3PM7El4Jk5wYspmNku8pbl5a5SxW1WSfLTRL/gIDSWCOHGz3Q2
EuJ/2sf9DtXDPsycRkhXfe0fyUgDi4qpofQwXPGK/c4LztdXt+hdjH/OjhaJTk6kdOKnUJDWaii0
oFpKgFTXoBUaXNFEwvtp8tpFPqtsh7MLzOVhznDf8heOQYQtY/4oaf3ds4pOFC5nJd3B39M17bx9
zibDgW3G4PIM9AvRcBO4zeG5B6tEu3yYonjNT7Nbk5wXNZEBzkS51CS5PfceSodNFxYGe1uHiZua
uC5OZqrGn0S7venENFkpvglnDdCSyBAnt31My5sc+8Qi+l3jKfa0KJiMcKMS1uaaXWxnkXH1pUrc
mcNq0jW3aIJTuN7EdvbanFDQFu4WJSpFQoTIU3M7uqfK9iJ8G2QByDJo3pTTgLhACrMFrWeik6hs
xe+SP1ScWjtQ2OXCHrfkFo/2lnLWD9fVtjzMRju9nSv4HXw3yjb4Qg1JCn45zc5wtsbmie27qmTA
W8AoCZ+WDu11WKSgtANvG16BC0mfAYht2a5sfndbIRLq44PsewludWnJvDGEDrKJG4XLtK+KU+hc
2LBXO8U1Rl9aF50lf/Dwq/o8+E/dWAzM5ROcmSy3wblIOyPBa20P99nzEW2cHAL8FjtGv1TQ7crP
WkG/JdFXFK2Vpyho6dGwWjIgp9Lm5qnTNRIq25AS6qVfu+4c4T1po3h/8aefOTr1VJPZnMcA1jgO
XJZdW1Uy1ghGGcG/hNOURq0s2CgjrVjEDjqipLim7cCt69YBlcV6gwU2Eew8p4fw/cBV0NzAZ3BF
kJbj/OOLDNLbym9Bu3Jx6YFl/lPKBvQtMRDMkWc3nM85ozb7fIOKV2tb9W7O9ZuEG6napOboM3zV
XFp68xDB/dtTJtz9NNET3JM0DH3UDfQGbkvc75FpAIEWmtf0PJHjr53JrsxVpD8AQxLFtTmsa1Rs
rSV1FrOWF55EdKqGhFy0/yzfeBdPN4mmeHt0e/60tTWwbX+Un76BmgGxF3KYfv4Z8AkowVU0X7D/
/BdqBdqnrWbZFCC/Q9ShaNVtIZZczSZ40tJxhIVLVPhoSAg0L0tE9vNlzZyoHKPj9EwKWGvZCylL
rc1zhFfPvPyiDyeRBDPw9jVcbdbclAsbYBD+ptpmAkkrZGAR2h3zmk2jTdmOqtFciQs8Q6bPa0R3
BwLJn9WmWL1wR/WyCaA/sZDqmD1TFbyXABpdaHZ69kGGH9lJrGYtkvqYGzGms+m9bIlY9lW2uM2m
Hk4PBwQDjHe8FiubzG7BTGGwUUVETHhpYCgpK23Z0MFDAajW911TVxNMqcuiAoecmizdCYIbLDUF
USir0GQ4JYf2v7Cn2ohc/huOwWlIWeGbszlxuY/SOobqQbVhVnCZnL9dg0o/pVZQLsCtarcZJwmH
CJ9a0S813wPdVqbPkhm0x21mDhLGCmN8QE5z+Jtu5900rgrx4JjZf6JJjmds3VOTT4jYfyTjydXu
gtf6f1jNsSGqBap4KAdRxwhiXVLZUktJABYTnbLMt/7n+r0i0HkNxwG5bORFB+IkxOkDbVP0+FXQ
5i1qbJ776b7dxPqHg0pMQoyUSQmS87WwWXos2qFHQaz8uIszW+itQM/WflcsnWkJkXbWijJ70HoL
EFLVe346MZK4HvTxd+z2sYC2fOwqRbe0whlRHSXgCpYRRnZLa3VXGWF2mcSIGVS6nlP+ncZZ+DFP
mnQXtZeh9PYOwW3hK/JsN65oemVJ+b9/J8ujmZjwDz3qyTEZZxadpWSQjzjrpGZLR/frNG2KfeQu
FqZfr5mfxKukSCLUVEG46uSc7C2cabioRtTuO4MJwb0IiEDQm5EBRr34n8d2ikAdUsxKEWxwcBjF
a6zq+sGYqN3aAWhMPFFM/Da0dChZ31J90ZsIU1afCxG80BuWgH3bUImFJj8ieiwM/IjoDmX3adzR
o+1tfpKhLio3M3jUNhx5vceQooXA2gm+4yD0VNSVUKIWQzjF2TkFzUSM6puTBKzMxOuLi92vPoZL
JBJuxN0Bh4v0bidPvJ38E0rEqs3/fkR7dS7KQy7vHunfPvnGusXMSwwV0kF4Eq1a15A6gJy5a4PY
uYC4nRVJSlhzNE2MQVC5e159IigHeRx/5LE6l4blB9Yi63eKj9kxCVmX++OAuzn/AvF2YAQd/uxb
lR+H1nA/TwRw74AWm9zOi1FRIRDQ2//OlSUbvhIH/VVSHRiuIYHxNbRfo911g3vQjuXJo+xijf8p
LSXiHDUdx1wCN91bP+wcE8R6WsRZgMkEsp/hcUcMbnVuexNBcsokyRvzy0dLjeHT14mTCz8BOTTJ
oGFn83Yrw69BOfgdPq6nqfH61zkc2AtGRbwRIF8PA5N39y0+1CBn5U4mbiUpagBjlpDWsywwTQKq
bAJhb6nvVxUYuk7GnHTnhqSEntAbbnbO3sz7ZMOm2p9fI3Mm1KlNvMRcsu9higno52FhgbIdDQJo
BPHjJcBIbMnIma+xvExt//YBbPeM9LjMOfsp9Hz0zg/rH7W/EXz284omuoXs0Z3cG3fu3/iUKZgn
O1MYuzT83f9w2orYJWSl7ZWAWJh3+qTlL2sU1O4uRFK0TEks4lHm+1nRGX1GVV4i8VNtaay8vOf/
+zmXVFyhr0wDsikHuzVf1T8HQJBxqia61sTBcZ/Tkz0KABS2hdFdl7xpeX+IkyBTzG+4YQ3m7CPQ
wuvkFuQNlxdP3q26NEbOlEwK5xUrphWrJOhoc2rAmM4VgB40w452GdY6HTCkksvG1F9ffKsebdbs
emMlMdlgKtk35vrc85UIk9+vnaqjJummvtBodvhlQ4Gkl2ZL1NzCyCuasOaUNg/3thIGX3e1VThE
MKa5IZ7hz3xi73YrcbJSvGOP3I33JBocw5wktrMwWtmtf8+3/Q9V+qLFg8FtgsGQYoBQhYVMw6Bh
lbxFiXpcbECDEgB0mI3sUn+8yw6XdovaOCMEnAQ6cb2nvrVkEPMcUdjSe3LnKHhlbhLN/Z6VZ2dc
14AjMQuEc6wE9Bo8gmTpw5sZBzD6DhAPdOGxKQyPSKhJoSVsmlV7xNlBeh7V9qSPwnUP2dsjDq5+
mucWimlrhzPWa4WmXnmvIvCyKR6DxL2zeLPP8RBlD3YOPUpXJVeqeSKtJEfvYoVjDwAS28lEqAwX
6IibCyPvSoGh8HQmJ94uDgEOjXK5NJ+Pa2Ts5i95R+0Vm0IwQNI+dsfPZs8wO31vncmPUcBP6+CV
7PoYbCyuPUvoUAjhb79jNHEmeQUsaXb/3WY9prrTXLqZWeSB7WlHuOLQtEZfrqhgk992gf00RRwR
DT1uamiiLYrCzDKADevzAC4CHNFZulyddzpWdH6YaH33Kct1CTM21cMPlO5F2qhlhaOgv2JgZNZt
991HWrB3zl7uZOVPMKczHQZrk9gDETOfZ9bt9gw6gLWztVFPPDMuV/+dFV8dHE4wNKa8HEZmCcew
dHF0CyZ9jtlwHSmn4gV6ohWQPvTJJi2DNFDzguTcbWdBc1tX8+G1WmUAv2HHPfcqsxxe+q+s4j++
qrK+1yiDA/0aybwjA4ZiDfOaRiT5XjwAAG5TzSFZraAvFuWh3fpRLLOCpgy9Hlpesno7oKWHRx4e
hEVDy9+EMVPZSgFkE0760PnLwfBuxXkRoGmE8e0xiZKeOGruJBGejCzwTDZ4qf5cV2xSnpZ1yFCN
OdvNhKs/ea42mVxDazjMqbBnXayPwRBVosAMBRFQ8sLOh2oiWs/ugi/4EH8WgaOwflrbYE4kNhyY
89fCIJgnYMCl7IgdPuxJ4QBoi7KVb5U/ckm1SUWBnDg03vcs3gSYiYaHDLwkLufv0IZYpvp7PjS5
UEa2dhYEFcJuihz4+t4WkS/YRy5BMVv01gOyG2Qix05P4BfJr907w9UeYutfWeNbO8cGrXLX2bi8
06AZPlP8osEtwEUh7vO9GiTqy6XfpqLRdFXNmj8stu/7hPkEyWeeCZdRvVNDsjond5a8xf8jk+Np
OVLVymx1Iuaqew/D3E2znU8ndLDouIQrUXUsjmhMrbKFCWJt1e7zqkAOR21yrEZIUxhYYuV0MZrh
1uo=
`pragma protect end_protected
