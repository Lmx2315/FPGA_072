// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.0std
// ALTERA_TIMESTAMP:Wed Apr 26 13:33:43 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
UZ2BrUdaFuIrKMIcmfs8xPOIGM0IYGoQgmInQ+sIJbj2WKozO056jofnIkeocq3Y
dfQ86XJfhPB0B638zE2fVyjOAAcQ72INqOcjS1Wg8Niwh+cT/eLbuX4ggul5tfLy
4kJxJPhHEIsljwPsNlhZlAw1N8F/2ky6lMnaJW6enls=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3040)
IPyf7PxPRh/nYe9JhopDfBIsvUKLZ4rH6SoRpXJzgt870estkUtvQoPpv6MhU4gu
EQv+LTn3mvhHCYEfBeSHRkOtX7Z+P7xFxX9uZrTw5hkzflYkmNRYC9I1KnfAKQ8P
8sHr8d9z1AQndGc30vRmYzHo6RxExjcVXumnVv3BUl22yjmtQ73zjabMeJdzKGg6
WUa9SB6K/2ft3Jhx/rRNIoSNvmej8YfwLLByxXmVzOkPtXTy3528xtQjaQ/ZZmEz
dIDPW8GObReR8MbPMouwIaQv22n4DP3EWGaRprHPiuP6XP5b3xuC3Veuqm2PChyc
vLIfbLSRkihTVGP4CT/20ApBzbfQgbVvLEXuJtQPY895xw/sDvcniGeJ63A/DJz9
SxX5rbkHUWigbSRljU8oOAXsqzPzpOPV3j9krpl6dPlzqHwrsJPM6Sbb2gZ6Qmmk
JvrQVDDqSU86xBKklA5EVYSBZvN8xqlLD2OOz0A43VrzCYNftQ4aLCmm3J3057VH
MVhQkvh0iBNYHCnGjskmmGCd/hPkUxX9hxilLVM971W7JOyLzfqq4d6fkD+GOjVS
j0aw5HNEkTehc+RTajM9TOs2qFWnohHd8pGKkiFKYEYPlLKrNz1yBqLkn9ggKMdt
LEJzURwTYe1h0JXIH7/00aeg+yUiNJDcVrOyMx3zaG6LKZo9xpJeTUFcN1tT2R8n
em6Thl5MgVQSwi1sZEzGjq1WQp118m69pPHExH5AR9i8v7OQ6z/IcLDQZDxQK59m
NN4bJAIMW8PGlnbP50nPmAXzjseBJzGA6k2hFq52Pob1Drv5DdYDBsIqumahjRYD
XRl6m4zTvp4dHLhNR6FwtWaYLhznZ9zRUVTfiyLBtTbHK6drV73rzKK2X/E+C7lL
c2U/z23ew+N1x5+pZx+13uUqRVq3FqaTBr1+DW8qvVkcGPo+Lzf4uGBIXCFAfC9P
O/CmhfpvzcmOXwZNyC6YB0GMx3uyFocSrtzaD5sRCC4qK0VQ3o8EZ024pJBElLh1
1TmI7xmgxpUwnByiTXjMSlFGPskRL2BNWg1EIoPZHVL8xZHxgu18RZWurStw7MMi
7GTXIxMZpLMsIcn+anrPLBng47pNvF1kPYYg7gQ4/d+EwMD7BW63G8+saOnsEO77
FNFb7I1S54MOI/5ySfvtNY+ygONE2xBAIgIqZnRxKD425LMDc5IGGMMCjv0ob1Xx
bn9MZhi1oQk7LzGXe/cPOowI68rOourmTHQ6ZJhAq3B9626z1oaauFiOr4UHlBPA
Z6KEq1YY/47z51l2d58qDBGCCUeXf8aKceZMjeLezlUXxUx9i06c0lmOaihuotsk
CpB+abZTs5KLYLQ8sF4JLqeFeJKnnW8mcsghEs4ck+L07MrOQ03QmxvaanZ8/m+w
tVX9U7l9iT46t/IdfKaGyalnXYQ6zLq4HOKgupk06KdFNzLB/9W0JehKwVytfqdk
OIX3kKCRVi8YlwKFDKy9tZ5sgIqX9Bj9psWdJ58W6v+a1SpJlC2MfjVZJPqrqwnV
6rKWfBmUZkLFYEEw62Vz5vmpAvcBDkdKOI7Z14AAD3ym82xkzlScyTce5K8wZhia
j+IHzdrN/LWgDG5emuni+2rVDxIKCHV0eIirrwt91oK8rWHR3yPfPDmIQEjbbAtc
JWus6zNmHli0peN3b3eoH6Vr6Yh9PQFgFh5c5wmv1W9LU7iA7/AgLWeAl9L4OrQ9
Rjfd75fYHLNfq6KiOpQ1yiUHF2gJt0ZD5JdRGIuhivD6gdvgsYNm2EoFYLSAKcZT
QbWyW4KOI4FY8ZvCEae22u2JLp7u1+4iNW1nLHTCdLMwAyWXsb9ruuNPrK7ER5SH
Wy4t16csLHC4KlF1pVsEvIqASutBdHx52uJwzc8uxd0Fe7kGCLI4MX/9Cn9PolAi
XrLLBIGDclg5Hr77LpeFRJefPjtS8BQP4LLkVEKtA0aMHK9DB018Dt3Ofc02OCrf
TbBMmWhh/fqOC5v45J3bYbcHxdlqy4+p1755qomllkONza2IBOLSB4qx7Paz8vMP
0prGKjn7FSvOlQgT9lAReT/FYbTYW/ISF/7ZOK9YkcxM8wo8qG4wgnB9g1jrxkVa
mX/HaLIZtd30M6bprk1+a/VfvCIhaaLzWGs3Vazg6GUBAbrHs5FMj7FaWb6sR89W
+CYIdVQ9XCHECzXXESXwO/KFHwzQkwy0DArpkp2desPHIiYi0wF3KF+gVU+ruUHf
KjxvkpU0jX5YQrlfeYpZKUs40eltATlh5ggW7uDoliI/N5SzrtUGZKGHgk8qBegT
nSkqGLKMeGDOwvHsWOAuaslsjtyc2PD8GEbMtBfAWEyu3wRzqISpy6dPPj192T75
+/uSi1i62HPRsGkHF4s2QXe+btEFRgNUoFzsOJJrDsaNVEY33Tg2LhOd5XanZquQ
Fw5XPk7MuhMBZJ6WDmbn4NssfN8rY4oG/xy3WwQ4thKul9PHFP7ErrdlYJiOsAdz
U69/6ajABzA5RzAj6gm/r+uuUmaFXiGtmK/phOsBvmtuvq/WYVT+Z29FweOZFp6Y
LdfZ+vRRz7BbkbRixXVdik9EEAfdcudTvDslDlTwuL4bJ8M/KqGkSLh2coO+kLa5
idFKDz0T3MMndgEO4ozUUnmFvE3x7GMxAiY+YJKtrQ9uUgneKwlzNHjcYqZrxQW5
WS8S2ASVjWp+vC4vGKN4k91CcVZhgr6FyECYHpLC3nHRi7DHYSTw1hXlZMCiNU0B
nYopHwNmW84GyEVj8dMfJV2aF9VTAL7PaPtayFJbvfYH4jvv78iGbFVeC/VQ5M+N
o8E2f4nVqCb5UZ4dSGYHeap+HOC2iLJZW1Wd8ls+jAvcDn2jHquoWFrJILhYoPxa
3JpwmZ4Ja7UClrlCqJjcZj0Y6QkMZLEKm/2w0S//kAEL33+AuEOnOu+djmEqreg/
Dd+0VDQH/lPFvXBOwqxLXLNrrULE3izne7yhL7P7ajB1fF3/ZlDc0rNy9vxWeG31
lauCmhzCaNYDxpVRJG5uga0/gNCgdoUf35WdvUmX5rmP/jRiSkcP7Zgj3ErisUO6
C6epBq37SdnApuC2ClHEmx5Mc2M8zwgnX+nyuQyISoBMYJtbv6bU8j+Lo/Zgr7td
54hnX35UevMtWL+b3mBWHze8pNdCE/JjEfnHKvaghX//LcUmkxwMVinFMFy6V19Q
456BGeEZdCWJNKSjjttCPqKIhGdB65dzdrEdtmWCQoTAx1xl/OAltHaLARPyk4X5
EpCmMLuZ12C0h68vKy9HeloGAt2Xjlt6JL1Qh2zjhtVHruOy6l3ulDgc82dI1G5L
uNlWHyqLmVcKHueLG8d48g2YjblgAr9mQ5Q3eu76Nm/B4u5qikznvN1Cjkf+6znD
MqzE571AiOu+yIEp/3NU6H0j7LRdi68gSbFC1D3nFiLSV0C+sSr9ieI0JKpOuM0g
NCa30ZyiSCCrdXl5P9EpuN/uGkn3VlkJFsVVXnTP4S9raZV55xVZgb2bZHY4Zr4A
LuF34AowxjrM5YDQ2PLh9LWDX2it6XOhUwIgWLgI3y59nOtlreqMhmMeXS5zy6Z8
MCxi+NTuEk0//zESiMSoLEW+6P009+F0B8G8h+wMreW5Tupo69vrXWdOLxcCjinW
+FVt7GQP9R2zbmHZhw+sCmRwbRjS8ai2iRvyUbRO5rkAaxECr78CkPQgY6/01Kj7
782ubvW6HizqDCLcoZAf+twGhi3F909W7pPmwl5W9NNT5Mg4uqTus6HuqI5H3hV4
POkf0DQBuXLtWDRS30vteZ/c8N6S/li/G8xPGMc3nfR620SodgOALkpyh2GLO38y
MTxkNky66pHV3n0EL4nzaescyFIfxlzq8iUNWc/Qt+AZ0W6WLVAv0jpvsLzjepZO
mP1q6r8+Wcq+NkDMqHPrxQDtOlaxz/NIGr0MRgwvYwuq8P3sIv0m+EQQUXYTvav3
oP/J/+rqjCZBxbyFqc4kwkKKLUJENovbcxFzo3bewM5bi06mIgPPydXqwLvl3NfB
1wFqcNVHnG7HDTwvI31+Bw==
`pragma protect end_protected
