// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.0std
// ALTERA_TIMESTAMP:Wed Apr 26 13:33:39 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
argBtHG9mAJN+brjpaNP7WKtKFiz1OUPhiTlJWNlBu1ciNeR9Rb0AibMuyOajK2Q
f/gnmPjUzknBGxrDTkLCI3UXeTpYTvagWqwvc10HSphpUyaDZqxvsqm6W/LrfYmg
mSH3Y5qbk7uh1nW8o1nrWvjMAE7CGdb+CDUTTggW5gU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7088)
AqaU8tYZuQwgOLRQC6XDgvAAC6YXK2tn0GZMcipNd/XNI0l9Oe42mbYgzM3jPCmi
fAucet9Hk4Cpi5FPHcs9CJU5ORpr1FbsbhJ/cubpdHZaYsbauqY+iMTR5MmavmLz
SMNiWF7L67ELawsPF0WwlyzViKEJ1uu9RD5xpkKgq1j6Got0wR6yO1K/iMj0uiVD
aUfC5ACDNeOcAR6zvtz50VSxUqPsSbsnqNebcgL8Kp27JfH1OjSFlkIHm+ktNODt
Yb6lQ1uGVY/sWRGLE96nduV4AvAGx6MVddOHD37APU23wxKxbpToJhYVCtelH4fV
Dkekkm1kwAoWoAjbJ8QM1YKvQoirjZRiq2LMxXvfD/e+KxsnRm4b4gJ7tZkNzVy6
MFWZ7uM41f3QVn94n5YXayB7SnT79rH7YYstAGm2IlO0mUEkceMkFjN67jeAPesp
0BUk3FALrXIbA0QLKls9yNQxMTi2F+r8PvO7kxyPWXCZbGtV0/wKLDQOmUzcLEeb
8aYW0tb4t77hrtIiGwYdMpQs0WKOUhBZ2jSBrQGuKr2naL9f1uLMLvHkvh+Huo8x
cleBB0ziCAJBRDNIzEUupuWuJk9YHJHuUqQqQRnHcOwFcEZ4/q+kaRDlm1Mnmp66
BsQuUxnNcRfNo4TznPgrYdhI7MDg/Bq18KlrEdOuBTb6+1rrdnxXBQyL1CuCCLZM
5QMkNq8i4pA+3YAWYrtu+xBhbreNdqb1sC4iU8eTZE094LK2SCCC1XBaHwkOgScD
p+NQzsJYZoEy+OCfciMzj6byi6xzynhoY5dcJu8KlWpgqZ78nriQLAoxu/KixIGP
V1qHURKuKEfJz7uzb915gzfNcYPjYrn4vYnoD4cXiMAx9NOS9iwEPrySGcVvGDuz
G4P2qmFYtZvhom9uDxl1+gj/ntk/G9ULtZ07+55tkiR5rs43fO6sPUdPvEDM/Kzo
+Uj4XEMUh4Ci9dgNynyCjLUTjnaRnPH+BCo4zz2UDrIsJNHCvcZii93J14ztlD5v
poup43vlnKUjaKBIbHVb3XBoVadlhMrm1zMT2Ygq8yRflRkM27Azv/BrSk49MOQj
MdPJGmtLE6kQ0dwRsw9z2gMB2+6sBpg82aon8Zn6yQnSJQ9R5xt6fkLJ4u0s5QSq
Y0jkJw3QmMIS5WKc1lIzHU2J8nzZ3Ak9HgovnokigkBhsdu5Sfa4UBWppCCBFfdC
mcs74bvzOgjkh0aV31wwVgLrMRAP4mGti6B3liZNBu3Myps79Ux28/w/YZhT68i4
cgGslHapkFpzfIsh6zlmukmQ32Bh/Fjg/z+n+ImVXuSDb1hgmYw0prWWjL1lqRWd
Uv0plgAtgjj1A01iDbqZOTOV8zRMYyS/1+f7d5xGR2gb1inQzIR6UKbE6YOX4TW4
EKIT2cuCNewu7QeyVn2ldOUNXAxUyNwm693lnLDTU7hkga7idYLESn++s9MxtuS1
rSMI9OW6tYZEiB0S2s/MdLc8fe05nWFlr4jBB5kIJmAGiliF/6synMvePXRk7tyy
0T4Uix36poEgKQ5BLEj9JTtIL8v/Iae75ah6HLULVprV554obqmQN5fjreso/ubn
ZRfODnu5eJbqy1cRPEsIlolMDnYV/LPYCAcdZkpu5oqwExtw4Xji2veyQkSVsDN0
nBk6g2tJIHb20F0Bh+pd4WTC9dI+z5S7mG+xEmQHxa0z8Jh8I01zUsxvNdjbN2sO
9N0K4pCcDDB/iYhvD9Xp98A28BL4XBIanc4Zl2bWA5HsHaRjfRa8T/+G93BPQcgh
RbsVI6NjAihi4qiNJy54OJTwFt5enRisYCc6pHzhN3/QtgSkHOYVoIq4XruzCBd4
EIkNXGAX+Qr6+GqDp9+xh3EhlYdL1FmjYGQu2fFfuJfSisd1nTJYpFaJlMSGux47
rtnOTQRh0SCXZ6Hk4ehSagUmjM/xh/HmecqIHbEcM/nl9GeqLWzy09x+CtEPU4gc
XA2/2DIBq21sbIURrAIX7lB6pIKt1koQHYXbZ7/xyFbt661hWcGeuvH1anaW6XNn
6nxvnypjjcBHw8j0o9lIizTcWaACsxtk4z22CTQNodIqISiEEhQMXQrCYSGdS3uN
14XOShB77Qkt+DliCh64JGXQ3ifqVO/y8r1cYXprZ1ok98uBvcrLfR36a+SyIpRZ
3NrTzJaM8QVC1bnJTyKC3SXZ1JGQWeh3RU7lYiVoweC0NEtKwGOu9aL+pCJjgHwu
6xpyqm6PdCz1PlwA3RQdrF29C91aIUSV1Lfcmzl2gzy+9wxTU97+NiEDGp2o0tNP
7Q8sdNSlWclWaPiKvC9tA9E6762qPChc43C63VEgRZDYPapj+ppZY+6a4flV1umX
v0MCt3OvFVYKyPCrQsr9998m3uHmy2Cp5FdDZWKhWbvRvNfjzUk5kWPMnQx4fSDb
em5Er0sDsaYhuAi1SM43JtYYQMvMT/KU+703/zP26rkpPiyouPSdLZIgWmSq11T0
qV6iKgDSfSyt2Y8Ivci6nO+KKAsh60i3MPJQXWN664jCEDraXYk6I4weMduE/zwK
lSMRlNwv0v417tiYzzVrQ2AhXr+yncGLi6iq2SR2yy3+VZVoqHOHfgzCusLl2PDf
1cpt0HHqd5oxHVgGFP8ySNodHqagzqVppst/b9/A11I4+9Sic08I0aiidjOMLmV6
fY3P6y47VU5OeU2lEgu2MAGc5rcQNakAyCxTUxITJUC18ST7CtI89YE31V8dwzvt
LdzkI1s2De8H7XLigVhad7skCubsfb2kdBbfgQaRvYdUXRFbsTuFwuTpf31T/0iE
E/8ps1g6SM0NhH9p/dma22Li7bBSUy0+AXHse7f881A975XclDUmhSfbNVyoIb+v
qndfD4Dq8ic/IsaN53Lvf2VTIWLxB+N0uk4UU/uDkC4wLwEcDWJSfIzSvUZv6xWI
JR3xTqRZCd8HenW9RzdhD0j6tr4F9/2BC49/RQ70g+akOLEuEcAw3b+NQKR89AY7
QIicjtlOuiZD8gfacUZGewpaEig+7ysHg6aMyStYKvEVhFX+AF3wLiW+vaEubL8f
xvL1WmwsfHPkChNKvYZe7dlmO8j3LGj/nQ+u2faJD5JQh6mqNrOBWkXIjIopGP1j
KhhpMFVyPyzMwaLAnbTmG8BGuLnKC0xw5VnfCePbFgsUdEtDXPUmOWOms1aspTSt
jZNX8/6qLxf6R+35dj/A1qy01RrayyJOL6xYZGdQ/3tTnwEaLvlpox9ohbX8A1o7
zWVQmoLMzUEvx4LDEyJowzi0Z2ykDIbZKcfvds6EGGTXUFxGWoDP5py78sRaoJr7
dFBE/DZbRIvsPpoaFtKs7ZPxrgARTLqxxDEQf1GiUrCLNIGbx/t1Wv0nArCEDzPm
1sHj/orcFKbWzNr/y/0uTSmFmha9bjqIBjOirQky70Tqru/G0+JQeF3WBiDtWWDI
u1+/EmpEW+43RP4kzWa7X00ig++cf3PZy8J5tb1OOoHR0jvMdyj57WJlAvX2q9tq
kL3JpUNlAkR1b/AFBu+u1nRTgJS/8bXXYoMeihYitvSqJifF+P/MVQ8WD1QZLlKG
rj3FVZ0q1TfXmdNNwoh/PD5WNXGILk+XgvhLbzNCnjyDu0brmpI0B6d/gHLtCUQg
BNK7UM1J3X0oCQ2rTQYJtvav3bDWRdGLVh+bePLlhJJZ3Jfp5pDQ0vR2JK/EbqEh
kTYme6Cb3wJ73KKJN130vYR2WhX4Vn7ZVVjUIZqGZdeWTP40RC3sIDXsRPGUyz3T
heOtw+BKPCn3gvF/D9Ohq93ChAdB3OKHUisxnrRqbgrBIfHReVu5RkVIh0qth207
E0YAswKaQ+hODn1FzhlRKiZUggr7nLcwUMqMY/Pto3//yYkjQGAok2wFUh9Jlyp9
feptCZ0lMPtKGVF8zOgMPmD02ZKMSIX8STibbLLSSeEsHLdENCm8YkuFkNgiofTV
7Hpz7PQWSo4VNqFx4kU8us2HIw4pewpexX5ASI6BlinfSXhpBMYnTDQkJAbsm5F7
xF5rPaDnTxrVb9pZi4LHisym7di3qNLhdwwTPseavExI+Z38oT3EJjVJ77wqKmOL
0mbBM9I8BagquGxCFZv+zfkPSfsWSG4Pma6Eu0wsvrv0QVdAEueZ02U26XqoFecq
40NAD0ECKaLWuDhNrOLYRfb1sxW7E9ZaODgCQmxrn3BurybFLQKw9y0a5R3vg1JL
kM5X1VUitzQTl4d6fwrOsL1oV4lTF1yMV6txf9I+j5noVhVdDcnqSEDi/vdTQGlD
ESwjrsSHwmm/YxIZe/2vBej0ctUdACBXgLAiFLJaR3A8Q45NHS8LcwMep/ljQff/
BCLJx4q5ugrz6Mo13HV6iZHR38VvuJH0kSCYTip14bCnIcnPhahutriL203TU136
fg5MC5GKt94mQBs18B49KERcf3KyGPmxbaSZLof8F8X+UWPho9pkCN1y5xPU2pWt
P374Ck2dmzj1kyi/daMsxHYw/v/jJrGZ1pihfT1sV+wOrg1LYTKtrDkQVQH4eeox
3SPNU6upHq4NZtwx9bUN0UaF0Vqm/8zfGkKhRyUuJXiwuvwNUIl8nKJGW5yomrv+
KYRTU+9Xnxc9ohDmEfY6m4cGowz1kaG2rcRj+86kiVgXzhBpRC9nh48m+ZRhi3YL
y//GTMUuoFJOfKXxKPAMQh+iCfFDkrgurFSV5ZmlhFXqVDHqai8znAo0E5jT7aSs
OwN1iYOE1KoU27TsQEz231N+cXSAvE+FIdSquTf1aPdct2MvyJSlObYF2kb3EllW
4yTrlLUN7Md3vh6iIw0ZzmJfHKezUiCR6jVXfT9FCZcvn+eWJObFnaGI3f1JUwbd
XsuzZwF0d6KDhIm38blMKoNOBdMyt0fMfgNg3REBKHAgHB2abeD/tDkp5fjO8kuq
yR5IpLJLRsyeuTIQjk5MX/CJKK74qxfGr8G3xKUg/Is4eu4ttjDVva+KzCNBwQ5y
nEXSEmGJUqKlOixKsnN7Yazqq5umxuWg0oZ6iUeai3UO/u+ZcCgoRuAjW5Acm4W4
msBOEoyLeiDt4x4RW642j7+440GHVBc1wgQADETsJncH4tDYHVtj0Cdo+eXa7zhy
/+5/JY/z6x8/cuMlN8egyqs5VPpXZa9+Tz0gVZXpvqGmcXQT1coj9+gcMFXngCcE
oJftudjLmaAKR2vokylfN+GW8uQ/PoE/MLP4Bbqcoa4Cg6JV8a70MKUnCHP2GmxB
w5albHXSBoF6VEKLNijTKwEh0SwH1++CUTMdYAncrHfBywzJ1x+mmhoWMSTnAOXe
/4Nrq3bOpemzBbzjthCItGFbPfv3fNQAR/eEsUS9yyzMzo4IE43TuWopIReuVzQe
PGZ5RNbNiYl+xZSzArHaG+QY8kqVBU3v8NxAkEMs/gyENZGdA1sk3c7eEH62bNmK
RqKxN6ch6RhJVc7iR1ZPUssFJgF6YWK/pITBcKRWbI3O4T0mzJtgE+C/DodTI86H
sHkaXtGktOuy/jBnu2XJBuowcLUWRjf9NydmyWHS2R7IVRDjrHwVmgV0voV5pYxn
tt/qhXDMnmRCnSNdMbudtgqFn1rbuzwOFyy/kvQ5tpELJNNzrcbkHmLJCNnbYipf
SVrsZ/uf2X7j9xM+Iq5ahgjjZV0C5c6LM1xx5lZMDTsoX8q6NYpDSB0b/+87Y/z1
wEzObOr8Ek9f3OSgUDloplD0Fku+hfdrNBEiiMA7+lFu1aAV9Sr1rwhSKjVKsTtH
HuAEPFNzYQn5nHBO37t4x1h/0LH8EV+CZ966/n93gELXR8e32yOIvVMobCU3KX1b
0dnnEo5GvUde6KrGYfOn8EjnPB8j6pAoP06BLGWJIDQWCP0wKkfaDh49h9yR6YMu
kmeetr5Z2OBWxxocBH1tyr8pHla3XE1uGaGLT7j83KO0DHtJNyEaCxX+qfJFweTF
f3+GjqhNgD/i8yAWNBDQaO/wWniUi40TpKn43MrfdQ5Hco5HMJVvPLUIEtmILfza
IIjru3JmoBjJQedyqbBBIsPe2o2JnvrMooA688qQdYqnzMFdHOCd1j0prOF+MgEt
5X4yHcXOYNz4xof85eAGZZCykKmL+zP1FVET8S1dt9fkrfMuDIz/FEplhxsW3+Su
A6efShWKGgyk4C2X4l13j3jHdm4T7spKVBPUGvQ+gLZMklrFHn7eQ3iMQVMYhgpA
IctSol1X364LZ9fhW7cqjtG7nIf71u18C1uJEJtOnLWPOtA5PT2W0lVPNLtdLV3k
6JkyzHYoDs1wzXHc22VtOH4BjCWBdJCnpSAVC3m7DfCTBstLrIMn5LtsM6qH3wJX
YIYXaX2VU1wN5DkWL42ZAs6wO5/hkN/+OOuXG3JbKaR2uVhZ0RUrUK08T1L0f4ym
LJWx03BNqWNfu1BVBywg5jLnLBgza0L8/Bb5dt4xo7cbwHsLpFtRwoCp3/UI4LBv
YyaN+vMM8FvkOLm64OEwefPeRuyfc7PbGG5rKrt3jfzuNTe+y/Z/xyeWPbR1WhSx
BqISoo8vkhyXViIFbDal54lxVGWVIK+f3UWLApbqAZlnBJtTINd4voBLDZ/MguVj
VSbeF6hpUDzwNYxW/ZXLKK/fyGDaHHyitDWOA8rOytCmVQ0QKS14zG2MpU8BfXgm
kMq2x17e0nod1z2tOLf8QyjwbEQZuqnAK4HYNI6EouRG+QOrTz676j1NZ+BSX375
v7GzxlOVUp9klGmrCd3jXXofBx8rqXVftD8Opm5tZoEgzlL2xtNEaommGIvvhlk3
kieEV2Iyu/TVBHjWFITNxvYoMF1Jv9aS35ii6ocCc4bGmIiBtGQtVJlvy6rtJvXf
iDzsM3JqgbLglRuCPvFo90EQq3hiC44ZrbiCgGtzzf3bNpHWDTN8jHMS2GCg/BkL
OZ78hIvkYyPIHoc0KVDI0UF1/YgafPSBiTND6u+vxG56zq8yPRQn9TrPmnphG5Ji
IYpQvoVs1CI9fVZkuxvLtP5BeOPRQy1jDGd4G0JVf29AsnhRT8VIS9aiMC9hlYcb
GKReglhaH2Wx6HJh8iSikdsanqoIOxRAH5xzTHlGEVmlTsaRtnhC7vsWoXzJsYFx
9C344/EN0gRNp6PcO1YAmXqkdSHF9pOqVvU9ZnP1BJ7zU3q8gl7BiwQ7JyozsvG/
z6kT9LI56OJspS92nudwKNLErqsMa7Sl85Nqwci9pYrT5HvJjYcaBN4QO9DiLxPv
fpaIZ1ZPy+Sz8uGnYgE1vmV+vkobzslvd19qfnnYpMn6qgPcTS2zKZcbWttV20pm
dofxbrJLByTi93XiMTn4KDTKJl6Ofm1whdh/whP12f80wyD0z09qLu7j1a0YcV0b
JZeO+FvU1zSuiIvxMnCgCdzu64DzaBfO6IKG0Dp0ioAxUHntdneoMMdY4NxteTzL
zySeNteOuYwdTQEPmqDvaYIfO8LdS5khR6Osr6BSRpUfd5OstXMOOPBu1B5LRZBJ
fSypBGsjF3NCf7f9DeJcotS/icSQrfBViokYbYneyThBR4xtphFLAYtMouOWrb1K
nDGqZTOPEaVxJuBpEUXUz0N9AwImPi/w98AlPHartZKhe3VgA4MlEFehVvoACQhI
10b/HrpKI183XeWdXb086ICt1C48o8msZJL4gQxW2C79ixGVn3rq0Lhcxchi8skE
yNF4xygeC6DzIgdZYAQplnZVrnWRUeRze/HEOyh0Twv+ooavyiedlXa4N+6MetEg
DMynX/VjMQb2KwVO33LNFUcO5B+GM2ubYvnCi75JXFaxgarQ/BDe+w6vUjBrNIsD
JuelpjNtvMBf9z9IAKbfMJsBkTDzfbpUTeSiqiTah4cHZAmx2OqN20fppbA5LNwW
zlpFMT10/IJPKN7bs1QAvq6Qz23Pbmfe0RUXFAd2R7OSoUoLU5F69YKFmARs0xPL
jDWaHkHC7r56YaOqdakuam4zHw9mym1d/zD6ASFU3h8zCwC6VEDL3wSGm9Fnfdan
aoFU0KkUk+NXdFqE1Ek4+NKULhnuZPClIdtI1XCsN167sR2m3UC01bG8RpJFpjtP
ttBDXL0rYQZXyhITGaUJqTTjBH+fyTzhZPlPIDsBjThnX1g36H27GWoS2AwMYS6M
El+8cA79ThuGYl+4B5Uk5nPS5q5pBtIDlvAxFszBkgFUGvs8eQeNL9AB0tUZvR7x
oWuUhYpjNcyylvTlM/Hc4Uc9Ow4ysArOlL7NIxkDTcpP4tJ7bhjfofuE39wKFqY7
ATKToy4SzlV4ZnWC5rGo6ssbnkE39mA0r7PBrS8hF1aI6mWjFb2ojg0+X8xLtsPa
OxGLv+mgiZ+QqFU45PHGo08+iY7h5ZoL6qbAlwQgMGG4HvmQDN3ganj23G1Uoncw
/KKbHulel4lC70uxXdnUnqwHm/OBdDaGhvyGSKJPIeD2XXZJ2UtrM56O0T8+WDrJ
UeOU8GeejuWExApegE7kGR4HrPWMAM4E0cqC1MUujwfrQhP3NJtv7BUZO/mamZ79
0lzFawbaKBvf+t7KCAjSuTt/pYqta9yYmcWrnkgcJUFW2yeN39YgcjDRPvL8giFJ
nAdyJuNPUR44MVjBckXI1CTucoGhin/+duy5vOGll/YXpoE5BNY8lyON6WebUT9T
x5Mil4d4KNV3LGQYoZAL2RvaMaeKmuqxe8F7CqBWAyjO5f8HJ4F1cn0pw0gF+BIW
EskRty9rXMYdKq/h5g0b1hcMAcAkD53/nbuCvF2ZG3awaSe7YhYyPCorJeSJhFgF
1dCUXs/d0afxMRi8m2qB+FdaHaIvnnC9Urk2ZJIoxou455LcT8gL3VKXr+tUNSAw
AuJhyP4wB+1BgxOIMOPKciixKw7PghmlM+WKYfm6T0sLdF/q32vkLU6Pi9grsmd9
APGdlGEfpYJEBCCU5wODrQ6YqIQRTDycKRisfhQDcdTGaOhE5ORiefBlVu4YZIfv
W1snMXQC9+Si2fFjjftLDij3LLh70wI6wUqnFc+BoCvBBK0HV6WfeG3TAvDYJJ6I
2vrh8iBI+1HrAl5qvvfsdN21iO27V0yRJ3x/kw7kC97/L8MWilezIsxgV+/saVzA
861T5fOFNm886cEnJLUIktVz7bkuqmZnfmhv2rFyRFD6YfDiv8I408Trgze1l+UL
1u+G9SBt9ipHEeOz84TFQW6cngHefCUbma2sb7/B7MKWVR5ibdR+PL9og6CyizZQ
Repw/SBGt34MPwp223K3YuHBepdIy8gIprXkmAMn5YVMaEpO+0KFoXYu2eCRlVem
bKcl+Bvvji+8F6zOqQwwnUgpSla/o6ZuYImOYUgRcjO9sUGGxyFgr1gMA8eSOREM
S3KdCSGDs9tGl42Xka3c630YmVtUnzhk0ENt4vQ2OvcO1gBGZYPKvZ0i7+uZKN/i
gMCmIzGowD7YD4mQKF89KF1uLiY27dKHWj5+SgBAd1k=
`pragma protect end_protected
