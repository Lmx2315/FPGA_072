// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:37:06 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
e7daM9gWhbGiy4huoea59pg1o2flomzUxEdbRESwejWAAQ460ld1eLKRo3At/QlM
AQdjV6YrA2y3WUmXsqyiD6nZG5Egkpr8BKZQqN6gSek5RKQ0ETzE6XTWj5WYVTfD
FZD4bu7Q23lYQ9o7hOTr9JpAPQNsy7i4358M2OG5CQc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9088)
GN++rvWLbtl6/qZoZyPfoI9EmQWl/ovVgrH17Um4Pah1b/m0MggMEQXLg3g7O+k0
Jr+mSOyIM56eDHxU2RhIrJYHpg6XNEnqBby35m5fs1fCDMuSHQvy5NbblKplNc5z
rj2EFJIw0kYWcf+CRkuHGs9Y6d/gOkUcOSI50FCENgADREZEq4Rk1cHidOY19gRT
r2tuPxpSS4vRi5jBjkxso7gArR+PG6wQFAOzDs105rRJjXXB3Sn4GEdz33YXYbTo
3WUuzaBOknhQXNEEc3iByYXmlpS1ojOGnLFF0nePndeLaYHlhFvuHYS/mdh12aHU
Ciq4BBzY6N+9dPIEp0g3wXdgsDuYcvk8ZuMufq56uClUty1xyS4rK6/EuYcxpCjm
t3NWtXeuij48bzLVUeP5/T1jUIo46JpI+3onzgVmwNCEB+YXUUnbTPZNNWriBCr0
Ckr3FEXKX4Gr6fA/G/N1r2HVwKcSx3INZSj+O03ZpSpqQH5VjDUMTol4J1os1pp2
c5F9FsD1SYOliMArGZE6WozvdM6icWfRvSh6b6c7bzQT+cT0tL4r19few/ygquaK
xvkXz+r2F8L/DfG6CS6f94jTHLrdCqieG8gRdriYyiCI+HycrrJI8fkagCM0p9LC
juDzvwG6M+HyE7tzw1aNfEgBfZKm1htEBL6ltOlR5E4xyNuYck1lieYMple59FsU
0sxxdpuuF9Hg/k5j/1UTdinqPhijdUa0TJM2VsyK0SraNHLSHE4sj8yuq3+1J4DL
Cd8AQCaGh5YMajG329Yj1X82G7QOopBMzlcjh3ZC3I3jQk/2g/8Cbi4LtvRZuW4W
DxChzs34RmtoBDliHXb0xBlsIqIyQRndKtvkFjwHhk1xfv6dAtCABli9rYdVzAuv
ujsp/330Z8X+iSHl47bV35idEvvXBb+46DptxHKuwQS2c6iyEzmtlqpEnNDQQR/X
2tyz+dTU6U6fBcHJDe5IsWJIPh+IJbwqmf3JOtQSGEGdIWWskLjDUCsGkAqp3F43
TPQ956xOfDW23avlcHbB7mBbaK8xwwRvVP1Ah01o6KsCb+XKtvT2RuXY2f4Eb/nR
yAZNzwnENGymJRZywoaW1nx6w+zMbp9mV0UYpYLEaMevilYB3h8MXkf74thUJFM5
Qhxa2uwVgmdwS5f3U/j5gfiR3SktUeBj/DB/jcdRYZIXGpij+01Sx083+74xft8f
ITCOmMHrbX91G6SSTHxwKiMEKT0+p5OVmCMrnYv8XO00m+/u0bk8f2DkGJT4Tmz1
kyDVyjd9uK/5TjpXmZ2SEtVzWReSJf8qEOwtpFBkAAD2ZQftNhxWOTny2hZMaSFX
m8sXxuRjjYAbPr5oVyI8YGXqtgzcavDJxwIA5zMLs8xhJ06Hl7SVStuZCFillFWE
fj9aFJ+EK4CMALNKyUzDC7DyP8mjxf4mdRY98GESvrKRc8qqjm7hDUfXsJMVWj8/
nn0CVr0kyrD8xUuSLs/ZiiKODUKQVFXkvJzps/1MuUgYHZTduIjkzM2/S5u1XJH8
HR5fEheqzPxHqLTeaXQoMnwEP+xeN4L228lBOzuXV+1L3Yg5RBacVTEAXf+K7YNS
Gy3pSh/EsYsR4b78tdL/1lPbLVHZHhct+WRmDAJn8j0R9psIthqaio5g6pHLPBSu
zTHLAwOe+oSjPMg08aWnSvebWwdVA2fyMvpby5K2pJC2HIuRPd97wkmbo24ZjC/U
bVeV1aX7lxG9X7cIG7RH5o2b8U+31JcnGdRMG5JG3efPFfcORKA+dBSBXVm2bOSg
xind6SipynWpmC8GaGeYFhdemjuT8OzxLVN9i0RKaO6L2lmBuNXJYo43i1KVm1MD
LRXAXCAUDBwrOtGujNoNJmInxS2CfkMCOhRHI/Lge8qf6PG8EgRZ6LqH6tjwywWC
Ai9nQco3Nz4rsJeDxIVR1Nt9sH8+uvCN8CtEIzr1h4eYdgkSSJh9LR/Q+/PTd0VL
qcY8U/gyo+A+EdCySCUzzWFTLa3KPUVP9JPrr94MK1tzuNDR/lQr5/Jvl5LWHCVR
D2RDULbQ9SZT1jEhPolXrZShQFA8uArP/SUs2sijEkU+sXB4/6OGyEzRFqPcEegX
Vg4I+ECro38Qcsjpx+vwsJ7egCaAA09fO17qaBw4vvQQHcFg6SnkAxgsXYqDEDeB
4GFCYcL4u9bcKFCMNsBoOhNTkVgxrMaPwGVGrBuiLfl+DoG3mRUXRelZjHmZcgyY
fpapzr8wXIUcbsRuMTs9PrvD2HjhNxcqV8ZgWBZjOgiE0oRztQjc2dey47LX3TC9
veFuDTRv5ny5OqszdTXDZnt8pgtyKzQvkRmVSETF1fQkUODnSw/MgfXXi52imv3W
iPdaXmxQ0PJfvm7CQkRtBo4iPhEzQdzn1URetXZA62p1B4vxcSaceZ4v0AYpdVfa
9oAOVXvuumFO+L+WIU+d1iyc8Q8zbjRsHvxvNHzZ14KrEDrFADsioU+rnZZW5CQ6
KzXepPNCR2Xy8Nrds+riPowwSXsAhUPRhnvibX4PnZLtLjP1LSlD3qWmdRWHfTe+
kqVTYjhfUqqXpyRLQtDdeug67074d5Ai3OsrAWyB3SozhqI8z23TrZ8dm7H5Npv8
Pj3KF+HuLUXXScrJ+GqEcBGU5jSvG3f8MQ0NQ/TxnrxY+t/rAW045gd91McKvLzm
xqPAEek+ykvm7ao4gIAksRo1OACuDqcra8CRzdCvJcBUs8g1Xi7VsaVquJYezwaw
LsfI+H0ympG6q3+yKvxG5R4tTMPsS/3F6gR85OgupGS+H8mX+9lvd4KEfjvE26Gc
W520XOmTB3zi+9J3Bo9p7+mqWjyfiBFlf9/du0hAThDAx+ssFSj3D5rjWQOjcuMm
oRrPo15qZ55ZY/RscpHwWFJtm9wv6LiNvkGzSSJtfWzsxunM8itbhOCG3eQbJZsQ
4DsOcKtBcc8+pPH10IPAg9crjTB448HPZZEPsLSh0s+2jV+WftnONNSHMZ5kg76n
m4+dn9l08gQQlZxNGkJaw//wnsXDtsQnseH3d7ScKyEQJNs8h5MMuOhuvAIDruv6
wP1B8odwPJSu6bEyQubgWlJ7wbSzfohEEl0pFRB8jKZ/QM9x64JMQL9cV67Z2YVQ
ke8jkZlYyG+iU81SnEADG7QGUBQzss7N88I4y3UGB0xvN7Py323rTefHngJcW7tC
ZeC/WcP7WVPe4ovCsUnIHnPTIs+FQQ5Dz8aVQshnCrb+whWHXnZzsuymTxoiTmWd
nzWmnVIf9ABZxHQZnVMB5QLqRamp4v2/+QKT7ywwYbsxzuvul1eX7mzTBwFhOHNV
ln8NugwfKx7S5l1//PlKEW8CK/TkORGSvZ3tVFEY3HSyv4MBqTzH59+2LRm1O4Tj
kWEp7qY0CE75ENPlpWZRHh46SuZakjpGrbfUqthLXIIIFUIlV/d6u7l8W+vP+DHd
DvfuqdHW58fBQ5dDvfblYNtYqQrDTklOGyf0ruv2loNYLl890DYrbQ3geTDQW3rP
9UyY6xij7BjHciFlc+fJGyhIqZuCmByxVC0QHlsACK2PboKNjwq4nBmoLG/y5gSn
hz3tZLwTE8qdIT4uogSwitnCJxZSzNZ/dYUaGgP4UTADMxJkf8QoV1a2/YPNgqol
HzvebvHTbuRpI4dE1mgG1/JT/juIFQ8IW6BJUwvtejda3EpE+4ilOPTKK3/bbf9t
vXJPshnnD3Z5ziM1XF2go6kU7QD5JWBp2AeaWeAOykO8VV2t6nXI8gkOgJWiOiM6
5AYeQNM/WHr8uKtdRrcGcXPI/qSdoX9R0b2MjpizCeXnBOPmeDglxMd5P17lG6Yt
4Naz070xfKN86SSap63B3ABuOQ33kkKf+Hdb2yNGVbWpRleEmpJ199+VkYAigh2R
Bkl73Eh3MDg91jk+OF77YYnNxZaoCv7lKmrJYCBssgUS+tPK65nqYDZNc7Ii20t+
cjN3mQZI54tsql4sm0MmdiRrXnt+nQGh/M9imaP9e61r53O159kKMRd8FnELhKNP
qwpXzR8jpjODnSvTvnUMRG99F2CTzSuk72Gq/jlwGWDjqChIW2pQxrnrzyuwtF2x
5WEHDR3+ueoXxFQQL0a35SLXs0j2PDCsou7fTBAXLbS1lWdVOmkAYhYbZ6L+X0aG
pEBRLEDHLk2V0yF72LpwD8GRSjZqbwGey1ZGIkKHVQXAeOntzGP1hDjo4NZrmbmw
zGynIa4u+OIGOXjccpoW5sza8i7V9pfa19yEuGDu3k636isSK00cQuJX5rQs5KTd
ck9nWBWZ5vQ7W5DGcNiNpafwDdCwlRvtWSOyE8GfTBrSYF+2kvA5boEEeOO8WWXD
Xau6CVkDQ+5MLq8vbttGoWfgX9s5PYRmWSi7z8cXKxvdTH68vXMBKY2c2TtNpFxr
sW7Mgibsi9WXEdvnRIFWW2sclZiMMhpWkcrb8z0zIvfrNYOkqEZkdC8Wi9B90I7T
pPAOXD7KWjOfUN+e/3xRoNOZS+cHqtlpJq2tF8ILV9Be1JHHl9kXEZU6KLbQgxse
3gfVnC1/B0NoYOYgsmIvtCWg3ITOqoLxaChWCb3ZfexqwxGGNyfbVycDSROV2fGV
GQziAqZCd8UnAM0OMsMJ55jSx1MZU2GMF/VNe7QaWnkULBYA61bJFG18QtlJO27s
uthZCyVoyCiZEHurX9yADpPyUzAiyuwShlUS4Pvx89OGefvoK24AJTNkT5VQ1hFx
6tflxV2PtBSYfqEvxfRRfDD3IO4W0oJB0FdbHzdr2MFoA1KRDJvhSgfYBLmwfT2d
ZQZeUZcRM/1UmaUxRlYMhWaZvLn/mUa09hQvpEWqlU+wX/1tBPJc/sFue4ZQ0Mm5
NqrDewRN7ItVWCdfCQkzejtl93ZwuBhObUc9UTBB4eYyKHrP/Ip9M41Pr7TGdjgJ
uIafyYexoetetlw3PxNBGbsywyDRU3PpkAsR8rirc2yNxCkrfxKyrQtdaMVYPS72
9P3zEVNOp6nwh1okoonc9b1bXtJjLTFAWi7h9KfwPSAo1bsHdCJSopnc5UFnDEEB
DfoAiVri/B/ko4rgJw7IQhqxQwtwt5JfLCSwVUIsRbn/4+a/2PZ4L62XEfCxtXfm
0LjMDDPP3AxSihtqIPvjmLxcPKzmUzA3lX2zq8UkIe6oKachXhSynapU1HyWbd1a
2a3zFdt1lbFd/AylEnO6WA78uOiILAXWDTStMBlqLqI3YKXBwEAaPkmPKkb/C0XU
rm35FZMf88ExOlqypAr0o8qiH1Xm9vhhY1hcPXODThUK/GgeOOufq6iUnRsHtGX2
Dw+3dJPy4uHEH3uMfPhWxx3FWeBuDuOOFbLwC4SWb74g57cM0b64Z+h4iwE/1XOH
bUjplkF9ZAiO57IMWXXe0cfUiOnwFMihDD/VUD9ObO8w3g8s9xTcpqHVMFzkMgYx
shK+okor5R7NY6kLZsEDojJSMDvgj0oLyYrMrm9Wp0TfmP3EJU7mX0L6eS8tPkJv
DahH/EYdrmqkWSg4yVzyqFQTNl+s5NHmojei2JtwU2my8mk9q+BjkI0w5+IaC3a4
FzGIJhRmHKYkUKSLM4d9ALf69S4I/AmcsYW9a+QaiY1Q+YQNryxP1UTMFL0Ix0bB
Ly4PS/sT83mVLFGMv7uv65qnZlOZ66nOSPTpvNx6CMA9txFfTs0yGwqV5ES4xQaE
k6OjE0i3CZvNxp1V+gO8KALSwa6sctrSFl0vfUYiY7wrqSBole+f0lUFTzEdRvKj
229RW6EcFifcaNogKAXU5hGv4aRnXMch8YAkUP/mkaAX+SNmR07dVw86rDVmStbK
5rec0perq/NNCjqNlCay39RZbs0fvYrEKF4W3QY+Ip2Ic7ynH9lu3NQOHxsLHe2G
fwnVLV20Ved1pAozwsi5/uhquWA7FESMcxgRcRtODsJFhb2qeXWH9T1UupyenjNj
pydqVLVQAyppud2my/ic97lRO7KjkxdetFtqhumjtcPhzCvdHYw6VNeQQ/Brqdng
QtAdQgyYJvko4L4jrv/4nfz84Qf1NokwDJP+DZ+iT8ze6DaP27wvuLC5NjQt5ARQ
SoDwQltSMGhzc4FKXrDUit0vxsag7Rn9nBHFvzDc8jUiweTT1OCpM0W+mDfthfFQ
vFBa+wntKtcSnvKpOtwB9tWdfE310hDY3uNkeBW2DqJ2Vj+xYnfx87PHGUb2xRl4
QSthYHlqqV62hv+ReY/nKTMV0QKq9OCmeIagVk9+XEIXKgZzr3YwW6XLtYwu2EpT
o6BWNN0/HpDor4Ma442OkxXS3HtAjLh37M9TRs5i5A2vtp1k/Z2W7bsru1FLB4mT
LDG7h4kg5/y3xqfo0kuvja/RgYs23jfXFxG7pfCqfVEEFh26VPvHaDrYVgWJsTMl
pZ8QKEywjJRmY884iypg0JUwbMa/oIpLc+G7ikEipw8Do6EYlIP4u8TKhM7qdJEd
K6ymv2i+CsTleElJuIFC4Ej9WDFcoke3EgnR9hxGAdRGF8I29CNO8f5rVSGbGhe7
OzmEBe2L10SGnHoJwSWoKOyUzfgFfdCA9eKXpkH4hGccSk4kHkYRCsrlOvIgXkxj
BlNYdHSc3+S4gSzBa/OG4HsHoJa8GO1BgA7pPsZBVxeLDXeQI8Vl76TWAioQJJJk
ctQSn/rm0kgiZOdBcFwiOl116V3vkKbze6HSt0Cj8h+A5VlDTevi1xuO9yvOcDHt
lnVWUElPEUWXs65auahSXI5YZmm69glvyuJmE/9jGaJbgfcZZ7Lmz+a8G1JXjYkl
0zOMf6oWbaLX9QocvigPKRK6y5eB4s3Xb8i6p9CBM4UZ2NwW0GOLmAWqLpNFhZ+e
oGy0IyP9lQQ5UqAFwEHOyBTS7oLIN2xopW8g3XfG3nwPkDLaVaWYEQIJWrLR+IeH
OG4zX6yEjkWbols009eqoJOxJeF5urs9GO7UfSRyKEiqxUKR6dd5/jGJftFvRXsn
JJJdIVnWWQSjjMwtPqzmCVtJDrCxMCFyLv5bydkPpbYUoCZix8PE9gExWAZimg9o
t9i7/fDZRvubkmiMBFH/i9L7I0Z8agp1BIkaKs7nZH1gDrW406wKO2+GbtRFku2a
druTR+O5hOM8bpxaCjFRaRAsTt/wI7M1uzYtsT7S1R3Lh6KRwq4VjYNv0m9a8bu3
taDZucrV3M0q5L+YEdPWEPMgF85TPHeev+v2u2BeSgd6yGQOZQRDWRHxsw7nbM8/
0DyLgvm+z5YY5oZ6YW2XfWJlCsmh9EqdtAF2eHUEaYZvk93+8oKYHEahzQ394Qmt
riGeZ2l1ZxCjjb8uW9HghorFkkk2dSGCStw+YLP+kk4i/iJuE+m0FZ3IJy4CO8yT
yla2dnXRzTg/N4QsnZCRIeebPS5T8xw4RaF1JD7vJN8IQe7J70170sXVa+AUOTTA
eIiSKuP1P/lomIZ8nP2soCVbE02vUGQvL4rs1QOcdv6Kf4RofOE0/NuPST1qMR0I
DytWYalOAkv+HLIFkPVcGFw8oOZ0fN9lQIGpfJl00htcgMwQ4To1yMcUm+h7GbBY
3uTywMo5AIPji5ZeyR+DBCVlI1mNkBwRciMvFqsZoH9ASkA41CrXcKAxEdNYUDyP
+HfNmDphz2xh+clurtAhFGMzGThkjlmviIOHv1IpruiPsIEzoI53MxnnT66T9DsN
Gy1w8KEQ7+vazZbRkJUk5zAl/x97R9Jxsqm9ge1ErX4QA8IyPdBjRVgryrEpkiQv
l2kek5IWKGXZdPSLE6sWLfkvUZ3Mw5JY0QdbHBZpJF9owr1DJtquDBfVOsj7Hk1u
Mto/j4WUpiYREc5gKc6SUz9k3HkAC5Oqu2rj8bCKUg9wb1CWeH2aICaP+WZAAOVw
KIPnqPrxTuJkA2JFb4YboGXR3WZ5cnmKUk8cWnsgVwSvUQ/MmvVgnU6IA4EkJU0e
RoElWO7iJZ8m3cNQeSuy1syD4L4Wwy9/Jj1bp3R8LWyw6Ep+/yHWOkIieH3JjDc0
4vXrF+gPUNTX5KB/T3mdRtg1KB6Kl8hazVAgUHeVo3/+wnv+eWN6STSBmEMT6rGj
Vh+7kJp+KLk9DSpfbEPpDCDkmhE2nsodLpr8DSsmHv2Nkv3LEOm4/aQl78IKqGUX
Nz2OPLXmkdRUhIpXO80nnHJCko9cVrhuE6P+w+pxDV+Qpdba4yF9hDF5ZigiTMuL
WKVuE+L1cLwctdAYA3VA4ZX5CAFZn6qebsjsoml3SjkAZvCRjMeEyP8FsTYHz4jR
3AI38EGWjLJtwt00arkNrKawz3xwjZpr5zH+z7FenRLAW+Z3MDrFMpy2rlWX/9C0
u/uks/TTs94WofVrX0KWtXd6iTcGKhFr1lEgEvXPE758ufXu06fUR065EljYsUvm
CnU276+ctWmXLsKkZ1wq0RsYSGPOIMkyrMegF43Yy5VMK4xDaFVbXiFMvLJxerlJ
FRpPqeY51CfvGqpv72xKrdy7zVgLoHPK4GfztRP0DX0ijL1TNowVIKtrR51UiX5A
1LwSF0pJWP/MZs2ps7ABRoA3CMq4T/71iiGtJLNf9HLXqG4dsr7PvtHEQwftn+6S
2VKkumKAsh4nzAN9LfAAHUlIaVE5BK6L2AaPvZYxFuzvRxtomfZ7aAQzurJaWHnZ
mVxW7kbSqkfinJltqpKd7FlcTafF4p3D5u30D8aXGiDI0TAMYtQzVWs9KhKl8egp
YL78Rf8j2OCv8KtqDo6PVEsjGguXQWoCHl6zJ5Hj7WnpaxqCz7V6KtLWLxleDsdF
5rPe1IL5ZiAha+fYtcQ+HhIRvWnKU9/JjP+kS85YpIyVzPjZcJKWovH/LC/9AOMM
uID8JuqLbopiI0B3JGy5UT0u7Hq4ixY+vXynwEqb7ltecofiJN1byZq+YxM06grf
BKZxtoqj3xolHsJ/YfgG1+1AavoQooz5fU2AkgOSlmca+jLy4+7fUd73jG7lgSdD
whCUGvv57RbLGzmmar7CNmb8X2I9GbkOBqHN+135V92K0Yc7IgioEzCQD8DLu+DZ
BMAlkrgJTzwQkvrDnx0qqO2zjqjQq8MVaAu1CfyZ6EUjKJsyYNziH6rM3PtLEki2
wE+bP34XpEbp9R4NypGSS53IU9u3u+9huHAO+8HK/c/BTIlPjZpZDfLv7iM/hXbY
4+4ujQhp+wTNuj2KJp/JqgWJIoaPwTZhPCuvzebH3UcjrDyUz0I8ganchYoetUge
oz2xaIArac52sO+mmWDLgxAzav1dy7r6Nwx81svqhfpH4qb0Wc00zsD/SteeTRzW
3n8f80Pp9JEGAPW4NtTiLYfHLH2PvgMtFAWEdjjGHEQS2Q4mBoIExjKfbfiPzaTy
gbNTXqUG7htkQ/N6mO9TNj44LoVMf2SDWn4WbIplbKwOVw1BI5p9jWuVhlfzDhSE
vbK8GjU6NEzK9IDolcirdhW9rAlVlzRqmvuEq52o+EnrTHGgyz/o9uH/dvxmIe6y
lucgTfp0MODEtD/EmkHke2aVTrFqm+BW+TjIIg9FgnKEtdfw0I6T4wT8lHy5fCF7
Z/SumcHLDG7bHZhQlKN9+tpi/ibAkA5OHixGZY4qfB5BiGaavHxlENfMMdws6oRE
9ctcQoCYvrDXZavV6531RzRsyuVMmmum8tTgjaMZhYSCL36SB8LpDQwfW6VuH1Oz
2Rfhg6al8Df38aCXIhceOL1+HlJlczA0Rz+eD2CkAMfinfTnkFmLTLmp01KWZ7pt
OI6L7rhOMisR7lStDUfPHV1+lJ318ysZt76XqQzL7b4UdpWFT8cqxa8nkUAhePIF
fwDRh/fNPKunGFPeIfkwS8vcE8+JeB0KpBL/MIep8/3qWyotJpVKSqhu1Z3cESoZ
464fmCI706pU7zMiIaW58HMTTXE/7gxJVA7tmNZoexenTHQL4bndd6/iLTe88jHh
0Tl5TaT23M/Dcw/fmSpAoYhIBEOaOqlvXNiFzmRepmZfCUuqagBhFf0TIV5V6KCy
OQbvxx9qamhHZ2CfZ0oqz/8qmsFG5G05aKJ2WjxzftMKTjoIeAbk1f2r5sRl/4i6
qeTsq4iBWwi+ZUto3H1+GZJ5AIL9DfhUaMtnZate6OiIqg6N+Rdl9vWqB0d+BDPV
u+7q3VkNy6YxreF3QGaRtHs+F9KjXcv4vDUkKXfBXgP87pjqWaDAzcHN/lbSQWvY
IkjUrBlkKZOchUPAE/kH0YiqTrJQZLR5Y0saSnrwjMDMenrDHh01qqImignrtcyk
TEzcXd/Ox+2eyCBJ09bOXetoIfzC7ruxgxHdL5RNxmAkvsHQCgGFiEQ0KrJ4xOPf
1sgbcTBxJgN3nko5ov4D5Nn1VtEna7ltDbXY6LU7LaY9jIR8OHfix1gTn6WxSzwi
uFMfmnfpmegqvY4bAf2aRo8asm9MjXNPfGGf+EImnwRhyULPcpdR1cxvr0JdWy1q
MEubhWSRZsb3pi8d1jcuIvjgt1vH3dQKXY3UHj/lXCKX6JzgyHEOsc5PyBpsKFsy
HUWcw4o8s2tcR3bSceXn85uUF1ChvK8PvtV2gM5U3eZRuPwP46I7QGdHMPne2Ttb
TDT7QBrLmuf9rrkh5vJ/IBM2svCB8D35lrqaXNNX9ZE61HWcsdgqpcCG8kt6aceC
My4Nec/cLBPsXdryZzJOKRliWOa9wLoEi+imWX+dF/tY1X27p/F3usZkn+bexpXj
N0eNdgEaxbhbQS2np24jBe4CZFc0P+HV/8CZHmi3QK5BGTYHitQcDAgtL394slT8
gfbthMDansyvkPaB69artf2UZcgz16CqPLQ2u+sMnb+K6FHez2WRckgMvTOPuYNT
LRJpYd8i1VZgXAq+HW5YuMu9+0qFYZoNhORFXMduN88K8+aDrvYTjBGCgMyXV6A+
vbLM8xV6DajV0Jubboibepfh8f9G7MYaKKbvn/PKlfaSiua1LSi7zSfXf0NH9z9C
uJ0ATouBRxEPSg3In/8QZfiVXIkhLGmrE+ekefhYLNBGTqY1ZawXQLEivutChpAX
v+r+ovRyqW+SozGf0UcOCojX5Hxln9k61OOVpIFD0VWnLGpNNZn1392xxjUVXybE
upOllrfHlaBd57/bOCRWBekYbXsI5ttzplSM5l2UTa59qvB0bJjI7jdEM3iwlEHb
jTUQ+gvtc/1Wanih4LY+g1UPlVs0WuxQeD0tLu4NSgSznK9dfNv0wSqPi70mefCz
3P8J99K7dxXiwPs/Rvj1BRaK96Ek6wxzKdYLp3V4VMracB0y5JXN7+hQ0QM3mbs6
nnMDYWXgH9uuNjhpU2FRBxXJzxfmZUhQzQNn+YDPA7/Zg63mI/hD2YaX4H7he5jg
eRCacIGXzA5KudJ+heHvRll6a6kyxTdrQf/41cKNIDNs/+nMIS1AwBquCcTJj3NS
PYPoC17EPwHK/JHGcxJp95HzJ2xe4hbmFsakR+6EJwLKfOSJwcTSjFrQZkVoIEi2
1QYW5IkhogYGDHn/NrqQ+L3B5UBZfAwf8RIPmPfgDSa4VxiPTvpAffMeSn0IO1dF
vybT0QJhnVQi71M1VrsiLauT+H3xPjF5d8uAfKx4vl30tbG3zIXO5uwrjGD0tgbZ
+tBY6u3b5q2qrxouUhlc3r5IpnLLaxC9cNdOF6tkZL77CZNH/mjJt93O/ukoZM2b
tBceOAdYUvn6ott8NydAZrgz/E5qEmJM0G2pMo/lwciSxus6J3/aI6DbU7aEwv/a
0e6xHoWdqZQEwjYKJEo3AIOvlyG7vOd3UKDTYki++z2B4iels+bn7ZcfKZrwQErK
KEn19GHbqey2BndDS0RBhHI8JjemmQKbwXev0GNAhzULuuoZliS9G6WK/2zyW0X0
URd3tH6ErTKC3qPURYF3l15xgoTG56rZOhR58TbUcC3hgmeHs5eahbkdpgLofZtP
NWakOE0qIz7LrhLXObAk8fbevLCPAzc8NYnUWzFMscIhXUj8ZFejARD/LCqBc1mZ
AucohZ8UFn46oTWMXQWfOL9uiPQSVGEU7SqhOWaY2STx2RS4iHKMXL558QX4tshB
sxgaVG2kyIwfBLUk5DrXxyq+fa0EWOnuH+545iGE2KAZ7ww7NpOOfJmllS6Gdp98
gAv9RaovA94XNqDGLwHHkQ==
`pragma protect end_protected
