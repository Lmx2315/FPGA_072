// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:32:39 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
KkP8oJnvK1yzctFvd/kRZM6QnH11LHVgUOkPdi5V0Ux+EI5CBNFC01SjlCVAsem+
vFbBCDeDQmSdTkaKE5nrULfB5bu0TAthJeAqkCyxv7+1Kc/W4w1YuOPeWAT7XoQX
pfEGXLg6a7Lk4TzynoZfhD9lwrw9OaXIkhuAUNnI8vo=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 19936)
K3zBXTUHOVn4adRqA6wya8D8dpSah8Z8yRKsI2JNaOzJUNA1GrKIYIJ+s6H1qDcr
V4Gc5nQa+s3puzirCY2k8ymXAGZxUVRRyfQqv+YgiKwb5rBAhX5qoXULgoEYibMm
NkeCMicsrjxgmwSAIHJ1LlnJzNOGdEXAUX5i7Xvyjo04DYYYhBCwSM5KUq79pTjF
z2zkCrvB6evGGSBf+iOfRZh845PQz4N3+UMda6weEy5V3dY1OU3LUqqGxKiTs/P6
Fw+DhI9eXlOuQbwh8S6AeMCRbfj8w2S8tRcHFcYFnfpkxgzjpiIHj0nzhrETt2fy
gFdwzXXhxzH5Zlzyq7EUogUNXS8GqEZDzBk/1ESiDfxrH2CvF9gRGuqK3nwf2+6H
y3jbIXw52ZBTXHk6EZp1BYPITummuz5712bpFt7PgIypMU3hv7AVwVOWUc7cwcGn
gC5VoUTtcZrux2c+hjrZbir6pfcU66/+WwGAekO3FO46xxJwgXyqc2e8zGn0DxV2
V68FsoqKXW39bv/6CxfVieVztkGmmw3l+BJHInlQx6ilZE+d7Uso0q7JSad+RW3a
/o7+dbInTFnzHZBLjAybOk/xe5cRs8R3wb9PLHxUUWLNjikBCKV6Oq6I+0SGxkSZ
S2n6iI6KPxljv3KE7tiJsOMCYB2fQmciRw15OoeNNdnwW1SinxZ0/eINH8haByun
c3clxn0KDtWrzqy47ILHPS7A8Av7musrqSMrAGgqOd9Hb5rzSXZ/Lo3I3aFZFZEN
9Wy28qxVTSspna9lErunMVzCGZygyIUCeIW26/lRrMQkSPolOUUmyqCDXE4ikOjJ
EY8TYY6y3Pv3JcEHqiFQVeA1nBIr2J7EcHaTVbABIwgqom4/DFLDkGGiiobBhn8Y
o8q8u8xhVVxDZs3I8/DcbCiglEsCeSwaILPrBNQqlL1IzhurUZGaHASIRwba6ulV
UZW2JlUxx4vnaR2WXyJiHcypYrn2k9DmA6W/IHwNXTB0mSi7dQszkvkiQLxLlc5H
tv0IuurmmSggIswu4yeKjYnbI0TTS/FKGDGb5OX48MlbhUOu/wBtmseAmmGEIu8w
q2im4OEWfSlTRCVlmNnJ2S2fRxRxiSbDDtpvO4qNOklKN2N8i2cPk0Z3KPcNXrHL
yYpZCs2QgxwMAMYJcIFAyR34Mi0nL2Mg6lUPNSHqWrhx8hT0uIhaNnY+9g7YrOLb
pBZhVL+Cix3t91znyaII1iMET694Ggzitw1bNtPkhsjpyUFY32YY5zL7HVz6EHRK
zR5a80hX7SfqSuRztUcsXU+M1sK1hxvfA196MWqvr5ylyH6BD5cCnkLVwSnfWE6H
PMv88qScPEIzikp6/TwzgnjlrrdYzAg04FPvi4jj0GQYjPOvv0akC9vYMve8LeMg
yWeO5ZK2mvnFpO2cYjfzIDwQpmSmn8QcjO6Fy+qCC8R+NiEXDMzXNDmumfobYhQW
pBTQB4DWq+CEdDkdKdF1JM1GwglQyOO2npBpOy/oRkhFGLerQFrWirl2G/PqMnzl
MWRkZI0T3YUWSFYSBg2LD0jd/9ocSuQTk1pKt+J/Kdb1OkM1vDHJGDvXI0M1VwME
MaWmNlwB98Q5cb8eaAl5jwL/hpn5di5EkxFaJcmfKKTJ2uwlFr0Rkv2mFQbig1xv
tRi3ae0rlKp7L/RCK+hM9Au+m+OORlA/728Qd+AbDjH0ogz/agFGbX+3vh9B908K
jL+Eb73e2brJ4FDzRaPgoT5mIbSa4gX2HrIzSjLu/nw76ih5qOkZlaAlzVxIKrnN
uD/RZn/equgG0aIXN5c2UvXFp+ZyPzLNnX1m8r4tP0lVHojn2acoztE431mZyTdg
TJqUqzEX96V2QwVIDftzWZRL+D3uzTxXXWun925obrkITWTUfEhnP9nTWf6+T1Zr
zAVnpwoM4TRh9I/bHbI6e6JDmJEtnk8YFgtNE7GL9cA6CYPNl5QTgkzT84CtmDXB
QVL+XMF1MZ5LxAAH6kIiR4nLZNE5uw68AWAUinvI7FEkU9gFZm82d1XI8L4Woyj/
c8M62Yy6dsTwhhA/GRuoshti4QAmqjdHATn24F6EDttD8F/dsvvVVkpOrwnCYnn6
NOtfB0U3cIfiheiLH1Qm620ndZMop1vxlav/b/1eMH1pezRsrB+OG+eNRnphy6qh
P5T/rjKPJxP15rlB1GU9T9l7bQt1LTx8rsor//P67ToAzh+Nil/B75PFKCCQaXlO
kvRwtw/tDFwHfQ8helK8GY2m7q6euuYZFt59xju0K0gCLOwoEhY+DCNphKTzZ7pD
6VSXuAkFO0bUIduSC3ywkMQXrnhdAgjN5Ne+eRa+8lXPwNUGmL3c7osct8XsYwfG
EpNZJfJ78ISieXITv9livnHIKuGTLjoL/BKsn8TJzymQOMQl9VKPHxR16sSdthwU
uI7DcIuA+BU4sJJRWteY+kX5yVROn7mrV7iqKiKh3n681fm6bQi3byxDB0sy5ez7
URzd2+VphVANMCBu8FS6xRwvZFz90j2sQQoVWPGWxJtF6dh+eMsNl0zHSfUuJHvY
AE5fCx13rE0X/Q2ls4ekWeJ5AmCwNS3Xxdd32MIiUtTQUbE52vKoRMNsBkw74TLm
QRb+a8akYkkEpK0IbA7vheq6NPP+B3rgLYtgqx8qLsB6AGlqFHQqU5kvGn7zbSck
hgZ9AjLqtg7EAjRGlnqdD1zNVmD5BkVPdR5wyxAQcX/naaCU0E6m1Jpp/G4WzuY0
uLBJmTJrWHsLsZHXsH6Ry7Wq+nfCGE+jpgxP41ewTKk3RofSOgMpJi0CgzR8XiAb
gY3VsfG9ebyx2MkEPNedDD9MAXq/E0D8hZDtQbOBbC6TBpyp4tX8npwKXlL+ufQ/
KlkXxCZSesyBCM4JAxPmFZKsPdFuKROh1xc5XAxB6LVtRExDSNyI+tDzo2SRtFVf
YH+JlA5pnKcHrTIj9Xv7norTlwaCKFPowsKzxkOwwoSH0sC+RSk7l10mi34m5pN+
OJy1GDQkgL0LfRMRIDlg4rqKh2stga8Q0SRVi3NAk3p3oj0Mj+KbpxyEikbHYQ09
Ooo7CExqmsnLinzyIPnk77e8YWyAFrVuAPcT7ckeDUziCZTOc/IVu8fjBqxhaOaJ
y4N80fa8WV1fskZf6Kw33LGyajkFHb2TOe9f+I2+xCer5k65RSRksZ7rppgVQGiX
iYAoVMsa+Mu+ED1x/2ZBiNyF3UWm3qLY36fO2uGoQAyoWKQnSZbB9sxqLmaB/Jtk
8ijjHGkzuvTc3ISojG+8iYkR4dvQ1dsG91AMTQagTk/4+ttIqqTb/lA/MlFMen3l
y8t//oRefVn6B/SACug4lT22VmV2mXv8v02QVF+puZTfnWE5HcKnpOQ3IJrmGcuH
nUJ61WZ6TwT1CDUPIMYel9v0XapeTjSAVisAndhqsZKE1Mg6dUChaVk/J3KB5GwZ
9oyztwTVVYRbakArEvc6IJz1CrKToKMBGVQmxse8pJISe29wPXZdQ4bTtlli9d2c
YlHISPVCJ/b9Tr6wOQ/7HvUMXYMKVTcrCWAm5soQ3y4zO9Kbil41lWD4inwVvDoZ
Kp/ljAZ8T5LL390iX64hqko0Dif4bHP/v3ZK/d3uamaqbeGYI5DEXbBXMnlGs09a
35n26OHjRyPIZj/4fcTkeXdmsIMhVz4tL2OEyJTpyiKYc1kibJpOJsjOcpP74zRa
f0hJIwVaGfo1FxtfIHvpIKEH8XskeXyzy94Xd4Ch9VVxYROa0bRsmQxDQKQ66uqM
/Us9gRLgW66nhTjcp31CklvHwtHEnkqaStklEV+q1KnWlCdlogbtXudX0kDN70F6
lv0yNpWYfaeutD0E+Z0LRkjudUUdanGvTk/DYsTvhBM01rqMKkwajg9u45Z1B+M7
J+PRhoTKzSsPmBlr6jTHX9YBrwkYC4qo3zpA4l2yxFbvQTXXKkDQkL6NkPvVngl7
zquLJaklIWsK/uW/JjlSpXEMTKFLUggqhc3SVXRI74/kXqrySx+jyFE+hScdNMbp
5MK2Ruob0MKS4mtiJsWX2ABBxdCVu6wlit+u3SJBHw5ZHNzfe4kuZ9v+dTvNGwkI
Hnrx8J1WVEacAD9EiLqLyicHMIsyCPVwTCbtz/0UEMl9UKnEmJkcXTkuSCz84f+6
3Ju+O+HS6APQUyPGcW9yi5QMK06VonQcmiAazHdhsukj0pPXo+bFZWTvSIu+poDJ
W7xRmbP3nBTap5tndsGcySlStQUCdD/PbGckzfIawqTsKb5zX3L4Sq5jGzTpv1Ts
g6zq9GiStDYvQjGzZ6QIWEdHH8GYQLpxo+AJGK1ztvGrg8F9yABAhKoKjnA5QJzh
Gux26ubw8BucjNj+F1Z7ASFusZzqgfnc8q91mT24EwpvO0SvafITgd1UAzUvtJes
yTWzv2k+3J9QlCK8NJUmZjpZAQIHJCQ7pCbZWgFOHa9ACPfQ2PbXlkvgm+cc8FzI
poguWKUPHy7rTDx+s+2WDFP8yQ5FUnroWqzraSYbSz6T4QItOb/QE4fp1jUV1pSA
ZDgNIJKfFiLWJIh08woJzeo8kRd6Kt9btPLdaEN2UafLJyAcOLnsgxswJB3paZ2D
PBJgAkfk0Nqtxx852youSUZqBCAtp/Z1oAaZgDwyd67ME4my/wTGdMpeTbTLa+yG
8Hp295eDdlW7c21MQAmxSaqURe5gYnudbo9Ib3oBr8jbSSZe8ARQl3tKzi9AnuiJ
qoezRISE2KaAYWE4IT8V6yajg33RUfnz5BhSAAjbhjPZco2EqzJRjtaUKPlwldtL
A56FeysD4B6DZdOpcxNczs5hqVDJwkdM8FYLzlU6pNSFuw/D5IRfxwLyNLCF9n23
9GFkhvhN5TX3oEHOAJL7BKmc/olOIRjz/+gaL0fQgRAIy1p5dprn1HG+hWOS8oRV
oXuRD/mizsqNk+WttdKqwq1pic3659SAVZvz8bCk8FyaYk9nXYwxI/5ijUJdq735
U3yWNqvmpla6lAI0U4BAMrnWHA2rOeM2Foaok31ysfrctDrSY5RqUmlf668acGMk
SZ735PesykC7dFuAgGUgtFCzTRpQGuSQFL6GMSAJjG0r/ddurvR8VToYm1mbeCRw
e7VVTyYeVUI9wIfpBe1mBBjXnznvEE/IBwMqDqoLhn+5jpYGZ6BJZP3oHO7+m7qJ
3mJOnmv0DoOrOEmLL7tDrR4LAfW0mnvvNWr0xQ10pLBwkvlETh780ec8ktZvKgBO
0w8CWs6t6fkSIAod0X9/yHYobcbrknrOiPfRC5/gjDVFptyKtrBY7Y2+5nGl30mb
d14TeEMUOXB9gfseJEwYwgSPIJDeHYOWBvVK9FYgaQeW15LtmkqtzvNwcyUlOx2Y
DIw+C0yOyIdm7GmXfUORRS2ClGfTxsXH2oTW2W0mdXM4EjBwJlfHIEnVUGMBeH4w
rhvrqOLwey1y2QdcKMOi0UG8UtnjZ7jP3LUOz/ufGUD/fKYjIMkQZDbh8VfzGAxG
fYFxlq8MA1YpgW4VqCZlIu+Ti78LxI+uLanIy98OEwjbo0JIsJZLmtUx7oQCLhZY
6THT9SN6bjSwwCqZvCdiNtpSvTPjYDIn472YQMJRxqbfi6onE24gaCOq2q4oLw4V
5ol6hJ4KZL4tpituV34Hz0hZcddaSTVgSniHBPZHzZ8QsR7pBo5sSjtuAK7UKr6+
RtNAzBeTqZfmlTzerSBitwwHBpeHt9x1MptT7q0tzNE61uAgjzMCZ5PUKCIwPele
PAHLzawUeifJqLxoaMi0bt/cIOjWys1za4lTqMRWpGPv9Pb4vLLdroTCp4qPY0Mr
iA/251XQisJYE4joHCRGrmeuysT/l2r5ZGhkHJP3GlW4yKOSfe5BOdNICIAqJHAh
nh059tNjZlOxkENAMILiKHBFHGKpbj4Dem+YTYIjFRo+dCo1XWQL9bPdQPjjBO/z
ysFff4ATGHuNrEL2TF5a8K1g/fi9HkPHG/AqIKXPPXdbekPlGDc+vlBJgdjV1Tu1
S9WkuP7c5oQBYtt2PvQt6Gauss41zwj5fcbyDMWJ8JyEhcoZaVBLdwNDGciOkz56
FnFkE551EQvw8PW6vfJ3VA16JHqwtrDJVfB1l1yL+IGEArXMH7IJfd6NrLfhyFjs
Ii0I/luWk2c1VOdyCxdFMYHCKN57bHyG3L5GkOH/Co7pEqBemtyHT9wjEp20/Ge3
DnmOoK4iiAXkFNCRiRm/SZ7ZrjXoQfF/jN+fS3tl8iC+gMGqxx/DKMIvoPF6OKhK
E9nb2bqeDjjRVh+8jhCw3UvRAO1HeLG5ThVmZx/I6yKGLkF9jRQ80s9NILp8ZL67
I5jSelopQu8FHHjdrU2hOeRrniwolCiezkZ6ed+lS0cyqWCqc2jQK50TLLIG7eqw
uST6S5PTVI+tt0yqoy+510+W9QTvi0/+oymRqyxWglg8KqkMl0qCVfTkhp4k2rcw
/dpqtzbgwlV6HIP84Gh7bmRGq0767+UtuHjvQWhPMd0DR0h0SUc+k/oXoa3GayGI
t6wcHCRBrfvM4ty6sYc+bQOXvUzjoff3D9TKbfEP2qpTtGoY9BRlGi0ibAcYgnEq
ZiHAmGXhvC1qwf773GpV3KmRUPvX0uLtf9Umq0RlUjimgpNLnIha1iMJiVCGBhZb
EAk0pehNKtLY9VELYBO+3D1K7VBnDuaZqOhJPxN7DE/yYrKJ7W8mXklr47vSY/vq
nOUHr/0YCkcKFeAH27IicyKjK6LIf4eADMAm4jb8E+iaumy+IU7xZux65UUBeUtV
/C8XY44ecsfvvuPrD3lL0YA9jSQILBuoNITJEmb/v3IQB8jDnPtSWDsDWjnsTlcD
Z+Cdh1J7qy70YKfz0BXB0N+6OFr9E2U2ILuSCixPtDeCcB37m0YQ7nrAZN2WJ58h
Yf1M1B606aAsyNUtIugIn0VOVsfkJL9y7QWC/i2smDsfXBfFLs08+Ult1ivNUvVl
Ce0LxV06/kYQ1I+UO0KKMczkWy/mr92XuiDr/cyWrLOZvAZM9XqTanqV7VJuoAc7
Qv1ZS3Xw9eWOCsSwNMRzFbNqu/pwmFVdAUjPEMS/cCofjK2n3toAB6Wec78WEBxL
Zx3lNz7QRbWCR/4KN+Qk9VS0cVqCLgXwhL+3YrD8Ew+OoPUEsBSmoFPYQXxhfrAN
JYq+VbC4REqhSJbfqFQd0//q1Zx0lBLfdx14yrAol3JhdpBVVmsfAxFveTdrt+IM
Dw8sCRdhdDakxHSMf8+O90HdLShVlR4OVke8x3eVpaHjAXn9EeIlvHyR7kikpzkB
iq/h9rWHckJAYWtv3lZEIKzxbDbfPRqKGpbv3+9x78ydlzYp7e7izcA3Yt4Ktf25
oOB2SegOpSPDf1WluJ5ni7NPhgLlLN+kYjqLFPUtR1XAQwFEpNqhnAQ02YQCLpfy
99bmt3MyBpp6lboxF9HueDn9PUK1bHI6c9qN0taC6SD30h3iyy/EwYEBEzYKEfC4
xnIqQPiMkmPZLoSwF7YVTOPochArFMRNXR0sDgnf4fHgWWc5Y3zFLpEa/pJ+BCR1
N/rXgrqnypKyzaIQuqe5ORCSRUuFMg/jY1ctORw+HEGzSIFDfAJjbMSg+QgO2XCc
NyamMPVaEJkMwhlWfVrnkCEhagP6tCHfWUIM06xRF7ojlN2PdErDzwnPZVVSkUms
y2h7kha6gGgy4HFVnt1YBX5ndNOmblJ79bKgGFCuH25YM+pd5Hm9JSPPHkIOrdf3
wxwTNVYvmC+YODiekP15g50HNju2bBhgRqSEUVVPC+4Aen6HouSukyUCQoKgoKMh
7FN6/6ry2/qXDy+RrT3DSvzaR9XZPio2BoGTEvQTB+9EFXal7JpuoDSvXTa2UgkB
27kIRLmTQ5916z4SVC0oxJSB1UcKEawyyZjJq02Fb0s76zzcC/fSMrZME4juvuM3
J+YBd236i0QpSD06hMfoQSoBqo3lHKeD8rLjgak5s5gKbqKdvLI0b8BLsyZas/3E
OqrTJKtFwiaM0JZ/uPLszb7Uoc9M0GubkWubErL7zxnYH6lXmm3kZ7kOTBkgeunr
z97LFkHgk1wldo9fIXrxqkPZ4uLDH4RZlHe1GO1NeEWNStQFsNkhC8kdzk/Tps0x
JYcEaK99Ev9kqH4wllHNB9KQDM0DmPcZLePxp+1wZ6WQBAqM8CRrA46ZsbPTc/Ye
iV22tXs8i6sRaWvSP/LHEKhoOT1ZXJ3Qz0WlaOM5XHSwu+C4nx8kNUptyygbI1Kr
GCoh/aOT8vKb2XOfg4A4AbsRNyWUQN+ggP4AOSlz/ieZ2WF50DqylixiPr9VaBEa
BF9hsyzAq0W3yjIqH50FNG2oq9pprDn70Ej3rcRUTSUp0xgrOnPvVxqSMsyswJp2
Oep9SenbNLD085GpzE8sZCUS0M3eFTgBoRpw2JM+ozJM+kwlPqWanAUDlvI0S4rZ
91B03nEkX/M8AfU/+Cli/RGNq0Nk4rc6YgJqkHP9IMAM7CbETU9MRp7fcYiiqL3O
4BU8AFQhKwqykJ08kbRsljn6inSqXePE3Q8TSnKs/I6TgoRZvuWBqvX17x77YXmz
HPhKdQtgwKlSdhcGCa/5LmYxdmzkVunXH46PuTQn/CFHRbW/S/auuRLDGuYlJNmm
O7eeFOfq+0WLkqHkkRkLEsRYIn4gOJyD6OZiDzJDVfrzkxkx16pwTV94Ww8Cm9fS
NSRBK6dYBdvTZ5X0vtRt2Y2jNnRTBtsUjGdaldafldu9is6ayRKar8OvNLUzG3C4
rvlwmeYdaXZmrIwKPAR4BG0vrp9tCLarxLg8RUq+AKKoqzgDQSExuMi+TACbqJdx
mXZuBSM9kuRzjP7JJUJJYpVlnJnkUyj3AikSLJV47zlrxReFf16h8TaKlqPW6RWy
gFHXrbt1TVJbWe8IqTpsPaR58UionzWLUjnB+Zz3FX8B208dWMRzO95+7BQ2zVHX
glEFjsPGUiN21BvpU+Mpj/0qCzMNpLC3y1Tg1V33Ie5oYDiDYU1Q92jOI0Hx6w4w
nC8mYPBBD1XBZ5bW8jc1xKVlrdllEF3G2vNzyVRsxYYzThgFPJsD9j4cJ2z4UBjy
wSuj+9Hb38aOWrPj8FwooDEpvDMAfe83LKi51NLKIii9RxSJq8SrGfAlBXpHJSM6
SgIpP3TWDR4qjrLMzipNevuLBPempIJnhyvlP+zR9o33Ed6jxlcgeLhM3Visi+eu
9DFcC4VdvXtaFVSUv1xyOWSiHGEGjdqoH4iUXYEPuWB0wjYgm2pBWi7bLbTfstJh
Ymc8MajjBGvK6S8ZKGURn5lQB1gJ068+PWvJSD6W+MImd5zWo2Z2EC3ng3tOmSBI
anY9kGPIcD/x77mIrLG5Ni8XmfOlOfEUE5tkpx2rBh9cOls+Qs/7qdqSYgYUtWhk
xrH+KcKMy1drbw9VKwlNR3AUawVZeGZhVUgsXsfp4EhF0UmfnW7Ctvlizpa9TqKy
GrL9bhGzuSbx1YqKniZojxDWaTTXvy3ZFWAbwTn1lgQEeIn/4t3KRsn5gI9vQty1
h5d9N3EvXbxSego3724azgTDQh1FMfcwQLCPU/jqmdRSnhFABvT72Piqcii8xQQf
u+y2mKBK/bMuWrC8SKC3RD/v1sfCkZ5PQpYsWj6VzFTCj74COmaonuQNFo27DZXm
sciISx8vne1otJ/Whug8dWxhaC5JEumNlYti8MTyHzOo2TXNXV7kRzYpRBiTUZUJ
eRhN0xV7GPqNLlaZwvOQ9I84yobBtxa53ArlwgXASxNxlkyCLocTMbBD9Ve+osyB
31sn8XOOey9YHAwkcWsL2nSvRDjJhMHIL1GeFQlZgv5c2NCF7YsCJTTv/iIqTSST
lf6bFW791tGOFbAXgaLB/V2He84mDCUoL1LAi+lnd6sF+su+gx/kjO5L0iOHz6T4
EpT/FlILgmZijYypLz4KLwtTO+9ItFBVOAqIYokzQ95NdE8ohJaQNzUo0J8/VaF/
V/NM8fJRMm70/vyZJBhkwBNzsigyzvTPT5uXV1X3aHWqiw5Jyr4VlMOZynZbuOBi
gDhJkVdO4JN5j9xDhJCZbcXjBXi4ksvwkYsIZAFnSjBq39Cgs7K4SXo8rVw85sGY
rFJeB/REGl8VSCwPZ/bEUJLHuF6O4fZJNJBfRMbJAbgCSFn1V8TL0Xiaj5rFkbQo
rhNMDgv8K+HGcCe7FLQ7qzKwbgqSKN81oetCL2iucLWKJzT3h7vayyo5bpu9Fw4+
ddLZQ9J1GMYVXjrFHEnGsWyUurejfAIGZANSqAxdvR1W5Z/mi/TCC7U7D49MVSiE
KVifAA++4MbCefItYk3Hp3cwBgMMbkqyXP/y5Y/JBxH8fKuQuI2DLoCiMm/87YTd
vzmkpHqjrUCMWpBzCWRMlM60vAx8/L3v4L8G8HdI4ohbAr+QsFgGdyRYfJDGrsAe
bxXe8HMiHA1FZSTxr8cXEAY8EMw/fPQM/UH92RPgw51Smddr2ftzb6OO5UhZRyP5
Lap5AgGZS3GPnM5bhEZqTWwY/LmgHT/+/hlwCEd1cP6d/72MUouU6+RcFLl8Krpi
pnPtDZfMRbpYB3SNJQsRYt8crgis/G/YmMuSaLbv352/fZEZzL8lauACDZzGhGsu
eKhh5NK4fQUXi+JwYW8AD0jP1FnOT5bQqgkb9pVau73Pv4onJd3fWdpy/1C7vdHM
5K8g37r2F/Cx9isqCMecKtROz1dwcVrebC9n/TLlh3iNS6l5QgOBH9GHdKvRbQnT
b/GzuAUNYMMbMRFeRBxEqrlOjfVgYG44U0/pm4r/hRc5AWilbt9T/EI/Z81VZa8c
EHc9AqNHTjJHgjJ+0e5dsyadGgjr0ahPr9EWJhtARerZJBC79z31G7aV1KmSQaZ9
jcl+XDdPJvmD+/VoP6OfGlVgYp3O4IAHLTK9Agw3XC9u740fHihHB5FultOma1/p
AZJJQ391PBlTHTWDNYU0KrqiWwBDPZQiCjZW6LMgCHas7v/SemC+o3EXg/5TkUR5
3/8iYDdizXh8H03Sb79h3zIlm+MZWe9VkGmQCWnyaa3ydxJ0Vh3XEEoWalxScFLB
YokFKuDU+K5ubmJpapOClUndym2eZdOzVD1qu5AOsiwkd1QhFH4Onrjd+bMcc3n8
ZK12dmIOec3Qp7XxtPToBs2PTBJdk8qeDJ2KyU+K8sXKeDPRf9yBbUYEuPLdEbVa
gu+8+mZ8SMvv7evpMczHc1cyU8cDQv0P6pAaFz83SY+5wPzI7iXKvr3si+2b5K4s
a8SkCgk1LKVL1zJgsm4nzQlttqQZ9iNGLS21az9EHK72VkxnEL1fXRtZs5Pqd+kX
z+T9htmLw5JDUtO9hs/jNbbDc37oyvp/X0FHsnlLcOH8RHuTRfIBUXn08dFe4Fyn
c7HbESaj95frz5yATxn4/AXNvG4GE/Zn85Qe+6ctNf9cRYwRSdn9GgNMwKV7J0va
3qBnmaINiEY1Am9vOaxfiyjBXSnimE6pNmiP+8qxuiwtu61ov6f0TV0RmWdWsEtm
uR8ysUdlFOU9Qm16wDx9iEG+E81r7OOphk6ufTC1OoxslGiLZwro+i8OnnONYPNC
EQCvBd8/6Dk2w7tkKLRYfvxnSxB4rtFrIA/WjPuPYIS4KvNQnEH0W9VkylKUO7kK
O2LT+TJ2wysmfCoNyrrgXGVofd0NeE7N4ZXUyqvTq3yhwHeDZWxf7ul4DMxVn5W5
PXPXhlHPXdapwjRG908nTwtIr0hsDdZ0CQoV7AHQ3YWe/51zlUrdDJmCiwCobgfN
+Odk/iylE4HR5H8AjFW3OE9lnuu1nvhX5BIK/blTLKYzj4WReALHeJAFKxtG3mol
LWrwse/boQG8mTtNnKPxVplcCpUSbyb23i/OvIHlBQPmvHAqFn0hox7I6q2Jm0yl
ACqbmjYWCcLAgfuRC6VL3W6J7hztbkCSSh+4zkcL80rpqN8Ncy9qXe8IyQt8udRB
zjbh6RWxB+1OGSxuZdwzjdaQzq6plF4ZWZjxxosJIidnfSbnB+RVtCGLxM+UGtUw
OuSS6oBSQcIlvgpkgNwGJIlFZu0H9GaBv7OVJy/+OZat6K6zJT4w69j34fXjAPmL
rMw/bZJ6Z66EjmPsgmbSCUoDvab4wlEhvuabvJhXyE4DnmhGOig/WdaXXis38kjW
mSKe9NSDWGGkmv7JHSvMFrXd+8BaaMn2H2amL0s2D1Hnbsrffc+/dxAAwQy2o924
gpFe4BcJKTmk/5lMWgOKirU3NnUCRLoZfgdbDAbHnO4vHBM0M4rCaA55H2IoV1B4
GxPwyQGhHK2U81Fd8HhQVnRxro8PdtiT6GNirK1q3W0CFMmCScQpCd/9lI5ucEbA
Mnn4Ok0dFqDlzQtM8yQJmsPOjpsK1lsBY/X9nVSk1rszYM+pyLe8yDCOrIs/eEBf
l/GtTmnQTZrbm2PR0tkgTUQHG7g3REgJw2kwFKKOZWoiqS7pxseqCiRG6wuA33EL
tqGNC9mIfrH5DmwhaYlVYLlnspS3iWRmxSbH/zSGI2+VCK3nSOJsPAc56fIiz8kX
x8I9DH55JcvDQENDymNkB73ckSHQumP7TDAjdqy/hdEDi3zTOCeXVjII3RXc9iZ3
0C9x72WugATCbJjTjExqB7ePtTmYsjahxf8JexL0QqPe6Q7AHvS3DBE+BpwyOYYy
2WQPi/wFkesxLkHj15rORMbTVZXpEPqOuaJ5X6cHGz17MwEdmTiZp1gJy9K3QQKX
2i7GQ/GIkoMDZBFYhMck4xIJz/F95CPlM2PMV8pvTiU2eENE7UHhLQLZNuZobd55
TLTL3yc08zC+FxyYscj5TbxPDa4JcSpzAF94LB5uFUrzuufZPe02KK6bzKK08zx4
1De970Lnch2E3++Z9FuaQMbP+YPbjuNZSXpNvgHWYG3sMA5BNE3vuYzwDuVoc2eQ
LTP9pdRX75T4YkZR7Pe7F/FBtw/MLMcd+SS44H26GSVUTK5s0U7EvjUX9Z52VvZR
B1Io+pCIbfPhPWOaWWoOmb6AYR9bWkRt28Ol/TOGUONlwM7tz2s+ipjYunZcWxca
YQkqlYFZ2ZTQjIDJALmFx7Hnfb9g5eWqVEp74+/M2noYkTvj3EckD+8v1INwWKq1
zUt9yy8S5WrJwogX/TPblMu3yl9e65KWGUoWpsIIsj7rIG6Qvvxnjp6qf+EiY8lq
o+blIPMew3Cn/tOEzKBEG7hoaBJdqLQXPzjhxez5vUK+RCpbqnhOZEsgHjPmZFZS
40lk2p08K3gv1yNE02rfFqIdjXhSGl4QrstCNV07KnvOYTlWg/1tcVaKExIrb/e1
HUn3DUGODMDXr/TQZlHu8uqXEnFiLEZ3oKOdrNJkjBW+JVNKN7ApvtwDUKciat1j
5rT/fR72GpUH5wZBM3asHzCEq5QWqPDuBlgKlF+dX4nG+sO3Zca2V2RQ1F8LY8rM
DrVv6GlRMw1AKY0kwOqfYr1puO6yLKo4gFN/jP9kF0Iz4/N3B/KR3sa09WuLAm2g
P5WYNvS/a/MydHPinVO8xJHaMoR1x7S5zYKUlUJU0FNRfZSSUVYdcaRG7LitKh7c
nbE+ZwwoIhBKMPUdiAs+529Ag3z0fSf4dpMOTSCNujdL1WICwTvA3R6TkIahua2N
aBezkc4Zas3Tz8OApnJiJNgHPZER81gnHLsIP1zGhMqudkpwlRmeN5XenCu5IBar
HoJiyFCLbkP8XTXqd1uRGtSY+UE3uNnP2Pcqx9zP6wfYBeJEGvQ3bFRcwzwndu8Z
P6WHwNaVKKqB3D4rcs9Bm67f7C6M6ZJAbC4gN/kNwCO/m7Orejj8y7WS4oNMqBys
b5Qt76qMw8QVflhtlIgLSNPmXis/WLahfwJ2pUG97IP7ihaI/wZkS/ZA4MOVovgT
1t+4tRK0mMx4xThzWiL1t0IbwIbNiK8jJvq0Bx9F8MOr3XUMZvJV9RbM8sGtQ1KH
r9VBvKw4xUSd/DXUhepfgnkzNp3UqMpltjx9iftKJJmL/vmXI0d9R0VyLwPcNYV+
/eeUxrwPt2CBpLy7HLb/2AAYMURhvC6FOyclFW6Wj/1NtA94i7As7HGuknTVAgyT
Z8GQ3EdzsYMwl/hSrSya7wK6bBvute+C/KPeqLWfnR24LO3CEijqr94vjMuhtxBt
ejqiW7ppmBWjWtuDXHIZr+oNQG9kII3SnlmWKr7DYPBnk964FDLWnbQbDd51yQOC
o4RjQpoCF8ouMaTW5mwYAQAmTXIuXCb4k3G9hDi408iNd3sGIaXYLOsMvGp+cJT7
5WIDfNOEKy6xOYioYpgzvVQYnZbp0A0B1PQNyKraMAjsT75xhSgkb09BAVntEBeN
1GWo0JIsPJKi1LQfw5ZKAfnkOvBXhloZky+HlGg3/cPdWJE9NZ0ncJS1WH6noxLk
ckn6VfYBks31cqmlSmT3wHqtRTp11cxoLuqmnqBUhaBXCYJjvrlTbzEsoPhT3Od6
ITJYhZtO3bW9FkjU4EOePVoV2mZW1vmaRwaN/QwgCy3qXvWbzdUNGqkB624aH/fS
ozXdvmJ3edzDhvM/5+2lIKvv+Qd13nRYyQiZyI7WQp1vHxHIkTNB6578n90lqKUx
IZUcBbmMzQ91InEf9QHzM4xZ4SpHEszPiq9OBjCDufDVE4pbsftsDGpGuEYhUGeL
ZADUjMVXW9iVQHMSC8e8cbRD/ZTN73nep5riXQxVdztTxyju+NxkYfecJZNv7p9b
ejbklEZBqb2tPwKR8MFEmpvYijizDGS44NAbgIJ84rsTcQ2at/2Pmqx0Y92hUFL+
EnA6aiQ1ftjCyxs5Syn3fJGiDssk0GzZcLYydUOp8b4w2U6KgnWsM4XMMJPNM2yc
UDVour1ILMNM2JQcu0BQqvfGrVIKLy8PUtTcXCpQleSkPvgUYfpQbVcJNGruQhD3
SfOZ5pw9r+S9lbeoUQGGNtyeuE8LP6FkDUDuesZTKVaZl5FrQbhRdAdRi0ue/I4Z
TXRidmirKhhZf7a+NmYQYhgXwtNpdUL+5wBcBwiX6Z3qLLqrgGitdVdpUaR1lbuk
PT1fcRJ59+yW/2Mva2QNrk+7cbcqBgA6qzh5cYWwzGQK9zKlbHlX4DOHNMIpT7jd
t3eCUredQiJLfemDPsC0FpVWWBdhOXmnMQa7bKZZEfdYT8JJsuFEPdRmPzKScz7K
5L71mHg0XXOHyv+S9H3evPd29YAebuhzy4EeBH4CJnYT1pAybw4dtlZmcEriDeJY
jb9jkgCwhETbZzRnPVsvcUcEasOVkiRmbUEINb0+dcr576qLw5f0GH8OXn8HkZna
9/G7F69WFY1fcvELfkQc9w7vEvLNkEhBupoyQXro74JPyMzsq3qBs7SBmUjYRi3l
35XzKLXm5uuo6f+XZr5SX+1i3kleqQU4Z/Sf7jI48yFZqdTMdkkgNnyoJnSzaOoy
mdfDN/dogXkpwRI61++fk68kyQzQAPc6aSOABQ3FUa9XGm73bBBqOJI2RzW2x9Nu
yrYrbCwqtfPkEsUd0yTpmQwvX0QOy6NrGVodBxG/Mb0yduPycNED8pa6XInprUaB
UM/PuRrsMMERxAudRArEP/X8pyzOuZYBkpvdtoeYN5cmztM1oKViRPFTDIWNlCAR
0FyH1k0vjo/MhfHJ3zRi1eaunlyCi4oEyNaUrulEDUsPHvjkhH2xl9HCF954U3o8
Uu+4m8iJwO46fU4q4+L2z5uzIMtPTXcsHmhz8QxhqwC1AfjXU9ffe+ubDaq0/xel
imSMkRIBYydyElo7EDi/2VjnskuI3B9ZQXOvRWQqsYw9sQjyN6v1/c8MQw3Majql
oYmxjfmFPfCW6syILp8Qa+qIKQ8BPhNOedTIMUsqWYDvKfV8/mstxGvdV4Dn0gKC
lkXX+Oo58adlDbHFpkdITs2mYeBMMjpElcAjeKIgaxgt9WGxwhqCFonBnMnFiXTN
1uVBKSNyBZKxfSozjBADGBCPN83lUxS2vXnd3tqUuDagTBK0+leVUe4kZ1dLDayt
Nmmcu/K7IH4uYVKQzrmM1edgEgXiJt7zwUTeHgCdk3/iqUUSsSEnKsLnagyNHJFq
DRbZB8wTRk9dcELZbmSj6MxSlmH4ncLZ2zu+CIP5EpXqiTurkIa/0nbEoE4+e+pC
Jx0GlVpsMDVaKIHWX6t3iFw+wDl0JiJXDlfOmuKkJcLgm8MDgY7BW9baedc6DAdY
0mKYQWG4xlyDY1SKBchb2Jtu5t56mWgFso2fokTi9YXFUmn4eKN2y2OqOrAR2f3L
8g+xveZiwnpatreMu8qR71u/yNeE7rAmQYBRhBs32VltxayaH1KgjHbFrBNNOWmi
LAp1ZUVAouIVYlVv+XAMGSQuE6M4BJykTe3q9ON0GFr77sN8aSB50H/K+9tK1l7h
Q3uWsyWi8wLBRKyOqIvJRBDX6gUviaXlZikETucyNyMAJB14gCD2yhlV8z+CGS2/
ak+2NANyexOwag+kKSyPHXR2ceYPP4eW9PK1dXu4ki+SzygaZ1Vhb75LOJ4ZjBwG
sFJyO8RF8vz6Zt/tRF0BMqtYR67XXQF54eQCTD7u9VXg1pqtqjRiOG4uwEweT7h1
yQ6zYgQoE8cku+7OSCxcZ7vVmvUoIvHqYXpaCDS8AOdsb89YVGg4R5OdHCbye0Vv
eexUavBApBvJEunbmCRSLaJB7zFNTlEaYDHIXedINF9L+6i6a7f2xvWTMjbhSmJk
FqaGBcbXkgIkml1+f3NnUraHlGm57L1ja+9PqDGNLYSaeg2SScTOTdBN2TXIR3ns
vaCx4VEMMqyG9+tTLnJqKzvqj6A2PsvROGSJ/5WpkWPe3xgGJRcTYhnQf/VipHTp
JY5Oe2wytdqUI4XvQWOaBhEGAmjy67ado81VIWPK7ljAFbR9sLYilPLUJoeL/raj
R+Ni0sihsIQYAbbjY8QAGUSn4bHWRE7S+kIPEJ0JcvJgFN9hhVN7wEIM3kNTOlT0
DweNwyzpYlb9dKFqfIDCQ7WiIeUpn/OrG0BXQAQAz+oA5KSBYypYmA4cmLkAfPAX
vIJ8UWzeSBW09kMDWEqYJz97WTQVcOd99wGh0x458o+GI2O1DPIV8ypIBxRgmNiA
M7ZUYiSMC9q1XNtj1nyyJ84IHtLxin5unHjPGte+MNo7SM7YMw2999YVqIFWfJbU
IF9gXPikxq8dgS1kXUjLbDL0LMi+TV4yn7qSn1JZgNwFeJnNTxwo63QEembVIwGQ
N1CZl6SaxVp4ZCwrak5dSqpJ43PSv6jSQxDaG75Eim38ca2GHddxng2za7tRh1dG
dQDvNShNph+P17krPWU0IXHzLytvRK3EYia+N5Btiuv21uolNt20OIC6B8kPHst7
SrCQbKrsKYu49m+dwBaLG09ltMerkkpedKRwlvfX08QjWmv5yCRgjOn8ZjTtyzOg
uUrGlXtMw1+gbGkDH69DQLd/7WiLSJTlLWAwOlk9/fJxjCZc/pyWgz04CO2/rWwX
YOaOOggCOK+Q+NCCTM4fgzhvqSJubCtJhigkqtvsoFTe4wXlQOHqvYbd3AbnsD20
kt1KLSRFvPR2RHrcuxGKWfBWapfXwx/60I7Z7kEe9FDhICQTlttOHBzlF+CBnPZn
2zcunLU3I0otfji3UDjN3z1VFIqg2rC12JcuJ8INt/dPhTuN9A6smaYVREuoZN3n
AqRITuHEW9I//uFpK+8A0tflgLiiTJV00dMHaM/OG2Xpux0hjBbVISf+QSCoFsQe
FJqEthVSAW4yQQ80pdQsvuEoehXEGzw3OmGQqCHOFrlso74uVuk0HhflTDQh8Aem
76HGj+7cIHrNntn1PxEyONstieLen6IKj0SQzw/tDDMJexQA8SPJWgvq5pXNaRgY
7Ey0L9q1ThdfmRCH3wn7lc/T/B1emldUzxoNG37hiWc+fYDLe8jIVfS1rV3vUbud
/9ujRw4xZyEe5UzDiVBGZpeU6ujLPp18aE/fqO3qA0/mXIeyWr/hurGbbOnL/Pjs
12Nz6ffOTrwjbeNrUHpBMKy9VEdxNCMC3FAbw1F1QHD0TDHKnh+OYYy4dw+9i9tK
t9R9IzNbQtHTnKX2ffei+j0fIqcaA3zGLPcNY/jSDiv8aSWK64uis34VpXpps6oh
z4YZGR8kkiMIhAqc1T+MVT4eYwbErsDC745pQFPZqE685dLud3/SQdlzHHdEAZBM
5dqX7oq5k8rVrc4pBUWSuq49JtTJXXXHiQ4FTZNWJp6c9gtlfgSLOeQ+1cakXIPq
pbO5IoSHFpdKh6P9dAumNDvKFqP4jJEvmfoqhXkBWJizW/ZYFn0HOibfyWflWnEO
3ZII9p/1LBmhmgYE6chenX/pINiFeWoKqkgE8tpppTlsCoG8RanBYDY01AUGm1Ze
Ivb8aQ6cdSZTkT4XtualH0o7tExYhh0+S/2fiwYcVNli8JqjhoANn9YqOmYo59u9
q0sCvHjsomS2F1tdX7SHrOQkrrvgt9LJaSviZwuUszLtB5k2pfgdCORJ/2J95R2a
ki4b1H206o4HHxSXenejngYqk2KRxDajKl3MtpelojGu75m3n4w5g6jcpMAlO4rx
yOWpxWcrQPRdH1z2efKJqz7FZXNdhnXM6Wg+bzHxXgLFtZYJXxWyHZBMx3DiME8O
CzRfvHG8xKiMujpgNrUVYLIlLsY11/f/JLR2XMEOe4bhu7JNMHwGT8DaLKOLhsUq
O/vwPU+jp++WnbBtHtxhw7SnPVJ2kiFTfzVjYrKQh4Vcvz4mkBJkbZ9MLBBY78Of
uf1hEwIQkoELJ/YxiXR2bHRNL3rTo7Q64UOErEwusRgfpSQbERIW0J74a7dWj3pf
2+RBtRnPDCQ0ZlKmG9Kow2NBtbrwY6CqOcQsz0M1DSQ60uHTZHWwUEOYWoJlDl+d
RWQ00s1SQPYNFdd+xnaV4iadfyAAo872JPtc1yZ1gWYKMPYi0X69ltvT2f6/Abi+
8ikuxdsPYvBvWyApczEeT8uqWDYj7kKPbpI5gv6zwdrBh620o4tFMKip3zF2wnwW
2ZbCMfJQwpn6HS7/3TPbt8bMFLVodQ9zvVWpVuBRPD9PRMAB+swrINQw7Su8tMsE
N9GN6b1j1q1PAuqyedql//QMgSYo0zI2tKus2gTRfVwaxoqfgguQJJTrKMXsBjvn
QQ6I7+Mtb2o5Rg61+OHV6Bo3HldZhc+kjqb7iuJNZIAypaUTdWSg4LAvR+QVrKHL
MEZBzZumG8VLfHoRi6Njaa3Edq/bDD4XqkSbnzlTI59oPMzFRWsYJ2SGWD3/KmCO
8kQbLfiKgf+THv1To4BGsogaccjngk4LFglmDA53sdmUNTadAN+A1gFuIWSNTafd
YgCdzg/yw+2+wSOXZlL23BSDrtvovrdEGMKHYlTAeeuxN5RPFkQRXiewvEgYdCWg
Oyl+MKcGNBHvgcfE2yMldOUtBd61jZcVbsFa7yJAothXVqMm6fP5o+4LHUh/uoT6
l8vO9zMw5pZ86XuZq5cVH4Tq6FORVDi7PbwtXuBTSsgz4ReoJCKjhKrm+xWJf7wy
M/OjQtjxSWe4C/Kd+v4OxuP0PIdG9+ksrJ7Tw/QOOM82MYsHBZgzYtFHBkTjsmJH
DU31fHkzLf7yVlr0sSDsxvwtSHFv2qVJ+qrazSat/PB/ufSW33xJjfF8IdP2Dk0K
eWdzJgEu2Vma07i/aS4AmD3bgjEzrYCk3Jow7M4P9ls1IK48ujH5NXZRblpTPVyC
XeSJW0TPxfSYn13J0aZqC6aMJ8/JmlbwUC1XHwkcln8hK4LWSKIQBpSlW3Xr8CF0
IUQWWf2UFeInNx9gYU/WlkRF4hi78yO08085VcPjdg/1Jsh9+XqDEQFkgPlIAarf
HaFZQuDhXZG0S9AVFgGCJWLWlFGt6PdXdb/1/By/DUkntK4tCnbUabMBTClvsjoj
kZge3qtVcRo328FD27mchKoNLCeCQZ/tzr0VMDrI+t4+5ui0JLhA/bYrestR4yT9
5PHMhYndiyxScS8AxwRWuIyfRE7IOtNAPZama6q331M+XFL4rNM1xO+x2FGj8ojA
KvUCCxf3oMUhq9TlP8iqsidHuOwedTvuNpgAuoJkk8USkfOTDx1hjKXkc24aQRAk
7zOab3DEIQtDzQvLqfQGbkfqd98bGlx04nfOdL7RZqxL38W47xPtd9RCRQIL+6LO
Jk1huOA1z/sqMGXMrEITWX69bqityMuf/M4cSSLUI3eAOSUQHp3t+rPh4yaDP+n2
M8eZs1cx16rT5WN2q/pfK6bylbMVPH579MJznQtEIXK+WTnCgNQK7E9ADXXJbNc8
Qml2hKYR3CFi3wQkh2fDOfSFgNclhLM+Gvd0WaEgRWopjECeXH0pw5r/R7rPUWE4
XWAuWaw4A9OtGdgTt3+BfW2gohZmvTiozHK6ahjAG1SHPcXLGVh/+yzRpivVRNNy
UdUo5bNzVBYL7TL34Tz7DUUR4qF/4Z3mccEhWx6qJsMRUYh021phn0dDsF089TCB
cTkYHAz0tKp7E6BBYdl1tYnrvHtsPqJaalIxmP8kyjsjewu/Z+FwmA7ZD1RJtG0P
mNccSZhDi/7MUaInqn9Uivqb1ocQMCFN7Xmfh3lRJYhGZsRkzkSrxmVm+aVf8veQ
W8bjhkfbRcc3ehtTQjrj/KxLg8XiU52mbTSyzS5vH9NvUiX8Eoq3m98gT6/75upE
1lKtSYjkqzUIAdGoKc1uQnCOfQymDPewHKFhnv8QuIRo4HPJefyqMzqfRtI6T1x4
aJUZCP7hyDy9Ew0ffX3DtI/oU9Pils6FvcpyCuyrUSGCwkDOndJsSUfJplKty0EG
fs1Ppn5IBcjpnwolFFVogSHs+4REnxejjxLOKvsCdhoD7gdF721dqQXyfdTjyf3a
VJjamvsYyvjoSFVjI7Y+XB4bDZf6cdGPdPcUcGqjuG2ZDW0acAxCJLJ/Hl8lWW60
fsAHFG8NjWMJ9ReLUFeRgSX4K1LIO8w2zMIqzxb03d9U30b5gVAQcVNSWdzFbX9+
hkCoWZLH5nVkXlBRc8IkMW1pTcmWbHMUrRYhDkTkU9XwWYYlVTyrBu2FXZbQButM
SZmzITWqJOXg8neOiyB79ghsFHLmzJkUCHgJBGFOJ2LWeRrHPL+5w/XQ2Rxt0xyY
PuxYpeBULSILp15fZ00O/PpKCZBjYKmnaMrCeY3u1L8acM6HTRgxegIrST5NyVzv
AXEKzY70Ot/ZJY+Ou7FwQysDquMEC7KGUR61tSnFwfk4yX+e2B854FnPc0mYJ771
nwsRpcOk1ICqJBh6DDtBmNFNXgrf/R70b/Njx7RPnxLkZGIpjLi/nwSzaZ2CP7eW
cZvTRZiQoGnh2uuZE7YA26Afox0nC6HM/K7sbTvpkw1f49mAV/U0oHg6uXblMWz9
4uzcsCXrY6v0/YUc0AyyMnsSUuaxXj+6bcHceEH9dItG2l2yFzRUy+79uOW5udN/
jXd9gaLwRiil+Usq0xBiRWxiSSKnsfaUBjp2b0WTyird8HvCXyag5VKp5DTc653p
FqltnwsBTpd0CAZH6DukmjopYvZvC0jtxwMe8533U0WEuBNg03SSZCm25g7vaTrT
vIebBY9kOV9ReRFvGp3N6g1e9n2LXJ+9SN9z9eJZQAAA4Rst8dYXJxgs1RmA+mq+
Q+j75OEE9F4qqVXudrn4kUPQiY1+36nf8K8JpwS4egEqZ3J6T/BQyl3eebF3R8S2
tiyb/6fJHwsGAAmztrf8gkOz7K1u4X/q9G15W0o7zXQrqTDEmcPrijSR+zpjWkGx
0Z4/bgl8jkClew3E6A9fQ6EHQ+vZUiax+sf6AanaViAW8QyLXR4UJOmlBUosKid3
rma6KFfzLj/Maqw+jGeEFwIfZDeZqSk30swQF5yiHaNSP7rXWcwe7+yR+Er5KeB3
0gqCdhKbMyfV+r50V6CCJyGcI4/q2VqM/rqUwoEn+lqpMJFnYWn3+sRtX8YnjM/R
gX2u0YqH0sKw5fbQ/Xftw3snI1VPhGDt3rxEKuo9gJ93PaO79tL2zoyl/DSbwgOa
WOqc7mlAdKzAhOW3eIAlvAUQvFQ3CwU2kIOu+bQvnbLeWz8AKnI5LM4bPgNOqeiw
knb/5NWFdS3W4gDv1c5fW/SM0crz3ReewwnzOicYoiCWaa2Ks5hl9CUFIgCYtrXs
4K4UjDFSvR3GNwxEI7VLOB7X297KopNJnSNauCiPFLU3SSQ9TAP7rg1DM/xSF0uY
+wXyiPGxnbzXy/eDyfw7wn71uvH6C7lwWisH/OpYjgMbHa53yYRWt9EQCbRxVyfu
Jwy+nkEcm1QmcaPCf+vf9xnyPHRUjjXGPlRQ8knVHElLsraw4JDhpxhITYG/g3sw
MGwPaENTLr+26EY4jLLBPgTKkAIIqvHF4jjtPR5adhTNm5seNg9WqOTvTMinOsO6
KWKSxIwvqoeaAJR0uSjJZdNUkOscFBhGnXp2aHuIjgvk353jyKHQjOPSnUVahCxg
adYX1DlSEsm5KPKRUdwwVERuKK8A+HumFaNQGPaG9ychWHu5P1X+9/oiueA0Mlq+
fPEo6lI5+3CnVB78cFF400AiLK9YriwRvm4FxDuSvRY3cFyHM+QcJGj3DawDkBbe
lkA+Exe/AqY0wFM/TifzaKpRWqA8+VXUwi7H+qCc128/yErUcbBr4RgEZsYuXfmd
XcVVh+sx4qOcpl1btfpY/Ye0K0b03IbOX8Mg0iXHgobt3VNyQURzWu33exZ10hKJ
0KM3S5MGZWmdcc0CluhXmPtW99BtZVdld5M2YevbThs1s+c7tND1E6UrIRc9FH/2
lLZmcSeklCehyw+bBwK9bFXIdQuCBa/cZBF9rv0HK8lP/xXA01phUiUv2DtwfVUl
UlShRV6XPOfiqFFEwf0wvCbdKDrr14gV10KkJr1o9F9DK1aj/b/cMX2HlTwvF2/9
Tz3TAtkut+kv9Lr8qIts8HvMaHOYYtfbJAH5VuZa4l12FBrd2jdtRDPqQraSz+z4
r0CPIHy5mbczYOqVjjkFg9AM0ipYZfTFh1W51SHP/hq5KGjGK+nsmbhZ6W0kjgWT
FcU4oUWPfMxmMeHB0zTRrhMuur8XF1IJARXTWWhQpHTZ4S5dEdCFoOzzWCDkS53D
1jG63oOEapMBJAbahEsEkEgQ0zASlpvmCSReQ4xNRJLuCVLRcb+y7Xish8jlEphR
KIcyGQBYNxXps7ytAW9eXV+OFdD832YJP6MKlATy0xFYgVsUYZZwcaX/oGOoZjYO
v6ut+fr8CDy9RkPo6E4rSdLKgNSmG+KwnUXxrLcGqEYjnjuzWEnCfk8YzePnhJCQ
S+dsV3CpK6aPTDBCJ2JRwhck3jCfDiI4RDPsi+D/JKxG+ZSa/dsyg/XcnAd+ZD+J
W3RN7GjEnssG6GMIQgNrTFCne+//LbO8Wqa+h5RQcrGf+xTq2on55XX8vugrnMAt
/IdsyLY20qpEC4qbdoIaIKxdOVvidKMuHoLN6ngyspdgpP0xIEqcN22J20JcHkdl
lqfuQXJHzd6gJm82LlayHYor6NwJrIQ9JiYI+xm6d4BI5Hdv9qa0M3iPoxVOCyEk
E8fvHEPKfl33M3OmUW1qKuCVHvNjpuXn+uc4uUHAgum4SDCFHvmEiT7LxtR+2SMm
lEY3glH4KCNFac+kk8cJ49DVPRfSBy08WiVexU5vac71WcrlAHxXm/SW+3MAYMTO
rE9b67cOlC5z3Cl9QWwXWUq3okd1kcMI94LNq2FdVfWPCuO7HKozDXSpT0jNQAOK
zMs3BcZovSUqrezZCKOb67Ouqq7Vmt8oSoNsj+6Wx2GXl0Iq3MQiFYCeyNSLzm28
9139WyJoIW+HyFaMFzSOXQoRF6Gc1NCeeZmhc2GVyt9R20KWIOe9xta4FOIJnSNU
zSg7LlR1tz+rLLpq5DkDw5UcBw3HoD6SeGNZ8FDKFs42t4vGQRewoaPY43qci2Ee
tWtIneCVBU9dUzisWA7KIzNgM3inepWJC2UhKh0c7gm4DV2/Wuz7R4H+nDHNSQU2
yAbfQhAwaapc6mWMyt19knk7BK7ysn3e5s2P7Ux0WbqJzJSHKjsan0lobmtwYv4I
h8u3jHhOf3U2nNC5B/sIuvxzQWRn3KEkMuplgGHpRyG4MR0FD4t7J3tix7TeL5WI
K1zPTG/ZDcR5j4lI/+lHiwRIRS4OB50qEP1uL/N7ZQXXRHCZhEGa4VHeJCbcYRNC
fbl23E4ZIdXB7O5bfCi69Q8jlJKOUQwLK8eBezMWwSQS8gOf9ooemcIM9+fge/d9
I7SjioVpZYlovfmSTjHNBjttfLVesWJeCo+GCdAqi1iyxxAKXZj9HD0eXVF09S4f
XSsO3TCuGXPLNSDSEi3TnhkntuT+dQ3XEmuLQFOv00Z+201jzMLCzpfLLb8xp/tR
4lLDfJgpBgW8a9DWJElH3qCwcxI+biNe6JafXQOBx8Xm0/nE2SH5mmmmj4NZ5NU/
2OqNZbofEjrNP4xNCsI4jItv3Sa0WP8eFZE6rLORstruOKJEsFFpC3XiKBWA2OTX
9EvMcQV2ZZIoX/GkwGtBTkEjKvo+AlPWCOY/ysO1PqckG3aOQhoC4gJQSl35MFc2
w4fbVXwWHN+IUNcww0MCDvHljSobE5uZyOW9ddgEQAVXu5mhLDs81x2Mj0Dcbhkh
IzNe8+3Qgk6bVklLmxXndYlRNIrj2+i6oQldIs5rjMbpsOH9orWlc3Uq5AU4tELm
CnKcMq82ZtyZvHjwC4RgZpg+Nb3QHQH54W3DVhrA4MO7ol5RAJpD74EpmCX1Rgku
jCQaHT/v4ec0pISFKizeoUlHOfCjcJrKOvZ1TRJx84j4uv+FqPfkwIKDJxvT3tU8
W7uEfXQE5Hb0i8YJWzYxVfAFOxJayBWaR0xEiK5R09j09hk7KqAEPqIYAQSvxcJp
LKzrpaAEXbT1KTZSouQSkYwaLlLzkGJzbkdEIIonpMD7Eo11Iq54N9cnSv1WSTeo
cpMQYKKT4eoQqCffiCfLIqyqyPRmlw/vzsBHwvpACt3PJEpq9zP+/8VCclavftvS
3j7ttfWLQw7R1vbNl0rscpr1Fbo4Ze0xxKfTjcFICr1krc6cC5AkikvbcVtuOA53
Y91GOHW7cWEl0NvVy67WrijGSdBeBJ+42f990VK/AtwLw6TclQGbtR7IjKr8qAGJ
y5KLMYGOOlHyeqgaO50CCYs/9jQonvwQjoGb3q6ddzwQjiZCTCFWTTBORhj5TW62
8smsOHfsnDk6iUofYOHHq/5SCBQOjUvepc9FaKBEtQWd+eh++XemowOEm5qgk1YZ
pnToI8dHZ1A/d+JVeMyJDlzAofgqwWDxh9aHS7CGp+DE97oMB84lsrzCnCz1ltuU
noO1CcGcV5RwhjNQ0NuoL+BHbPwH0pE6OvU7P3GE6fKgquT0lrdzWXvJeez6qZcI
PJGX5Bb2osfLezO/9AA3BF67A8WhdlvaeT0OV4InBUVPaq3EJ2iUF0NEWhe3HvAP
ym5F75MP9YtAAFV2wPXWZi4AiI6Si3vl3AJX6XMfweOSAdwrX077ioxOb0cV8zuB
R8owpyC+5x7QvSumhv8twvtmZe0kB+w4DIbdzVPEy3eyKRPHeHMRzuDyDE0zGMvB
edidZk+i/Jv4BqvdI77NtHXnQKOF6YQVwSLXMvB6t/PxZ2XB0mOAnqawf329rBPb
ZqeT4j5HUwkxLOf3Mpx/azPgJX2gnkLGtdRJ85OqMCNVv9aD7Bzo4zytxGes69Uv
fZNq2Dbpf2qLU4+W7di5xBANroBZ/ODUKwRne2P8H9fKGFpsGx6WkGtyPHq/7mq5
VC0x6mj3ODt3iHpS5cVKKg5tStSTaLCsycqHIegGwfe9P0NbZj+OrimSjdY+H34K
HFKdJYEOafUEqxXUYK8ngv5L+AvDQMbLPuI+hHDLsZL/yNpaQKeT54Gg2pz5u+IX
Y7WXY9bGppcmMk7ec2+bsQjRgpuTgCAaCm7qxeNtgsF1dDkbq+yWgcE8D0mQw9eP
v3XxJN+IaJoj+tDn99boK8s6G+WgMvDjiJSySX9ygFFBm+raG2f+vIO0i5XTfI5+
cBEeJQLtAIyGO0frNKCshlBs9Yw4zYBmHaQlBK7d8xne4aVfnWb3pXbWcjzzMui1
JEZ/GMl0BhFikMlwih8nFDXNTouHOWjcOilfFv1qu7aL4CE769668pG2DTVCXSLs
4Ku8/eK0RXRir7FAp+Ou9/+dLT6iaA108Ves5uVQ33pie03/RxxhtuYl4/Vyxm3J
1ZDxaq4Vr0Cs0ZW/5jep1ZUwStJS/ygSqwWMV8hyExpbg8VtWAO4DJ4qs6+fiDSG
ybVQXpYssDLdwILG4BbB52p5aL7bEahK7Dc/7RLbYTX83cLhaotnPwl2+WfanBoM
p50+4LINwQlzvZktaG5VfINM0bOSu3LFHBIJ3mzPCoTkUcM4SimRddX5QSV6/mxZ
xVbkbpTWhftvDI/t4hTbGYjzvosIkHRY2uLdMwGLuxPkoiL26nrVWY8VWEt4Eg4O
nhO2L+YZY6besXd8TBu1iFYsNceCMlnBJsk2fyAfO6H8LauqrP8nwvYdodXs4XXb
sdjTVHawuSn/0HeYUcP6oQ==
`pragma protect end_protected
