// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:36:54 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Y5fDXS88SAmYzLKmCS4FW9r6okgbvaYkwXtH8IUydvBW6L578jpeU+yEW39kvMve
oY4dvrYoqZPIURRsgyuaxoaqAx14pSYchwH8wy8PoC6AnSEFiYJ0MxSvYIaB5+z8
BoIg9w1ZqMosf+iIzldVUSGPn4x6MccLNVdcYv4Iw9k=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5200)
gNd/yawfsQY78fE2cTFONhPnQG2cKUn+vpt8CuP6wV2PXcqEI4cDsBaoxDt5SdNQ
tgywYLAsu9RnnkGnLiVel40sY/tjIiIRL/KekbPEJFQ4cHnWjnR1suY6x+e2zegb
02Y+sqr3H2fpBZRyJODuJ8D3+mHA2wCC7cG0V8jzal+77WKWxo6Ot3JK9sCfwEKl
zCdTOH5SvIfpn+0ou/aMLZ6CuCzVBuxv6ds3NqE4p5xe04NqeyeBpx5uBxF3XXVQ
MoRJL9vu+pxrLamasPiL/NJS50Y6qmq1XA1mKai/lCF3iqoDGAP69IGf+y8jcrCf
SHvYGzJoCuZFwl3ztSneL1bKy4T8FoQc+boEM6I0cZARstKHVgjPot8qf6feN/jF
xVf9/vQ1vqzposBY/i5+UJjqB5lPWl99V5/3B+O8XwJmVCS5tFr1rgxHuArciEXM
DtyoVE0P8MOmOT6pLVV4WyBFwFTEkanGYff+000/tf8tD76rKlw5B2flkv2bq0Br
hMJf2C9xvUi4KjyuPvhhuUUnz/qJx1bm9oTdq6Pl/dybq1Llqnu4WF2MGKx18HJR
RNP2qBmQa1A+yFQplhs0viqiY/QthfsJJMZfh8Y2GGLCBE8VKXqu+5PpRirCBDwI
qy5kvvdjqAm5+jLBTK1PQsFsD18ikstMWPB15zJyb0imm/EmgMta6HfxC6kQeLAS
1Sua9A5Uwa4UjanKNgdEgtaQLf2WOizLgL7IPGia9nf9vTB5B/CvJRsC/WJacGLF
BN/0glS04bHNixpQHnwqlxOiWUlM9AQoZJT4/byG7xQUXfcOeLiMuvshvOS9vozm
EHCDRCTVlkE0FsHI7D1jevCF6W/zVI5A00KHqX/PSFpvOURqvF0B6zEHaUCrXf/s
AYwVZPX5gV6GkkKwrg4z14EtSDgbO1gpkOt2ePChuwz0uRZesCrEtKXReiYqryMY
nZJah/SAhYSfV/PK1z2KFlPfyp9G2+598gdU+1tWak1yf/4c4pNVtyUKGi4Z4iq/
9qljzCRNEH7quUEdYSdV//Lb0cCKL52zmjWDczjC3r84ZRDhlUoh5whO7IhvEQ84
2YnHnTeh781xzrjHDHqrsuoNs4GSdCtL4gv+HNvacmL1WyVFfmVFhEqdV1G5oBD/
JDjwzJo5cV8iDVcPFHFs7SmR7EOqbvSAv2wcsmZ++3rOqfH3qwnfvnko5e1m/PsP
Jhzra0tleZkKhIp9ac7TW4Z2B/ucNS94JL+bpCmZczfAkI4epqAgyzUwpVVdFJe6
TY9DPc/SIlZvEQ4jybV14wehUQGM+r+ImANaE1jCfwOaiGChFFdYlO98tGxszMJj
UtKOLEdStYIqURwiMi68vUkgRewY57XSMiisTmwiUM/Xg39mEmJPAMCaeFpUgLiz
QIjA5PcdtlErCAGoV0Zs/jcY8tfpUpLTy9BtJ5CERAn7JBQXu5/5+FJVG/D7nFcm
QulJ7Hji1BICqO6UGu8/lpJxgJkP9gMLtP2Pn6htUSJPi1ZY6PdLB1O1mrfm924y
qWuE3ODfQhXU3a981DhZ99npScvMqfRtdwolHEFTBQIdlrtblHMeltz/8RSD7XwE
OgkLZKuAF1gy6zp1VkmbO5JOKkMPo6HCe5NijN68iOxfXakjL8Te6WuE3dpra52i
z857eVZgQiVDuXQSl2+3cL1yrs6tYvTxMDG+yftdDq+2QmPf6i5sWoe/o765Yf7b
HTY53KwrGTGDrar3VpMOOc2FiP4OR8szxV2TvHhYY+NqaE/LJKtlmBC09DCa8rrW
TsfnE3mPDtEhoDSNKoRwlyar683tZVCK+v+002KL8mnCYS1kSqBKCsTeGS9roziK
Zn+cJcLEODzFd2C1Lv3xlru0AMrnpIUtSuZvO6NJVJj98OMOAEBDPMhZzaFJQhvD
GNgMnJh6awjBE/lWWY/jvh2sHoUTTCXHuRhJZ9Hm/P2poFQxB2VHqSS1S/LZT0r1
lcrVaSKFon1tkyznxxOCWXT0xsJC25DDDr2rKcLHVu6INbfw6UPXhGURDCJuOYnt
p4WtaEKz1TQ5uIqfnSbB3YdEw/0auj4KQx0BLinYUdurt1Aa+AsK95DB6uq7UJsO
+1qoTGpeJCHmELVAac1Y8t8KbieQ6zoYEkDkpUXAb9d+pgSzWZEFbMtqC4r1ZHcC
cLp43Hrw+C+70EqCsQDFylP+rpW8ESpUblPVR4RhTaO4feW/7oeO86WBDuf1kg6U
rG0wuEjecQdu+MVTg/bB9FBYsTTBFZb05BDXCNB2TRCTTjsTWEob11R0h5AOoufS
rmKj5LzcDrzcA/WgoOu70fDl/503YKs1SMyV9M9GqqVUQK5zWRmDrJPjSmcEOtfX
s02J633LKvhpsbNbZqFKJvSiOyqiZklHFbaaMPZQOFqJqBsdpga283+5+mwAXASy
QRqcbpUZYLTR0kfIpskXzlM7bj1LYzG8ZSNLQgRLfjmymvrEisZ9vevTOXVr6GrQ
VIklO1Wkga9xz4h5eJUfPZsUG46sjdAwzPJYslp/3n3Dj/3/bfbeBPW4R5ouW6RG
nCfAxrg2B/aYrv0UytE4KKc6e/MuiGqSC6hfU+tutA8moKnBthWGfSQik1PH03wG
QesHCw10F6s4H5qfCTiqPyU1s2TzOv0f91G+ckl2PbYGdBIRJRFpJrS6t6iljhtr
5+MsfskTS4aRSmggXUrBi71ap+Cg4TGowopsest5x2lmKxTSN42dKJoyT2Ga2sT+
R8/k12FZje2900I3BJ4HRAaYLjTXzByLNvwPc5S/KXXJ6vE330bdni94hv0gxBQY
f6QPrhSJ2I0ueD/ORfZkciD5M/EQvcDTr7cCMvezMtoFTOxi1loXLE1HWatJU+vY
iHAk5NYpZOBPzlQ2laNAypQCYGaaZ36ZJw0jvE++oUzqUQyw84JZiofj71hgS3IH
9tI/mTjk5W2U+z6jHS66pgSsl1p58ungOCy9jWTfBKIvAqVICjsIoJtZYMWJDb0C
mL6qX53NTHwxEhuQOiNE6MD67Ai+/bVvGfEMqY6xt3U+gkdidhz/3VQRoy3VuX+v
NtZOJizQZJDAAb3Tjr2iAjvqNdNSRnSxsNUaFix7QUcA4EQRhlz0TxTXZRA10gHR
ldXrty4+mh2S7LlPfJuhBJ6TReA9A4IvCA8pu+hE+mTnDeUoBT1SZL6ZC/zqQZOD
Y05EaKCkvsrWDy6AxCmtHyLw8j65vYX6r7CSg7wpa2LIk4g7E98yYAFr57JH8JZB
AgwjcE6YCihAqe7p3rBTlv5IhyFrUsc6s25VvUV5ymRPO15L+3C2FsUYAmGWPiCk
i6tUgWsDIHZuCkAh69I/k7tXz7Uk8KniEVBnHdKDctQfTOpZdo4Gw/GiACr2i+gK
Si2tzp8P/ppRAVCaUVxG65e2ID1s0MFp6DfjsxwjUKIB7mF+hFVn4LEg7UV6xEQk
BTKu6XkBpecLiYCV7LTNp/jINa+FrI4CuKwA1SfrtRGDUoK6R1/tZ10aIfMrP39y
8vdmgNCvH58zW80nZ3jWCZgh4urP8D1KIThFIFlwzwa/5s6frghz5Q954FW1cVTr
WzoorxkjTSgm18T6iNcucvzWU08nzhRTOhmgwbNG5OyVkD7u0bpZNjR2VZkQ6MPH
Qw7dGxDFxjVD1Q4HERR27BEzNSH8/dXzRJIAqzh+fQ4Rwd/JYam5RzJbJWewB8x7
58COXFDcbeSjn7bSmyB3J0YVYYEeGDQFYePY3TY3ndPucynq+bLJ9ruV1eYQlvn/
MsaEDwzdpupWHOD8lI7wpY0AbgIgTo02zKLLLVtRiMiz83M/zj7zIWJvba5k4kbL
XF73bkzd6BJ5Z14apcI/Vo2Ucp7MwAYjZl0yKYmoGjaDu4SU8mCdcDtPsPjCqU2Q
6RiGK5rEHPG5EaDkpnUEifzwINFiDpO/BcgNIBYTl/+erD/2NUO5tVTkh21gp86P
MUQo290ruQRAZC4ERLxyrI5vTI+GYy5EVBW0SMA7+grsa5HC65w8PxNKKOdD+p1s
+75f0wXmiXKrc1tjIhf3vf2dHfjKA1HvmNYO3EBS1vyDhk9PJmTIHFWYI9wyrlwp
0KywQKGGE2hRdzOCkRai1GxsAthi/6mp53mq4eRchc9u7I/s+JZXk4hTgQmcb1CY
eEhrA5YyVdGndl8+7uvbZXmpk5ZLttN0MGJSsEbEccGrNIfPXGcDbHK9vweCUDqs
y59t/OvJV1fQ8My+0XYaj37UdzVp5+w+NdB3IjoiLDAS1hC0GEgngNKjluzE4Zzs
tABHCuykj3sIHDyAvxPglpwv/bEVCTAHi0Ze7ZWH3EXsNLTXrBIkN+0+Sz+LbGoJ
xtooia3+BhcMgJ8SKabUhE9EZh1pdmBrBkMj3o+5fL7SLOGHltEtX1yKVkozLOXx
1e0xIA4ZAL4dPJQ02Dlflt6OEwxOa6VsIXD7OMG2+n6h1sxJB/gafVQgYoOfmDVd
tJqbaPso43jcbPUtWhAVSNJw1XBh+b1PnS4sawHEK12U7FgdXM8YEOM5YEFc0aPb
9i8662/Pd9ujS+YvGf8vtpNsYkFhA5ASAf1muUwUkkjVGKz9trTymZtBhgTNfPeX
MV8Ih9CPHt1BnKbPwlBY/TI1NHaYjCLEQ2XK0MaZimWMVga3TgwlsW3a0DTK7hAV
4ZhlPamq/eX8KUqqi3l6w+/Ou05pTss7TUbhyWVjDI2VDTi/qNciUW7sxwyoWEQt
S2zLJCbVVJEr7ur608+2cVgGRcz8oz/7C2IyMr8V1+kpOoHc43BD3Y9UHARc0QIF
1zctotwy6IlIezhbllU8YWofIompHft9pKPpwmBO16QrjJ4QoZZq7o/j756YRS47
CkEwU9ZMmfIJtxc2FVCAtxd4Xzk+0D3LvVqmv7BF60e16xPDRnKQ0igBBuJA4vqm
NxzULHedybKW1YybGv21bT3USfpmqTAoKhvViTpr3Vl8RoIbL47gLVUzNV+y7J4U
/7vjDh/fPzfvoD/u4bfjSMH7ly/hfrJtEFwOvTcns8DQx5bq0hRYDwXAfl6IjAH1
6AptSAoJa0zMkO0iPJVrrGvzjo7sRuXnM2xUvz9IqmL3J+epv2w2Zq4E7yAfhBVT
P7ckTURGjmlgDUw/zKL8ZWkGdP+88phfUzvOBsxtBHqytLZnHtH0fE9l+G0hCWjX
bx95kQzK5tarNcS9gfU1oNF18Nai8hlYxBDmvLLT4BI/SlCnohSP/37p57fWDv2h
gAEaXQn8ipyteVtIcJhvifeT8ZH6FLwbMWG/m7ZoxGP8GNHQj2BKzrH56kWLuBZP
RBbCMepkdNdzsUXr7mePWauMbBuBbCpcSxmbgdHYyRMw9I3sHCV4grOxHmZA6iWZ
AwCLiIbNx4WZSxJT2rC7TL2QrVPlRn5pVXprOnjHfRle+nmQgGuJ8Yq0vlF0kJoA
pNFodyaIjUMYHD5UrcW7TlwnYuoJlc68eDWufBYaWnRVNStrZphBfHqhV4PmkRmC
/ICPLZkH8EBVCRD2JXg+j1XaAfRF+v8gsALRglbKHFYRdVAOA1Ots8ODyoKym2W8
YcPnvA17x1cQIBPQKXNl8R8Y444Gc7xWlOVBK92//4DIlpxAbQDlIz8OTzNt6saM
8zRbv/8hzLIJn628Jjoe7lyqxsKKDsDmpf+NHiWzPNo9ldNl2rrvwsEer8fkv+EE
4mpiznEovVReeY+WOpQ+PPi+Wp2G4mKsgJJaX/M5qZANn6gnSRnjeHyquI+WDg9U
OxhB2O458tcSWg73gzuL6kZxHpX8tCzMtOfZuc+X4G/esn8fDDrAaR39W61SIKHK
Mbp1N+18GL4YkBiheLsd33vnEq+8Z5zXNawI5eAeebiHiqp2bYUggD9w6knl7KBv
mBZarnzD9KB3LpIit2o9gVj4DLEP+3CX59WRwutC3c4SqcPLCeXYMjTJmA16etRI
ec6pbQloujisCe5o296rsESxnXlUoz3GE1sexYnq84IezKKjN2sBNJW/vSnYqs2P
IupjpHuzOCGdlULDZJJyoL3itILeyALF/7VHez3yBfDNFNbGjQmym2cXPexjuA3/
5mMAuXl/7UfTIp8H9dgXj5UXIz0cjwBxs5jAAoJnhoi8jlSXhgvHFaLSrPvOzRF2
k/3mLUEKcPMbb6X4g7NKpPT8Hpx4BohzTZ0GOqbxN+1Hf+S/9i7zd2T5L6G1pqju
puHfX8x2o45fUABhay29sX2NVXywPB6TW3I+o9Y1quD+d9Po3+BOxy0RcTY1Royd
sACKNUiJdImPkb7u8PIqPTbNvD9xg56QcsXYH/s03GFjeR/fheMOSy/6XXpgGwyL
Zj0f1KsLrv3DN+SI8tS6EP5dtvQZAFAFqgcBKT+/AJeTh1lv1So2ZawpaGpGqPuq
gcRz6BmlZ1mH2gYiHm9lfhmAnQM+JDi3mxzPzA015h+0CKiBRv/BVq0g1QZzhC3S
c2zEdt4lhOvFy8epWD9wJMQ6QSLyHg78VyixTg9A7qAboZPpeehVMKDtUrI3MTgT
vjqjIZ2RmHLTeJuGnPVKYsFmxjnRtfRbUEg29uttBetqoYwXk6loYv9CMovQQVrY
qVX61SryJe4oXqVK0MV5y7YCMgJTvBtYRN9EwYK9OqnhqrfZO8ieY6H9COY28aDD
J1mR2aH1/NMi+meXS3VfWYYgNCvr6hpJUgl4rLEITS+anC/KpiQcihl7EjKjD62F
XJF9FUKbGTQdhRy5EQxjAdFYSFtwczDyQ+x7nxLOQpKgL8EGzooMlRl5DxspuZXn
/NTPtjzF/p861/tikl1p+wHkLpAPGvFuqBqZxXw/lpz7cCKi4tAdph1kq5LJbMNn
46y4Lk95DuNSDdZQIuTP2Zp0mXaZYfnE+/Tvo1wdPRRbME0F7s5Q/jH326V71ws2
cLc86gz0jkYjeLMUGlX2/A==
`pragma protect end_protected
