// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:32:41 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
t6o7cqvQLudiAyQIjQ5hJWde6Z3NWSbkU4Uh/IvfYQRFkWkQyW0aZaBreESGi2Ul
Mzl98fU7Ghwe3ntKW8WGYoAOdDiV5TTjol2wBu3v7XY+Nt9i+l1hMMvQjH04zZbR
SWJqQAjw86f4RTeOMDKpiwLoJPSKIfupNaYR8ZdSFJc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 4848)
G3HbSCt/6WCv69kt2xm2YtzvTtz6o+nAIdJBaU3ViN7dLwdnC8Xze1cT6kbG6QW3
G0/T3GTKYOKCVS1frzj1Rzopsdu8APgNjaBwVL3njCapS7Ayzgy28Hja19/Hjege
NfV7zGfae+iLHrxmkWT60HPefuIjPv3N9i9d5qW43C1OhFhES0KbwP+4yHk/HtCO
d+HPWGmTqLnRHk3N6oJbahPpI0n2wlvXgTXlEw1l2NiBK8bg+SRM07Q4CcW8yNwX
jB6CyC2PVYYP+eo0WLBajrW53VA3oek/SHOHr6rUevqgbx5UfbcGTfSK+mqC9gak
iKhrI0KtEsdwpHZoJKV0uPSgrVLXjjfdV/PT0EQcHKmY8B0lgKW8EtLUsPUQH6cl
P/MVjBCGRFacFBIexL7YtpyGhmH6g68cA/Z6eJ7WyalVKZ9EdnxsxHSG7q6my9Qo
8OeBiCXz+yzeXJOARMaqSrxPedK/mMqwEklcxFLfDtqn9/EIvIcqEbcAE/yqhxSz
qcTmzi21zm3EyOxCoGC8YjBBwsOheaGdA1wfD5mQvkIPggEiXvzKwHdUXVKzrMLw
DC8P9fTdqkxlBNftFgCYnnwP75BQexrKRSsqCWswN5NJMCZJtY1P+zpIcDd36Wd5
o2kcWrbv/dEznEvbcSYw11ZdUITTGldxr+ZJU4fX48ZRYTj60CrpqSdMSrwriGyf
W6+j339R4HQp7DHQDnZKuGeeXFNv9JjEmMfsI+zOZ8pFEOfmrykEYERGcAXSRDdL
oDJIJmrMwJ/gcguPcA32hw1AjNKFEXW4yVbjmCywtI+Hs9se8SwsPE1Vsen37+T4
cRn3kLWTClx0PPcYyRNCLrILP6bI/IJLwBNr51Hhn43Tp52BXlOffXF2TlCFLYod
izbQ8lRRKZsdjreXnLcHdwt3amDRSxJDZEjxeA11SQOY5jbH/wXjfimjXNg9He+H
06Zm1SznHX4ifG9XRHMFqu8tVd3gSoVZon82vB5rUSlGFsozDXv7cbuxB0HGAKQz
aiGRNHv3jsn8PcrkahpvLT4FjFP4Vzz7C7b2VRUq152nbKnNGKHcZ7G6iHMqlzbV
+0Y3+IkIzC6MA+HmuP9Pr82EBpEqyyAJZxoPtGEq01Xy+cmo135x1ckoS0g7oSuw
PPgQ1fN6m/q0yFw6Z3r8wJIHB9GQjBvqVh6vU1xr+4nJj7Zzvq4Y+rZTpXvg9ZiY
y9KoV3gcO6PyUkyxMqxWIaVlBjIYL+gSDXxu/4qNZoPeF744cuuyCTc7C0sT57Y8
ALJoWVtuoxp/rtvpmN5oGSJ9dp/9Uo4dQwfhT1Gyd0sii2lNzECXa+VZtCmdfvmL
/ejrr25TeeuCcqQohQsNQb//UMUWo9LzkB9gr77fBiVzXTmmTiq1bvdua3Bh7OjJ
2+WKaZbnc+h+nGPNt+K28Zs4d4EsJghS+uIQr3Soi9riwbLS77spWGhvPKvLoVow
eGduui27zE/+o+8f+g8M7bEJorCv5hEPGPv9xWg+ovzOGRV07ui8pRtWLLNo3kLd
djbTQWEK7Qplgwo+KOKfO1N4fDKWFpzCEPeRI8jeurUmYkpXkAEjsSpxA29izQlG
P3jAZ5Z4uZzK/90NwvrUlhItyCAmx5/zJbkirn5q5nBrtK+Fc34vwxprroDmHflC
qd9meOMhMGpGJGCwNf3+vAD8xVWoFOuhVVaOUlPYLTleY6+aZ8wDUHQRcDQrPUVF
TN4C1edEhbTixQyAEjZd5LdTYvYV+g4EplWB8W14Ef5ZaCD2lQpy5cWw3qMa5cCj
fGAWxQXzqF2/T+56m4UjHnR0o2PfyO/AbNYGn38F3W3gqRcslkEFVUyALi2+Vi+D
davbEpCnV1PQYPlYv1E2Olj1AA6AgSbt/f5MHpcrF82iROac5lCoq359Z8ug+OrC
PDa1kQFSQxytY8L8akbQrl1SZUCHe2ai23YG8y8uqyFD87+QYtB+4Al9FoHd8OIT
Kl0E/iSPzlw7vXxGxT9arlqZVgFkpJKf04BWSxqyIgowFnPHoqpUPuXVa+m456Ir
sRrZm3pKZh5Mq6h6OXhPrpk7pJT/b9eBDW2LT574xcusRq9s699aQFHSyXn9E2Pm
ib13Hy29ejTItb44BZqHKdholS0DegP+j5CeaBYN8rdVW8bmdX7TZpjLWpfVD1by
iJtpneZ4+Wat7qBi5SCF5s8gJUQXQnU9V+JfaJpGgAArFZhd48yfwRd3BzIjMdY+
AYNSdLmIlI32cYYQOF77QbtWAsoTec6hb5iDV2qlPEpLt24tzq7eMOU2eo+sgA+q
d6oQY+1afY0bqrzeFdOVAgQgaRX6A0t97RUSmOQa/PoBwUb2VJ62SuQcESYFLlmc
QATptNL1pEEoM6mvuUiR6NZMvJ6tJzvSHO7Bz+3ew2V6GtDOsVqmFnZtkur0pIJ/
O4YgKLJdB/1xe46gybIIfNqFe7OPysr41xuv8oNB7EG7w9JCw4FNFplAFqosgAt2
Zisasi6d4GmP3p3D5l8pYTBsWug9wifEhDL5VbV0hX/NqthwbRdU++KjPQiN3BJk
SvLmadQyennyWY70T6G758e6mOa+PHjN25LDj66eho4q7StDG6MYl5hMLC+Dz9Tj
Au282vfsIDmaKYkO99IZeJWcG23FVc8LR2+AAXvxgJAn008gEr/gITg1vIOJtW2Y
fh8ZmlzxaQ+J9ZXwzxaT5j3glXO7D36Ofjvy2+6i8A0MZ3YCv5h3CdIbWB8/qV2q
EjD8Wxr6vnToBcrZ1TnSM7fj9MtlrGbl5qet/2RlwJJB6iJcykX88Fl2yuFgR4Ta
7gjMle7qzuFanBNSIxwIjBSBLbKk+anSHhsBQ2jdIxZGuk5UfLGR/fiYCRX9Fksd
U0PLsmw1VXktEFEYUXW9Go3v88p8m0eAlHtDR80FLNsFJyYxM42YlzOWKoMCgSHi
CSvc1EpOeSuudWsyU9dxz3XmbjkThiiEg2G2fRfdyZIdQP0LFkfGDpi1XuCMpUE/
w/Om/ZV/spimrzcAU76lJ6izydwRr14r7y31Pux00zWZApDAryRbVaUkfNniTFrB
GrghKjSH/Pwpv21mkqATsRiLL0JoosLkjhobB2Zf9NhpwV+2mHRyqtiJciDaVck9
brUngFsAGdGyUFHbKyDd/rZS7859O7vLBpdE3pmdE9OjZZyadWC4imNurW+wWpUA
uSiom3DB42vnwOfkZtxBku+r+ouHId8kcum6qnsdKtzYD1lYDMQ4oHq8pc7hXxUW
tIDbDbcAJr2kZxPORgTcRV7GqNDRvwXx3asd/jmpxn1Tnl6Z/d4eWFxjaqe5OKHE
s6QZTOtkil1hZOT6bPofa9TA07bBoDn7roQRCFEMKTxzG3mhU9Pos7elJti0gUEN
AE5Kxrjy1JSzT0xHg7Hy6jgNxAcaAHsN8FVPYLO9RXSbDw1oFqY63lGq+diwIbl4
HVZKEPeHBw+Nn3oJcQVVN/sSoFJTUnOo6DNJnpJ+bMbGg4LeEGUPonkGbq8IlWBt
MnkDzn0ngKsiVJKXrmgUzYleCDHBu9hPldT/pTsDe2q2WwLj79VhC7pDg1IZXa93
zW3BRk19X07K6OQ1sBL8w2ihnODB36C3TH9Zq8nKaMos0AqkOVTnTkiposOUPYcR
/Ex3hqcIIQxL5rYlUv811e+ioGbJdo+gbha9dVn+qrmOVg6Fs1cMk+a2fSwIIj+R
rI2knpQPHdnbtkEpisLa1d2L9sufvc4l05aqkVH9wIfbknX7HIt6GmccKP0Qcg0m
//Epxb5y59289bZwuq8Zdp9SQ8Lgx1zi3Yoqs+ryD9VRAd8aGVVtdxLK4iRSe87K
eUHiSeIjtg+KvgM8FmXllok41HVWmSEljSPfKGQBuLchrsq4PuTNxVfekipqE3K/
kkU1WFkaWMvStgWrru/q+1EPaW57J4OHR42UIl62OyOvEjnN/da1eEIGmsvz+3h7
Qay5qle5MEwWz8GAS+H9i+ynUD2KqGbke1qQwood8dbEy2Ri5jKDifvnsKmdZ1f/
3IzvMwG4kz07z+sHoQ3gNI/l5LDpxid3PUO+fnDZJIT78SOy5fBXjnAriBWY3F5c
cVEa5cIZH5BSfBf3jwyPnryMwpdDlVdn+YijIHZuM/JbNzDW4JvaUSlSPbjv5Bks
KI9N0ogURMOUG7jCG35+OcaubxVSpWww5Huq4DdeuFt0Gz/Mytn1tuM7gbXqabfN
1LLOSbif1bo8qkb1XTGwRW09WNzOgs5FAT0zqOK+cHS01XnJdTHxF6qnvYeUNcVY
NP7fb4wgKbWbooFK4c3LP6xX8VSzFZPmTi+i5KJuW5Xm91nSLsAzHwSi9BGYVDiY
0PmwCj1LeCs9CunMOsoiyaRjFWx82GUFOVDX0PCndobC0/azw6QWbLR4NtVTseLD
42Ei/ux3FwwFTeuQft9U1HqBXJA75iw/WA/Lk1uFqHqXKSqnozyDQIFs3X9+hLMY
213dJt7JOkxX4N4+8dtNUWmiHM+fBgZMDT9keRiz1ikekA1cQmxvR9WD4czwBB1L
LQTk3TQOOox1CLD+rsFNF/PVWIpQrOFAGOOSoRQUpFG/1vtKJA/EYaUziKGKXufe
43McGAvr8vDqS3cOgQunaqmc5o9ng5Luw3H4Lw+GXIUcle+918JOqghxWIJLwdkO
SvX/2PVaZW6i0t7Lwg7x8+LiwMd4qAJsjIKTGu9jIskYBM+1mrWD32E6VPvsTG/t
Svv+UO0SLcF062ySAeQVXpzL8QnFUGU/5yLW/OEh6Jp2V0J0m5vyLcdUU/JkGtIb
78lVlJT50lyEzBhpjhwzqhxDK+AjagA/ahnggFSPdb4zEIag03T2fCQBDhJm4jOX
ve9Sf7wqvxBDDpYPPpkKohBBBv2EeQEfUjiQ7tmY7sXPKkVjmRx+q6NW22eGzJaP
j4Amlmnw596Zq55npd56lVTP+WyYxFrayssB81xP7/LVVjGMrK4CPuSIh5Ek85XA
kTwji8kloPQ746d4mA4pdkkVBZ8wsdOwsYCn4nZsZ9UrzZFWF3jaCQ9k4d0pbC4p
n5DPWnI3nINvpQK/Rc8Z2TC3s38c+jgIzhDp07F9C+MEpj0VdpIzHW0+PIBqbAfF
/FBNs9Ka5KvXC6dcQ/poXA1gip2x5xHCnKZrVXCLUmsLsJzLWPE1WLF4FFD1QkCz
TziP3DY+UoTqU09rsJoXpx+vM5rSu+wFa5ZkESHlj1rVsp2odkThu5Ldn0imDwMv
o7v+cFKzvdg6nsAdUNPTTyZZaqyx42VBSScx4B5zO+QYrSUlTmFHiOMV/vrkKSX3
FEVQeIGQn86hDKDS7uSDLw6bL/nJriTSQxe6mnFPbpWdcnbO+17VkBj0NMB+lUJS
w63haKDs7Ytj/vQ84kfvte4Ki6Dy0gsqDrv4nu9gH5svmTjzL3KbhOxveU3ls4ep
X2JE8L1UyW5eeF3rjZRni1OVoGiAbaZ+tB5deb4C7sfQNlEnh4FGzlgF2afoTLMf
vNhZHlmuxNnf6XFPPd4cOIVPA1UhL3XJeqoY+7ssW6y6DzxhVSZQCq6tgViPVbz3
aqZLFrMKSdn0k41AJBv7Ok0f+lRZGK8J1fHTSb4gNgGpJ09bMMw11QznDx7IGBqa
ZcFSXCa6ZO1rL6gK9N1M/h69YPYKDW2XHaPRfWyztUMwC0BehVZdUUv+gYhNfA8H
1mjRp+G1JzCHKobidgE6DxN52Cx43l6OaOXyBRod1v3/V3BFelNDANskv1hJGSHW
KNvs1YJgva69id/TyAyFzSet/zQRHiWtoz3FizCaSKk30uQl8os0Ic0Xo8Y44dcv
mc4FDE7/qP6artGLjdrI5TBUPz8iY0L1JSn2C4xYFvWsN6iu8qg8BM5PY+RM2fYp
mkVP/1bk5fvmw+Kj+ok8c5fDGAIXGMUp15uPBHWFuQG0KsnmwR9CJuNpdS/R+Tqo
1JUxIIEIu94QP4Wq4fFJX3FraJ4jpLyr9myGjnGuzs2xK+kabjI6hUUivH31fYy6
MsAa3ldJbflNtJzKmQkduyOwoXCrlcAzUz/q/U80pXu9+PpJGfuSwZBWfGacDlwe
FmPO/XHwDSGFeI1GHC9y8kYoPhOJkrDe/7MGHsMEHz2/J5KyJBfd8QPKhk8CZXih
vqMtCiXBbrIAkdD6+Nke2hLkl/GhgLvvxucGHci0XYDlP1AIC3VyShCFsQmk8kt/
aeKcba5RyzBMwQwgpxM/Wq0Awv2iq/IrUVPBx5/BXoTX4DFC7uwO2AwTLoxWCDvL
BVDlMCFpre294n4kvDfab+dtTvl5MEn3e0BEIJJSdXbwYH+INQvKSIo4xROWk1J0
BGZ27T3D2MM2GutJqJJz7F1lGLK9439iJs8iaPXjXxdpi2qfD/prAXiUU/vZgjF3
eHTGuzQMIRAbEwD4ZUPyRIsydfFwnh/fkWD94a8ZCFYZ5sT/y/ianOiP/KFnX8CM
`pragma protect end_protected
