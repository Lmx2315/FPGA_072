-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
IarF4JKkWtpfOP4DcTpeUXNss55/XCdago8bZXT7N3dkjoGPhiYBATTxFIMV4kdwBwmZ1L5Nvpo8
8wOHoPtnlCLFCPsIRNy85bBhkL9FGTV6pOTY1FYTlLzleDwX71kq0Q8+n7TjBw6sUu6RBBJQtTCW
Kvffp5JmuaDTFiUzR2S6lIasJ7UBdHBKgzK0dvvxhe2mXc2JkNHRuMFyyWdh5Z7ktq2rjlFzszqk
BTquhKgm7YtrtNLiur+Nq+7zAXlEfC8KwJO8f8WxOe+oLBQwKP+9CT6QjfWCkYYTAK0m9KDBhI02
uO4nG44u7WV+WimULUrbqc+GB7u+EpdY3L/Kfg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 8048)
`protect data_block
ykMB+XPWA8xoiAvDHupvtw3oSKT7nvQK9YMjfAkKmx0EOyH/sj7OXh6I7t5CnHCuP17gYeRuqEsg
mPugj+1kCtZoViT0dkNG8Y4wAj6ogu0DRozaOBfQtcuaWTrZiOK1zfcBK0eKRGb0VwdINxGMbR5W
9E7gCsPpnQ6WkNUMnvI9yicf9opldkbl1Z1V31sKy8r/llBI3ws1UZQQ4l6ghcyDtTSgm6JuiP/t
yqXc7GCAAh5eztDjPBf69O0pdAhHAkZQ8UWkjcyjEAHoxTFKULMEQltGsqDgO553Ve4S92zzoXDz
8Bspn65yjxtpv1g3Hh93YAd3D5TjPvxQs1RpKtx2MhG4RP74dfcylKM3FpZuLNKZe+dT/C5B4aF5
OzpVxOSXJsN9eSW9JmV/cW7KTpfNt45G7T3U4cr+RB+aOutAKf5AxmxyCf4f3SSnyx4yCd4xpEhP
1G04/c+BXj5PTuIX0aQ2dfD5SFWjLk4/QN3FkZrMeipR8B5Wb9kzAi9xzduVn4nNy7jnkV4yfaYv
8L+RsCJqlssy9ava9XYLqd1tF0imcZ3v9PJlPkR6H0OcerwWXNyNvaEq3dFtp43VxRkQv2Ew5CYP
QlOLVwbdj/Co3t/Ozfd1DJ5C1z9BHGjhPVxGng+zUl/k/ryEH2+pVfNFRMVJuq1pN1mhb8O5RmQ6
TFTz7ICafDLVGA8HuI/6ZB+FMgG3Rr8Qjqs3TAoaaKYEgkq1Qh7tahk0pCX5r5PbS2EaRSHNCR8j
EUMukwOz+MxXuAWa3RujgX4V8LDS4bLN06RKAjZE1dW4JomVhx2j+BO86wO+JNDO1QeNKyzB+tOb
zCrE8RNYca99v1ep9iPJhy2aSvdRFr/v/5FtNuwyoqBQT51qcntCQsEf3EIdNisIjgG3jTPlnoa2
uEOI/1zTL3AQc29exh69ZApvGIG5h+yQDQ1EcErNnZR0YtNiL0qieEvncGZWfc30yA6Sma/s/MmB
03noOK5LoSvpeTB8J6dFLwvVuKTcXSt+IpCC79umLzBKn8xUU0FSEVskCzrZ1kLduWr9WDDMoLLG
2Jvn6gwo1eZ15GyCS6gR/pchD+3rbblGfNh5vR5ndl0O1XSjQgHYKzV7BH7ehzd583cFJ42+T5hz
+BI33Ve2l/V2QmM8dDE/hEUhQGsZC5i/lTTDUayk4TeWAWfTLuEGEDANb+04vQ6W3F33VVVmpDYT
Vi7pXUNPVgTgsmsMQb46QYGlr5j8GPedOQLiIQ9Kpe6WoEpYbreX4XRCJB7Wb8FXtsiA4TUM4XqK
O797aCWDC30BfnKFKE4NGdNqUj02jxFsVxkR+7mYARpghYEBLOBfVJbavcYkdIImwMuS8vl2LBoL
aTMjgbOZscvigDaQ8tjZl496xuEAiBSqLARKl7xzxV/UX4vtWbGzwyz+wNig5g9Z+T4eDucj3QuN
HkMTUJX0o45G/pUmZ2W5ThTYkOmoclVBrUYOQDcU0DAa4ZUulmuPqztWa1AxEfhEttxKWyuuM3bd
korPIb2cX4UB48Kif/72UWUBMCzflkgGqwAMb1bsoqObwo4rAdGjPlZSL1SdiUsrkUi8wJvHdkMx
5tQrebnOK1sDP/KQL8e7XzZw3lXOWq/91gpvsyziv7g5MQiA8qanrbtn8APymLU1Wr+n9s7M/M5F
KAUjuVhKO5JWgOWFabjyjdBbKf1Xbi78z2uG31AQuROF/ywrMy90htZQrKGepFxjlL10RLJqK7i2
kJsk+XtIYMCRbtD5aw+/GcbZqiJVhc8RlTbqg5EtyCkuclSYq9DHeA1s8/UMb3vurigGjJJMKMEe
zVjDDBsGS4FofFie/aKk0ELm2CWgq/jbpJpqKBpoZOEB/rxT3/xUHpwb8D+F/w2cojTU7/2IGxn3
eeub5QtVf3PACLWb1/uetbLdUWjjCRu60UozCDD4/+YSLM6KtURcDd9BsLiCGJk1+5Nh+NL2NJSB
uDeO1O5DfGSEgpB1NgLelBdoFc9PqqoyB/oea4TJZwDr1SpDvBfwQC8nOr5Uz6Om3Qpcw0rmAWYH
z+LqkcA8JO386G/dqtFdT1pjr/ygU9x2H6Jmk/qWz6tWVr8a1sycF0kn7MFllMW0Z7lpP7DrRdIB
AoVGuBvBx/dvmSheSh1nSB9X9hPsnOQ7Wz3M/S22bxBtcSoT42zGEqZGrEurtGws7HukUF2ilFyf
F7M4D1v2muUsIclhg3EifKqziqPYo2ORmjzaZI9d9ggjfvmmBWwJTLC2I46prsVr6IlHF2o1LTrW
Y2eR8gfcBxKy6kflrHKocrCHawfov/k3IRUEAEb+o2H57OBtXWZe3vv5axoRdvpiTNTqDzqRGtru
YY+Wqo1skiLui+EWmQO2TQXeWNQigwh7nLO3fWH/Kk/LO0YgGLVkQik8/qE4C/aWD/jGDinluHlm
ayHUuuCXucAxR9l0I6Z26f2Ey7VFGR3vSYgSjiTUYw9oB0Ju2ILZRdA8Q8SrnJY24fpBm5ChKuct
l5UNJHpoLA7LX5AsJg092p5gNNyv5ydEFmeLXkKHwic5FqYJQfUl3wgbdj7Dhv5eoDQlLiHVN3Y+
/RF6PJ6qndHcEarcW2mR4p+tFX6FII7pMhAj9y7wRbyRnsEYxOnK1cq0gj1eaNWyj6AWd6QRcVMW
/yzz/H+rjVd4PiFqlWfI8MPh5IY/2yXC0Zzv7UUWAl9dn1hAC2NJKPB9mjDd39j/ujHIlVw+nXyh
XD+6Tiyov/NQWEkXOqIOiBX1TBf3zQ+akrhw+pm/S9L9ZBkel0CstBX6Z/a6dJLMp2IubixjS7pI
rbpchL9qDkZp3sHcGWVlunligdKPxw+Ak2NnJtxihroH5FvmcIv4SsV6xs7e0wKI78Ae2Ceyw/m6
4ZD46O2tVLrbjv8q3gMmhnOr7ne444vR6bnBDjt8W7nSBuU2odxHegKTnGsEyau5Tkq9sn3v0MF8
TQSKuQhwvwamCkvxPsR+5jvHP3GK7UriATBO0W6dcM/Mc++/nrXpjMYoSW2BeCn5bviKJBhGX9F/
UHLd5rCPt0XxLOsglAHLFIR+QbV55XgZ5ZivcUGvVwGC46H7Yst3rNbGztwu6VSBV7+ZbmUGXJZs
xiFI/sF5NxgiqoJSLb17HoJCl3EVnpPRIyR1PFwBKiiVHV8KWa/KeBBotlieS1dlzcvv3GRnGuyj
RwGTH480pFp+Mf+O4o5eG68IHePQ0EN6H25S9Nw0KGUWSC/AAVoQ31hJQ9cHBXkvOng2GqbA8B05
07iVEBI4SskcRrVJ7P2Mvy3CL4/QTJdJ5hSSmok/fxGMwbsFd5iigmvN6OyP1eyCoxOOuD1t1Yhc
oJQUIDfz5VFc68qGPBdO2DTVofHIHSZit3AQhJI76ZAIFNu14JItv31sQQ1g98NzUjKLWx5MaZ8n
dEASc80DAtz6toiTYPOFnf36mRDvFCHaBedMH5Wl+gVkV5kXDURxkUY6LY6pxJrpfsWqZbLKg0gl
M2AGFcC9jSU3oj8b/vymktAOhOl5SOjxi3pRZ4EVfw2OQtEzdFMEr/FJIo+iKQb5y9Ld99I07jWC
dOv6FHVx6yQwlz4O2oy80Mf09QMpBNpEWSE3GfD62Sh1oJ7AXCWcNKRmiojgSGsWilSDdo1dWX9X
YXzxcaBn3znUQuoWYhuDX7zzQ5oYcRtEt8OmRDAabM8GWaCDJotqPncaqHJIiQQiKNmf8jJYCC2w
Pb6c/x38/61JQ0EqfQLM2CtlFojGAYUi9ZSsWs3rGcBOLK9TcJX5WXS+TCW23/5vlR7I6OEGyb4N
FwmO/27/AmSfvo+7tAxFt/zQFH0GB7w8zF1Nn2TlNVqXZwotdE8D5vDij0uQMXX/KRAM3vy5Fari
R/eBJ79e6GK6BIHngfiwmVpBzGJw4yPboVd8uoA+evqzjX1bl2rM6UWwr45wDp5CICJQMOCgeoRm
IoBJ+42t2bVeeBf2xjjwpN+WG+bqBC8LXHx+mUhymXzKaRQc/nZNBNfDyXzqpcQMAh8/3fl1A3wQ
wX+jIXVlLQKNG7MulrJEYnzwtrWWNOzxvoxxXstKDmny9iHis4Xqv7/utNOZNKVFrFfInhNlCzOR
3j48LChSADUFDh5VFnyWREPwa1r1nzSrdNtn2yz3Q85o84d5pxCoSokETMV6yeIQa/ddgBJzHcp8
dfJFeFN4GvHnQbarPhPQGmJEPJroHWClRT0L6lsoF1t8EYmuKnzUmJ7FoFNf9gdgp5bJ0ZZJIfEh
aye0UqO+zvtbZVbDwunTVRwxzfYoCuqd+RA08WJc8P8Wp/TTXdX75G/jnVgA9ArIf0/Jr5hYqn4o
mm9c/Ivl1b1ScSMNpTbXEPKfJIS/JuIKTr1nJKoqLiRqellgEIt9wQ7KbQ7ZLKczeQz/kh5A1Hxs
6C2nTnAlEEb2WvWynp98mZx/bW0VQzfDflqPbQmyA0u3Ev7Co+z5BBXBFXQGOFNWe+tu/CMHcKOJ
U8UUW4pj9bSfmMUe+ZaEcpd3R7Vd5NZgAEDk+TzVqqiSDbT5Loo57w9K7zC5Yu1xpqT2TvSEtAPT
tgthF7indh7x6UvXrrT9Seh0nBBjWn4UQIzEd+OZtdCr8QaPVC41zv03C7/4OCUyCMDraxZ9UpVN
ycXdHN9VdOikcygtG6iZhrqhMx6zcsJEoUw8mYXQTKIOX94al7sAimbJHLTPnVnt2/MJ3H0qDHm5
syz/ef7y2rsFhOcBGLuTVIVagBnJEVhSgqyFf+09vMocNX56X6FHGcpEuI87QLmoN+XRkQXYB37h
J2FywSsmFcn/DY9DxZ06hb/4FF5SnDRSOkBcXLheTXOmxnM15lG4KCLU2RP+0ZgHqxuZM6Z93FxN
WegEy3tey7PQ3RQf+jLGYRBiflUr15fEn++45o5lpT/RIXJ4n9YQ3UKn+YeojKtrYBOk/mrTaZYi
jUhSEV0287XEiOt4yXRMtoDFoLwEHR70ffx4Fmg+lLYul7DgXE9w/hgZII4A4z8MEipPjuHlxYxT
/7Ga6A4AiZJ2P4U+Keaa1h55FMMdFqLpn1JZx6gMcsqbbtwv7fyZLK+PEMT0BilgwgoV428ahXWY
29PAgiPfky750HfFVVzaquSVXIxQb2SA5yWXOR//z7VqW3gcSDPBDPtKZO6W1EgANUvQE6QBG9ki
bDO6DBuQGnmqWoIY7NJynkRpW7UQCa3zQJA0kBZd6PwQvBI9Faxy7K8oy2RXF22Fgw1LBJ68yMMx
cimxYBdRI9FbIPBoi/c2MxiJqkaJ1YjM7hsii83jMgjDdYjHKt6+OeUzh+qaX5aCqornyGuicBYv
ezDdpikfJ47sLtG8B3BQB5lVYcwCS+uaKCaBfLJfhmnNF1dNE3ZyNkCmRz5bcA3Mi3HP5mBRbXEn
Um+vVFOuN3DyjV7F085lvEIj4I+zhtnRcPffpEg76Uxfg8w23HmacvsqFqPh1dcwiDJl838o1GQr
4cP/XZT9K9Bd66bfto34954qhg4NejlOSC74sLMbhxc+3dGHPOSo9vETjSVMkPbjWjpfGOLXkYbK
jYVAh1Exx43uZq+n5T63y+HI+XfrbajH2FNZhPm3UX01v0IMn1UqQLQCx13ZsT8Ffp1Q1pZBuizL
jc9ELBCxsYexOr1f15WpqyfikEX6nVQFPYTZqOMDlzM23GbOc7fg7XnPDeBSRjsO23ok+urIV4Ix
qXAP4xaWUivszpK3mRUI/pIW+3rUGHnahhalPp+48cTEl5Z32pFDIjtayJIevmu8uVFwU2fVS2t3
8Kc6hoTJlf8f7VGKlWPTZDO5fSFXhICeh5RkZ/ZHZxZn9ffzyZkWg5YOLnKkH1gDDB19wypbng58
r+Y+td6F2k93pUc2/qka5UaC1Z6lM5cUNbv9OE2x5cCSMC526ey0846IdvQHXAtxsdrpqRQHsKGJ
dtBi71AuL6bhEx8qah4OFD3+bRtr7v9LgAI1QSoSwFcTlGJuVC2zfsWXZgWsiWqIxAfIcmHqBlx/
MNXYeJ/+Gkxlxr0eET7F/jXYQklv9gmvFYeDSI1C8oy4KyEp6oxBjjWkCwjX+EKtgBMOS1DFj7Ux
INB7cKedvPgbkwmIg1ZLSoPf1ylFH1yzHRtOuQl787I72rV7a4+D0g+ZoRX1Tc5SoB5SEDb4yDrG
ouih6C3hn0Dtad+Dm7wavh5N7NaWY4JxFa3SQRGLPpQLRLvGkzepg43ImIJyNldji9hpxqxUMY6o
uLM2sM1Wh9eiyrVOOy3GXtmRI5J2kPYVtQoSQDEQffnASeuM8Vv1YdlPjyATevFL4Bu8mbMCFC16
d3TRjcaP2jzSlEJ3SGruNfmJEHM3bYybihtF5B/m4IjznYRA6/X9QfE7xI+Zpg4FvAJAVTzwZSv3
/x7h++Gx8RKb1s1o3IcEJXEhQr8qz5r12cZeGdDC+/nPzSKqq8y/PQZ3p/+46LU6Mdnx/aJ0vgu6
AVoaNyNsqBsjxioSIfnt9W+XlP+CSGcazt6m4JA6nfNNkyQt/C9K7mB1S03R3nmsr57btqmHAmQ9
9anYQVLUzawY91NTZ6fwFaLSOXdi99qkUtBDIzIo4qYN1hNecpQgKF/zCQsmoKYjnJpi3ZVOwxqo
cIoG0+OLZvmFOUtUmz3J09wB3WhuMIm4Xf6lEREjbiC6Yth5KghP4GDCBPR4lQX3p9p3eLbBRgMv
9kkt0ZXKp0kfOon3f3SkYzx1bLpjeeb+QJPvU7rmAtOW8rdFByaw8vvTqLFrXpoDQSOB5giAQSu+
ZbZtck90Ik4mgg4fFen1FyUsjRCsMgXZC4q+/pOVfSGAueQgV3b9H3DzrwueCXl2sGXMpYyfmf88
Jy3wOMYVrl/KkKVcb1rVpQjEW7vJ23USeVgQF/ZLXK3/gZUqZzqd7iWpoDVgwRp5ciPa6zZlxF65
sqmuY/506Q6VKk6xf9v1Gpa0H5d8TGl3MhU33NnjtRqr9qHNZ4YyPkwLYGOkPJGk/m2YAkDe5nC1
FTynUZ0ed9oJ3J+yj+M0xHsFL3TLjyiLT9Jbz9f1G4Xec9djOEISkF9qt7JaZKBRtXkjU5Jza9kZ
ucG0qvyyVWuUBbmVs19JZEslYv9zwn0HxP5kw/1SASsrBIERey95f84dWtNjETXZZXmosFaESVPJ
zi0E5SuvKmax/uu1s1puYZsCWi1DYyJ9aOOHkPVfzZ6SNZpwISvZxCiEIhmL4FYzBYecIhrYxQ+a
fLexfhDGpwyR4fQEMrBe85V1SxlQ6YIQOekFiyKj/bZ1oL1h+XFJ5qPd/jGPUiUN59g5VT3tOLpa
nzd3V8brRLOXQz/pWku0nTXV3/qF0FVw5DFT+p1ZSE09sIJSmcYxxDXoegWBGj7tVWxye1ohUhWW
SVzZ/vJi+CCcyPCx/oqVb8CANpTy6zCPG2NVqjixQ0KugLxQGnWEdZ4PO1nO22DJFS/24NTIGkPQ
7/wXgB9ABe1HHTBMF3fm/UAEvE3MBUt7hWqtE25f+tetPeIRDjH8buE3gVU40tptlu8R3NzdjOtY
d1h7RcRhk2hENPS0VlS0UlPypvGQ31g32Damp7eNuTZX6zttWhtPKkKs+T9WJBd47rtq4cwvhxJA
fOEJxx9/Pv/PSRCX8alP1stfMbLSSh/sKpLXq2Q//XxpYa4gsbZy1B+wYFfTsxjrUOQ8NY0/8g7N
3JpUNlwDJIQN/fqYiQQ16zoUfQWJ5sidA7YkVmioxoSHa6YbOulhm4Vn2IGgBJpZ83zTJtBxc/8Y
NZpLL64VILCQZrzTdCcsETrKN2hG9qXLNJYZv1u9xB54S1ZLN5P5gC5gstlXFePKpAzWZIbv8bnH
XklRgv3cwtZvv9csIXzGsUov+MHXtHTTlXxtmlXGWRJBxCovwhHDKDYut2b3zUjG8eSNhvLZTqm+
uLFqB0TYox+QPUJWmkpjf0ABJKq5dIyp4RsTRUh8IqGpfgk3WqCCOF0bpwMZvR20ZsnaIPat2VSc
chml02yMMFjBAbK4jUcFMfJ9VbmsKNInVL61ln4X/n5bTDVlQc7+ZfarHECdJhp9AYOh8uwSq6kP
9lkYg29sHMdbVr+GR3Vvv2JdO/UjrvzNrT9CgESzHUkeZ0UuxvpQeZajKtAMB+gV2fksXd1Pl9Gj
5R6KNyFfBREpEMwbvDup2MPcA55kRI0iViEAzQx/IjJ5/ff6zLqhuk56ILbsrNIwwmiJZws89oon
Bgfv0WQvI09i6ICrnJ4RFFOp1EO1RbEqG2/DHbdxDjBhx4to0NcdvJLDrwyf8FToKv3S5BvIsNuW
Pzq3TkcEv0KghrA2/IMeMUC5PUF0GF4G5EIQSp0XjF/U8XtGEH5H5OZaZbQJB8Gzq6AW4YqlsRvq
qQZNaAoo1BpjT/o5+c+FQZeZdLv35lct4DJ9uFvKCZ+77kYqdodW+7mF/o6mW7M8a+1C4HeuQMIM
bOfN3JcF896RVXExaq9iSj7OdtfTCg7GS083T1tNc3hCI57warVpeYK8nKZNpaMGX3mrDzltrRKG
0CAkmCTfPr0BP4M/PboYNbk0FHxJ5M/fdSNDfzh/IiRTyLEpB95xxpjb5iVmyzCjWfZEKzXp+s1+
9Qn4IurGgwGSu4P2JLGJqMW0Ck4dOg31MGcdOtSJdZckVYeAHsebU5YVlyDvZlarF0c6ULyV/Zty
QmWuCohrREfuDvdmKJm73hY1lAwQt4NQcLMPtbx4i4rDURrVOPEH7prqhuO3qNe44CIKeQfk+M5c
1MFUaPerwLsCZNYFVFGL+blGpy+LORa5dHrzBksTm0Kqle058yi+CEMNE+t5kXUCL+xDopCmAilg
MOAozxc6Aa5Qt6iwl5RXd78nBOvZ8PPHzUJ3L5wcfF6nn9B60KCTAJBTEMcITzAeaNKahw7Qo3r/
uExKrZ1NjB5MGKZk383z7ZlMpAsmB/l7B1J+VUsTis2esluCi2hYFtlp8RGxgQqA384NNGRV8Az/
qbJdM1+lPAxyRbtDE5M8CWzF8txjbFXrumcCINji6nLKvTMkzRSiVxjvQjo+8xSNUdb/t72Ua2v0
mQOi+86cmffGhxToYq1zwoD3H2bpLOFHT7JGjjIKjclnM2yLVHRqya6KDEbjD0y1eXTG8a5cs7JA
hKd5UYkBVX0Uvd9IL7edZUSapk9csUV4yjZYqRU/TNZIsAYxyuH6dSVsiC0hr6lTyRfyl54WMzIC
xvZl04FrJeET0ocpzNvHDGwKGrlg3uHOQ85EBwM3GyAHjQRQhZ/ZTHY0McFJFzKlkpVjVVkAgFXG
K2a3/eSxhfTsvq6QGk+vjsPDHcHwWn3aZDs6lmd+SYz1QuLLUyhgFCBTqYwiuCnpgOo6jKWO9hSf
y6i2e/ZHTVVHcmjSfxCUZ8ADTKdRnE9BappwSVjeP+RyJ3L6CTIyit1TYrJBQnMXbkFVrOPOs02l
9Fzu43kLLSbB7OsYFKTUsZEg7AYmlWaNWx1yo4GxP0U+cjEueKe0lg1/K7kw4AH4184Z5i+PpEQd
mDh1dW51WVoyobYg0vnsVbOk784YEtNy+JKk7zTumwmgMXJ6yH7n54GhH9WKWQ3vkIxShzKgXxYm
pz3L1epujamcHXo+H6fqvGL7gtHUsA3RAhn/vQxDdKRMBqx/wtA4hZBlMYKL8Bq3BGmxptvOfLb9
diEFwMtcwIe+zddaGwrfwhzfgfGWpQEx/jsY3ezSeQZ6UGPvg1HTedZcxtDn72JhEb9NR/gVX30K
k0VvgNVOAmdD1ShBrlGHzmuRu2ZjOstYqK91DeczaEu6z4pC5x1+TBu+3e4fFodFfsvqu4DJrk1g
/wo5TfteDDyjmIJHkHQ6RMtr5nph3oSdr+mpgVyrUTn/K5bAAUhY0IUJVz/QcJ0Lui06lVtrNSIP
WcDDp/34TnkP+ZMOPJN4EJkHfFtPfV6xZ7lJ0pTOPodf+9p2TcSW5oJSZ/dexfS0PKBzfC1mmkhz
o0tGBl6MGG75KOVNbWvMUZsDA99xid53wD0THIc/ZlIrnPewpqbrnm6RP9AlTWwcnAeogwrykxkx
P/WypGaoGIN+/3NQlHj3udH/2NWNVFFsR9RTwbBQbGpRZ8RnvVxba7+eAlw5X9t4qd1/e7Ph2UlT
TdLDkaez4P5p0jW64wumE2DRMbgKWV6dtXALPfAmCwm0noXiSir8Y2+ONJyETx9Tzy+6LrxhRHdm
dkwNBRB16L6hZPMcpmirD9MviSaAkbF1d0I1RjjN3jlxcQBXjZUH1UZZTVa8Ark0ddoTgGmo4dxB
4yf5BBcg1xESux5vourQNXGBl+/h6WWsyK6cR1TEiOMx+GfFaNT8n9KE9gACxW8zk1Y7w2De1Wh4
Td9BeeWyczqyi5YOcKW0ADLkv4re/iEXxhTxozO4+9q1ZJYk1UiggQwR9u83Q42RLn/el7EiB3pq
fR17oY4r1CWVFW5LXxUSbCkhfsU+0nSkGdNSWEN/JGYlzjZLudHmc7gep51Qr+PH5gSnEEzxAxOo
sCzY780CysbfJ3vNxCscQ2ELoBe48G/JM3prCy0Em4XlmTAznzjF+XVcsuiml2b8EVAqQMMW7dPZ
+ZOCL5CN7OLBgeducm7f9Lnwv8c+k7n9MuVvUuNVSXpaIIZ7rk+/7cHAds8o2mAnUBT6cUzZG3Us
j5CG2mMCxc+cl/kncteJKWnzK4i+vqDkrJkSc/XXDsbBD0WJlF5mshY9h1SVLW5rXUjNAOGhoGVl
6eF2jGxvy72Gk4s=
`protect end_protected
