// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:32:45 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
cy5egp1awDuZFWM9AgsViSu/bFJjNLemKAkFYwQf6AoNA+2zvOF6Q9BnLr4+ej++
yC48HWHhWXUPU1NCroPugyOsk2OpoV8iHnciX6KwLoX5eEYNqZS5PWBUE59LzDdC
wt1b72ZdpmeimJe1fFOpiXZcS0nqLZaPDsnw66FSk6E=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2272)
0NdG/j1eLUENSkblBRMjdXK3/N6+XQnOToKDLF8jDmjLY36a3F5R5j+7B2tbtR15
olf5IqRoaP4iP2ORnMVHLvADkc+DQ6BDwUUmr04WWXBA8NRyIu1MRZaxW1a9t0xz
ic0eZaRgPAa0YpoAakw0OvnBMeSBihXcRUY7+B0We6vId+X4BOXylZY8w9RTvXI1
zYgTsUlI9UQb6EWZwatxq+LgD2ZHjLGwl+3D9vSQbXYxCCW+vs9hywRpFbfQm7sd
MwvAerPObFCkwK3xbjUiTYKetLNmuJwP5mLZfMRHi7b+pYRxXfKqlnNk7wXf7AjT
xLwpPnGwf2JAYaVUqfsqFUxpgvPkBnxA2YPOVOgn52+MqT8TPf53CDsZuAC/QGrw
pjb0Cin0PbiLx6yDN9uh+/JTbfNakcefrIHGKn5TJKu7TrWkX1bci/PKJlu1hgfd
ZZhcocVyr6HS8enjFNE9vjLjqivkPY6fWS0oq7WdKyzhO4cK40Lx5gQPnhbhFi8F
BTUW/i/9pdvus5bEQ2ZBDMEIbsHKEXxi2XrLgxLq6Cq6dmRFTWEbYIIcGbRb7ySr
B5IDuE24JLpebIl20ZTFjzNab7Xx4Wnl0Hf2o8XCBjFDjccZ2vClowATobs0zoRw
Q3RbBWJjD7u+SIY5iFLT4kJ+PGg/bcNBN7QCxyNJOwDDEXvT0jGTjwxyAY2o7G4U
ST4LUXpDM2pklD2vd/1KgcgevgM5m65jxcmGAoNQFYhuA4jmt0xz6Fe3oWC+RWjI
emalgrIKrI1dH6GPSJt6BBKxNvI+pPO7K1B0f/J9B1VZrfjD/Fq/BxlLjM7npQMG
VON2uskdFibcbuK3d3enbFHZb7+bjWR/IxEWglAXlpZWRbYyHjbbRu0CcliN6UrH
lzfDLueRF5oM6wn6Ro9IFgNbzIlqwLDGk61azG6AVns7WAdoDE19/NSJZu4FK5u9
raC9+gGb7w4hqEI3ULIrciHq3wu3+Jdb5WuLni3Qv+BIxbdTgqXXWYJ7Vu/Z12kA
R3+jeD09zHznE5KLSV3EjIc8SxeBO6rUttfYtL614dSbpHP98FLPMDevF7wrMHRi
HHEzDZtQwcPaBTjgxPEnoGgRn61Gztc4wHoAf8MSQAeGVj4pcR5BIzazSZ0Aqvnc
KuccRQ8CUS9MV/6hqqXEfrahTPJiDVLuhNW8iimjOQazJFChSavm958beqjX3Oak
zQdLsbAgTqYnVFZtvl28zeuUNtI68ubqGtF6aLRoNlhVjPCMYTM0uhQubwaHK/am
aAKoHlB0GmYYxVdE8eB2zMk4yL/NAwBmKIhSDwMIPRmhmG1vU5yk/vkpOrBx5gKl
T54l72wEjvK9ai/IrDbgwXEtaE0kUz3dWoudD24rrxq/2PTBc7AOudlhjYf0I8BW
x49SVOhMqfW34YALH2g7NGwOGh61l4n7QJY5VQOobrfCUj3bNeBB3vqHf6mbfcOV
J9j2unQER8l8JiFe2y0slzEmS/1rl3ms8671j3h+MMLekNSAJbb+wCbp6/YbpMTI
dz1SqtuskRvz4jobf15vNeLqd/fxeULem9LjxFNvOulnrN6XDb5HplYjqumWCnoy
7UkJfDwAgpczTA0rkaZH0OkNa6kI4y5DOA+IYi1CZ462zXPVD2Ua+A6dFMC288Dx
iUn4XZX6wcTbb3LfsxfvpuddP3f7OoyebVeB5V2E+3TfpeVcMGC0JFbX2K9FqvfB
r2+7+2pBLjFQQqjylmZBhyKMiJ38vcbqmUtwXD7xJ3ivrfI0NkyRkzZ3wVFPjrNb
ggM/74J7Wc+OCVibVEbJiHQyPOathn0+9x9TzYX+qNLvx6py/7MrV1lWMpI1dT/R
NdfoNgyls4ktxYCvv4ltppUZe/82FZdnblYLqpF4gDU2Uerd6sGV/4nAJwPKfpPG
jLGxJLTh9wmObYdwyR4X6Zn/0zeTrJIxvh9IwymHWIK0YOdh4xMHcKgwUDd80cSQ
fSY1Bsucbh9zMPy7Dvw+GinzLlDvmkzxSUnMoeWbAprnK7ArAec1dN6A8QR7k+sr
1xHvZTkKagatwZdgstnaJFLVw3QNxxEk6//94K1TnonwWk2kLEbwO+/1rZEOL1cD
G2xsrJK8Vcb9ZXTfJwFTocjlzoCPzYrR/tEFrIYChnidLlnxtgC5fsa17Goay17f
0B0haIyJ7hLWe3s526QDwzNLo0AlVCQcaae/4ea+Mf3Bem7v7YaC9+w7Je7XXIwE
OaludYLcgpK04zcUN7GXxIsHkfFT2qei6Mfy1JzH2dNvojU/iIAOui6F4+rXTp/7
IQG18Vk9cYiLaqU8dUtJJ2utBNtwGRzR2TYx01HiOQfkLUI7ytlcfMwinZw/GsWs
ftix1GyTCU5cMFn6atzwknlT0+gFdwrnomow/H7iIpkV0xeHWo1JVZFg5gGgXW1J
BCfvMCrILifJYd6jXIheWwrBEuTTMt7X5N2wOjpvG+xyxRhs++dnphVOAkFXxV4y
kK2Ms+bI1RguQ+KXDJQR656zwDrWdCJ6eosFIrrKvKTU9MNSlEgQs5DH0xsdFrQu
aa+xM4WPt/LTCEVdNaCBDA5idiJxeddqKEDVrG05/djDnbl1VJuN6d05IzwCPlEI
JKA1ofnFeHqOt392s6CR/4uVVkf1bove5TTjuMQ0XXEihYAZBotkdp8mWAidm73p
pJkIU6p6Y3zA6jGupNaUWCtG8y7BqaHbMKZt/6noL9HCe7zOi4aQCP/cQjGQO+t8
dN80jfXi3W+Yv7n3PwIxqgl8Mo0h1PkEwP6xmaN6ZOmq7qG2qrMDZT3ZtRin4IN/
Vf/exGg0NOITGlyColhJ3vexxY09wtNjRLiu3UTZPwJQxvq48dpnFn5nuNWVeWXS
HHYal4dNnfvUWprGF1te3EmpNGbNmKzG1FU85Hm79k49Aa/ACcymIzc87J1KCHxQ
2gEAKz9b7gv0HNDDzir7edEEnOjb60YjyO8epjGrU3e3AAoIpzYEsIbRuU4eD6JC
XbKtJMV3Lb4ZPpa82f406Q==
`pragma protect end_protected
