// (C) 2001-2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
L8KCvNB+VF7qvvgFs9SAAjKZFBL3xVD/lkWXn6zAYVi87XmR/CHUZzbQb5BcwVxR1PSUhJAgHyi9
XDA91MdpYr/HB5mtbVIz8+iFPbDKyMcOON+likrZM3JyBRAuudKH1IsraoB2eX4bDAOHysC5wRIs
SXEMkDoJ+Te/Gn3KQoSrWlvIvHkNXEkaD9vqdNq5tMDVut7o7qvvEMa6+zVgi+42P61oxfMXIn24
4ynI4bvtuSMmeajrtHuaCnDmJ8xMGEZwN7qcVMxxIbj9SKdiWm2DTyHhGpcD6Psr280j+Vvhtwc4
XghgRIKIKuYCXJ8Q64CEDQ8Z/5j2Ptag/Up6Ug==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 21216)
+mc60vcj7lAUAHkXjVW3tLhRtr3WdfQMeC8+S/X3NkTZSmc954XhOBupIEoPz6ALR37Urq99XMFQ
9IuVUAiUGfcAZhfo5S8lxhYcnt1mDCojP8pgNZD7P2wfbZD7dJq7T9/datgmB7zd1tilFQFLr5E8
NXEyKSHYeF6g8diseLXJgvvdnbPGd+et25X+nrp6mR5P7pD81DDFIRLWY+/g+RsbumcEK5w92d2H
BYKtafBUOpJri1vAjeR+rxfMsibDpW5lsvCr6CMKr1bP8gbB0ct5bbUelF4eRsG0nYgIQsh7e/U/
SkndK4aNyEXW6W96XpwH3mU2HsFh3liDzdazbHtt1DntMKgQHAVe1oCgljBPfqCWnCLR/nD1kcn/
gzKRjJ8DmbR2osH2K4pSCLiasNtuCf6mnwoDp1BQL0NVqATk2eX9hOVEZkXbBN0Tfw6TnIjdRk/j
OOlW9RtnB0glgjA2KJrwhHF+x23d5CXCQ25nDloZqJafPwGAGVhCNyCDTOpHADQckMUnpsj6vTPf
qde529Sr9hZ18EBB91lptwO5LhrchpjYQhCMkkS4ld1I+xtphjcYCiw5jpwXci7wVDZJjiAayAZU
vG2cnp/LlpcjHAA5YhKJwBV5QUwPLodWNCggCP0SeaTDV3gtPMli7XtrsU037bdVJBAhG7aGI5bj
U5tv5NSbXy5P6uyQGEohlfOghGiBRZVjoBFgqw8h5jiXBH9C/+/9fAQVTqun+vS7KFmdxy2ESEVk
g38X8t1OFeqPUbxqMi+EYxVRccHDAy5doXJWdTORYnR3g35tJVuFIot+mkNfJ1cRdHSiChsEaPOD
hmwyk8XIAK5mWhkm+8ZS0WHmTIGXC9Eyi3q7kVJJkuG0O58ywqNBUNdT21Y8g5GkJOWJkbbvTREl
j1pd1AUUeciKjdrK48MPHzBf94eBe8quJPBu+lUegvXs7tn/6S6ukz8nCdDYoVH+79zTCF/HDhUB
Mb6xI9AnUmlX/KCzodbQ4hmCoUNd5wjg5lRAk3ijEUmpt5OXFYFUVJvEuEbM7y1cgxex8cQNtZcr
1WyRi3QaxNojn0KPXx4A3PKycjBB4qhoAlIoSqHjrD4rWhwnT24yGgS+A2BI4Vml3cKnpdUXQHYZ
6GTYZRCTSPKtB8bZHOY/Es3IGL21K/4LAy98av/hNPO1xwnaIjX+ixZQkxQ+iPbtd4/GIb9RYCjm
+/sEG7SjFhmxQkDaFhBudf/YIHNa3rN49xNIb/IbKNKzjs3s9rlyaMJuDRMKzIBYMrq0tyzXvCY+
IFYGUFe5Trs0+IbNgOfqeGBAe1/WIq6uEZwhyTHgRYavJa8xkWtH0L81ZNWTTLgvk710wc9yGZhB
fK5veBk4YjJ9QFXwcej6HlIivQtljEJw8mxjvCsAkHJaFev5TOgekEDyieIFTcjGuoY72hLO0oS7
+34vSmpnFFAQIPGrttjZrjO8eL2UZJM6xmd2QOkJRxKPHV4icW/fM7cK+zcJgFvCuHHppLfflV6G
T9eaOB11jVqe/zLMwYrc/zv7xY2c9ZgLFNFlvm+gzkAtU9dMWChQG+LXW1GJAVb4sD/2/B4DkwtB
4Dwp/adoBBSewOsYEQVTELIp/t65BoYlhYh+MhfoV/cvIonR5cf1NQxpNW6ppxlCQw/8XPQ3RSMt
TNrIEjQpTZJ5t4l72I29lSBgsS3/CfzsncGdKf5Y4C6vjk4wxlSf/vcXeYJ7Ed7HX4Gg0sfizIl4
CFLPE+DlSO5Xx4YWhE7Hpqy+ViqfBkbHWszvH9iZwPYuPgTiUM1k1LPOZvrrQQsGt0OPeWsQcEEn
6R97hk1qBdUuGLWLFGWnraDh9ct8FS81Z545WG6TQY8+iVaUjluh53g72uUgrV/P6EXuBCqrUGzF
ImIBTXTnUyuFGTGARnSXY6UrUz10K9tGt3k0KscNJU5Mc0LcOcGVYvmRUb4r7vrNDWk9kq3iO77j
DmZQfqUsOMcbVZSes0PqSjWuM4gPCHBQlk049TePFdvQwtmtg2LcdKqhQzps+PZ1xo2SAHhlqX1f
X77tJVi2BMPXJZ55NyJVLc+IJ2/VmQdRTgvuAjvlK1wKY1f5EB4vVSh80NUjm8+86AchUIS4FbEw
aRY06YL07xFBVR+FVlKYAHfQFSeADpaOL1Otp2dJ9XC24P38jjJfczvrGAWNl5beYYJJfy4Xb8Kr
QWi4W7xD/EbfDayljeWUnR4Uk1dz5NXc1E/CzqIMQ9TYNEJpkxPWNEGkfVvT9+2HG5TuI4pzUsLc
KWsj+bL5qZECGHBiVAOzy6z1luOhHj/rgOpt8y55BCl9EUssqsxzUAH9YsLECop6ipDcfwjgR+ZF
lKUK36IvJcnkObMm/NwjrJIsQB+xbaidKlgGCIqwmUBto3y/wCXYh3ddNv+/9Caar/53m1Yhjqr8
ycT7xzQxYqSSRRU6aBLV8j5eltfFgZ+r0HQkLq9fOOREC9kUTcjvKRn6sLkMIun+Ht+GgFfpFTYr
LvltUgGETU3BN2AuMZsSkhyGAM8TPtPL1lHRJQcB+FWVeeFns4e6fMzQXDvakwCZbDhSYCFIpmrE
Pnyp4Cgq0hAO1bUCjM9Nemej8R1L5uT+0rz+pOB5ltaneVqo9NgwZqak73ofsa1B5IWw9tRTXnQ/
kl/2P8jyAtj2pgNmeaIMhDMLMh6gdZifD8CUybLTvQZ0v65aMCkUS1XqtW32fRHsYj5VE0V9ma2x
fTsUE1MDM5BtEU82D8lbwsJYIcTtJEFHUWyHTiEzx/tDDj6uw042gziyYmMAxQfiFuC9ZGSLN7yT
bqRo4n9Yil1k+khIG+IOEIO5wYMK7FXws3qRdy/eBPB+mtj6tuS8dGxNCjXgITIhxXXZ4akmRXBu
JV5vVzxRDKVjiWSR0mHSbBl+M9Pm572x29TXs/Yu2oUPr+swt6/wCU+OQgJG9EKjBwnpJai1BE7Y
EG5wM+GbPaBjtd66i6I7E+BBmndlMsOk1nlfhNtRCW8BMONYO974ptudHxht7tsMpDzSUkYfvrH3
Gr3soptLJttVi0Pn/B9FD1/8aLLNj/Z13RIsvXZMqzsW06x5WQguOe1bBTS1m2VLcu2Mg/nRBIsP
dG5bIrUFu3nxurDnfvzMS+rcxkzOAlQjmTw6Q0p/VMnHyFNHVKl7u3q+7qr0cVq6uahVRhtSuGCv
CsUo0YJDXdM91L5rAdfwijCGumeF62imP869S9+zLf+SaebYOpZvzUvBsx+Rc5NAKaKKx0bZhQLB
TUWGTPKlrYtzT7vrH237+r/HGv1h/kkFTLt2eJk7NVRaDhHNhaq5L3ibfPjVwknUSVvSydeh79mX
wxOFzsKyNPBDHYvRbeAde0uC0SwgZXL2/dyOn3ZkZHklrcDGPW7Lz6LX8gU9s/A0vfslH73s7dRp
ZGBdOznw13FX5KTJfEYuMQ+lFhtmMRFpcawF82R2Usgfnzv15ggSN9G3hdO78U9wxgjSs630qi0d
5mmQ+lkLYmfKikWqUHZ8qvA4IBtXDUC71D37tzRqRXXI8kzv/mUZaT4R9irHKj+rg/lQdvPqK865
qB+ihhWUzpz+IuaGbgBe8C+hUsYhqBWoV6BgnstjtXoA4CKVLECMPNXBGp50HZwvf+dZZ2OdOoiv
gnDvKrExErISe78iTr8uDpu7tRZeHbfIyy0o8M4pOanHh16S57ZwrxYWhBmahmB7w7vvU+jyHRZS
sOtPY1lDaxQ2nb/cR6qTmKvWiOujT9x2rJb5g2R8kAt75cQynJAI1vvpZJXcl/05YW29GEzyqSQU
2aOGfIEs1x8+DbcfgEAeI5L+FKs0zPkbpfM/TQznatw/WdD15qbw97dnKQJ1TSdr5Nh35gl9X7GE
GzVBiN4MWa84QyRcX1AviVyPxmBBEk62hptH18Is/JmZQWWUmArcYynVevvbFyToL1rhzDP3IjIB
bnC9glEIe0vGE/KKa4hHrJewp1VFN/8AIa1/W8EGEUpZmWi7qUlZGcim/Q04labFYOZh61098Teq
bbnSpGpwXyV30xvdx3Ps8Ovq7iQxa0h2ms5pdVa+wKcKpaYRLBloxFgj+zP0rG8RVoNKUUnmjUr6
yqIH11cq5Uoo+fF1XOm+KsXeGh6KQPmLPLwpY0CfHqq+KIxiH3pURP4wixth2OC4R8OJs51FOVMX
Izh43ycxlyRxfAVPk+CGfWbi0+yzBQEdqXZska1j4sWOoc1JCiSwYeTO0Li1bKfXyebA/kqU5ome
TunOI42H8/G6iYFHSW5ChwbQ2VwzyuFx6Qd26oqAadXqt3cMD6L+0xL+atIsXQxzw4Rpjp8WS79Z
9KiXw9Y8JYP8dVcen69P2g8w/MDE8gP/mwLn573qWnI8VEm19vg8Kl5ehjXo9hOrzD2qhlbti34f
8quQPCGw2qNOb1BA2kvlhyMMk2OEFTRSqSzUWM0Kzv5AGaVozXvvCKIgf7A1+1cObqwTiUqtQWh4
5cP2O75u1/28gmIHq5cyzV2S7As9QXssddCKKANN4XfJsHOoYhfuxFSALITtdsnfIHk/TyOlHJLt
g21kYlL3DL/E5uK2EGG9FLfwQmhO8woTSfvcgBJdzH8cSeuHEXCWzJrQpHB47RjTlL3X9NRHh3w6
Wj7y34PLFfBInj7SzPOFRCdSFQzaRvlY59y5B3S3JgFTOZo8bV1JH8zisnpxP+akPs7INi0Yk12T
L/iR96TJy7b0uDGd0unuXeKcQ+/H3V5UGkrOKYWXN5LVo6n/EckkRm0780ye2aGw9aorPkcNzjrZ
ikdu5ruYnTF6PiPps7onwgstPI9ev1SizE0oHaD4ceSOR4Lf5eAE0YPT2c8acghL89CwCs2Zldu6
W+kWg48dYiQUFC3YGE0dwblcgTlEa+znFUgzo0nyRV+d/EHWSduVL/LYI5MDeFuPJfPHZzu5Jopu
XzCsZm1R8x+LlIx2DH+FZvi8JnEAJY/cboL4kRVwRrLLHoxfDgZwnYzJjKL8u4cmrAzlSHEkEvRd
+x1i+qkCsp+6/kt/YRNnjmq9XWE9QVXiu1tjSbEWAtGN/hsN6eHdCLKRI/4WYbd+oh8saXTBozC1
lCCbwNHx6+kBbyeYwQexj0Goby+BrQIBaewrbsA32uvjrbDKnE4hO2+zKREdhxFdCdZgflC2Ri0O
CqeW/rnax1cvdbRG9MSK2b7pdwG3yqFbhRO5MKg1DOujo5cvB+TSeZxSNL+CIiZCz3ENG0teg1/I
szo3X9Ddon90P81TJ8xLO7/xO/lzr1BX0kXFBdkFX+iU6CuMdeVY/2RIqekSG7A4UKYOJkHD1eVT
Fw0DSRVW3ta6HoP5Bw1WFuVrtyHtqwyDF9+0dqBtPPDvkpl7cw1ybsQgRAff0NMQLFusiVlvIELX
4AV/nwqK//QeMu4faVLpU6ZR5Po9k79MleRBSxmGJ/+UpSI4zZpkn22y4GdoGxYF92FtW1cJkUNQ
8h9keQB3VR/AxARKEJxsQsTaN9ScRCrJ+qX0Fy516o1WmzucHBvUdgRqtL59Z1CNEQQmaTqqaUiW
AfC/KoalG16r4d4hqLXbGxc6tmKyhpgKS5S27CoTIhnHL1ewYn2DrDCPkTeNnZ77Ags4vIFHMm5k
XSdILBkNLBUN9oDwDA//GPpxWWml7cRTc+gqPabhfwVzzzWmqW4xokmSYhgqnEifcu1DX4HoUMqM
PAbe3dDSFHvHLsq8LQ1xkYIPL5jFqq0TmsqqJK6UqSNkASHkDD9crBkkEM33GvaUY1jx20EJGCxk
+rMOU2Q66OtVZyzyzmlR92PnYaMA9yYyz3iuObc9DGOC2JHbeT+aCRa2X0kGsSa1WZM1O46/sG9s
1h4tCLospdLSbN5piO2hBWFP5eqJx2ZmFQ62S4BZ/c7Nsi1cGI5dD7s1NJ2SvG6NgtoAKIZnWjA5
AERMOwPuOLy/ntzksluJetuMz961KLdn+WJR9cpgGQKi7iSvq/hK1QmayGhoR14sWSJI0dG6sf1M
VAoYJ1ndq1L3+OkR21yLCt7ZoLIsUat6Da9xzVcbWgK8DJeEXuoZEo5UnVSit6PBg7hNh1eyHSZV
tLX83Xh60qCh8lVGo8N5Ds0SfC/xF7ZznsNsunI+qWIL6kDmH+HudJC5VOGBoTly1v5rK8gApnh4
LtirQhSYm9/J2MHRpyk+345wc+j4KsUgovoBBcLb30/arkhFQEHR2DogKUYK5R20hcHhj1vYueyi
iuTYeOjPcB20ujCtryXacFS+FdFMOYm+uaqrybSrpU6mcFf6NU/GhLhvnP4cXO1uHY6o8tFaS/eD
zmnZPVCWdDEfMErqe6+TZ+MdKzeH/aOr3P83Pb86Hzsb1E51n0WolM5pkgv4D+/8hsWwGIJTthWT
nL+zwd1nutDqs++/SqajzqkqI1Q3Q9WG1tfKonYbLId2q7582dfN9w7ffMklvlblB0CoAQZEdf7g
7lwTYvXAo98lfNS/EPadwJq6vHVf9svHYNH2zrKwE6MnsnWl26xJ8WjazBjtZtdlRVRsDWd/MK64
FEW1ReFacMC8EmTqegYUpCN/fhmBxaHkP9C4U3mSTblBvXDgIPKCjC50Il0t8burToaWC86PTXrr
OiazRwMwJqSTep+/IDW1qX5rPcXfT9EPmr+I+gFUHc2z7ju5frbGgt4Dl3pCMxjl4Bc/mL+HsdpX
MMeI6DCRc8JJYmyZsivZtJZ6Im7YqucB1Qkmw9s7prfvdMGUn3m4Skv5kIPkXqukIx8GuNPYhgpY
sRXMJYLd4lMKPIUrInePGQZkH3BtTKI4H/7rzyud5HHkN8vaVXX1zOznvcAHSJL6EJ9SVvYykmSO
QhFKZCse9EaB0BP43QKt56jJ01Hb1Li1jlxgEo5nvo65VX9hKpyNY320wwrU4Phu55kODpCSMuSl
NSvE/0qRrH9IjzRNvaHFWuTd1DNUvYrz7j0/lPPw4JzAqccWyAMArkLM6/bPlksrJajDsxmZzmEX
ZA44Pq4s9izH0e7n7bZeYGz9Sl2lslSOUOQEwNvUlRLfpYXL+7/4N84JwGdy10kLNRtWxe5TXpIB
ryYBB+cU9csfXkov01XtuH+xIuFt7lwUXekJ5eeXja+UqYLB99b6EfcaL8H52Ouz958C+ibff2h+
hvt+myyianiCXMxPoTSfQtR4G28zSxoYGBPppDT2I/kCkCd5NhigM6KEGdJ8J6P3GjdShxtjqGE/
qcRiaVTFY1NIMLa7RqAnOJ+ekQlBKLbgeOr9TT+ju9yq2EMuLVVSeHGZhzbcfkA98g6CW171TBlC
Hl/gmBKGN0JI9MH3reyEMT4Tks3KFiqUeG00YjmqjYmmm4PhbpsisgJGnspR/fMgfCRtYkGBWIFg
75eJBiit0AJDXqgsAk1acnFMXVJSi4098Tp705ATM9W0fCcgfiu7sw8sv8QiQ6Ilbi7K+amqYCAA
HrizKyeV/fPOc/pAqHJkeJSmUHue+7fBBKwOWy9KpXX3pYPJvwmW4UsdGrrHP7owxrlPCl7y6wdx
nhxOs1BUekDM5clBteA9O6hye3zb9G1Cx0WwJTDvyHBXqUTCXYL2aDQq6e3Pq73k0TbzFxwoqk4i
yLJAdIY+F1XugB6Zcz8Vo0W/aqDyFRF0SCYzqD2/qxGpEn/GpZKIEIx7c97meNmWuWZEp/zwtvJe
2x/1gfe09f8CDzhcScjVpRuAd6McE28ISor6lwPiBgqZ+IUF5eqdsyQUXsY/hT/Z0jJ+in/fmRHV
WA2+qvojm+YzCFwp+SR5ojac6NpQhHwNbTkOqF6TS2r4ujxDasHGkK3ChFSAgCLorHYxSFsj+0KE
q0L1g+MhYITXhA//q45b3y1FZQb2LNQEC6t8wIH5kvlN4o4d1eGYcRozJZGgZrUUIUUm3ZB3k4m9
LPXPwq++l2DEi11bOih23jly8zeutYpBnP0ffpczyDAgxEIxWE1tPMGZSqiqiNgd3FiPxh2dsgH6
OmGYNE+Ga5Tp07ZpaEMFFNZQBRMS0AbwFcDgzunyd2UXG+tn8fBXGSWxauONPAN/QkRlku1Kv35Z
DRx4Mw4QZWCnHCmyZApCXmgNtkj1Yb0CA/NgWkbl0EdGROhz3Hm+24qN+lvM/cfhswQn/h65Lbkf
JvBKWJF3HMGrNh9OEdIFYwzLI1x4zkvSEOLG+stldi1+YoJrPsAVuuzivhMmzLzAhysu8PDfdblu
oEztU9bctKYPmNEYYFT1uKTop3dVhX+THBVc479p3rjf5kREXqgyg5ziy7TczSyKOKFPzDtqSOnL
AnwCA700aRplgvwS3rcZaxqu7hFfR2iSzFzNhP1zOx+oobMlJgl1wM3Lmtpe/eWhzR7EhfSFSFL3
l+vhy9DuV+vHaxQcsaLo3xppooP4fcNuOvcauWCWYMy1/14dk+y+ZVQfDTERMKXVBMf+aTWmEjgT
i3zJ0N3Qhcwd8Myl1GFl6RpKMpQSpkUenvekwQBE++9t2yXrv1HW7W2tZ0wSAgSqjR7B0ewhdeyR
xgtZA0v+MT0IYMKzNG0SWG+xMAyg7JbzVpaXs6L87V5yMMbuOIzZLrw0ft8Yba0nUvMaY8u6k0OH
9pkhdbT6RDE7BCzcEt1oIA3lzAlOYXincn4rp04psB6SmjHC7DqDg3h2gNDow4p5JWAMa+TeLQSw
7apejcWz4mlcSev0HeC5viGGE2vCCSN2Zfv6voEr/lMW7XjgbHwTFoB8klWUYEXsTnfTSAnMRla7
Z/nkhvHbeDSu7ggIzu+WmYTqY43N260HHvgFliw5p84vHLosysviBTZ0j+BISqArn8i3XOBfkUSk
c853xpnJnS92zS6rL3eLaJ4Re2DCIWcBFOpS+1ZerjZdpe37vOgYYA+hAswYxLwBcGkNnZBHXaqP
G2vBf/yEuUVXukeKNqRGYNRUGfwASUFelo0LmX8nB9GgEno10I9zb2VsbEytzQTaWDkMpcRxD+K5
S2/wbMDZt0De/2XQrjF3ZcJnLV1S8pVsiurvpIhieJWCg6YLfDm1fu/22A6DIo7HDt+ol1T05gwx
wbGYNhkYP7nLFsENky5xZxND7D2PGgopGfeSa4fv07XClJikHh5A8jvxmHdLojVcmoiXD0OMsYWL
dUKYiA3s2l+iK77kj6dTb/efS6Z5HsMSKrDt0nZYAxaoAZY6JLdaEw08Uw24zenz3yrUpVq1LFR7
jH+NATd809zFXRoiwe49DtoSHHvNoN8Uupg6eluaOcznlpJuzbEI1bVCuK7+uXmcP52XIBrLNF/Q
WcGxBvnnpwRY+UkvvzTNl0Zgcv/5JabBs5zpx0INW/TRsKLjqN0+N+jcLmxGd98teAtOt8OSBGDN
Nkqsa7KMIT9nyX1jN9ZlCT+Ik5Inud5jfGQZeDoRkJeyWerju7deDgSwCC34LMJAwjGRBqUDFFQM
zRIigN/0+1Ft6rzavOZMo/qRj4D4/C+ftJGxfCdw4ZmOzwJHE3vQeiiuQYt3LQ6y9fUJzyff8VY5
X7EboOBBiiEsDSZLCAhzgZoOPQXzfPaBsSlRfPPi6XN4NHET5EunHDKt+9W+8IEiCBjZZ2TMWpGf
vkNhXHiXPD87+svwhrFstblaQVbWbvSlNgXosr1f9Qs+fftxLuKyfJ2sp7sn2wbpSwZ0xVLmgA8g
dwj34D7Ysa5sEYHzIQtWihsQc2bJngZ+hrQQl+0dUyNavYKiKeqRtlKPbITdHzF9I12WiTTLddXY
1SOgczOYOkonUKIGcBFktA8GEBO/lJdY1DQvMAAqLWxDV7PAinkQkc1Xa8Vcm748aGHY7G7KDRNu
MsQFHJ1UyDajBtgZdf59t06zQ626hKXRhjl+36SD3fA03BS0pZr8Gd/clKP+gMZ1YCSCXXoB6Njn
wODRGht0UzVUERiCc4563krU82OdagcJ3NVecVxNUACO0UR9WTJjGxJalwcGiiaddPN1P0UD9KlO
ZojmfUAxOzhnvl4C3ml3m5AIVBqvfWBgGqCAcCnA93bgGA7RpSRWf+O61fFeQhhoeEflYdzNewb+
NqCMtokT9Wj80k/13zydAaDOfnCq5Z54/oChJ87Kv1Xtw6yqZFz7IU2VS3IxuKdFrfYpp1WbGS3k
wVhj9YH6H+Z9jDmDjabnwoiVCGY1MCPKF1M3MAr88FAEsZE8uiK4bR9DHiOaniCFQ+rtOo/L6A2K
NZZhrGnYZg8Ail8lCq4lyhpuEaOX2hjownP+UUd//KHvTem6tIo4T8OOW/dZRaGo5wPmJbRNmLRP
8dLf3wwxKmuHWTo9yOyCG5SJqK5yhpl0H9yldrAGre/f+HwDzowWb4P/58Z5lHMF4Z8SqvWwEDyF
LA9jFrbE+EPYRyFlMxVT9ULcjpGzjOmbq5lQQI+wRnwxwHs8fn3iNelrhmBHJMXwJrGTyWtrDO8q
Qrr+ZDyi5opGT11/MUlPlh+L5oauM/NF4pSHQlndSVlmaLUb41rJj6t21tHDcKx68SeHcyOktyFd
8CMPp/q0FcXPctcl7fKHOko3QoxoXdplD3XLFFTMDi/VoOanejnB5cdqJBbNnRTveO3Hp1gcIKaC
jJORPhE+ngOwtfxjM69IS58oIOrvaHW7rmaoniGQH2GBo3aVIJxwxUD6Y2zkNpqPgyC2R52ccyLI
L7rZYQ5bzUxaFXbfA8BQ8UyeYq0Z+DGiUWBc5i7SEZwa+WnoBNYZY6VZXiY+DhUWoZf8q5uC+LAY
YARfubzwJVTQ/nzZ1g0irMJRIgx8NREXbJwAJcjLSVtFt3zPz7amjUhkUhRXxOCTiXJxfgXeCOCG
geainO/UJRByxaQKVtV11M4PoMXKH4uhP6b5Z7wQyYNngej7TjkRui4poW+upLTj4Gu56tnjlbox
Nx8YWATzuToa3eok2n0Mxqc6tyZdbwjdjN2WagIo+bIAYrce8GYV0xjF1t3YWCu88OCxADcaR9uh
EFyuT6B3V5rXFEIrE19T5NDIEMV71TZ2X8ijhoJDUMYCXmj/0Kh7weZRWmwXJwP50W151SNjoLCE
lwGvaL4rIe7uNASKszjfXYlnHvxUBGvOSrFi4XD++qaRr9v/169i8qjDHLQzQuGtnkHe2uOLeKZ3
aGuj5Uo5bB+RYLJzsB4dcVTBn8C5QyZgOY47c3M89vY4EvwNo/Ci/bNO1zq6ERn5tPet/KZflXjp
JdCARXoSdlBoSeP67/d3yZSxd6oIvGdEUv6efC5CT1dX4qYStLFD7XjtEpXYM7pLrc2W7LYxvQdl
q5ODEDljJn14tRSck+rSKYIPbivFFKdHSUYZ486W6iCjU/592lTX3j9krUj01XIh2ICymBczmNDh
jXOwLTxV5RpkgnMZFpHkZdVmOLOKh5y/XeGyEYuQgCHQdl1TOKmNwJPGtSatrYlRd/QM9T0voDM6
dCt5n0nFddJOqEe51hIUGfZDxFWJNOMHCxaw38ysYMpArDTtd+hnC05r0Rz+w718dS6YHh5ePwoB
dy4iDvPyEjFrcGE+T7hh8lLih1mt64czYGGIlmOuHhUP240cVNxR2gx+MPMR9tDMKRq1LD9BTbHO
B64cpi6ZeelOAPps6MiyYaHBPcIIF3HRkXxJxa0dPIg87kJuaAuGF61Y2A7e+lbpoQFYc5UvZHOf
RBAeN6cJ0qnxvi9hVULrHO4Wrm403dKox2cZcJSAceV9SAt86cSwN+32YsUSKVvJxDVd3jHKV+Hu
FPEk+ytrEKqRZSkpz7ZnlxFw6LG9BXAKUvMmOIn8kd8uTLAWHAcAt9rGItWvqNT5JPgbddQ5jjwo
V7vgBEEHpgqvoIw2zCMaFFM54NbhFXm3WY1AzTbUUDQV/0gy1X2gL/WGiLY4+uHEqEnEk2v8gf7u
F4B3dMTUVaGyC9Y6oz3sAHWqLUXBMFxQMTcVq59Rynn+hXFaraCUzMLAvt9obxrVctBY2zZtLkCn
nzaLocP8A3shmrIoWIqIJ/YMyKcupdHEHvcGZV8Swee31rxfhXFE1/9U33XOABL3tWd3kMJRAmY2
iYLWAdva9a/yzvuR3yYQSM7AJVZu56Z/4jodaSqfqAie1O7CCZX0kE12YEcmQsOZSFp5zbmXZEfB
oKKOsgkYLlKSWZd4wwSRY0PEoLdzXyh+T9lIeWxqAPuCLVNPRQceW1/G2bhUmqV8NEPCKEk6oLkj
p2cr6sR++97/eYTIwQ0/mXaqwW8NEu1DWrUNSiYkwN0gpR+rc+oAR4nV3JhbXU9m1wMDp2cZRqTL
OXycEdJer2X/1Z9Lmm9ancRkhMKSetbesZhgnsqJlHnHryRNyGLG/YDW4iEtR+68VpXBLIaZPRn2
d/JkJB4vdTDgR8VPQKZPWeA282m4iZtCiirXcW0yJVbvXtmC7ocU1RWJP3MkXYAetmPRiy+17zjO
jPXa4auu5qdfZoV/+zr2e5+XR+AcrDClA0OFPbLwoR3SRqu0NAHptdxC5K8IYRlBHl3dVZte1/nS
EsJ0OL4K2l4S2i3TKJ/do+lczoc2Eq1V21mKs1+Dvipr7fo1hH9ws8aUkPWwEE+aGPo6/hg5oc0q
y0O/jGpAhPbMEqvUtTyvS4ZPe/2VXy8YsUQSiRgO+AKjlE/P1ONuLUjpR+WZqbOezs281eZAoRJ6
Ul6PF9bDQNo5MWiyjo0PHWkdvUW5fkmEuDzkOEBCZgQrRstNihsBfmJ5vbZ/Dj1npqjeU6z2EwWz
MLHZpLPfjdHaV0UaAKeSgln+u6xvySxXGmjyw/OzUlE0yA5EqLLRYp2O0g9jlzrMieiyYp22qEfT
95IVaCcMWAR5XyeODmZHNnmK6/ZHXWEbBnbkEOcJcw0p3CZRjUjM8If/ZfDZFZW+vDUCHjJX7V5s
0FiGvoAs3gb1ni5g6IVLtbXCdqIe8zs3t8dvjC0GJx+n5Rli2fvkbcbXKzwxwXmV1I7ptZPY3ooB
eIgpy/rED+g5HPCGKXirWFAiCcsD132Kt+eilL/yI57YI6auvoQ69TeL3oENKUbiHYzjBjqqOVXd
HWbnekN3//8Kuk8y9BLgjoor5WZkx/ke2WzqJvpJkYfdgIGhA0XG8acETV5sFb0JEYXquldZoff3
KinwP8yq4RrqmBj9Yh2W3cNjbj+dOamErMZTBsIhcm6Hg7qC0+FWd08pDAW/BYcaoYoyCHn3PWtM
7sUM08Y2n/nmZomOGm9LAOSf5P4OR13CPoYFDePZwm1yMVlGv9hM320wnxNwHAhQIJWzzDLwwn0D
rziA18PKg6+RsPDlsnQ4I+wxdRCLWNJSccHQVOdMcxRMX+tu4zQ2Hs4nltTPHhvHNfFc/b4m/6Uv
yGrEBeDr+4GgEIXKQo0w8WR4HiwkE/h/KuaianpwCbbHbAqGS3zzSiB3uVJRNnQ72oLZfZnR0DXK
9diR4NKfa2KaQ8XrhTbD2VumrO6Ofm/L6sP3u854qE47sJH8RQOZT7GajCUnmpEITC/s8zgQRJ7A
b7I2xjLWVsMJO1sENxzgqj/HP1IgqW/Fxslj0uNdeUtFKwcQEpNNhBFO5O9RiHHuVdl506yotdH+
PCijOfhkRRMQjpfLI4Mmg0tmUMGQHzLsBjw+t/GJ6MOhF2aD1wzN94iQ/2bAUfE73gQuWY0+ZbYB
HLYHvYgxiD5qT6sBrx8B/bD0nfERw0T+iTPHilYRoUd7sUwoQ8Yq8Dq2SoF2ks65836hQdJj2rhS
X9Z8j2hR6SwtvI+IgOupuBHq8QuPzQWVrVZJ/thPPpQK1XXLsR7y/sny2G5sWvewlQV1EfhrI/QF
R1wx1+ObaOn9avLxtCv2ghgjVrHF/8dHVIQdDsCriw43QKN7dpCrj8/IBqov29jJbEVEGNDRM96D
utDYCPgVPq/hqiGZiatvUGW3UxlOQaa0PHjVMlvAssU210oZI7QifaCjEGVx3z6v7jJUXkoEBi4V
RiYl17BFGRgd/LQF9D7vHQXg7TtbInbxJxHym4sFLEM8SGlMX+RBw3Esv87RDh8TimMbGOVVtHHW
j8ibRN1Yjm1+O8s12nkG77XvB/fYSTK8Vwi6t1AHAR8/MQb0fnwxdrF+waRJE2goccIPbaK3nRbj
mUDwA0OxFZ3slE6VUjxH48SPoLlwdKCEIbI7V7ILBTf7jrtjv1SqOzf+VuVFO97tU2jh3Lb2sPAX
5+j4BKeQd5YsgdpfiRhhaHVV8u2OfKbv12Sv3mDvi09LzB2hc7dAysMNa7QdkcZWdEyMlsiBITEr
fJce3o2yGKroRy/9hpv1816yIk0Mjp0n+YE+qdu86pwDyxS7cNDVSSOhPuCx5KrdBfda/rZHE8xR
9DfGjZYLHPX2yELfJ9/arJAEcRIEf3SLhzZ1kcCWbKgMLKvpYYRgVl3nhwgqavwIrMP84bPhlRs6
kOVBSX5KRHRc0zbBD3ctr26nEi0ik3K5k0jtO9KVlUux/fu+n2iRRWbaJdDu2cRPbGDSACMHiVE1
pqAo1K31p04yGmIjVKZxwY6XPDETCCdlBPvBmS7625EhvmJAUR0/Q97TMvLeok2P6cAE3SG57/TL
xqFH+40TJIi/U8c178e9PsLCA8ZKus4iY8RBihdBTgKV8LVAxNZWAJpF0X5mbQNpqUt6JPdInj52
ZvJHy2clsueLu/4PGYsotuEi4J+Zu9OCxxJkGOe9Ep3QkpRmums7+R3gOqID3PgSL1V3ueywHn7I
b1d+AUjhsN4XeWIHNJAwBavwmTQj1FHTHJg21gGxjhQPH+EzBdLR1tDFVslf5SBi1eI31b6pZKJD
Q/kbR0jZRQ4NbIvsDChW5PIAytw8bfkAnsJrHkFq2JisleQ0/6hv1G5ALGk2fKRRkxBON3ir75zV
pqFeJYZ321uSaD9wsbvdIatgOQolfwBTorQF6LRy5Y3ZV3xCYcUIkF1jY5ggsejmSnL0O3fNH/BG
fBHc5ucNBBaT3uevsA3G2gfyLl0xmR1Mfu0op8eKuAqH7e/rzxGdmPlxiDejv/Eq3JWCD7wehHC/
rhibNS2WqEy4Wb4sMtRswzMyB9V4vQzGGqnpIk3pD6jcmCc2P+kT8insHu72SH0qpQqFj+cFPogZ
Z5igdU64aijRblmqWqqHtseIvZdfhfNNj1+2j1ByTc88RsDoDTb28soFZ8dG/FGqyINO3mTMMo4f
VeDj294TkLL4LVNdSRFb4Z605J/hqj2DjU7L5P3ZXyXtuH3O4RGWI4ZBCy2yFo0UhF3BFSQROW/Y
kGrS/osqVkqvA4x71zMjtGZI+Ri2IH/CAAuO7wIrPuY3LWiGATlaam2j7Ze77AboydsRpbWxEJHy
EOpX2KBl+oubp+TgeNwpTEKSD0NTAUug9g9fvEZEt8T/ebQFokj1gbjoPAh3G1cbBTQxgqWN9kmI
9PjIb2HvvuMT+spleNdHd/Hep6vrlT8RFUbj8I9D8QCZOsglS74zazyNVnSe2JZUSZH6s3hj2iox
aThkgC1ER5Yc3vNilAyPLLxFzCnDWmn2F/qs5qamAv+MISpIdvJVq1CPnfTOXR5jQfyvGOLccpC+
MUSnTbHFR03Kgk52ajhclNMPcmYAu+egbxcCa7O3ijmDn02JmoOb0REtYULIit++u419pqrwXedV
y3wFYatFeJyDxWVqp+c4ZVbnuKEII1vjjkaSwmynkyPi5PlHvth54TIxZfSEUd71eatZ6aEegTmM
0ikmVTwR+rMvzup5JJEbOiUcl5rQyIT27ucuey7he2+DGST8Y4E79UwFHR1hIeyRm7H2fxb2k5Fu
cQW4VcO09RwCevSC/qAbDoQNCaOJDS8RIF1mVxebd3TwIcvbqX2BCNSAkrpZHg8J4n0cyWQCprvq
Tv4n1xf+AJm4QyUDqjK7KwuiVEqnaMWt4TLiojVyROZmp25TIxlFWfP2vyC7uWiem7ehOXOuI2NK
rLa7Jq5RK+RYVAhrFzRTp8Y2FurDU37Ms7U9pGDgmXfEtpRznLg4Cg+iOEROyc0/CH4B1HskWr9a
WAQDPbYtP0B2FP4gnxVni3EZCO+tPslXIzvOhudCa/8mzw+ByV7elBbZOITD/kERFdZvkGzQ38AJ
BZ5X2y9DqfFPbF4ei1nRoiA1xE9DMy3mGm6TUtQ9ne/FVQlpbGWN0OBJ4MCMgXxAhTw7pRIHAXiW
WVANNGx+2gIGZ64xvBKDHIcdBFTaq1KbPkS+DfsNjF9FXW0+/7xMGVFm3uo0lDHoSdW3EKciGtvz
X41R3KQ1IGhjqrPv+agJOWnwgBFSVzH5nIGR2DUWaKW2OnKz6MhbJPko9ui+Om35LYjT6to37p4/
1JJyKA17lNspw0SKPBQ56rPoBQGoLdiyTGrQBn9DbVTUMYFq6/AFv/IbdCOvexcETCezdcuo6GHU
kcA/Im9WJ1YfsyB0feS4vnuiZjLG5octUML4/1vBGFcd8+16Q258xCDOLCVi5iSJbdQY3Sb4TPQj
6BlwNNsYC22Ad/4TU7i1KUy/lMUKdnsulnAaK2lgKOyVBwLK6FWMWe72DXN1TLOK/zxWj2oI1rnr
nVS5HEbK2VfqVIYtSgUBFQ41gwH9qL6KXV3ZdjJm7dOQa57OV4mtEI2vO+B/Dtc8aP2Q0PztJq7v
gfEUMOx/KQ8glTGTxlrBT18HfQz3Tk3jBQpbEflXkpC7hWUCTv9UfrCQJEg9BrMme9s5zD80/x7U
fbncsT8zkveVfohI9QbpbSDmo0ZT/Hq6AYAy/mTlb+6Dher/A/gjp586RscKjw608OVgWG/L5VWi
YNXcuFvEWF8Rll58SfZzunYkP1jLlfqL3YfC8WkXOo4BvIsVi3TXnB5H95/IsOR8eQfuTO5fCpjr
HsOFpW2MDprOsIPv17rca8TCijs00Z56fVDRUYLH5HQFbNArVdjPfwUx+HXC6d5onO23VngpdXSw
ausRujDJwDZ9F9YLuXiKURR6Ei9Ljo5CCF6fz95tLQfsl4vSJgXonEq+Al53xLA9brIYii+Kx7ns
riF4qSNmZXBsWm3R0NBaHZ1jbJIqE8YtF5KLjeEUOsXrsYNGQn96DM/6zTIOHaRtYx0+jjiYmxWh
MoT9AbIs9tjHSAhEgVE+W7o4mBx6ry66MD4GQhtKPAx9hVRKizPi8rCLnvrSo6m5/4GFCrzJOqCU
vDrEehz/OyQmkfVdKjCSNpU+J5TpWVzGuOPbUnFMjO8qsg6BoOsz5kjhhM0jtVkfQBcPJZGUjE7u
M/pUm2X0qtlKiKKUf+5Xf0Fl8jifO8+JhDGnMnnwPta2MlXIPj9mpeKJTAmJ69e5ELP4iMuaQVVw
OQgbm+iW0oiavp9IAZ+vap12IDs2nfpCXcsWHkc3QXvM08gXEtLSkR6Zbomc+R1Z0rFMhR5u0fyr
FeTboFycm4BPpq3Qc1MfzNUzwSYQ42FX0lSI7VJ+KQrNQjGOeAjhMzh3AzfBSVduhx86AlBh8dzY
Z8NISf8dDD9lLCRgt2e52rBVrAHui7a0d7nz1h1YwMXMABx6PjuUwrIzVIW3+BED0d92Owd3OU+G
tve8L5c0Y1vWuC+28Xcuk1J8hrbBmchfyszco64Su1/QP4LfdQRPqvg6XhQP3iIz/DBZO22E0Fsv
En5QD9+OG5lfyJBfd6udSGlhtQ59oWeVd545sufgn/BG8x5IGGzGGb4LarKWBSEdCVAr1KabTfP8
mYZA7nJyXo0XyCfPNTnzQSXZ4yLK78MpJUK+jb3KV4matHif/oFdpBRsjgaZGZhyUDx0aPoI62/q
4sqxWkU0deGpsVVRCSNiI9FS6xx6qIwCAnokJKBggDk0rAucS5L2XoWN1Hp4hcgFHU7SFkFMiwEs
q6JDIx/HXJ8QO1z4ZTkvHORt0GNWj3a4mb/fx86C3XBxiDqcsRmqp41ugyJvE7XDcj+BkNrkm7Z1
oqtHO10cAouU/RxIIExjB42Y7r2cgMo1uT+ixPbzfGt2p9f4XyPCmMVlFnaK4J2T5odUOTDqEr6S
5XkPUEXmnwBZULJ1fagFG2i0Zhnn2/P0uGZt2v5i+ZuWXTIPYUhjMAkH/wlEdILp+ianlLZ2n4km
eEZ+Xf+MOfkPiEoHaaNiBTva7s6f6h4r/rlELfmA6UiksAGuDOfHMGZUMlZnQNs8z0xLpYJlWxNG
SL6gpP5bduNcXcEfTrW6bb3g2E0KaCwX6gOd5OVd4nJTiXVB9TY9adGDFaOIYc1JJBvce7k9/11N
GJimwvCjY+Ciz+9Fvyv7MQ6c4/NPVkCEHUdS1TT8vSO2N9+CyJXh0CJ5UPaPZPGNt5GC2jTzJu0W
J1zsbgBRVMVyNKC54V9VeRDkncC99nFZNSYcuwpNcK9Trp3ZijkigRsXheHx+v12BM7zlEu+yuT8
RaY5g7jDLa1wsgGlhDocdXMt8rwAeaQp8CpjdgT/AIZ9D/TvnS+GVJiF5a44wtkNJl4CiYtKYM4D
VxWrkRvsk1mPLiUwSl0Urq8uyqN0xtllBaHJvyFNxt3fR3VtemhXSUFlEpjSp81ra7QOQkwObVm3
llEwxDXKDe26BkpWwyEsFD9POxCeEM8zs2/+rdeCGs7X0eyJWstTjYNKUwpWrgSleYPUoDJ61KNE
f5i1snWBnBK1SizHEnapV+MSwurFwq59Vd9JMD9zrDPDM1RXc6TuVB2+W2oxczPAQwmQ/rTyLJ9q
t4WeysmipHXsXOJ1ZbDlZdfIONbv/dnNB1bg5RNF6NKWo0ipOhGnJPTHTMbx0Ro67a4fvCFIzl1/
bmmIfHqATKiXnW7hqkhxQ8fZza5NDO2IO4ofVhxzW9214dJPnIzR5pNCHWccyw/7K+8AF+1YGA7Z
VZ+RZzBlZILBfON0ZUArjDMWX6oB6FYumrR8n+WqiqnBjR4MC6PV9OxC5BEJLF/XPMvfKBbSMu8w
AK3tgP5IcgDhLFuhnM23lIY0qOVmkuKmD4l85rKEHoI1NeuR0Z4Tqv8y5WR0xJj6eeu88WzwETIA
Cp2w7Xz8id8o/uASL320x0m0zkk3vPD4HcFaQyngHR42FX74igrZZv+533FQVOX5WQTQOl2hVXe1
nH+FMbbG2+NPYw23Rg7pjMkMXJj4Le+oWI1RjnzqoGb06I4+UgBzYkOfYA9g54hecysZftevTk9s
oisleLpc2ZRNcf/zfpa6FkDQ5mUAAfKNMBL5H6bgAFZkOxate5dj/yG5NUjJhL7jxtO8B5rgG/XT
6ch9zW0O1Rd1rkY4y8bl1fNkmFQXDu5BRPO/2h9TZv5ARkPgOwsC5A322QcBNWuiyRlGv5bQyTwv
i8m3assECmG9f5iR6yThFiVYszkkh6tkDvVefYexXzIAcp9+XqhAFBjeZRjNUA9ekl8fBgdBES9h
6mnR9hRZ7Qk+phX9ldzr/pqdyukIseyofitZIxjZWskF8e+XYiztgPBuf5YUWbyRfg/aVfizCSIt
s2sW6M6BVbU3P9wBSk8WTZhlsG8Ymnw6w2I4BZez+/CRhztsf8tKgbnib15lM0eKVmNRlUK/1DdK
VYEPCJG8T2Txir6pRINogncn6XO2OySAs92y8a1vNW8r/HZ9/Cf84EAybP5WEGpmtn51PrRHDP9V
hcTLMVB4SbfO94GiXoh/zVOXR6m6JQhs6jwbT5opHhOxcrV/x4kRvDVnykTlNIehv5sSOZYBqZAR
zWPEyhY9z1h216CqMoJUAyCerv21maDDm0qasykK4+jjG+CfK5GCv6AYRyjLhB8nqIVj2/Bz32pj
4hwfUA9TjJngxvgjy8fJY5NCIlAcTcNPUfgoq/u8eAPKOCEQN3VIFk5IOq/RFE0h2lNgZfGfory4
MnLWxVv65YnYlwy//6c/yBZp43h14azc9s5NvyfPTSmt9Q4RrnI7Ob6K7v/DrHo8IEeQ3S/mlQOP
U1spdgG+8zW1+lBP0lgMyijSAiZUZTZjO0NoLoH8zAZ60XFUfd97+ZRfSvukQMnmPLb8UGjeaH+s
zGsKLJih0KHTJUqIlFPthgm6XMaF9TO/Y6BKO2fYkaBDeCiN1X6GacYRdxebHIInSeH7aRmScgZj
RZ5HorMsXSG+D2fYFKHTt5we1Rk4CDXvleSqM6RCWWOxdIlly6B2l0sLBhgcpyZH0V6MXkQ1LsWz
xxRvmpgQkYzthTFFW7nEyMfkXchAv0BvzWIJ9vwhqNUGHSChKa65t+lOrJ/0C3yX3dQYeQSIPZ9a
6s5gFeRmD+1AlDwnYMuhfyG7wZoGKgHVYO5K9+mmETKYntsEEWn8So5QBamzmmcCVwPEgiVv2qHI
bjcjpOQtIMyP+Zi0VT0WSHdn09AZUV4P2Mgl+oO/RAzBQApcnYxtgt09sa4I1+ZCalFhvv40WFI2
YlEu2Ewq89io8inBsGfbgun/EVuDus5/UJHu+ESE/nanI00R7RBOY/YN6z7gInTx/3Tk8HKA6RqE
gwny7WU1Ivjk8vXRVBy3TYG+fFu/ugJDnaf+IF4sQYFAWtTj17bD0bDBLZlMONw1XDsgUBT06LFH
fBwT6y+HsJxzqdFtC9DX4yPjL2Yb4ubK+TbYp6wrBV9EF5+TWwnLMfRDpWaIIq3Bsb2EVBdy8rl4
WXqxfbZzKT4DJmJU1vzLskwWkC4wBxFS3jthrJIJxqC75aDevyuQ+0PrynflEoNjzI9Ow5lgsnF1
CN6eRWHcR3d0qkL/cmhDreaTZZbZpfdqvskOEQ6TSIco2rYWtMQbpk9R+qccWPbvdpk5e0WoQyJJ
Iml0c2WeR7ROVSuNEpCsfcevxZcyAH+XphppmzHmfTsrBOMLWeEvwW1/8+wbp8LScfVETmxoIHLU
lfXixNfSGjMVvv3OLBk/xw8bmIeB27/LqRE43eXpZaUl/xUJ91nm9OgF1iQEqJxSBkuIiMc4h768
41nmo2VAJKuA7eykIQ0833x1buDtYxIz7pwuyrKf8Gvst0hp+2t0uFQq2hPoxNdZDvNwg6OEGygU
vVZNLLbq3WdxagOL1NPXpXVipknuXNO2M0Y+V0BKF6ts1UExgnTNuBA2mieBo5sr3sy9lrP+Vneq
KoKpIguFzOeGVui8Gj7dL7+HipqgqLf1oG5sZ3p/yZ6plhlqc242Ul3yksJx9vtYG6nWO4wEgZeU
rB6uGAbgGixF1adwUaciQz7uDreCW+8jHzN3b2OPYv4W4ZJ1a4bCXgCZiUqJsQ0zF7y6+Gyl9uda
wv1neVYZDbR72aYDeIA/HWEZg/Pie3hSd22xqvi04XOG6gh1Bccy5NSOcNOBWKJAjBCIxzxciDTY
B1SmhtuWDnCo26qBQyrWbf7FPvswBZZFPcaHSLmO4cB9adm/3ASUv8bqtKntQCNCvpRkuTM0EdF5
QYc3HTFpmqTPGuQtEhB31GgH7TGawkZ2u2TP0zRH8Yf4IFJkA525hLoksSuTl8tlb+bi+KlmJ4um
xgKYbc4iOKA3ZmXn+n3Mw4gzVNwE6WrAZnYh4fLc/ncpBIFobqUIh0cTvfw1jcyNVaIZPgYWZz2j
XjLgzfXuvQBeoM1nfh7bfCQqQInGgtxEbC9ikRI4O60bHOXElF/cn7z7y1toCfjmcC05isNPh5/q
4H8FJaYaUOtfa9M1/M2sryO+dr2kvn6FhR5RGALUXyoTeWskKRYwMisjOh45vvLxqUvOUQR1WZOp
MgIR4u25vUPbbZTALP0g/08Z8VicYxzanTbtpxHiwaZaJQVddJeuCxRk8/iWbmEtnYMisnWtyPC+
fngvarSZZEI3lv16ztJFLwLcP9XfeQYBEX+Pc5cwJDOc/NvTXx+JIp4tfx0Z4CJ5Z02PW4sZY1lh
eCirZDDd8xxxZKHjVcP4xOQtXcsdygpVWBv15PY2FYpxqY5psYSe3aURYQ1RVJBnX23P2ryqtZP0
t6knmbAG3y/k+cCLXdqIQQR06tYeOYeVkevFCdWnVxKIjAwLWnt/l2btZuh8tz/72o1/VdMATjSC
3CLut9bZ3Z22Zcx4unlxidSqQVmc6CyDWd94sUnzcUGblUI1HV/gCjGUvQs7BuMEBUoSlI0JCWXI
tnd6cGTAf6LoF4FZ9ugLryKuPYDbZ+2E3/3dwvXmnbbhHdOCzpqUEo+Kupn77fmL30pP2a7L0l93
9ejZqgRNJtZG+ctPqiHYP39musqa58Pfc5tKNLDdqYicv/r57ZrGPlNWrzXNMiuZCztLKEi9AmbP
WkYTH9wZPnMpAk9sPhMZAC+skle7aNjddTRKq2/UuFx3FwKJOOgJkxMYffZuL4T686rGjI7/qQQM
KIHvsb5jVYW1u3iJsRNO/Hv93bM1pwvHIwNMpY3aev0xgg3Rj0GnBwlYxWtFo6j8/zkiBDW4uqww
Mo+UzjeMXj5jCCHnPzCi2kX+bE/oULPGMhTzt4MQCHMVAJW11bePc2h5N7jcEqjUN3dZRMOMuoCA
Thv9v6y2AwdJaEPSjWZWvtg/5oE98c15eNAt8x8hHSp9KAt2kGN1bxHcgXDbTg0tvgfe15lnQ0qm
YO9BuI/YQyZJU4Vxm4gC2+SfDSrt0ps2+x3UAFNcydjofrr78/0zXbUnG3vMK84b72d7YInC6A9A
ixikHnMjAHl4HcEorypZ+8Q+Lw89cfPoz87b3pOQLDiIBmoNbA4TdMyF5xpJB2f1UplrhJsYqijm
HF9BrL31gPEflyjDhLSfC473EaD2LpDwlmBQHQCCIotl9SfwN954RI4EKXf7gNsq3q926YwnO+Cs
dMJmeeC5Iq5/VLO7Uzxg2xA2vMzKAKWJhXtZQqx1Ig3sb4q6X38Co/cddwQY+D8DPzN/cIu9HPEA
FW4pFs8e2fxxXIJCk9cAIn/YJCJI8IhEq+oydsh8eBP6o2c8fzUvjfPCtyyGQpQA82jXOkOf+M5Z
D7JnCudGPaqxYv4tCQmIxOfx0xX+EMZKu7tpFm5ERYI/C9Oq50LT+2C4PIW8OFoCrM18h6x4Flg7
ftHi6iiPHLrlNwb25gw10DNYdEi01jgP36rViFDEeJuPYiwEu7BE7kgMJ67EV9V91/i5k0PnYBIm
oyEWrVHWkPpmou5l6qmZHchTUCyJfO0G8c/2AFeNEx6Z0aNXieCMl3teak4LDKR30m1Gl6QYW1EW
EZZXiSUBs8dwavLr+Pnmjr0p91ZjbyQDEITBbJi82+m5LirUfOTmtAt91fHCePJWH9h428ynG6b2
fJWhGIHtTeZNuG6aXqFl0VC+lojyIyFK5qczCF/4tsjQ55eKt7+Ex7B4D+1MKFMmYv/O3d/71IsH
Uuqxyx79EKKhSCx/GIPsaBhsNoRVkkOUtOS3CZxBtMbScLpzHtpIx4ZN98nju0qrhUNCfgQ+QFRU
z80aqkNNMs7S/bad98jElB5Xs/KAWQNvEqZfipIcVfbPfneRr6ImkDMtkZnaZUdIRJMcEb6N4zWY
5U7OMALWnkB6l58D289dNGbPhRNhf7yuiChgQoB29zZDd4LDOfDwShwK+MVtLko2Hl2Cdt9DLV/9
Mo9kONDZyzD+83+ZFv3HKcBrchEJD0kFBornFvbHHpJF2yoT7UIS5ey4CFK/Le2UDgHNyxd7BDRs
BlPoa70+mQKOesSy9dpegXO70E5i8FS2+meODLzZaIs9hYNTI0lSggnK0B5xl3xC+qI0CimeXIyK
e/ZwBIgJupHV3oVdcWw01BdMNcsaLhurVqwbQ+yiv8DM6tuSmAsu2j/lLQwlHp9PYy9PRhloN670
oEiAj3FjWsmdtMJ9j6IyVyd6RcqGVGTHK7HxqLWTzZ8QiUcNFNOORUuhcuFV1BPKCfurjXv6SwKh
IImSpY8d42PT9tSrUecofI8OzoKQgj2KgkcqAscgx5dB613CI3Hn9TCa2QXU9wqpEK6zLliOVZxC
Ao6SLymGncRhzjXWQQgiOHtWThl8tidkNzTZ2YFq0elxsgozy9rssrnavwyo5LlzeHENCDxchTiw
bHDRr6izH0W1JnCcB48iEAbgLVWQJZQ4ANWPy/LLJX2I2wQO+6Q+8HIOKOHjzwgUtH/B+8enoFNn
c7193q5+RuuUh/HH6yZiaTWAQVL2wkj7L8yuvmJuMzTyQ/EfwJVg2BYKfUJJbWahAahLUr+AL2Vg
F9oWVHJFp/TJ6Khtrs6w4Zlziwec4OObOuL2Y87/nwNGA9qtpFiAMdTvUd4ckkhli/GXgF3bT9uE
o/iqKeSkR46FbPTF2TGNlWLxyQ8p7aX0XHBwYcWMcrwuUiemoOQfUgwgyNaSWfHMU6NhmQoEc4HD
jJ7ZOVkzxkJMB8WabyWF7XGP7QyzOJX9c6gGXbYGA6/ynW6JYXv3c+RAZloGozqHlsuo37S04a81
61ofgCqu1WpkQmtaOG8IMyn9jJGV8UultvUlEQ/UE7twuQRH7a4eLXgOrH7GpZwNmkEwacszpfMb
5dz3JcGJsXuE78QnHOa0awd3Yvax9rzDLzRuRCcLoUnIaO/0rcZidhOScZX2yuOcmYxIrWPJb3Bd
txSYoLxkiXeocfQ5CwzgizDTGT1MSEuw0xwIecsV9k8uo2DlXTlrMjUkuPFF6fiuquiOSGUPvGf7
Ck27Ccvo4S+bX+DkaBUQStgLfXxoJ0wOKpF1c3QU+KjcOSvGsrE/iS/YSmf7OiUKkfDxq0yF9Cow
umU1JGONFyUjqIM3Tea9YXflbPIcHuJf93TV4o51pIrujk/HXZEaf4KVEi6OwAs4EMud5X3hbBTl
kds0dzk/rRO2yl/Ko3YpWxq4GxTbz/hd5KRtpOyu2xHq5FL2Fy4065/12SRAmcVdtxcEHtMX2W96
zyHq3yQSyZ8dE7ZuPMZIg6Q3Nxz701uSV37jNA6cb+HVqj4gmtnxJih+BcwH7ZxKNNK3Ndog3PLO
CZfcCO231dVr/1WJuRZUJOOaTTWZOT7rFUMf92peO2dcOH5AlcZaSsTwaGI7k7VuUUo1uwvpO1eo
zcBU6WlBWvjdEO28Ood0v2izQd78339S79RPed++TPv6lpAQ8Fvw9UCquGh4ueklPPNN6Bu5LMLd
3gmjAnDLT8LxaQki3gx8KNakAcT/dTAJvMpdXSK+7wmJU4+bI0ERMdlLLgh4KBywT2BlI2UP0vSF
nLXJfoOzlpZ0bJym5qJmVfoT9CneocMCyn1Ow+/JjLz0eFeSh8TwWRAtyxfSasjwPJWlJCaWKY53
jpylUMpbxB31pbB1YsZAUcg5M6PPRLdFt68RfEkOWqzAx/ta0GcNrof4XLM/lhzJrVDoNyFFR7wY
LwjYd6sEUrFIozeVNs2YSpsYw40LqyxQmzgfJitO5VzqA0HAeQOZbmT2x654mPonWAxtJyCWirzi
3CwAwSCHINFVAwGGboGxJKERAcXXq0uVWeY3iV5Y6rkgTAF7+b26Oj+wAj0P2lTTiKMRpEFzJsqq
QOA7uV0t8J9rWeehLBsOEef89gYxDLCS2IBEghT9catNU/4H+awWFG5BL7n49Xx/R/U/iPq9wy1R
5pYUXUf/OfVCyJP1YnB7FzBSR/oVLHSyppRJCEci9CjEJRSxcy257Zo9mCtfJV1zR5q6PPN5Q/wW
Nx6gkaTS8LJt9aC5PXXA7YAMj6IYVmYSFe3WEDbMwhRudjfsiBGK+7deAUcp9V5ZNX6GDiP1LMDq
ri5XTWgd3xMg/rxBM7J722AIYVydXEhVaYz4B1ZF0J7nTkAXNaZoA+CtK66NcgYWOfuoTo5eCSuv
Nn2yWWJQDUlIBxatk2+c0ykut88tZ5KfKH9U2RVxcXOqM5ZVLVCoLK+xf0fYgwDR2tZr3RlKLtHQ
cNLhIm6PDK6Bi8XJHimZeTOC7sDkFempDyNiBgxeYud9TbpgPUBKCExqmr4a2FRp0oRFZgFUsmPe
z2AlebgTapSz8NZbK9URFcMHNeTJAzJuTn68gY5SB2dS3hKhBAXQjygA8I6GyoV7JGu3NFaL4Tcd
H77dbGf2X1xDbnJ2To8eg99BxDdiuMXMyP/nsgSYZaa/ZbF+vKETaFROqonWBB/0t0A2e80vvkyt
8tqY00CZnQNrxio8orYjFcoGDUNj7BzvwBdPssmRIwx1viNLCx4KaIYsgLBaMWWPl4wK7CH9BYOt
54FF0UPHTp393I22d57jt6ArNX+uYHdPojxd/LyuMW1/hCm/YJzVXZoXQa6fU1Zi6t2+xgfODpbS
cI9cA0F2OVOxsoZ+llpIWur+kcnW6tXm3pNnGxNnJzR8+tFg9HvS8V/LGfjoZm8st/opcwLJEzdS
xOVW48UIqjdrSnZDnlIIOdl7cuXQ4XwZ1VOwISRVPF5crUoYSwGEFW9Q9aR7cnn5TC8jWfS+kzAc
cGfvpjddlfSkrV3AmY7bimrBV4xD1vt+mqMwKOrTcOX6wTmXZkLkDCeUi1UBNFUJg5IVCxWIrdPU
911+GcZntgRE0KdxQPj0llXzCs4RDtWWPErzuiMjHVtRqFAbCJyBxJMr7/WjSTlnjFAILFMrq++0
ISastTQkxN939kfMiQFgI/s74zFP4Tp3ecklKQvIasjjix+z/hgUg2ZyX3eFN8YYGeVXpDBMHEu0
uB8UBCPjc2xmG/LfBJGPTd8ocU47KT2YIULu+zZaZvt0Wv3wZLBFtWqnwVbqNOJOL47kgf0Amyp1
JGuunSGkqQFQq0QatiCszIVFKqRnPvBQ4GyXz56AeS6arp4XxnUi19z/s6IzvbGATIQlaYScNGRz
iPTSDgilz1tjlw62zynLG52hGdtmTDFC5lM96oPidbFY+szqJjgaf/0edBOTkqJ4DMEsKS3vy4K9
aWy8OZ1u1kTsgeK+9HnDsFcRQjJRxMLIfC5xoAOra2pZ5ZnHEVpZNpEIYWGfagkDOvCCqXo171A0
ArqCuRdfInUx71ZRg/krcdihj/4Ujeq0e+C1RC3YKWN8W7UNme9nDMgotzcqgjzfKlHAEC56VR0S
3rOqBEkilZw3v+AOzpagQ3CDaHyKpbogys58GrvbZkex+yV86DYltGvTtcM9wAYhmDh+LpFh9H4u
czRxxF9xAujS0ODMVdqHkMgqy7XCRMIY63GW5hrZPa14WV8FZT0GtChxbE4BpiomjpxYiLCeZici
YPOAN996yMeIAO690zHTg27zIzFbLG4RdEnpOYkwlj25DZX/m6LoOBBro+C48YzVNNNjWWEIrjlc
yEtITgyZlSFyDWTLL8e8ylw7/2hZFntwL9nlX+9UxFIw8Eg76PHopY+rlxuN+fdl1xU3x9UDqI87
kYUW2xECjqISWM5jCH/XJZDnc24jL3LqUV92JyXsJXQo56bPKgLobAbPRBUEngPTqjF/9cO/N2GN
gXSVBPqupKKS1CjABoFHKa0a5fB/2CD1y8JfUCzYHYpc/BTaQ+QKncXkqlJ8WLDJkKL2tPFNwiCE
BhIalnVorZHellEmq0m+OvhguEyVHEp+Wdt1iP6FBu3xsAO7C/Sy4GEIE9wudICvE5BxSP7uSvJ1
LYR5/LCixk2UodukMvLQXbIcXI2BOL+BfpSKMYOaJMXX0VVYVgeMA97Zc3RJhAp4CYSF8btEd5/G
8PBqcmWBF0i1/BVkLs1yT5hrapIB0rK5+hQVSym+ePd84K+ReIaCfYB3LZ/bYhyViQyia0igPar4
PPgLfSuKKFj9wAr3C6rIbdfpISFAenMtvkpjHYeh1Zqj7X3sq6VnPC7ZRhaf3pnvCowxDiDAbbpf
Hg/TrubCY00HVvJL8L6JPfoKd2Bh9RVfW5/GYY6JsCZkHu1F/Qs3n5oudV1nX568769phOQXuSh7
Z/HVAzEqTRj505KxUPSCcdj2ZzZDt+GspaZUrminPuWp2nvHvjNoSdp/zDZtJB0oN9uhCSXELncs
ynf9CefBdnEd8KA/eGSSGRD7tQFM7Y0qNoqIapOB7rCEMXzxBI0hgbtWUPJ7LVXunpzyQsn3gWlE
cQu/b67J0+ue3dRIP5psW+eKcd2hlN+j+6mM0cJBPPdrFm9OmMXCvwyMUhXpNyvG/JFKw3ZyzhNj
2hals8ydqLUSU9YIM1abSe7yTLf8N7T89HnxZm/I9oW5xSd/u7yoU6P+dunNVo9MiTmGg7TM/u3N
svmnuM4ae1FBs7iqEki7z+Oq4MdvCYzqQr42zG6hlEXppDfmOW/Odrp5s78bL9ZgFn0HVe0GMEWy
RqTjabKaNbXzHUjXd3tTMwUijCBhyhIjeXMCdLP55ls16gRqGd8IJida0gVhuI24yJPYr4nKvf4A
Gj3ixjHgMiG7/0uTp89SKeAQgwYsO2cZmX+LejaBrvI4CC8N2wWz4aJxiYQOEWbtRmYgDAwyOA6U
eresINSrAphgg2bWeUCf89KpH7H7ioxxuPDA8LiH4WGtZR4akw81bVCOIZsZVP5a8lnxGc+asgsh
LtZpxTTfZGG+22+u
`pragma protect end_protected
