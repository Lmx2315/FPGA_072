// (C) 2001-2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
jpDNjrUJIzE8NMuAAJpSa0d1rgnDKMcw0lSepNmv35sSH5Nnfnft5wNLDSm3pnn6DTumqypPZAnf
KlOJPv7TqHfWlsBIw8ZEkddwAhae68EaxcfSGSxtMBsDs65B0rzhiauo1WzAaYEBy6CyZL3IxO4C
WXaKZRMo6ItS0N5/l4PrPb0OdSeb7gQIXdqcN9WFTjz39hVd60FrHlJQAJ06JdJIR5Y5YVSj2Q+t
79UEixns0EOuGmyMbPH+LQctDX0ugcf/NVB4IU71vFEs+kXanBfvpQ0DnpqKS5Bqg5RZmdLkYSo9
k/QNjxJm3ipY0TTsko/UlvXFkz1kVykhgyW/WQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 22832)
RvqvhmbifG187cJTiZXuLXKYkstDoOGUvWuoQvmhVIPgjEwV8411+5JtbCNuAM/CJz/42mjPGeVq
8AiazNyz5D5ZLFMDurSpVvQ+NEj2ACJsPDZ8ZrOUHWvxYm6nlCoMPpYkNJ7+BGAdCUf0pWpWMS89
YlhckrXhvjbI50v6JAR2LL5FUNENOaYk/x8EMo/2BVvtYyxGBQgcqKX0oH/YjMAZ7ZIYBErmx3Jh
MYkjrfT1qrf9JY2tg2pkZ1qIZheqH2eFmJ6MxqbQQ7wZ2M/ljEdA52aw0ACGrUuUUaPowJpkhoBy
atRQ/ggeGZUXdhnDhGsAWvp4a/Ls8IRKRf/Bw1SEZlfoo0g/Go4dGdubIWSf21g8+jlwkU62VxV1
wLesDwVf1n8wuUswSQYS6lKpgZl2tIGIxowpYLJNMS3UKUJzttEu5ErqPJd2Co5ufFO0WYvqmSx6
u6u4zu1Nn8E6jVJEtURXlRGltUI1oMtxujNMQUiwd6S2vGJMv33dIgZLFMrHkI3SgUtihduBLnGO
FJ4GTVnR93RfyrFY1k2HQXi7m0md7L1IaN5XFjbLmR1nxoUiFl1kAlEvdUhARaEeJJBvYLfJQZ90
Cp8MtGhloMGGE30gYck+7wTvcsjt+vQuyqQhkgZaLkiDADhxbwD2CVQC/+HWJnW9bgJGmVRysfy8
QqC4B1laF5Nniu/V2OTTtyz3TpUm4ii2kc20RbvSfcwkCqT2wAgSkgTWszdbXZ2PNQZU5KnIqV29
bSwVAUbDW8UX+PBsoVqF9bc0z6e9Bo079IdxJeZXq97OkV7hTmNnYkFAW5XEyyPPwCq0T0iWU3sC
ZjQtD5d9SzlOE0E+jP8zUurmrV7mqsqPX//QNuSMgJPu09gScRdzdV0++ejTepGRf76xvwip3KjM
FMIiA0jsz2Vjjvik2JQ7sFnUKQ87KgR+uNqaD6E7we/dfcp2E/w2/qQ/H8xRMqb8rwd3dsYRygi6
D9tKE0svXy6hO/af4S0rs6UH9fSyx5qKQtQupei4Dkwo6YHyuh9K5FRpv/SxLbCUD3WdVNwcmxNQ
7OFu8eDHSAM0kLmiPNRLZyrpCh2+3VI/F2gsK450KcZH9PEnVUUbRSqIIg7BP+hxy4ATlhiBf4dn
gKb4yFbcPPDZdDsRNT7uoYnyiXif5pCAxpwh5JjCYCZ0y6Jej5t0RmxLcpSq6wy0G14q+dkj3SS0
TM15AJSivVjl7XbPd6FomWPWE0fghUkWM8tuV9eOEokZQOUWgvFES4sESUi5zZeRLr01ySc2rQY7
STd5TpnocT2vYR3AwqZ6tdlw4UN73La0NhmCktAZpKOyZ187DhPn+nMw7t8cN6CeL1zTjBcm9kn/
5JzNwZAamARA7LbpVoPIm+LhcbF/wSZP+GAGAysXpApSMJyKcACxinLzGxGLE4y7cWgUaNp5cWJz
OOMxbD2jzX4HUMzSk68vmG5hzLGSgrxGtEgovIIHml6pWmtVLHB2XOM+/lOuvswDeepsl++x3v2O
ZOYOk4Ku/1TX+7BWxV9QsdWtZKN2X4QAWYAusDyMVZfy+blpo7C0cuj5pMc/HVqt6ikTV696YdZd
cp1NL1Ga3+4JC65jTFrAjH+XYM+eqCXwa2aofoTBm8JsC+F4Uv7vehyJE0UCsH8cc33rpo8KVW2V
ChGUSLe1mnWAIsWoaWtZFTXghHZj2v5AAKgP+AqaEiYMC2Fn9HcXoWIHA0hLyMDJxDfYCu2NkTs2
73ijwW4bVYsJ/lCDBubQbW5pyVpm2JaUq/cDJTk2M9cNV52Sd6qe4pZ/0ekFl3fcgpo/vtxuTC9i
KmwUCE8L8vaBkxeijolYkcS42ZCgoRIxktJhvNbUPSUp9Qh7IJakL6FwF4FVYaWH/7B0IG8sy/Px
Nkte2eR6LbiGVjwfr/Bu4rOJNNeQfCjltoa+IbhSwHLNLCftzBIEd24m1Fz6biY66DG+oSQDnroO
RAEsJm0UW0Pp+7/0as3nzQJOPUhhj4w7Vll2p4ghwovtRLzFZ+ZUY2H3oEH/nIDeQITwNrDhE9rx
mhvX6BdAW2uVWhHIWU5tlfHa0p+gsHXxsjKXPRX2RiryEQtPhoHa2pC/WipU1Ck2RWNbYc5ADyo3
NenGjJ3DW8jrWJGHwWxuoTR/f1Zplp0bVTakRgZzVbKWUSIrfSWKpSAUa+KpRnOZ5QvoRj5dXAE+
hAj6AX+dNHKdIFs5Mxhbuk2lZ0faE+H4g2mG7LOhmT2yUX4B681uDre8+brgTPdgHXrlPSmN4YeT
fJMhXpoT0ATow7UqtafjRl62SyN8QAF5R4T5CVeNKMjWvc/t7yvTWhGC/4rMnJILoSDWXWPqyy+6
KTr6hCbGS1d+VBnE5lh2OXGQltzbxyAO8/DA1AIlgOPM3m5aOD6A3PURUCemMBpSoswF7sk1wuWV
MD2I6QVYSliLB/qvbTsEEBY4e/E+Z4THFpVngxgXQGOe3UjhGGM++vlVjRRjQmgr2vwr3gzV2kI/
N5kqbCjeJ2XPZKahfJKeDM54bn3J+klHn1c7nmL4993x+8Js5rJolfNYlv4qe0dpO8PlpIuR25lE
SCS5nsrn7qwAzeskqKxcIUIs6aayE1cR8RIL5gASl8KGla3aXE/WQdO/hKdgkztu2hXov0f4raKQ
oYmvkfhRlitRhiTjDEqNMjnKbNs89yfxCduzHE7YRDLK//keNxPQlxwvGHj1clmI23q0o52nBszP
B04WF4JspUtnqc3W70G6AOZXp/A36QxDd9xqkgtUe6VvUNANTUDuwTa9GPEN+DRekONhiXiP1AWj
A4GYJvxAj5d7/moRbHrAuy0V4NfqnHgRSxu5ZjNBQZuDQ+5kcY+3WGzHi+zDMFgtA4tnBSDIgxMA
IqMjirVElRGnx9gbl1/rOzbNJBtjQUcgtmUgUghJcSJNeiXDlVqJJw8y3DmddnF7LR7tj3nf3zzS
xk5aHMp4m7o54b4ZszGPJJdt2NWpUkFNiCBgYddYrPRNHKbl74OvR2RwCGuKpUfPleq+7+KMKQcq
QK8oUPRi5Va023oq0WNCpoBQ5sj7mqa5pZV6tIVXuHKELrvQooR+rZtzY/LWjF8Y9aquUE90xH1f
uSCvePBGuztJlnHtTMOtzQCn+WtzkEDdgZys93zntoIaAaFHsH9xiFv4rvwUnojIlbTrS5Bh46rJ
AVjbswlPth80y4a/zt2ILWKYEncQzkITsGxuev3G0So+CyOuFsRhr8vVkQF/7Uh+fiWe9JQLruXT
18onKxE+bBARTjP2DeUWmri2Fj0HQxGkhpUdLQhk2c8irVplj725SJwjGLhUiCLHZqzDDlCJ7DAC
7XRFjIHJVPBbMcllkE2VptpSwMRletqLItekDeviQD4LEWJ5RRC4wqwnskPS3dTqFdn+8X+zQiRg
3ahwaeSMB0k23837cTk09vvrdn1ilqGktdDXXf80eLoP+R6HzuKDUQtzOldLUuikgn01PtFDvNOw
ae+bVULuHrwCpkd16juL5LIrxZUBfzXun/R4tA+Vr9WfLUQmR6cSFr/htbOMzMcc/CkeAIDYyzb+
PhtvJZlzqzebbmWcOmUoWwgf5SwgMILXbrHU8ZRyDPBjB+w2szLNtWeFL04BsD4rYoB4gz/v1VSe
2NHF+AhRd1cuoEwjblzf7Xv7aDnRK/kktOGwhP7ZpZ9VDaPLmuSMmvkHkaZDFPFrSt0InFLbpFRl
EB0iYZwZEbORErOb3QxOryFibP90t7ebJp+IL4Ie3dPl6695PrqWUhZo4WfM2+OZtQW+rLyh+H/e
bKLnKPIWfGFQYHbYmAmdFj3wq+UzIW75rorsTQETxlpj9/GosZXh3I0mCc8bPSrf3KvE+4JTHGYu
+8naut9snel3Xk0+tRf/AMuLfqUE2JxN4xogoVRUE5ofCxPzRMi+76yxvVTKUVhJTkIGFF7tLWuW
jACzeXLHP3uv+3vFfg2we4nheHrB9mBEI0/4Yp+LY0FtSei4EfjJnZTypdSIyrY8RufeUQyIv+ND
EvWXt7K6tXwpDI0N9Ueld2cCuY8y8vZb3QazCW8uSTx15zDzcbTgnAZk0reUtlKCYemApUfhBuCk
r/etY8crG7R4xqGKaLpREs3EMnyzjMyhrWxW6i7ygO/kd52aLjc4qKZjy6l3mECwEvuTrAROzOje
nNaWfLVXgwZH6JamA7cYCOC8UPP8zrznwPvuMLuBpHAZ9fEb9X4GN0YpTI+5sPPfzuHK9kpx3I4l
1zaCF9sI0L3mbflCNQJfjzxBUANQfQJp1yBbuwUceZIIHs8ni1ZF44YdBl1rHKTC7GweoiEsUDsj
Y7Fcc6O3D2buh2/FDuYakWQHznhf+HPcvtTp/NwWU/COag5vS4OhAJIJrenjx1Q09w4iimtfDgcR
67VHcIiv+HdfrW+9HCHc82l2awMF9dTcgHlQFLYUGbGt67ZvGA5fOn15vPTfts8hVPfKIqmLtpJ/
6c2m+6HmZgnv48NHzG0Pzf+WmUbDJ1KrqKoWmUM0r+l+tasFkVgKEzht5WdLBeWRlZUZP1XfufyD
awpilua914jPEdXO0iH9wDaHrHg6X2Nwv3+gEd/EmB5DaH7G4aNcFWqFPLQM+YZxWpQsuRjiOzRp
yoOpmKIdfMj5Htcz5aGpSBa8sB9JySTRrSlXPkpKmtI6cKkZwf8Gh2YpIKTusgRuwU2Oz4RegbBL
BVYb1tToE/TgaT/KuQ0cDlXQta65Gtk8YsTUCscCuGWhr1OpGLYln2DtgwwHwiklQsdXv3S7e2/j
JaHSkR1+Lr352QVFrpvNmj9bjSVO481V0iGx6MBqmxQrfX8Og2kKYy2QiqY1Hlwex6UgB/E/pwL7
7bVpC6ISzOxCUqxkDpgxlqxqmImc2S4S04MgsoOpfYcBWwK7kgFJzusBqcZLtuoADwU+Ye68ZNhk
WXWr2xqPtN7/N/UJG/gR+zqFfAKoq+HuxsaBZb/TdR0QdvZ4X3HcefHBIfSG7kAeHt8DT+NL9L93
ks8XQEgp+fQXKnCUtLDl9fwmiJ05sFwbkGaQ54xJAhxPZdzVPx85XqCsnOI37TmzF4mViXHvw7GX
WOrU4dBHRHG3TnKqU9/knh/moVvtvYR2ML9uoP3+IWKwak8yGq+mH4xnPzBvzxYRrnQpdLKYNrns
QVk1mZkCZKhr5w2iOJ2wo6PsgkX2WGSQjkEtSrYcI+rHXKtZZjbyUEFjE+sJpRV0ZfpOIbBIQ6iB
lS1GAW6eSN8yNKedGc63sbaoq1EaSfOHZE52giDYN1a6rFHQhQha5wkZsu6O5M/jRWU1T5QzkkR3
QkeOWSWN+O2SQSnrdJ7dYDyuT1J2UuZUpWkBAtK9MNbG/i16X5FXxxz6LooOT9wNgonhAnQcf6S9
Lim22/uE8foDiIwYt2zdjtTaBF0ZO7leTXZebL6W7PPhCInH41eTdOoSXX+SDZwrWVazeKJClObu
lkfC0UArS5gk1+Yrx/DXdsDLbjRWttFW1JHV+CZPO0rEWbwoz3t6CUVXeBmVjToK50ns9qrBJRM3
0iarQzsdCGWBJyrcKs6Xkjis1TqKiRT7UIKkNbgdmu7hg79jgr6FS9C5hTGcYSf8x/g0KDkw4hcB
bgiXdR7NdQCU2yjA6TVJH8PXeItq5LLjlhFAgTDyDLg8kwg3V71BV/hN8PuwUSYfTurekmgjHBwJ
PcwZbQV9K5aB8hLMzcqf5XS44aFG22hJX3k3WzhCvjGGyKehBAYD+3gYCdZbYzDmxcGrsFoO7xIb
FGEIKx48J/uMqnhInhJ/27DpwpZ5W2HKmgugMl/gf65y40rwKLJo57hn8ma7WZIQxmpc2RFMhbLa
kwKs8rD4EqOVaCo1VebO2Q+lYHiBLLmWHqBxpOvOeDc1x9lewDbEocynXvrMwYozoKfLgbZfaokD
7J1sA/hBiJd1qL5QxhCFVpoDFb7u9q+ubOdm/Ww4e/VIyhXJZByjCQDLbPvfr3l6ALVopNDbBXWx
5ZnSgVtJht1SUUNREceE5SMzX4QPAkcRzA1ObPuS4f40S+YtSAxLEN8KbL1eMKtjH40h1CGtm8po
qhTJlo7XSdCtkPOSSNL1gXxyyd8Dx3jid+IYNhPwaLYylTlwssMMGPSRyIDSyQ5q/5w7fy07ZaD0
WguPXvYKUHw3GXwLSCrTz9gQ1H2rW9eEMjZrV8K1TpJT2gAjuN1wsNlyqJEYHTbCr8/zM0UyosUS
oWG7LFuC97fGsAbOpKauGWVmaX2ar/x7FAaX46LAndnGX5gT3Ewe1C0oeLqHTrxlXDsUfMg+5OYO
PwEd4Bjj3XkyW/ob5ii6MgbvRi7BFOcx5GAt3bdXz59YYmmyngmlx/h530cyApKuabYxc0QOmwEk
n7dH0LSaFXNk4p9oHLNUHjlGKf0tb/jl8YGxkMcWPH7Fqx25FHUhJHNkKqe1kAROdZ5Q4ea50mpa
Yo9tifFEWcQBa7hyWdh7A0wEO6C56nTq3KNooCGYqf4T6/3TS8TGHkmnVO3kKHLy4LbeqcimfuKq
ml1J2rUj3Bu2KqvfPfVmYhx03PH3lfKNU9ZEadDCBZvh0l7Pkz2J3fN4LxBZgPOmIiU4+chIqt7e
X/Sc4Y4nNTinx2ZWFMJI+7+trWp932ahLbxG+eFY03+3P0WwseWpQq4jap6reT9bOVdYZWtyz6OO
kmiIfQ0AXW8Y185KHnwiG9OQ5eptLGCDZZizPEjhEsuQI24Jx/p4PG3csvd8JnlfNDODCJECslEX
CIyoFdPUxJQC1EhAytuePGWgAS7o2iwNEvxuNmj2sSSszQGNZSwZu3VxodLb1QDMQdLZsHJMhzjT
ZqdBthWcA7Aqk1W/ZVKdTdaFtzzyEz1+ihiITkYZyA5elR87TVREZUqrNfouF7r0B1bBtgbBKh6F
dY62LZMrOubA1LrgQzzWCQ+luNSfU4es+G1/MHM3esCuw4QLg7f/jN3gdks9ARBeYt0hyn7NAtSj
nmV7+OmGfCJHfHJ/7THPDXRiRBcEC8AjeFHNCGPL/n+rSCD6Zn3OyJGh8lR8MQaINGO3JuZGhYAf
Y1BBLSnm3UAnV3PEiaQFZBjN7nArhUvb2adGn7hNuSfibr3unBf+ihKuz9dZ+uyah1oFeVXnh6sN
4taQ4RjIIp9Y457MMKxkycEC3tW4T5HQCNWzvWrjQWoYE9q2yKaSmA5i78aDbjGA1hL0mRykGwyj
yUpKMYR/MssTyDA1yEz10M6I0A0YXxPQvlKA06L0qQ5AzBPOYagVSLFlQdQtE4ORyEegNPp0EJhw
2WA+B5q/R5W+tCrTMb7SzSm932u3H9ulKkFz7eRyiBoPFSlAO/0O38ZqxVPHu0qmKScYJKA1vrvE
61Wrt/DMIZAWKVD4HQME+K/vVNFsrHAturOeKddbqCFzC0LnshB+Zj1XbfsmIrV1UyxAYUHMh9sl
XlZNBmyTNwKCK7WEYkMFIUYIPQNykG8GiIAJXDXktSHNZ3RHI4tBQATe8b6/JNb9RZfhFYgcAxJk
+IGqZjzyIas5DdG2WvLGMyQ/NcNbz7RUJSqmRBIHdQSsBKfx9H5L2+l0spmtFnFkv+02tvgRpCEb
av62TNMACXlJxj5n0W4Ec7phnTk/+HG7EAToNR6FDlZXV+WpgM/wBoIoIAp4yWLvHed3Am4tlGCV
sIpuuS5gC849ud3JI9M4u1f0K7rXP1A5uHvUTYSIi+W7EVww50TYeiaoT8egxeEp8YErP4ErNJEB
cEvAqq+UR6p1uFp7qMBBUZd2aj8e4IxQeijWS8cp36LKuC8gx7Qo5D46xy1t44hMCjpPyLkjMyoT
iAIBo3aNvJH/kGk/ggmVIhWX1DM11g6htNB+/ut2nmolJPbIYjcwCIHKnPOMOsDpQX4/n9QTbzbT
2vYu8mtZYGQJHl9V4vIPDKodG0ZzRYAMT3v5nrOJl+bfCMWgusXUFasn6ifcs2MpeZQFAr5tr4XI
6dFZjkO0Vi9IwsWciIt6PFp2hnGXqryOrtZz3cEb5H/ZughuSMkZ8STEGTRu3qD9LnY581gh6NJQ
Y36LDR4gECr/DprZGUwk30KiQxBeHVFAi8LAJb4JcZHH7RcUp96XDxgjkGHGHG3kQL8c9TLfapcO
+weMxOLcPgycnamlSPy685Z4PvJR5bEV9NX3h8KIvMfLyEZaVKabGpALHLID34TpETyOPI2SRq00
1Y6xw4BlRRRf6Kp3bXOt8UTQxf59m0U1b/ONz0RjQFLNRINYLmfyLHwrGsmIqWJZaklmT53SZunk
Vqba+BSmxKKL3bHMQT8iYAEr4/SrkYf8xD4PbIQPYqMlgcYemDjpa8bEgCcwQGzB4RxqPCFnUwjb
LGMUqsBgv27JzeBzYonGAO4jdM1X3qDtiCccj0eIxz6hABuaZup6VFHqPsu/8WzJX3/naXDzuqEb
snKMrxcR07NdDlcqWKGRhpxhJjf67ZWT5LlhKiCps+T/gXKA7goHoiIvINcLt9IbF4o9jzlWUq1W
wSXcdEZl7qAcJwdnGu6tvEI0CsgD4M+qhaDQ3JR4ClQt0geW+CvmKBfbTHS9htAUWo/zJRlXq3tM
TRE4/8wJAvbCZZ8H8ifcoxhuGd/8VR8GXqUYz4KWn8+Akl44pn18YvD/rMFixOyDX0L0NEpH4rWf
2UkYp4KMKAVv3br/ij5h5sPafzgg/hC6XZ2Fe2s/QNzZuZeWHYlUX3X7IzghzlmTTH9iDLsWGy9i
xGHDcigEEAK86NZ6z6k1nPEsA+Caf06mbeIv7nrFFmf9MqXd4uwBgx0X9yqDNcPYGT5xgWk823XA
Uw9284Rq5gpXpXkMA3sXmNW8QRIvaAqenLC3XtJ7fSSKTGjVzgz2cFs7iTKDLjkGd2ve5tARbCKs
JYLimEPuRIlKJQEgvDHq7NWGarW7Ci74+W2udXH61LEvLEScMyAeXhqSq1h++K3CJ4POWYFcWaJN
LghG3Grep8K14hYmTpbQ/IRYq+CZvW+u8HAB93IRTnx6MgUAggOZx9LSaSq07qEQl5A6f5PjaQ6I
eEqEU8iActdC9S+ebnuToRVV8T9q90mO7s56nBr/9zwMpFatZdoLRjtPU8JMRLmW4QdkZ3x5iGJz
TzXw4seewCmEW95k1SDDgs429K/kW2EpKoNtFLH+ZWwQrhBkLukk3g90wvPOu49nlKr4NFvRGKJU
02Jum/4nWVXY7nDaAuJsZRoIf90qkehtHbs0/k/DgFr3isYfav3JO94fG3E+GWhB60H9TiOXKJy4
luCvQ5hZ6ieincueMdWpKfgUrTShMeE/3hwRrfOrehmyBcjcqkz/L/eO2BXDxpWqO4S9HYTBCQP5
HtXqS1U+hmOpsvUicSTAPmJTee9en8svOCHTwF4HG1IaeLNcgkoulMRRuUGTEktZGjiPwsQuaXq6
T4WTEGtVe1TFs+LCK4VSYo7xG0CbRuRKip6YwQeAWAgkdqdh7zwqEbCX9NcOC1ebEXpoVBCTIEZB
Id6iOhE7d877szjtp4UJvkkLGszZpSdNQRr70Yvbn1qqBbdwzwG96NUtu/qR2cTCDCBMdHoUpSv/
cpSGsBayXWmzrsP6uzWRt+y1Q0DTZH/XODVM6HeLAvujWi3p3zHkxJuUPQJ0U9h2toO7uxFmIg1G
F1Cvs7TpaWnOg0fzr1RkFTiPCkykiPj5zTpVBTFTKDgLr2Yw4+4clOohCQAQDdhps1u8+gbymFLp
ns3/UVgNVw8eg6TQadszkDPD0yl2D0TkzGE0W/JGliX53rihlu5vzl+tpoq+B5pgNYINk1abCs6x
XWn8u60TAiu6tJIH0zlhrzfaxO/k7RuBUYPEIy89OIj9f+42E3mSzg4cGo3j5/AsKl/u0sGZLZKx
ONgVSfNL2dVkji1I44nvk2U2GN3iWo3Wv5kykH91ry/hGRHFrBtykWJI4g0wkyhu/zB42SjyD7/T
ehbR2p2eNxQ1PPOPZY9AFf7cRVsNLFa6ZOTGJBAjITLs0+MSgg4JHnHLrkkyfzu/6+fhY6EiYNBI
WsTpc17qFBJJ6vbFoNP+p6wb14srglmhbBJAJb9A0l7uAtuZ68qUjiWJ1qFgLed+KiwAio6Yzg1k
JUpD+kyCUkUdG32Bl8S1RU/maXmLPzuhWJMPt0HyjFkVg2oc4bFLpHUsnStzXya+botJtD53aG40
wxiM2LtWgTiJ1VIOrA7roXgMUxh4L9sAooDkBATs8TGSzzVJTq2DenhuiVAsNEwlImSyd8TXji8E
SxhvG6D9bYKdtO6UUqacJnAl/UeKmM4T15MtVcd/oEXV1IxdT9Ys6TD3kEOvjvnvg4pBL/Q+J80/
MlVd2F/1Gy2cMUdMEJHhwnr8dIQHqSebsiwmO3FaUZOYueahOzL/gWrQ9GvHrKrJRVjwDpV1mo7I
yGD0cJlu3Hnr0DZoVEkL/WCu3KCUJclhJVDpV8BmGiZPS8zmW/xLubFbbtIUl0UvtQxElPTkbocT
C6X/xN69RDZbHUEGEcsVum5Pp2grtutTbx6pSrbrFSeeqTMnSTXXm2NCRZ2Q8z3uhGyV1ihLe1gc
rIdITLjpcmspmmTNAklY6UrMEydhJ5QDAQLi7XYRcOm/d2PUncMtEzQ5MBsfw6q324bLpdVuvwXf
SBpYU3WlsUUqUYzkznWLuM2elnMFJuXEIb+9Xrrno5/CpnTcUSZe+MwM6HRqQshoGIyNQh+qseK7
vNRTi6PFy15jBi5vHh72bpFJvXrkwxgPHl8PVnDSHACa9FTwWebUDVbyHBjdWzDH9McZlpqCpMRb
tO1Z4Ao4FPAnCGL0MIE2lkuovvruhgoVIgvAXT7bVingYhsaSurKQdyN28/ye+DntWsDCR1vvghW
aRw0f6n98iVn9X4zhFBF5zvReSD3Z0/bztkcfZet9TWFQLG0IfNAKq4R+CajiKfVaakg56Ozn4rt
1oLJv8a2v7tDJ3un8NbmEqnCABoKAX9HftZ4Bom0vygF3Ps9j4/Rax//ZUt7IWBPmnP+sa7KaxF8
px90Dr9RSObhvjhHTbwxFoRro/OAKiXvV0jgpQWHN9RZMcsAZaN3eDbHC5YN9LRFBqQlnY/MeR+h
CIjegMa9tWi9z3sYF3EPhD72DM3O50eHDTKDIy4v4/YI0nObi8gUc0TQ4vlEy4SKUgwWKOP2Iucq
M9WwGEmaN1v2wPu3LG+zLgfjXVXmsZOOKeNt8hIxON92sWm7gQWAvC0ux2/EyINjYRxbE7/Cz9K1
nEQU+wisempl+wSXlz2vh9GeOwHRMfAWFhceL66+ht9chP9UpoxTf/KQdSpjcYTUfFoAVR8X3jsD
glvF55gCcCDww+nlqO9lPpbGKCpAyNkxc5H3qDyGSlWPAH/WzMOlPak79EQn/DjzL85phnA0JKD8
ra3MqDrFbgc1of0WSc8r4CotAjMUDL+xdHP9xzGHoVUdWjeAKeKGXigWZ1wTIRoiwSxkBPQAuJTS
yeyt4ODABXxAO5sExsr2sZtx70+6ogMRhRY4f6GeWECG0r6VyIVJkFZSxs/uvBULMNmqdT1f7fux
ZKKQ12jEGXB14CpaDlVYy+T68I8gdMn2SeFeyMUHMgAC0RKu7+s3A3FlRXNPkNYzbcSq7T1LwUei
J8ItftLjyWJJ1r6pXqjcxBGAUYbahtAofRepcOohgxw0Diq/yO10fh97QARIzsgS3JMRz4OgR6n/
2Mjjksov9KSgw/sPN85mLmtdZtAYkSpdDk+NVkOXfwCpiUQe2W5+7DnbCN0T+n5h1kLlOjYU0t4S
c3pgzWD1w/DxR+k29PvrZe8JTIJrL2hIOpn9t5Z/ubSeHEMIIeeok1SmoOV8FcVGWgqes9jv6jUi
cU8t+Qqj5E/Y3NnemyuNP3uYD/29iPoziC70mDUPLnP90qQqFNX/VkwTynIchZPNdupgvTbbM5qv
1DGjvvW57oo0ZdD2z3zHY5CNUw4+FuchiSHTe1NcPD1Da+aEIKJPclBHRAHYW8CsJEQaJlKwhph/
e2u85Yjc47Nteg5irwqWpd5DQyoFYWnj6wRMHbnqAdptmck+1KXIh5W3oHF82tvkYJkogU/+8xjN
4wrXh0etBxb6VYH4F5wkpUhLlB4BXtDgvQWqMbF4Yk8sW/OOd0G0i2/iECuKxFmkSXSDTicZb35G
pJt0/mmiEYCHBVTK6ndh3KBVQxo8CaVQ9TgTXO+CHGwlo00Xhb9kVsTzNzIrZ8amTelJzXWSAybL
TwMiTTXx8Zamxa4FHREjSk0u1XNPA8DY5j7jZGXq3HoGURSFTFm1MAuV3x0JWK5B1Ai7rhchMIz5
m3JHN8gj7uMUEUZl3UjCNXgqFUvxpvB9gda2T7NNWebAZNIvtzKNA3wGj2+WVj+KA9rSOSOkADaE
x8RHqEVkPjhkwOoE+15pqvKdMjpeHKZo0cfuWXQRy1uEMHfVOhPWr7M7uKkE48yy6+NrPG8GZQO4
wXZPlF7D+aXwll+gHN7cd/u55wFbW+7uaEnaL4k38ddJm02xtcYyU6tOmeyqCykd2Xn6lCZ8IFfl
iA/uuuWBZ66WNnzVG5/uRgLCf9hL6zSYjOWBRDIZUbaU35biH4sFCAN2UHcvgh5NuzmeNBu1nNK0
KzqZRd+bAvO000lrR/XodNyjtpaqnSnXO/ZvssLtsJlUBXi1xqi+GkaNVLW7qtFs6mdqF54CRTAc
3qoClOWjH3Tvu4WAKtYFArjHkE0k2oX8IJ+Nfwfc+B1S9pnZr0rvHjXeS2KmmoB9T8YY2EowmUft
iSC5cKFoLFWQt7EyYXWVrycQmgw3EIvXRJMVWaVAoQecoX6Uaa4E8IQiC8b1EeL9BkO2SglhIeks
bSgZLUpsyBM2mv9pdeaEVylL1cD7yoH+KadyYVLsoX23oKK9ZLHnmkAX8Z/PPu0dXyaeDhluneu8
pidL1R7QVELeq5mlAQVsg3j4FrWq59m/hnrvFOfZJ+URgHo79/ZdBNWlk5PJmSGs/iUw/0nyK3+3
R9gPAZbyjeYnmfdB8LOsqyn3g5CnP6wxdwArHOPXfmc/oKIqRSFQgEtbSyeUCt14f5Yb7fb0KRQK
sxxfqMpTsaV1zfinMU22WSXB5w4YYYCCx8Hh4hVqMZ/dbshbL/9/YAhkFGkIy4MokqOu0WMTlmsk
nRqGi3sCB14lv7FmjI5I4aACIUqqybZBXX2SwFrcHr4EBLh0msGRE7ngMMQFcq99OTDiAGi3kNRH
9aI0yQQ+WjBgG7knln/EYAmgty9YbPiWOYynUB2FNuBt6COJfFMablj33QWfXE9on0f7tmC4H0Zs
irmDFf+N2BcMny4PiydOzxJ2SJsu2QGqGjJHL58JmHa3bKKlAha6yysJKLF+mzhy2ALkB7oXNJxI
enb/QneOQwPqBU0A0izQV1S0X8F+CkOT99F9ARjFVBJM3c2TVoFiQUYtu+iViddyBbumWSwfXycC
XQX/TR2CahyzkPvLcW01ml74jgVhCxiWS2q9YPvB4FSWUamFVFWuD78+vl5rPG2XjWjNjDBewb87
zsKK+DWLZIWJasNzEegfFC6LGQGNdNpkI+x4iGpQJwN4UOyyUuxxVihS620UiLCYhLn8LDB6eRM9
pjgSaJSsh2wqKoCO9boBmbMZ7a5mHlahlHIE1LtRH821Y9HohQIYyeEldaE7PubfqdN82r+NdQYw
hF5/HMJ0rXWbFwrejUwlAYfRnlaSkO2JoGklAUZEA5AFpf4NJ5HiQtTCEbxwTXXzB6atJ9n9l1yO
5yFGx85n5npzceJgpqsde/1wYXDvDOLSPhbFZybNNgVbABaINuOV0Qru1umd/Y2V+HaQR8gjHX5c
Bnn2HPG6TPIpwWBLPSXWrBDvtuZ6F/xlAkfUCCpnOE3WKSuIKbzEUzS0wWRq2jFDKdDnnFimxLe9
1WixuLTbzhefXnuW0HkWoOt2fCQui8GgfmmIgTug2vtgqZfZGJIkWi6slk2PzeKCmtSupXc4OEyD
gh4BwP90NO1f/H0dqxeBW2jjVxtFFZ3+5/zIU3ENe3BX85WLzCET1VzASWB1wl8YxekQp+LvmQqi
xMci1o3wY7AQJCU3L/hAokI/kUpMwObD7egKk/yLbjpdXWz1kPkjFArYn5JL2OlYAS8Eu+e0gZup
IZGV4kxwuVQgRZp0BdBjX6uJ6zuQAHc511ID384c4tdMdhRBc1Dc/g7JHGtcwltjf5BXDquIf8Wv
FT9enei51tHgKIxYHA6BRNFz2fzg9mWwoW33aVM2Rv4+nQOoBFLxPRxaY6/ZqwzOTNEe52e3x5Bp
SJ1Aqi2apSIObygIkbZl3+XVCwtIFIzixPxA/qo59RK3zX5H7KbnLpjO2/Fc2CtOfmK60yWBAfwG
bodrE813mq8/jHBf0r/CGJ17SOt+LdsWfDH5bg2dj4LqPX0IqPBxwp7dRaHibv9KExGwNrp08JVI
HKBdhS2f4T2jcLFCLoBdSq5x0LJuo4ipENU9AaX9E1bCYcn2IblyNDpmAC3GDGH8R0NBuZCFEqa3
ps138lOK3UmCRdGS7S2wPHkmKhN2XcQyoTKRi+tBAyscF+qaen6BvSjdatgkBc9ld7d0YMUyxV0L
BpLSJ4Yqcv/zr/L14N0yep/ldp0QPIJ8VkWGmDg2g3+tm3FiO1s5jAEwXl5Or1Cq/jCheYB//aBH
WU8j8bPXuADbDA0aZ3zqFHgVCDvsGelwooW1P8i4fjoA1JrjuUqu3kTIO0k0j2AbhWEtI3QDHc6C
D7AQvdICRvlJHjtqW76Pp3FYdcHetcoXYlx4gObiKsyUB49IqW20rO0MzSseu7il5QOYBvhe9LWg
MMu6mKkav+Rz/3KhEIfuzsvc9Vd666VmF1BpPJcZIjgLypNO5LMaWV2Q9abtAYXh1xXviZwgSuBq
Wm1ia3ABL4LGu3FybuiX1SksoOrhkAovkUZuZmoyYejSv5TVskA4F7hR6LGNx3MPMCrl2/rD12/P
yfIQAuDItaCffjqDFHpXxzl64z68h05dEpiojh0/WM0u5bVT7APO3+DFGn74mb9pMfhpxILm0+tw
nmMvHULeKQCtzEquVV3NQCvKF9Ui0gv1Que/i2mxW9Ekus0KxwgmDwfUX7EjUsRt5wHco1Rx7y2z
TgEUtPOgSw15OOYYjhLPsRXDCdvJR4V/TYEZmA+gciFxR3pZsR/LlunP7/MSQMh9HSqvlFUShHpY
t0J0sBR1AFh2cXll5aT7YZSSQ4PKicHyi2TwPVPIRKUa1jkJ/QvOLHWFCylAv8YPK4xBmX1BNNHW
rzIP6zGN2ckW26xwMpTtqGNkv1csvyER5L83Dp3IW/ypSUlCanZ6OfTDmYsPZof20c8TlhGQIwCi
Lxkv2pe4+0VjNfSYHbuozTVNjwUwjLH3OqOZvlJHsTSSKRv75OQeLdsTqYk8ljeopBtX8gecxpCR
gLnJvPpssf/eQeWDXiKy8N+Z4YaDgw3QGtVAG00INC7qQHoDCBeRGWIfh5GzAxZh+JT6yCK1iJ7X
OwSC9KGmojnGOO63KCd8naPIqyiOZjetmNRshh61OKKhKjYSHY800IymsgJn8GlN5Ao19uEaTPHm
gWVpyPCw1fTA9GPQtgxESsVw25CzLgK9eQv+WzrbjnsWVEqTpEXokKjgZWKa3sCEoBg3xa+a6Ffk
KhoRfjNxK7+sgV5lOSivw8OsNhTXNuee7tE5joXdVJrLvjalhrxBphm1vYMbfBM6j2FNOQyge4o3
NdAGFY9518YHXwybU9SnlLm9a9PcFtoHgCJ6gTFk/LTdS/nnTseMB6THgw+tslfEE4u6h3J60Pn4
N+a75s9kUmXmOG6HxLUIEfIbstmlwf3n1I0k/SPm93g6SBYJxsnqBUGuNzWOVD6oouACipUvcXv2
0LKcEXlbLt+9WnPM8FkbF7M+3gAHnAxrkxwJjW+ep6ff2MzXDCkL4Gpq3sSQOgyei/B+8WyxDhNQ
bS8kfdUIaHeGJSu1Ztb7feLDvQcMmSJVlsc4eCz8L7ejMDuh+p2l/nx0g4tcgc5bvwqb9l3LGiCv
kdEgd6DTl6vUPsJO1JL/CmpHARjTnQfXMOJpDE8L1DtzCfx0QeoKfP7jmpFseH/W1J7VP5bslueB
cYdSf80vaDQzOHtma8kCB3Qyps5C9MAmkcvHCBEVcpBoQOwbWyaJ8PXPIlQvHiLZaL0Cjq8Y2NrW
eQOBjAAaoi0NJkdXYUkW2m6WV65+xjdJUDgy0WwqoxDon67rdY4sn23XFnD97qmqaMhgdg88ug9v
CbfoNsT1EwUqszh8FHlQrTCFHVs+ravT7uFAmKigU5rGp64DU8DO6y/yCBf49DAtxGo1fTP9hhBt
0jS5R5qsOHcvr5jYMhMzkc95cTFi//ISR+m4b3NsjVDu9BGMGp1RTdoeWtaoJd9obE+onY3/2HAx
3qHAMNbp6CDE/uxatB6uKMmwdRv8o3hO7CAX7UyZhmABPAiCLqFdveurI8FUcrtAwsnJQfqsMXX4
Y+qDRTzSf/lRR71L2LQjQ5D0lhOJGaAIV0ioQ8ByvOLPn6Nuo4fLok2DygEKExiQBrfa9NfWj8rk
n2oWwYLVTnJiJpNyI88fQOwpLZ3P9aq1VOgYvbzaZKWJQrxTabYFZSxTaL+My1qghM17qPCyUXyZ
bIfPXwViWfDrcXr/oL/RY/ljvS/n1HMM0H5rzUFOWLFxUZeQYNYYpgN9cvTxsELuHSwUyHutQ3o8
jin06Lwan9JwWES9uWmzmxAxYPt/OrwhLoQwmcui845OrJAyotmfP0b4C280X6eB2OEQZ9EB5LOB
bkjz0iEeT/WEiQayYiG27arvnU7u7G1uSXbXrWN1p/lv+4WiHTMuWWlpEYew1JT7LXv0kasM1IdG
4BGJrFGBAyrI7pD/k6xCA2te6K/ehKfbAhsV1kM1IDP+l/F5RZ9cKdmKM5J3Md2HOaYhQFRoNfpF
Df2aIA50GLdtc7+txF7XKRO7LKj0NTMmmx7rV94jEr0ddpOh29sg6WJZKS9pPua7XxEXcZMgIYmt
bd1phgZho7NdoTldt3D+1Ipdl46zBXURCxQ7H8fBx/0nm54uRXSE7DQMPVVbAn1790C6mRaTdLFA
uznnGOX8U6rcVObfdwr2T++kpeV5Iy6XKKsyIqByBDgDqtBhe/gg7ZD3AwHGQqMb4Ivk674Hp5Ra
+0fHjc2j69DkjKf0wo3r1PR2KsJgWraEWRAXYJSQ5lH19/oWLvh824NpyTDoNHRHclNodwQJCFJ9
G2bK2uclfjhWORzCDR76tqRyS3SPKFG/He+iE9oXVA37OP/oyQmohePWrYbX0CR2kpOf995VgnN0
GoxUkA2HISP0dWrvZRiwbq24tHg67vFQj7NfxUHIs+re8Uewc/2lOuIrNrrZeY/JjYJNBDQpQMZq
208y94eG3PBOZCYUVEwcaBDTLC1HJKnkbEsM7V8Ei2OWkPHj5gKYUX2rFwwO8YjD+gH3K+Jt9DuM
rDhAjgSP0eO0+z6cogVdOZ5ALKzmgj4L6Gn1+sO75BqiD8XR9Fuw1naLuxpZ/EE0ciQq5EzEof+l
EFZbdBw8KdQQimpQkqu10oVUcxcMb6Za5gz+uNJDOBskrZzIgfjSjynz00G/R1zehM0+ItKDXGkf
FJj69u1nOPK2Y1uTsSSVMRff0h4bAjL73mEDbRppSmSPqH2VbqJXgrXkjNW6b/z7i50VfoCzf6PJ
sUbpXystutq4AieOhaHLzJw64eFuh3rvylocbeivg6jXpFnavBZDb0ac0HT9ga1nmRRA2H/BFupl
2b6kGuqImnRpBmzGNhK4jBx2gUuoj3THJ69vefNWtzn9OZThqhkGhUAhX/WvWgwk21o1CF8UVLqe
W5Mjpe2W1mxobDA+dt/3hM/DBYL/yIHxuftVm9CMyIO+W2jOzXWFD38T5KMISNVZZ6mFYXF60o5S
TfD5eNrJYSBWBSfCcPOmQ1Q/BMmXl4CIwqXkeUjsFy3YOtLSQSbq9j7jSWXt+BlbFcqWwJ3toJ5j
tq/tABA3/vKkijLBe8zqmz1DZLAdTHhW7WlMDtvkm2AQLriI5vuthW6XK9G47Utq7h07N3DSprfr
rQIO4US/xd39K+H1KkecXCfn7+yC1Y4t8rtLPGZ46/xh46qFha6Ja6pj50YXkMohLZBdl34sLN6F
A4B5tPtnljzU5fUrIMWJDQeXrcVCdTqZDIOIPTZvvA2k1tdEs4yIiwCUovLhHLDIwzXrFsy9x4cG
eQXESHoVtTVL6HfoIgVVFBmoDrzkYpvNUF3gQbJEq3tkYRoVRtp+iSEp0P19+2wqEm7me5lqwyQN
JsfejdbvDjT7Y0jq8Yp3u2ztFeu8ABcPQ9fApAQCi1wOwTTB7XPoefmaqY9lTNfmDdNhmLVlXiAf
dt1HQjRFmSYqHZ8IkRINNL5FikLei0PaOkUlLAH+h5mK27HJguuiUPW5NWhapwU0XpOkN5ISFUcG
U7OMnaNy+Jx0/cPW9Liy6bqP82j5qh3g1TOrQTRf+WxeNDPoMqbj94KI+0qK69G9i1R9nUpZa91j
psOCBQ8Yza7wa5N6YvqY1+rkOxdFMVs39iJMuQOs+05ChK6DIPFdLPNMp5/9+CXQPl1Ptvt1iN8q
kQ5+YL1BnQvE/Uh5b4+YXMJtl9S5Y9ng4dHrjL5y/KsYJhitYhIMzKk0ApOp2fKZdW1fuNRqvhDU
c1oYq2/SrQU7zmBqzrrd11Z+mak8S2tuYSQ9TiXfSRvoH6/CntpKQL+pYU28CFIMljDZFMw0Or7m
fN5Bed+27XrgOLzMi7EGlireOrN8p9s1adU6qkDm3PZdkaL00ahdp5B6plB50SYBHE9eaVrx789P
boyV/Sklx2wLc2dArT+ke/NTYFMteZ6vm8OuZWe0BTNc+lzouLcBmEpuZJhlvcotVJZ7Z2nf0SXn
tpcG2XuPCg2UIkoR8wxZ509Os0VPt6CKD1YVCcrDMGZODtCbxOXa6dAqe5dzHYXaAsKIwMtKAm47
CuM1LLsz2Nc0Ac/DsDEt+DW0/vTGPiKwkletNdecNd58U9HPKmqnZD2FV88YUOlZfrpNvkVQjRIU
lvs+d/4we3nBxJlrfDbDJUQ20MJMAkUHXVwaM0Qu+nNK23JpqSZomoyn4hckb9Z5rX/NG7b2TEdT
EcHp3MrzN9/LnYJUZL3Wj8sSKUiL1r2nMeHGn+OAzjAw7q9kuNGlx68sdfxfMNh89SwscJ6lvV+w
o336Fz4gfYxyc4bzGf5LDIHSiX5/katTxd7+dQaoox3oY92hcJExESWrh/EKJS+e2CmGmTFJIdtj
gCcvS5tnZadYA4IJd319qYddJlN9qKS3C1z2xD9Y+ObCtTMhoky9CpYdyWLwcJyNM0ATYtTp019b
RXQ3A6EZ6GVX+2bWy4VfRxyywSzNKGPi8c93OM3+nVW2A5EYziDwxgE1Q9908F03Il3d+Lsemzcb
S8kRaayxvu3tENCH+Q4K6mjqfAI2lHFlZs6rG9L6gC21A+Kuj7LJhLK+ATQOhXXICBL8fK0JcvvU
0gRcS09L+zGX2aCkGz3Cy4rnIXw3Osope2OTvU1zZWblSewlHjhsx0XBDIAaJWr9fqBbo2+CXDDT
oX5CZtjUCMZfkRkvj5At/aCcYKAmHdbR7n3pWqCiWXIJAfSGfVrdUrYrqpgSgss98AKQ5YIkG2ro
SN/E8pSU5e8YH9Ob2OElq/Lidmtcjvoc6nfLc4wcRnHyySRTTdyFd4CMM3yW+y/zvAnlyAJH5kKg
OhCS4IWagJ9MVMoO8vr5Ryjan97f8NioA9yFHbmo+lz9LEguIVX8BIK1MC7RPoSUMmLLhCMjTrA4
nxOhTsevUtFZVqKI8gCIVO6jIipCBZzPq62JRq/+68MrD/yFVUZ8yy9rIy1wn1kKGWBGhZW6m2U8
HDneGL3I/IJXcrDr6alIyYgBpolJUblBRH+14nBmTyxRppiiOnLDDd7eGFL5YJHL95r5RifPw/gE
nsTCbs4B1pONUhX1hyxEFhcrZbd6lIsDo/XNCu9gOBQFx6Qh3cp/VMSA68b/lNd0+bjjiWZP7h4c
Y/Knpza/uzq4VHoziRIuanvXia4qEGl35mA7a8dKfWDi4q+0L+DCpUvk4Ve0ct0IEJ/lt+zbzaPk
+AuI41/02N98pOkHLRqfjo2vAyY6cMZERE6WCtdVYaPREDo1/Cxcjy7t3EyG25CFYHXMDE4vqBax
GKRtbFV7e5hq0gyE/dx09YzXMf8UqG7YAgRS4qZnveBHOhIlcJ6ov/YawX2SIMki2JB6Cjyw5EuA
wNliHkc0TZY8TinJ1HVOrKorbVUN4pSR3QYF1g9py/gPo2jh59he574DromzvCqTAkl0PRBxKVg+
ZavR+5fMsJVHE1uTwh3TfAtWP2PZt4Sq99zmdeBtSfeEDQJEdHjnuGLuSmnr2G8p8iei67+/2jrq
sjKPdsQxdQU8qT8Nrb9eY4eAFbtrHGTOaZ4ha10bSxHQuGEs4X16YHoilHUQYbMYx3FSiC4GeS2r
vPAMIUUbJRmn2yWCXiNtJ5h+w5g3OZ2vkDfZglsZ8SLl9+y9kWrG8Y7zZYJn5yFwt6SFbVdjUCpN
dt1hBSa5G9/vW+AiRC58bdNdCM2aIXeLKxflBCrE9TuUYOab7XEFdNdbBnCCsLWu2R77ifAhYyE/
cbiAiDpJjMjNbM58CoyVLvlrqg2xzTaSSyY1RFjUTLtjH7KjWnb8w7+fedIQm86raww9g/j2gz/f
iqK1DE6HrIDFg7Sn7gCPO+iYhzDtiTmDtsyRvmyfaBy7yDnVHS19jWFCLnaOBCZUFxCbhVBOkgVq
kyLBKUuyZtExr7qCG20SbKPJ1ahM1fIVu2WtcgBFz1O38I9kpiyrfkwDhp+qqAiwQzsHADRv5U5U
D9Q50jIMmEDetIqQpxw0AVsn+9b8TOr5U5KaSbAbcIgXXsK2AEdgYLTb0uYGwAO64KFSclzzZaDI
Pc7BF2eW/o4OHsx9k3/gdwkAdoqnihlnxPLGlS+YlR6toDFaUhaBM0nqLYl/8arYpX8NzFgaXNAY
KUHaLdWh1pGorAu0xXgyhbeP6YgA2tXaPJoNzuwy1nfd64r770AegDAGl6yAUE61CH/2JY+Sueoa
J+hh+xn1UOcG1Ombx7yQAcDLkU3zfMbDnJeUOhikmji1b8rtRFKgkSQ972gYYynUj90p3kL+A5d9
kte2TXUCWHJXr1q9phA3w3961axlhHMiPjtjF7IAtw4ZFmZ/OQduathJcgPLBitcMonpoqtG8a0J
5b3Ag9xJaWcp97d1JPOCvmxbwJhp4Cb1dN7v9XvIY9fGGZ5Sw1ZcxpIbPwl/zZV6HlvlVk9+Jrou
PvKyanvRI3wPAZg1QtRSUQE4C0FTu0HMoMzVjSjZXxX5TeiN1zINO7fPfTafXTujVNKIrFfBY/yl
cWe2E24p4Z6z/YV8JkcjtmkPtnjFOpnQLhR/7QraijBPQSq+d2vwHZ695gTROLFC00i8RjyZ6Mat
Sb2r6Z4gbVKZJrQwGg4r2BjZdytPgJRvWR5ZnYMhQT6oMDo2RiCk/gW2gvavZygYUY6kihcje74S
tsStUb+0g5uMRhiS8G3N6ODHLNejtKjpLNpX/+Oqv46zYKr5E6aNR3rvdAShneb+8lG5jbf0xW+s
68RqBuPpnSbXCdi6q9n6WZ1gWKdnggBXN0L2tpvpLaWsUz1BsK99rW0+7Erol8m3HZxOtn2yGSsH
COigJW9WyOHHN1PdBb8pQ62DTRHuMcXJO0ClD27Cd85lLp8iQCfMV/9o1A0O5Y4bjw69qndk+OJK
icNDLnaowpq0wOf7pOkHF3EviP9ufN+na6eU5CGDijOB6XN1MiOvBYGFXr3osUNKAGX5NMlN+5Ex
wEhC6XgpkU5hNj/4M+VMLBSRDwPMeTakYyGrs1UJMV/e2KvMtkpXN+G8kYjRlyntpzYQj0UyUEBO
0Il13x1MclNrqY3L+qW880FX4KX3DX2KP1qwIlYl7l0VTBLS9DaHzDzbIBMiA79oXkHZOT6o/4Wa
oKhlkyQHdMJB8DRRYDjB3zcBAkm8XJXOak6r81Z4GKDx5XXx/nn7xsiN5IQ3YG/Tzt/vJS2MCeT8
5ADsOdthHng5254kCTJN112VUc8lXtGeskVQCXRWkfPPSh30CdN+aydwx8zI7mRGjiAEHT2RpBqv
e7wuvtEDNTEgdonZ5t68ZeOjZapRAFmKgS+1565MQ9zMvSEEe2gcglQGTV/SS+3ytJJ2xoGLxhBc
dITgEyxD/I0pSQxxfUfSOwyKiDgoZymirBtVleeVyoGSsqYBS3CBQMcA+PSaDtXZf/5/jgPIwJrA
ubHcif4PU2m2uchph1MEdamRbK4yBD9yqx/+xk0os9KErqdEIURNYIOVpWmtJXlCULhHsrZ0AvO9
/7Vfa0SFt3kNeJpzuCmX/5FLoUB/O3QpI2u6mwvDoSkBb5hldQOCjiae8Rien58MYEg6JxcnUNfJ
qI1ZYVLdJMGA7RNaqNm+OlSZZef5IqjNh6TAKVpsYDwtqwhgcNWaX3BwrqyQ2SmkwGFwPdU1b2Cn
jVTNc0Epmr/pKTp78fjm7gGxXRVYomGe6sIwKCoqpWDiEhQKwspwRozIsJMX9Qa7X81YTlBKtVSS
kWkEdHsLnwPTGVnM7IYowRNdf8VwcJUn+go1FLcLdXhUzIK7MHB4dJgFwW7jOX8lFksbijo0MUab
jRmbD6oPnmqJ3HedP9M/md5yWPzTZEufYkaVoXU8MVQhl+2bTERuYCByhaHDZOdnhJxxdI+exq3o
/PzjCEc/NlfiwyfmfDwLGiTiEWr+hhOrGhtGnSnKkU9+3nSsk2mkzgVYVhI/nMm+RtPsqxTmu+4d
w97XaaBJBJhdnGqbxx11GcNBqQdg913sABNNfWaAqCVf4oN5MvEq5AMxG/CUAtwLyiKzEaX5hRoD
z2dLO5yQmS0ehKzUcGsMvLOha5xRWP4yUBo2Z6Hd1sptYLfjpFQAiJm0dVLykXED202j8rK7JHyL
i77xDM4F3AUUFT3cpUhY5XbvqZy14WirGRt6Ji6N9mFS8e6U/OjMjKVVaR6pOt4XeNWh/K4oJz9Q
zEFeGLe0tgGjgXwKByDFfeIMIzW4nUutqqRM6RpZ7eF9zN2Kc1Z749/uTeXDpVhbmezO1jvad/08
QdAFcNCGCHzQw6/D85TogRH/L2eK1ZvZLRkHYeS6PViOOhl9zT5HqOol9htJpVfcp6ZqppTWuGg1
lEnaltosYhTiUVXVQr3rGYGxAeClnPPDYLcNi1v5LoFsKVc5mKQlZmf6jZryak8sM4CNGTK/cKno
DAHf1zQTQJjEQQa3r0OpFo1WaAbpZL7wHYRcnSyOb6a8ntT8OCkzsu7bX7VcnFzF6DuIEmSU3vpA
rKYl5kwKVzqHm3ysOZAEnZ1Khqs+7Si3Z1ZR30zSBotDu8ed+UTo6ESOICxRFJ0Hb2MZF2PosNqv
UomuwWRLPJ6X7csBEK3zyc7PUIsxZXgxFZas3gmxHB8kE0FJNQHUh8ayZXD+x3O0+THHYshhoX+w
ZfExORM2lf1TiYpS6OwtIY8366IyzZOsNVun8PBNs1giprbKDfF2Zv8DZeaGjwKVXa7tmnz0w7Wb
fPv/T7fkveitiTBLxFzXRIeGMVM9qPjv46unb6LWwoZNl/iAhZ4iYXXg9PAScDiAMjj614ClLzB/
zhWYy57TyfGR9P/TG4wob9YtJKgB8XtXqiE6bNWqMKlhcuUuHdsfhUfcmdL6fMb/Gss8qZ78m+PL
5b7pkSX3MCIQLIGahqcuVn6xVC3aD0T5EpHgj8ee8Pr+J+dX20G/hl6IctZLXjPkMiDwJ+7rrgMY
aTraekqe1b/kTKYxFtc79FPlYhzvWvRvdwc9ww5Q5QE9ASeY8ZNdBLpLDNn2ax+0OJ7cK6EZ+pi9
94bkRLZg6a0n3Gkh9Qj+dKUyMJTnUP+iN6h3B+OpMBzP81bmpTJcIanSBwtrlqfCPFXCobTx5N19
S0AToB86/mcjfAaC02wJN3f7p3CxP87GrK/ugxPsVY0Pw5zLIIfSGLl3VdL+C/7nRFOOwdkVCKdH
cKC4ytCEdGVEj4hF503XhUvdDzqUWcIbEO69GssfaBC6VbhFkyi5fJxarc9W5qlVTLaGW6IkFD6g
hv989rqEGOBwUOzzJbLrNeu9zXjJaOl2K6MgJ51532GVHp+SlfHM43DguiZjg3LvrSk5VMwATdj9
fGvBUP1VrM77toL4nPDm2xTJot9/QolS5asQ0+OUav9IBN+Q6DcYdj7P7XQsxHgU4LL1VL9zvzdr
UPcpRYroUleECRPVw/SWDSF5eWLijyZFq8wbLbv1Rhf7xeK0h3wbWUA1iQyAFk5kGLPsR8P6ig+i
lj82TR169mQ7Uf3h2VoA934LD6VKdVhxpyWlf/rX6XpfcsnIFMSShIOclTaxmg/kYJ59iVipx9Bi
Dua/gJd9HqR4EsPHkAZ5AzxeVZzivXAwH7q3IPlg7XEF+Eq6i8bDuOIpwJavknC/WyWiDkWYPkBu
F5u+GCbeijPO9u1tGY7yjwLWuiFdFQB+MPwqX7whgwV7E94av4G8hH6A5lTELUJuXMfLbkXF7p62
L0wpVw0FAU8ioxb+9fAoJASqPIBwMQd4/ixdCWqtMvIbKFvQGvdgXUPvBAXQoTXNrpjvXoxF/kXJ
+Sif4NcolRMP0S4r6YDDCT9whjuITxN2QHMBt8SLnu13gwM9Ao2XzGPiyOQu/wYtpMbtgNIJdT48
8KjEuSrzt/jI8IuLhW6AWMeWEzXhJa/II5P2JiIL4JFzyj9rk9ugcoHT7zhcnNArieeR+/8Z5Qlh
VvwJwzv1DrqlyYx0W0pTcZXkxXQdcDu4uGc9gy99hYS5Ca/aQdeOcJfWQGTwbTrFh3OT7kfxpbT2
QhLgsOPm8a5B+C6ONq3/57Olkygv6AG3VjWZKbDL1F4Q10HR6mR4CuBQyc8mSYlc3baGoNcl4dk5
nbCzCBPG4WAYWQG1aBaGbyRElVllV1wRKpXS+dXloMTy+S2jKnPHUkJMNCAEiyqcA5148B4NFzdO
wBAnJ3tYMLe/C4GbRGv2Ivi/IdOk4tkT+y45cFnopH2LHgWcjFZW5Tc+SgucdD9AZgxj2Nk6DEb0
MSAvepybMmp3OyHMTfFRdy/CTx9tBI3O5WyMrjGSC9L37Cc6M9Bl4BHIqa95WjlOlWue9Pqea1oT
B6JOQloGDl8Z5tWKD4NjaMzYLjr4fSJpXP58iBH79y7NciCBQE3R1c3rZ3Fvbu8n9wfQ0gjx0UH3
QG/yBMdZLcZaflEEK+MbgrbgpoYySVE3UwgxkCshU/178fM93beWIsbzqdk+rq5xDhjv2e2KJIEl
UdvXmVi7tMtgiQFK/2YqViq0RsgOH1TqogvilGsbOoBozB+Bgz42E7z9M6qxXhrgEBkHu8bnzsnT
of4ID8hcsLG3CSLn41NsoW2oZ9AeIR9riQqyGb2je6rCHP0rNKfo0XfU8W/xhPNElBhyvUG45AIU
oKbRGqVyFCrjUzZjDRtRN09geoFAhfYaidtIVJyF6h9F1b7uIFxxfoMLNNHmZ+UHVVRdYELr2S1C
L0ZlHq9NNdmyjFnTbNKGhj62oM4/slCjdxSpOvSUWqgp4Bw64eI8WaRo5xVyHFxfcj6/PpO5ikXx
BjanYCqQ0cM2Sa7r4UkzfDMis0TTr8LjthHX83b73pheaxv/C+ea/a/KxrjWfa/SUwEU6KxTGVwS
hVe0simsYz8s27skrvxDvYDJOoCW9+7XdXFtAX5sdzwdK6/rT3xdz2KX4H8slZN4reES/I7i8ZnM
Gwi/NwHSttz0KrTkmPU7AJkmdgBaaAs/0xcDYVjPki02FrMOTeCfiIUzDrd2bcEUuczYlOErQwyF
zC5BcqQiUdZewP771GV9lcV2F2U3njvRrjyRhUQRvS7RfDCFYXtdSrcZb89igrIuyPI7l2V7C9rg
O5KHl1PsyJOvWgsp0haB5+/pw8r0v7eoXRuFQD7csHqrfu/c3hL5Xyco+qfK6xMKlX1cp/kg3xyE
BVnwd8UnaVIaJb+UK6T7l+KXVgrqa2WHwv7THGK/hvNGDy7fhDDNG8GB/dbMhg7mZkbTHkPgbeuu
fbDDNp93n+v5GIa0zttWNeGZXAXCOD1xH3a4EjI85mJqKWIuA1/Bs+4lrv6JNT9vZNwJUwERMuzX
FW3+WhFkGc6o7dmITXjVAsrmJr8F8V2vUJNPagZucEtErynbbt0Xu+q1OrOsIK3/FjTimeBEDT+k
GO+JDBqMJuCHqN0Dt5BQKCM3DYxSgXdz3STQ29rvX1AhbDdbMcc59ZwvNHZY0lqb5+P4YjH3gL4B
XjHr9w4sznNBkB48UElE09C3UUDRF8FE0fdRjwedj6Yuc2FdPhFpwobTU7XkKKPdid9IlQsmD/GW
lm3DTm88WnHEvYWhu2qy3V5bs+dHAa3yO/rnLoJ9KAJSpb/88M3jkOrfHTiGKY/MYT+hVHKETjbF
NQPWgiQGRtax+bbr7YzEFNSkI454IlTpUZPLaZxcTci38EZiehPR0uagB41Fv/L2BaG/ycT64InM
Z2VFqGbSBPpQYnRHu35SKjxEhYBqYeUcoeEnnC4Z97XFkRR/f7K1hNvRFCXE/M2WC2sFK4QFTC8o
ePsX7dTk0OXQ3x3zr3Dsmvc2j1AyFs0tU45r5SXrRAx7IU1oCGUzxfByOzk8XPgWRy6PVhR028Iz
yzhewPxaDlYSSi0exR/DEpxPRFV6k51kSKKvjrUjfvQ8ahPtPRkIYCqtAkg1SFe6LYaKu2Ju0lbC
8ZuxYxglwqNYRIJUTlAWivnh/mHvYNDrDOx+AwydYNHCkh0+YQv2g0Jjstuy+a3UDWek14uE5ssn
fa9Yi1hV5hlG2vqnfUa9EEviIKw/+PjWswz+6DMhvAEza0zkFmuYGNmGOiHshnv+7ITZaaGUr3DP
4gxtEI11qdhNb7XdVA6PRAi6qKGs3C3hiM1dm1JDpTr2Uzdhbtp3PGu13IllcpAQBsdajkWjKc8x
5VI4MrL/Eb4NVDFexc67pe5sOKx620or/8obTqOEfcvW0Uagk/cl+Zp1iyUXaTMmGrp4pCR7FqIe
YuF+wiyDmov6eQq67m9uudz3UWOy+PLU94MwF1LIb+q0j5vTF9BeWZKuLcqmpTPy83rWu/H9DZZI
l/eWshyjahjemHerGvvAsNswz7aWqCL57QAp8+secrA19Qm/5Ts8CckTWosgWSBBG6Os4wEJBtcw
ptlLphvn3fyVUt4H7DIoIMcOfSzx58z4ItpJbdubnDTs0oX6oZQRoTEVwCcT0qF7Q/PQbcSMLJfZ
HldEMntWUwUe6yc2XNGLGy0GyverHXd5FtdBKv9UM66zDBYZqtpqBt/thBr3Zeo+QXem38a9gafs
dkcLlYP1EF68vJLDIXsn88Gw30ZyaXv0Tqyc3KwqVBNjGN2Jd5veLhjG3NzinZ6JCm8zPt/X6kD6
ZXytF0sydlb7J5/IkJW9gegodjs/77axnZeh47LRt/hzo5YX0vAL4aVKbKApX9ZRWlXU6zecI1yR
x6Gs46Kiz2e4mVplW7/KpCvbP22vOMhG+rd4/gEGtGsDWJwqjV3BF81ko+ud75pWjcIl4mPfagRz
f/6og379eE2TVFM72RvxgD2/0G52GF8QTBtSxs2NeB+qqifeGXTqax/LxAMXg7l8JplAlPnnl4m1
UiFcFSCpm0qKcvqKZvW8jBhbB9/bghpeo+fBz+DmYE9z8lrAODRSV1U/lPqAr1NKP4fpanGE8N/S
CHAAV0WYB18bu2SfD+fUKPC5b0ICb7NxG0MQFjdKYKxKCwVMheOglniSL1jbA5sGTo9Zd9M3VWAn
p0GmUVPQz4q5FJxPKljsXVcJ3jwTRVmZvjU4hKrfImYn26tf+5mTd9EnO8T6e3zJTZsNmH5XQq5h
JtNC08vY20+kXUJII65Az7it3Gtc8BStj+JQODs6C8QId0HGIDfoaoIHe5thLWBpm89CN/UIJSxx
+SwV5zl2njbGchnlhYyeaNxVnbXIdnBv0qsGgUuVW+g4jVbX5UF8iXm8NFG6cjcxpj02Sk/WCp3c
rBhDOrXgukeKpUEDUbQtl28tyogwrlfTT1b6pF5wQZYwna4TPQ8RfQEBL0fZdbazUiJgJ7CAfH2I
lCdReshj9dXUyVLBSBzBuLWhESzl0JtYk1YeLwxfW3dA/3+zYJQ1bLnuj3dV3abF+sVuvkZ0kxIC
TYk7lh/2oZfsXL1T+P0bdfnTj0ZRrXDfH/+WYaNYVd/FGBF6bqV9cxaLkr0nsX+qgYozfgfeEb5O
DPrXW/zY3CeOm5cZDU9jxwSXdppp1I9mT7hvx0HS6jNIU+Ygntcy5zXInG6j5ef6zQHLbpza/OjA
CuH9PJ6KuuFAzzD6dTEffANQYTXM7/44LciSjMbrRqUmriTmM3cXm5Xx5mtdkG+atlAB/rZiyAAA
qnn8Ip8xchP7UuMcPiks1dX59klCt//4eVsIQtZGOxdl27HZro28zVCe/OvnFS+/3ed25TxI9+HQ
gz+H8TKEHReYxBUAjnRsIDp0mFsUjiYGgLfp1HQOixFLmLT1OHAQjNRjxhgDVV7dJvY5bH6igxo0
h1hHPNezyxnzu6wYdQFR6q6mD+p8qLVNNqYjBkFQHbz57OEjzEHB4a3YyBomRJQt6RzO1SeATKm+
/Ktca35VDvVDukAFZJjMyPtXH18HarGT0kNHl3oAcOUJDYT6yySludCAAcfuZanUY9zAhg3sogpk
b1vAcWYWraBQruYF00uaQenoKCtEoaqbzn/KG9uqIT4tEfmfZOuJGijSgklZvDzSv+9PFvdnIAhM
6aoI4YVRXaePTmvxWfxaMC9XuJHd+0vYcvzSl0m9vv8Gl5fZER/wuWRfaOClu5t2mUM2QriXcBdN
nbk24oi1zm+LTEq1IDhsYGxPYOqrxJ37zfNOmRJjWms2yqXSKYtpYSH6+Ynku2HB33ix2ZAfsH59
CqLxs65h1K1pabUIGD8WQotc9QI+tTknoRI8fKnHqKg3aoIhaCxT7fvBYt9QmP8GYS+LHaQiTv/v
9Ccwg/MVJfJahXfmHdF0eXlRI0DYYs4MLWFpf9OW42ng4YvflS1W68rQDBrAe9jFiSQnDFH6sMuu
b8Ov3jSDA4UAtrQdjy/mvqrMXyAF1aTzhv9wiMEzgQiO7X17phxC6tjPMsj2fAF0jmAGYpFt58ZC
5KRqrqbFxblIfUlV+T/0+PSS7z7eP1xxgDCmjdmgp9Mc+yk9g3dMstNLvHj9Oq3axrfnkqpwS9dH
ciX9LulqF5OEnFMIvI7fkmL38ZfODJlXehzJ4V3f0Hj57SOqwyKqeXVyp1DNwmHJuysgN8EoVyCW
Q5ZQQbSB4tXdNMoewy6ujZsLMUy8L4a8x3XXcHVjIL1EBvET/qgqYmjWkFQQndnIwlkitTB+2u7+
oNpRuGnvECjsDwrU4bTgKfXEiYgyMgWGgIvMvM3XNGYfH7vy87lqGG6RidCGBUxadvwT7nykPBic
E1VDKyjfavEFKzCAMWn3ztkHeL+b68ZRJVv3aOdfM1DDaG7YWeytRHCPYuDZKdNF9fvJ750PNmc/
l7FOZKOPeyW/jvUT/YRXNX52iq+IYCXOBDw5OSYNo4zSzT7uYiCLUYJiCvx+mxglQdT/wgmsCuVq
r/MbdiUw3pb3cLrSvoZA7L67HkoPWZ38tMOYiFB/lOHbWEQ9/bKoNrEBKFLEcfKmeUQsfuRSUaz8
Z1FkTvUHHa+M6kshiIGPDz5KbSY8csY78FvKiwt/xnSjXgGhoNywtzVTgqlhxJwNN2fnmQEsdb+c
sbVSb0gUyMDHwPHsky50ROA5QBdMC/lrPrvsqPKzS900/2EYr4FjXw3St7bvaDJG5X6PgIkh+O4Y
+wPVeAw54qcCp8v3HiC1FBXxfqVqeXynHA0g/XCUxNAZz1AiyRYtr/uxLPddW17WmR5MHDwFvze9
VjBbrpD0OD0JMM5i4fnh/bYgoW+KSpcNNEYfEOEYiSxXOFMdsqCaGo1L76+noUocO6/L1EfvNUVn
4FhA7CJTLnusNvkgM3CRd3vvykZsgKoRWgcu9F15nS4suwJ2kLX9h7q8a9NKuJGwb5XrWvSCwbdJ
BVxNBPD3oWR/dYcgnFWaob0mEKBPcNb/XaGkuv5jx//LzHtd4U3HHapvUG6k8tIM7p72ViX+LyJ2
66+W3IAOA4Hl6Rq5+JJu3Cvi+Mqooht9vx5QX0PVKYkkpofqBPxl7ChQam4Puj5cFiDQ5ZkbGWGE
1YyI+WvxbgeWghvMrM/+WqqMqBJuWUXfN61+fgdUAklK48tr/mqRSl2HX+bCUumiMMoIWlteQKAL
neyZJHc/2sRXozpd53h8AEHnKouf+USg6pITahLW/rk=
`pragma protect end_protected
