// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.0std
// ALTERA_TIMESTAMP:Wed Apr 26 13:33:37 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Gp/znj9yXJLcYm+0QWxX21QyKnoCilJqlkXDyKrcDXkBy3goAu8+91yCtkiviYa9
MxJccv2Grdcil57pZueC+TRw/JGmtkQCEJL+zqWJAqWLnxe+ckknTk/xwTp3L2xD
iN/JSLgNKrDSuRl+/7v0OLbfNbP+UjLXYFw54ZjmfxE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 12336)
Ns9EH98gxyjXbufLppqef8y9ORtGcIAzyD39i01NM695OwLsdsrC8X8K2ypUankw
Oc4bYi57xEFnUzhHrEyV5+aFlsFdX10WSVO8y28yDkEoMoxFUjT8Y/4YZvHPnMtq
eGChXrj+WGLNGUkepWzTJRfQh9t4YaMHdnhPVifszIbHcmdsiD2QfTtjTHV5SYUO
t+cdnBVlmjolhRWSy5f05fDeX/krq7BTuNbOrSBEhZsdH5ZGqJvJczwBiTBPrwVl
dkgDNdsMKrX0GANhumwve0BvCCHpDEJsQfwrxGZyhRozo4n7/pMYeOC392J1YHEO
dzJCOxKKzWKhb69RA+uZUFMVzYVyQsSpOCmjiCAxNbV+QqAdky4HnRWVbbbj71Dm
Vzam/kr9uFx2LI0Sz9kbVpy3JsUVXH9HC8XeR0QrJhdUpJTnMgKCtit5Zwnk4Qsn
wkk9lowlxj0gfS9aZVcO0/SN0kbN80NQ8SV8GMi4TXkFm1v8NgsJD81WvvsrRo5d
xywF1wue9N4zJzqDcvAb8EdauJOKFcKiXKIbmqYaF85RjtyfcczZJcTK03vEHQDh
xNHGZysx/7v6nzOs5FUo7500EkRMz34nQMuJkrvnLJ9SWDUb23nsa1EaYumDrQNl
dj8wtqAu8vLZhRQFfG7BLX3P0uA/8pPbn6oslqlyJiQ7hQvewU1ul+r3Ug2Ku3NI
6kFV1zsNrHBOHZDf2EST9ofneGmtSFW97osjnZns2I/PJiZd5XELI0Jsz4Pe+AEl
s+s1Vvy3jo6hb3AvNEjXUCaVdSv8NhoZvdLx5jzllMNolXg1MJjnoK79T5+7QiN+
yVPdvaPrPnb85jJhub+3LIEAgJp+4ks8wpwLJlliNvxw6NO3/eZc2nGf6PMt6enr
/0z3TQetjGC7HDHYUc9m/qYxjFOTSx50EqyrcFKy2MD7cMPWfFPZv+yz3mFkUnyG
KTwZEiFjA0o9/wmmRks8m9BzNpy8PxKq7aMfJDtFceJbjAGDod7TgON4zAm6AnUH
6zsss32zM4coB76arQg03V3ApuUbek0MYKWfH2zHMDp5ZoGUNosjY+Y3snAtlzl4
cK6qnteURvmwUz41XMDy/TojL3noJmM40cQcAlFmGQ3iDqpS0xJyUJBGLUX4McZI
NfVoE2BLniCmX6fL/W9AqTZxe34MiRe5eoe6UWR1QOvPEGfpmJUbLTdK7H5dh1/9
TYR00KfaM6MTfGpY3YvDMEeYfJGR4mZZYA95yTr82qSBLWGdm7FZOPPr30xX4hyb
skfptRnWzU6aGOcIC8L4yDkF5Ubis6fTmvt1vdfxy4jFPMDrxJkczY7dZV8d+BU9
4eGoiUNQIJjnJT+UhKZiWDrRMNZAkUR1bqknxtXDKXWdBtAgVyVIP80/fi0oFPcV
FKZFGWnbpGtNPusUQcbS6d7d9S2wPiXXMFirFRgMko9KwSbYR2Qn/HyhwBaQHByO
CDezWBabfnuv3IfJNuq8rnbpGHsXrCshe3LOtxQfiVPqG1agwL4yiYPO2TZkr52v
xZk8j+Ifc5p8TsKXUA96stvyosAlvPqVBiwh7KesRDAf/ghCJGEH7NomQJD6+hHm
eq4T5eITIY2JeKEoYAH1P32ERRXMkrHS4EFUQpCFse9OE0IPsrSk6NyVaHm8TT+4
JOgOGJiBWJW8+k0CnPoSjhg1B0KPzeoUn6eD2NoK7T+7HvmN1FWtTeVJzlnDXJad
wCQ70801WV0fGGmwAlphCmNuQ74DKMXxPcUCR/lCmGU6G9SCNfv6LXZf32e9kxQj
SIzr/huA9OLHoXboglcQZwD+zoO9Zuxta/PoOFLmfZmJCR1WtIr6ZLdnAuICwHR9
qk132asYP3V8UMDKksugt6MAPxMX82T6fcHhOe97tIf3cJMTYNZ7VRgLmXCuJ95u
55sCE7wafXcCpsM+pgLdcApztE0rqWniOpwFmauOR7KqcDMVGTPtWDP1ot8AAN8b
bDa2JPmy7zmN5k6vtHXtkeTR1itr2gxOqt4M0QHrXM5JNZ0Wx9o5igQC/5YiB0Hw
nUFmF/+26y96S4clEy/xmDP8gpzPSHTMTiSdzP08u2FoV82aEtTETWnA2ZiTJnUy
s4NeXep/5T3iAALM32qguEreM9apE2x4SEVcg0pAP4tgwSJ4q+56ZzT99BcpYJYB
ByZLvlJeC0YUwg4YemwXBrwT/S7hmxMfvVgKKvSnPEw45+VU7PUg/6gwO8P4ur5P
K+oSisMgtwSO00kULkoad/0dQwpw5XFp6xaiqgIjyfqdw2h2UGvoAjx42e03EZ9j
63YcqvYDAbCTsEWQKN6DCiz4Ao5+rUzQJpDnjCd8uffEDfsUFdjRpR1Zh6Db2ta1
SimcOJOBc5GuhTfRC1YEc3hs+KHy2yG/M4fQVAteS4SY3ujEUQqQlWFOpIQjxobB
cw/JXSdwaovxvCboWh4+dkoQccW9flnFPy+RxAuuynfKU8cSZSTTILHeuWxanylW
LFnk2/32deUYL7oolGqrlWuGiFc7Fpz+pvZxmdb5JXhkfHZTq1r1KmVRjJgdNX/0
86PSxsAHbPM3tgJRfmElFB1n01J2Kz2U69QciE/SqAgiZxjA5kvO8HEvU2MTX2Pv
9Uh8mioKa9zXccebzPSPDZ8RZ2e2G7KFzddKLmsbmR0mwUTbKrnCjVhnrIPJCbhx
2mnwmBjeFyFOxgdzu3iNSSbcRqqYiYtcQqbsTIPI6mhkHw6QS0WNN59lK5Mage2n
oaI1OvFV+xpbO3LN/577SDjrldA/jqdoQL5azbma7ohSU12CHY8bKJFl6UhsTEEC
X+GLNrkzSHEK9HM48JP8sLwc2MdHsk4ywYFfJDyE2XOhZElex16tkj4SIDYG/Eey
swtw6RhNsEycSov+aj0yp4RR7ue899/z6BFYDebIBZFi1310yirQzhvCrRcVjD4g
QVVETl3ucIt/qCgRDd9p/bSOePRTll5tDonUmc9kDWfhhMArAhba2VAjVfBTZbmD
N90Aas1HkwuBdQFLXPkcojathr8qBtBM7pxGsQoSeZMYnnaUDUYZMh05ZSyKo9QP
ZGKvMDEIj+/6Tb6kN/t6y1HsyD1fWaxq/MYBDfvAsj7WQO52mMF2bBAl4FcCVNkY
BKGqioPgyYGmxVHVWGeRmD3a1PRu9xaj3LgEHOrY/FCulTev5h7RPd2WdagBIRku
QZvXXJzLYzXazNhsl+XjTsJnjRSJmSnQyaScmBoo36on9NZTkXUO5gVz2H2nM0Xr
WvwITvN/rqN0wr+MD5wO6G2EsCYQhy/LBYpFVeWi+wOpfPpbPW80Z96hzecbaXzs
xkPpnAS/bRalI1Sm1rajFx+yq3bB7N+y275NAKXz+bK8UUOVETWqf9hWsYW2mN2q
EH9vdf3DGqDrVedKeqBzrvnzuPiTOtHa6hVZlaEtW80Rs9e/SVoNk4auCiGY+ywq
Yy00F4JFTvefEy/qVYCzei4S29x69deaXHBtl2DAXazimObJJJ6xVOKBSdRcLWdI
pLQ4j0mmUtrvsx9sbpYMMH3s+38osQ2ByplhX2H4os+etahoElEbl4IFFzcdSsLu
t8F0RUTwniyqo4zIR05/P6sFB910vVJL75dhQSdDstVpL+Jj2b+K86nn5FJqe/Du
5dNysngLVVuLHxKgF3+gqz0vOU7g4yGR9uguew1+1gwVYxa0Imxc5YWoyJZHKyZ7
PolG9ekisu6h8vQ8/a1gqL355KYGV0PHMRLsjCwMzRCiXQaPthL8oGIlF7LwPEzm
7t9Z3ujB3siNzCXhNBdGsJFJEYW/eaipGq3IULk04MQKJQv0GsbIHwc67kcw44Vl
SLyr7NYBMpzDa3jZ3/DwQ/Yl16RcH9/EJLUu4Co0NdbZTfuPMr6O2dIxjCANvsa2
P788vqmTLb76iLDOpvygDbFMdnwMeAgEgFnDCrG9Nx29Unkv4c4oLnOOhjvttEcS
Woq9Za1CJCRI/PwiKR4RMGubr09xnx/9gz2uzV8KbLJesxuOJJ77uw/Fzx8S3yJ/
oXsxLw9Guyhcf1JKw12UVpD6syv1Ieffw8Fk9eitjE9uo5ylNqp9qyMw/UCZVvPG
Jzyx6eH5SB0K02L1qtHgN5UvwlMKs8qFDYC8QYJPVxOyZrNZ1xMGhWxyJoqYehWY
lusyhN7oK4A/vEGOItdxuhvZvm7X+DRpa/lIyacQBepFAaxIZv7eGo36m2bghzEm
I12uDOafpXgkugMfvK8b7xy2nP+DoEsr9jbP+THTvbVbHdVuF0/9AViNVGs8382i
JypUAfmgfwe7lu1FJtoAkDO3ggmk4M499xzrTbdPt/5RzHZFH+SvfGGeUFh0I5U6
QA8lp2oWuv7jS8hk/SdNpA9huZ9QoOef1ms91IP2uJjBVrAOF5lNjbAbpL+NIQmL
g4F6eByek7iuiargx2UNGrpZuArWWgOZml9z6kYIDQi3E4KwuMqkmDbL5rFQjxxu
0Y0fpIh2/JPNlbvib3+QTUNiq81si7WplQEDlMkkvMSBkgY3dUsEhPPJKnI6sacO
ZisvepVW9z67uZw3Ex/vlv7aeN82Pnf4sGDX8kpDXXhQocu2pg005IqzTlhdiFSA
cWANsspdLJAuj8R9DJpC5ss4lXDtHy1UM07aRcBJR/YE/fKGreDT9sL7/+LBfFkb
hktOIePWWo4TsJMOBl0gZdCwlSLfro6cF6erlpTumghAKSikWw7PXZ4ZuqSe1gTt
rdI1L7kpb4ZccXHu8R5K5cJgfduqRVNkZmKdYCUcV/gTC3DWs2hfBYYppnXnG4EO
S7aQr2mkxLFOCeYG/skYhRiNRQERCj17Rtffj7HmtWfVRFOQQqr5lza1ld+p5o0G
DUBVLbM5iS3CNgr8S+VKdmOHY7jxEqpAAHOF1kVkp//7Wl/N9WshgNH4/6WE4Bwm
EkLPNxO80Y61EnhQBcesYsCpbVZoTlUJ9bF0CUxPoxE9T7hEcHTGm63ty/qb7kwd
/kgPqeygOCa8yBx5XXxu3FLzI+vtVXsOTJ09jAcIddVlV0bROIyDpTq7AT89UxqC
odhD3RTsiAZRbCcb8g/4Iv4QsPYBBg1srX71gTVvh0yx7B7BaAv6plRtmyn5FrIz
AjAhsst9QAIe29loLlXgTOTayln1YTPFhfOb5KwGzyD3iE/T/6Mq/hNs4pDmZkUv
Ea66mZk5RiAf2Djv06jS72YLk3AOcIXzCV3sWY+zn4uYYU1fswcCSFYkOgcMZRgx
hK0D4CvKYpvxsUbUav6WSrWg8n7aU3v9kIIFCgfaY0PA9SGGimHIsrIzZTAJgQ0f
hO3CTYbwluKLdAfRz8EFdO4/Bl7w0tlFYs3jJvXpNEIpVNDDgRw56OUO36xQm7tl
8M9a5YplN6SQqXwpROBmdi9LGNzsO/GDQmIVQr25XINEVI9mtKetdwg3qoKxI3Ag
R1lzysFG91zd2tePdV/V/vl8wPTeWa7rygdyr7imYeLLzLToFzHpJ7l3+mi4Wl1W
MENVawBvFp1CB8DYQ8ASoOfskDLQ0WIZ22IQeW0Vze97XrzEWZD7vH7eGgi75AxI
J9BemRI0HwH3VRLUVJV8ifWJVHWS8IyjsSvZNrcJkoTZ6tLYFh9UvRnb+T4sPK93
SD458qDosfGf8dZA5+mNmvmuPN0yzGXSrC5TcPvYOWsu2DO7X2hoyrf/OBklpCSe
Jnw+Vy0OU8Xe2yRYy96WE4XmCqgVxaQ+12RgA6gmEMDYZo9cCf/cu/R0xdtbBVkm
tSJJ2zBkV0zE2t4JaX8w+FIuK28VSJRyzAa9TUKv9uX2zLwqwnhF0M38HcwoGkCR
NcXOnj5Ed2ajMJT2lDmNteK4Pa3gCR0tlC54jWJPCNMUgHDeRlAtusfs421yg1ks
FuUx54pDPMgZJuyyGKPbNbHsXKMbsgzG5z9Qb43rsZrucG9oxI7YAxt/UoVzpMr0
pH3HHxcYEtMdQ6dyV6QnyohMlFbuhUCwB+Nw7w0iP31ZRb8zkHOkt/o5IAbkCilt
t8VYjGQ0vasuL5u7WgIBGcIXNaK/7IUzTsOj5kUQzxdAn6sbFktWK5mS60v6Wxa+
Qszbswd4LkbKB7pePfoiSzNKpHa9SGBWg3rFlnkIxyaV4rQ8ohpaUmcmNN0hvtGU
C5cXch3MMBESXYugU6BIsWT7IBip1ry+GpBs+q1StZEW9LUPwo2qeXSaTjmZSWji
E8Pn7vxeMer2epmQmzmTBfzWKRa8J8Sy+vu73iznNez+8fCHNw6VW0Igof/9NZBQ
f9NTRtQpfpWkkVy1e+bt1tawMxvjk1xwY5nPyBvWKNmfdI1J8OcYM5ZwjRgKPuzA
refIkMPsIdSp3+7AHjCRRboSm4C0srVDX0q3TK524K9KlYoWUbFcA1WIg3VJu9DC
BIyKM0Ky/YJXDewwobfshtLzQmExoPie5M1y+PEmTiCHwSvLzgj0P8xMNQGIUHn5
chV7xuTubcxx1LLwWtS4HDGSIl5m+rzSuTh78LULrC8ijIHkUVHRTRrvF1OhiVNU
eNZjQZQn/bwttvkxCxy0UsG62Tcx3gXZy172aXmnGn8BYAH7V/+hhY1MUpIuWfg1
zB6Iu/0m8CJNyPt32S+rRuFNkJNZvFlo36bH9WfoYIPXlCSO4oTlFXWgpDC2i1Y3
wX3oXEAhktqQGCfzUqayIIzuEoY09kBPTj7gO3sIY2q17oPCreDAgxNw3m4OKZxh
N1kMI2LaI/Y5VxlZTvs1BWRfPZiCb2JL1xZRx7kU/OoCOGXr2/HgXb9s2c8vG0Hj
dTgdl6qoOVT0YB9FXuqAQc2fUiVvlFOASZb6iUTRAhOinm0zaI4OGyXk9Ag7rNzU
ijdcENDv6CyRAmCYgrDGEmI8dv4tF4Az5uEvVXW0jvtSII4DLE+ag2+67sB9m7RK
5d4fXO4+ccqicGdRU0UBKNl7/eKGQlth5Rr6Fd7JzCvnUVz1QaVnZ6cCg0LBngfU
GKEr/5YKoUWOSl0uDvxF95Uyd6NMIwUQU91Vz+NEGNd9RsCosGi4upRtV7Duu92n
vAmiTjvOreanDt1ZHaUvp8Ik9qu/Ujy0dZQ9mwV5rubLyxvZDo7Pk7/kMq4AWa87
ymeQ8cljUhgp+B1GGkpNS0WdDxD544koF7ji+IoMcFT+svJJZeZC+ddw5TgUMIOa
VIfinjHITCowS6L+8Csqp0sX2Ih6UKDQBfs5L0+48wfWzQJVk89a71TBq7WmZyqq
5iWNyS9W/k0Dtbw1y59ZTr5ybYps3mvVB/BGDIrSbyJzEn7ZSFMyt2awkjZuClEH
dIw8uxnCc9rZmFyyXWGX2/+FBwWBbApm9sGBMqOE/hVnMS5sA0VL5QSJ6/+AMQg1
aBUpTxJFEYRpS53vDl2IYQklCatAaupwWnFTOFEwLZeh44f9A+L1kyUxZIN8BMHZ
YEZ6FjfShEa4xAeproqNhW0ex88E06VmqEr4QIiVxaNX3Q4dHkw9wiyQGnmJ5yvT
A67Mdi1lr3WdTMK7hGMxfjB9kTrmnY/o3qnKow5at8E2MSt1RQZkRH9ji6A/A6er
SW4of7I3oWR3CPJByZ6bGT88VdYwN7RNrIsHGWc2eIoFEmIPMLckZTenOyxnZFt+
x1OgeykqbaTUp8fybAaIODBA6FD6O8HEIz7uOpRkxkq62BQxp5QrLg9H+LK1aJs4
ArPGz7GbCm7r4mlhAK/ftieUXOLc5ctRBKTDF1yVLpy2wztpeqJ3UXL0Nno2OlGH
BrgwmAE8p2igdcPNpaYZi9MVml+upSxAgk1QfMiLlLny+ZuQtne1fWPus0r8QUCQ
QJ4trlSX1BWEc2dZSvmYTsHyjvvwavc8l6PqsoV/zgxYjrssmDUplGgV2IX4vJmh
3+UGbA7eIrdZqyu4vxeki0mmaA/d9G1vPpsIZs+wZzF8gGbAeq/1/sdVCLWNr3ju
ShoZdLmLkT/V2qWgHwUsfcfxUzjWXjDmdip919Nb9QRwEJ+BH0gHllcVw8Mojj1p
O7Be9cl3pbpjETTWq1BwJREqcB6grOMIlsDDUVM3V/ITY7l39z7Twu19NLzCHekU
RS06j85xI0/Z6Hmt8oTRK/jD4YBHTu6Ygxwc2OKNjmmOVkOr7BFx+WcjqhqKMYRx
zECuhhPpocgXKBobQxWHf2TnGFfADomgmWG+E3bEmg5npiJpsTSav9bpaNJOVFd8
mElD6wojjSs/Mmq6KWMwKvZdT0WuBM5HyuzRLrllP17iFtmuGSvMg7kz/xQlcONX
qAQu9bXwA8sld4YFDFYthKB5JG1a+mj1puJeGmB870i298RV3B8KObZGJUIgs2SP
Iv4DYMrNaEd5zVX85zX1Z5I5Bzw0EpTO/vL7WHLM6DH4tTaYG+LWR+dkNETzqHmb
TlGvp1LH5oGaxAQz+41mdfhIP/RuTkHR/U+MklPwxzFXrE8kWLTxrVBts2BJua/B
yhryT+rJy5ZMGYPiAGLJSVHT/+BfpNPKfXjxKu7C/8I/vlxkB+yAt64EhdzxKrEY
pSQI3uP/p/QkqI/GaS30AGeB+NP2hqCtBbkKMTGerVYGZG8Pfb4yCK9LudCKozjj
E5y8bG51q0YDKRmEZXXXWU0B0vb93RjGQF03p+C1AMrM18NdUKI2QXz3uk4yA/Wn
hqTLivmcDEQrqwKklc0nJLHnzUoFoOGF/pRliekQA+VhfZP16bgA+gZlmdLhayIb
Ap71X3WhjC/5vDlcetAjjXu+K6ETwnQt9bpfu8nFIe/AXbr3BSdt8l6ermn8a952
a6gGwwivN/rb74yOKLCFEQR3iCLewgI80JlCm0GSlh3SOsNgrS4l48TNtMt4A08m
rfWb+BNpXhA+Mv4XvVhPRE1CrdAuNA2+QMMXa0hG6S4c5zuS/TXdjVjt3XoWp5+1
KkrpZBndfaSFDcsEJTxmVKOtzr+LRxCBwQJCE9gN+h9HtRxoH9IG+BLvklmy3VGh
/uAHYMonO9m1xN+32WDTRwt22+vjSjiPbHKk1d6D2W8AJIgtmYh4PI7KJ6xOXp/Y
xqoMacbbHIzC8OP9iFu8PI2mPcgURat3Xo9TFHIb4TGUXp4eHBh6s2D3NYJ8F8ZQ
+wG/oy5X1DID5cNkqGnyAJxtuLPRvvzhBzMkAaMH6b26tsjDoX4Bg1SvMfmMJVoj
M2DqHshjGuopzctQPsy6tqKbuXUZlMyRORgIPyFSzAugq7tMT6VJGiVUigE02WZU
aP5WadaaPCt/0mVExBIo35DbNzSHkMjl0/6ZHET2uE4PE9PzVgF44K9uq9UNbgHj
Uvm/ZNPqTykNs5BGNvDBQ0bPtewmhmqCTn5P9lwFruW04/Ywrq6FhofvPF4G4frS
VLe+lmE5Z7eo4JF0FWxteTULLyDNUt5aFdUbKFvXvAGmZeKud7YRGY8GMRvzSkUc
3Cl68ceULtgcpFXXN4T4R8F/eEpJPZF0r1J+bdPvyQNHyVq3CEj/JCZuo4xyI0eW
C1l0uYHN1oQHPmRyB6vhnHtaprjmsAr/icSZUtCAZC151p+twVAZxQWsTjRIN4o6
ewCy+/6bOFM8fTbKLkMXZprhDX06wMVJC7oaQbkWa8D7LyHJkG55FFyzE5o/XMWR
6RX/ljpEIt/WBXgo7EGoRwtYyM4/f4vJ9xzo0qKQMrvYajj1OqWVlDze+GWahGZt
A6gzsuvgY2MnZN3iB5SbFCBcmoQb0KFt0l/5G2gqxeehlzyxVIKTaovR5DmlM/Lu
zKjae3p3ecVmMA2F5LP4+j92KZ8xRXveChz0hMf7DTTEt2KU02KwTRWkasRo1RC7
vi4F0g4dDNrCktqQJEH4qXMxE1k9c0bCtb0LeHdUz3J0T+wsQ2SgTRUtQnxM5BDU
+gK2fBLVh1/9d9fRCovpiULBQTeswQvJ3lfj4Ri9Et2sMZSzCMJtnQQ/WxA6dXZ+
4lDKZkOtY8Uq9HRRY69Rt1k5cBzKH/tm9SXYH6amdIfqg0RdEXx60pJqCE/UPFVa
1gxJ7GKuq6deNHvcaxwh4Lbh6FOKJylesagT/Y7TyadJEuNhPc4prJj6l061x6FQ
fAeKYYVYVzIIArz3fooQbzQJXqUbOp4MI4FfHkzvI7tGfLzxgj/m8z7r3ZaIDlkn
XMK4a6JOB72g0KIiRX8b1pW771L+hVWanFmNTCo9+f4MQ40l47zZ6Q1HjyVFRhY7
0gVmcZHrGZ0l/RVXFX9tlVnMVsZHfZrgHihDqquxgjd6PtIegXD8De8gO3W25QWo
QidHiX2YfSOWOmlxMbez7FSuDKmVo6TzdvyYLEG4P1/PNW46cGOGLftCJo6WrvpG
g5zFlLkHffslN0KOXu7dcI+nQVIgpVtfuep+nIQ5oBHDdMozNSG11yBfBoNsCLkS
iZ/7ufiI0UsRfLGQCznbO7JWCBd6+HSdkW0+aZiRhWbmA3qoA8+cTkuDV8EePg9e
QA/nEmYfUMYE/5X4VtY904qGikYL9bT0pA9HM6dI3CePY5YwzmbZDx1Mdwfkt9ep
BpGUGFELe99F4zIILywsDGt84LneeXW5YNgr7hWLPGxJveIhTm15OYEbIF1s8QUn
U9Dnscz3WmTcI5usKLTRBBBG4aP6TrW4bztF6VKcz9a9o/FmRMK1+xei+ZUWaUil
guB9k/5jDLC6NgmvXqIKK0sMfFq7MKEbyU5hko+ytGiRaxwYI06XCIWJVDUwT2Kf
jEcAzGHfvoXhba60NmCT8Sqtwp2Z8q9xw3a7NDdV6IlsPh3V95npqdAuJu9BETbE
xxcGvyOx+mPjFPPhVxH5jb5oxW5nOWhvH9sBuvhovcvE+aCeUKO15XYrMqbsy80Y
yeZIYR+UhKurpFn2euoHKSZFC8vDFdJ1T9jm0aV7OwzZlxvZPCQdsFUFx0aj3arE
cBDl6Ry9lByIMd4nTDOLwzA3vqhkoQdypjvmaHemZ2EVS6LIBAAUwQCR/4tr79SA
xivZg83/gChYFhQYAhKGNggnbwHHDKubRs2MTLxKSoymSKopJ9UroAtzv19Qz23S
v/NbvmQ+IJsvL/a6VS30i5aCdT3B5dahEO9wLstB5SWPzaVXHXasmqMhrWKorfCV
SCYk6T2epHo8BeufRwHGgEXO4gn98GHoMQmdg0KzPtg5ZbAjmQADo2l5g5Z4zYWd
9ojHEMQvHRO3Dhr1dzinY87jTkz9bzMSmA97YJrNTj7LMPlSH7nlZmesbexny0JO
Fs2zQjuLDd58bvcWrtni42MQ0Vp0JESbfTALSVNqgtXQXYe6OLc9mQqdNN7FQte8
pLSYPd62bNHEwYKMV0cwtorn7/5GVbRgWqVLw1pE0jUSdM1vbWyo7vQjOQlophut
ZfWybW8T7AZ0GrfShrtAAG4anVYLPHxTVT9IOJwQQbfMK6+Jocj+2uXSL2qgcrw4
Un9SDXw1XRiwaXpE2l27b9f9SeKZ7SpFhOXddeAkKdh1vRNCUBrxLXAGnUDJKJqD
qwN9Qm9Jmau2b3NoZ/FWCjdNHMCYcmDFib5iAvhyLOfw9cWMdcCoGyxx6H9WS6GM
nyHK8FJ34mr30mGpmhJBWpLlnk/+/VJHeBjVA3wwblJrxqOOuJ30YAIxwlCZGPVY
gBTrsHy3Q7iX2SdKoIDzbuSD4wpsC/yFjyMG3hHIMMGj10nmHavtq7WIZcAfJMub
TvjQfL3ksoMQMsSK4dXwx8ACLj9g1bZE5B3eS5uCx7A3kZlQo22AvJV4Sdg6Lh3w
JzhKbqGuA1mJJ50vx6aLvjjHmwrc+wbr5G2fYrnXBS/PdfdDdfqrobeZbBnOkz2a
Qg/UHeqic1QjUWlWMO4042Yykz6GbAQHInfIvcqt4UgTjpetgct9GZGFkj5VRkE8
tqsNOWxxAQeSxrFxbFcslTbVsiHujVJUCpjxxVLrzdpixrPXW1FoS1fDSXyXf+YI
Z3298b6DmIS/nGr2QDTILW3VFLwtC/ae0EBpcHI1ZX4UF7CU2haEdiF1VwkCQZcY
irH051QjiR0fZFUclOdmr6cRPs3GAkfgj3dn+/tqCzxhOtAAjQ/FXaOBRH2p8pfI
1RYF1TWx8CEosELYhDYzUHPsT4Zn50UWvbkMAs96tk3texCfjDXQ/kR6bsag8Wqb
Ae39MbiAT00AjBMvt04hca8sC5R8evZKlvies85hXEJZUMB5eRidyqQMCyNxX9N/
2QB9hhslSmghcFyZL21+b3KkwwUYHaJnmT0lSDHSxmzqcBV0XFNYUkGXmgRoYUrL
YlUzD5h4AbNxd/Tm/Xkgq+RXFFgCxeG8ntAlvHFx9M7Hbuj+QAnLalAgopBDo5P1
V8Mzkdv7b146APo+qOHsjykftYgALSHyASCb4Zrl45VNC8g4IewBqnDHED1fkb5K
j2w23SgMIbDdh9F+3pPVocH17E9TdydrNIX3YvvUwKMU6qH51+Y0Vh4P8IIq3ZSk
wdjSmzJzMWCFn9YsQ2r4+FHgYJ5I+6j51xe6S5tzVkpfMHW0JAcXLvREFtbr8HHN
WLWWb5LiBuWOJFbnCyDExM0BfXksb3d3jGPVdLZTNATsho9k1+2u+a8PLBAONzhz
cRWQpsA5cFmGVlmO3nldt+9n5VPIL+VyAbMMX+sHJREvowEGI1V7h+0VGbPyOJ1I
40sycOF6FnXf01mZD5cylll1aZSiEE3eJVNtSoezvqIW7+nc5Az5y72C5jABs/ri
JDxr3L2gzjTs0BLf3ZqMPAetdPmmt3qgT2AlK9agZ4NOriYUbeXcuHgXVKO/2YqK
wGRJF3ZWRkmL2r0ZTnTKP+QoEW5ChG5w1bhiZsDQAnZyT5sKSmC1/QX636/dg80D
u3QDEeKNtatVqyJ2DarJTHUpvHgYobpIYav2yBkkae2+A3//dIsQQuTLlIWETWSW
kZ2xPH38+xubjUFtj+ZIj/RPjP43pw+KczJ0zrJfe1qvyqCkG8JLn+392fwUfw74
Q0vqwdfVRDiuy8dw8DJ3sDAFGbsff+T0udxqxE6aS41FYHwaiiBaABtDXNR7PALr
/MbrFKG5JLgK77gR9agEIaVWwXsXvH3Nmk14HXcnZGgs3l6uDz21QpXyjzEMe8Ss
Ji6Qtog4QRPIh4p5iGA0Wb7KfYqpyOcPPLi1ko1gfrGMDooxi9IzyR/tSGFlYWs8
KnOrlU0uj+06XAnCQcmbVQdnxDSm749Kqku/J9filAgTEs/pm6LNbgKUbPH3TPgN
vG5bycFL46TJZTP88OBpHOKCKhKFBoAwTwrWhdoV5S7JzYxI3VyFWNXwi9kkD31q
OWIlu439GmqbeWx26tiDLnrdQyK4TGwiAF/5sCk3eCIbzUbAG/Qv1fw1irQYaPM0
sloEQWx0/551eYX4uxsjXzfjI8RrgT/2xS0+kZlp8kWEoKc7gLniJAc8HWgwQTSS
3j1cXkqkSm6kak7Ghj8kEz/f79FAJThjShbP5lbEuKjiuL3nAdXUp1wU5Z6HdYMU
JQO02dSRNg13LPc9a2bdqKRiPc+UKinbJoX8XwhVwRmg4UUa3BFpS9dpbJwcndBc
so6vn4VSKYUT6xvnoy1oGZ0n/O5AnzEse+Zx+l/pxW3LW0bhQMcDPcwTsv88NUXN
2WgEpDuK0dTWPEsfPlbhiBkD0zW3CFIMDiyOAgfvXJFzAfu1CR2S73zQrszTYRR8
yRA19pzA44cg/LvjfWfQduSKwWQfIyjcr2WmjhvQWlRpVLP3F0xOCjzMWxh2U27f
8dNeLuGpQyA5JBU3H5P7LN+3pEN1KNi3Y14uj9tAfZ1bn4GNOLKdbFaf2MdnAgip
khG8odoK4XU41marlM3dRCoRlNtpiz5/k1ElQh4IiEAFyFj2Q93DSAd/mDOZDpQH
QeiZpXqFz8nndwbuFSwhOzZVAUxrx3F5VxtWtbbnqaKRWD6nAIYHtZnB2kVdEjq/
01vU9wuU03KrrhzXKi3jF09N+/VBAJQ5GsZstEsCyB8bTQ0FC0CLXyeOobsyHkNO
H9rvpOUH7pNQx04r7zLDSIBFGk7u8n7E76Ekith6//BPEKy1Cjxy695zPwkoKFPc
31H7GOmMNmwnsIbK5PG9DqK1Uw6+JcS2PrKzLea3kWGirTw6QSxf+Km0cpmvPJv6
7ZRCyKx2+GzrRld7Lh+8gx/+ihPiVhMEECzQ1x/hmPydOEk9Zlv8l5sZp8gEoCPd
shppm23/ismTbbes3LmkhUFcWjbIzIZRASU18lpc89lmRrssekTrXrPwOrtsyWo5
JC2tJldjhOIKfpWkiTF3wrAVnJvmYjOd3iX3N6ozjPpFma+zmtQl4zo/BLrdTw9v
o50ltgCp8pEY1zXgt57SwwXlZgsHbge7qHpcM7Qb4viei9LYFaBzbObziZVehSuU
FNpw0b736bqXA0o7m62JehO7WCSRaeiTKGx4yk+G8bDJntfjcaxLTgCFiGEFPoyW
pA1foNTSoS6SgjlXbzkuV82GD4GLORbbflPasgMj0+AL2on17QaD3cOAZuNL1BAL
BFoKL+n4pfNu2p61WOxMLkqsZrjq1O9/89i3KfLw0u1uRaeKD4G7xSrxg3AGAKBC
STAWoIS0JBdtU2G2DeD1lL+9bFuwAtM9Btg/GjKCTQXNRTakIWv7WKa6TjtOhXAU
atwMxvWZBMwmAHOZrq9m6PXbHSZvJvUKmqr84a1f3BVuw8hreRiPf70XZdx+0inM
eU/5xP+PLqPJxUxv7NjnvKlqxnP/Dw2A+h9eGvK/aPdZU9og9LbgvfCmDWxsLVp+
YGL5zVhwa/exEpgY7h6roz4ysV/gMRDCICbnA1j8VMuPwaOND35z1hE9L/FPWzJF
n9VFpp+f4suX6Z26Aj4vtrq6KW4M1HYBPHq3MFcSP4YEAXR+EGKBzbnL9kDsfFzX
KsSXxH0fIV3ft69P53qYAmloXWVvE1wkIZQCHFduFjimWKC18nCzhc78taDppWDq
3Aw3BkMzusKcHRmxaTG72FRfsEITp/9OXqhOZf+Sqj/f3QW3w16BJIf4avHTuTFd
LS+l7BISCmVqh/JiZlNmri3qufPSjTxBWhuxxTNjd4QV5Qtt+LcM5aSAOkyjVl4R
tEP7VeW825JQZL6BtVkNDRiyXfVe7QcxYQtOS5fGwaIYmHDLO7kM0KL3UUCOK9nK
+RKv3dghONQTbWvpG4GsEWqHIxuK2w5vlsvIvdlrjQs4eMXvAN9OAVX/DczRlskD
RwWhy4D0EFh3kxtrrC0j0xFTYgu3v01GE89UXeIA3KF4XOUKTfpnlcAXMrsZVXu+
g7b6W4ympRzMCVPC7mkZUeB4zBgzVD7r6KoEJZtU+VfpH4BNywLMbFk9ls+5ch9F
sfUHospsMUyYAZ56sLnF7g/oUk65V/WKEqJNDbeSh+s1C5yMl2PUfTKdxS/nS7Wq
3g8qxZ1BSKLv0rER9yShNrulNcoe4oVDwprp4THeCZz0lPdYjob49hRzfAXym8rN
6X+BkZYJL1SgkVRdDArdY2Eo3tYNAUEDtQqUtFNhaS9L0Dl6hsQz5fGGIRM+QGKj
45ly5t0lrTMvPkv3OeGoKun4UHl0vykCJw3o5NuwMn4T3cEHjuMyJuAKRPi0TdRR
PGbcrqMSzfhZK8cjYceF7rcS4i7DRbrPc77g8qFRRQlwFW0LPI8fNPDSlCBUE6zL
iEfR319YF14fMvunZ4tuoUDcfWJZC9V/NPZHkD4V6qhNVfjMfLFinDDJyQ6pgsl5
BATveAOZRTZ8dppCxYWiQuy2AQ3p/F3IJnvuz7IVE6Y7s/dZfGvlceSCzI891DBa
fSRyOl8Z6laDEQY+c8Xuv+UNPz15LYb2F5o/uxQEp2er/qe3xy5ZFKRTbXgC/PKN
2GjI7I9AAon4sXXrH3y0D+bKlAFsYmDHC3XONcakHtC9BUbSOrtlK2ys4XdaGpiO
4AAIM0Udn/hhq/1R78fiLAX3Zc+x1ygk71TRPAP/n0TlQ/Xg2tL+JChzHud9Nc+a
jeH01yUx5lhj/gAElT+JxtY3qug+FJ3N7kpf+Bn4eA6O6ApHrB4roNRDbqRTE5nK
w5bzAmFhoD0QaEfE30c5AHcXIsCINaNpUpHHegxFZdeC1gn616/Rpf6AWbvou1hC
NbZaiRaKJmnCWZqDkAKtlfTioJceqI09o93DFI9IYmyTPmFhrrQ16B2JJVI3t5ee
RT4cRAHpPUjGC8JBApYSPY1jyh0u8X7iZwRyHtl3bt1OnR5wVQl1pC6Z0HZ0quL1
yzIExsf550XzN0qsgTkUOj+V7I7i69dO0UpiCv67VWeMriEYR2bNHOaIky2PM8xc
J5W0R4um1IwrrHujQaVwReyUS+H5xWucYEfiLmgr1uLt/4WJiWIWCh+wfJUMvUQg
owP8esrG/Y8NAvtD+f400hkI2jO4NFJJsMhOlbVV/JFaHkamm+Afsd1R2hMRmU4+
qeZyvxaJgwdhzv8XPl4Sg0oQqMsbqwRhayfBSeBa91FW1nuslj19uoAuZKwYs+fi
`pragma protect end_protected
