// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:36:58 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
rUpQVQh7tPMKzuUTOBaMiQR3JgjvfuPmFDY2qwPGaiAlVnbxHLhvw/KHpeHwT3wr
Av10ohqy7CvgLzYW2/utMMDre3gQqWlDKmzY4CI3tHLZy0lErIUA8JkPzR67nNNV
MO4rVPcNi6T+cUm6+WTUGBIuvhy7Kr+EnlwnsgsqBPk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8256)
IAzz3z4edTS0wrkU6bBruTAwJA2I6ERFL5T8k30twAR5OLxVS25c5r8d6TOTaM7u
bPHV6S+JYBGXFihgJg7vnILgyOgnX+5VZKnZSp3MMlTwlqFHPDbqDiwA3gLIhuP6
2wmqzpZb2MAWo/1BnN78xtVBjCsx9g5d0HugOwm2UkzLSPvIOgsHoe0rdTqXoI/L
ws4d+/w4U8ftsRA1Kg3KT8ndUYDGeI30DOYJvPrQqPhtL+XN7JbqdbP+oiAYbV7V
EZYWx/Vm6W5M3X03KXMkHukglkmIjyKDkvfM0xz0snA6qhL95bpIZ4l68J0SX54F
PdzvArOYC0b8qHBQtjOMpxVSaHNPJCb2oQBOhc5xY8I9dQnUu3L9GQdpB9oSVqIr
T8lEXHzPrK4gJ1Y5FaLjrghS9JmyK84zxrIRJK+hi19WxivWbYXyJqtspq8aThfc
NvDLz7qlx8ThcvDPS9EJO/QZxTT9uEbVzbAm4O6ss/0j5mN6usYsuVkVwQ6uJLfz
av16yUlvvTnXlckbdjoDMC7S9TAOOvClcwjkzgDgGrNJXI+5cENRD0h4kXfQTrW/
9POSdCbBX4EgD8dsmAPl6WZEq6eI5Vqyr9TUZFbcwLiwRVhlx0VjVrIK+1UGX4Nm
L3/CgtlgaiPmV4iCq+ASQ3bdQEOnvYrls3mAqZZZBP8I2HjsGBWDAdS7PjCk3GUp
L/XcuN972hCgG+NVmner4DLDDH0jVcP3geFwcgFVXrVYC1pnopqavQO07KelT0ac
P0+Yw4s7aFwLXUSLHsYIJA7UB3UfGsEqrYFgSDH5ZWmZg6wqn9XXCPkzy2dBfC98
y7HnSk/aJY4B6cVSLMCjsGd6Rs7/v85Fisa/cc6oz8swvEuXbc4RIiSz7I6V9LZq
QKrxxFL6UOinW5i+XXQ0pb/a0Z1KN7BzgxAiRAYcIwc7152USfF6YZktHRDh2WgS
pcH/henSATONE3UGFLs83HnFfFU+F8wPStZqebV6BVN1PDNCpTdEIQV/qGbQrfKO
5oJjZw6sSB1IxE4OuuFAzBeaJTrLYMpH3io2cR2O4OvvWBvanRaw1gsUmDP3mJVw
W830upl1u8OOkcTeIC7zsb/AS9wt8apVMjxpMNIhr1SLolgHX6I7j9FKFazYCRa0
snuYgAmVG/6BYoFDel/vAIq2OXXugvIoXR0VQw9GDtemdXTjoO5EaKnoC81Sq+lu
0sGwp2JJlBWNBvCaXz/WJs6Pspkob3XyUJHWfkgp2mzM0HojDConyZJDlqTtqsr4
dIg6aL4Mw15Nlrd5DZEGjrR2W28dDyEeXuCu8Dfv83c1zhnoQ2/CblljhXIMCUVJ
/S4fASPqVz3PKDrZWeQVlNTVEumNs2wIBTG8es1VdolGEJMKYUbg3Z6xE3ThJZS3
Vc0/0ZXY7FZDWWyLSMPmicUJby4oh8S0EiQlD7c9ae6Uk1kEMSV5chie2OlsEtBj
32cxreuk7q/RX4WUQoMl9D2q6kQSzzOwSh9ssBpmYoknb7aGmNKHwE7rBgDU2Gl/
VFJ0CGqFCIXNLaSqSgEVJSFrTZGg/BEItEIFP+CbJibd9Pibb2QjG/+LCNzGfipE
0xNUcSRu4ZB4CNldk6q1iISe+SlUV+1DOANsV1687O2KRfv55Er8tuYgm96s9nUv
CvDIY9Bl9AmtTv6KZ3MyiMsNwNmbEKzIHsV41Iw7QdCnjy09qa3AL3fennL+xSxo
hKYzJtvVPkZktxGePrfMo8QsG6Ma76vCMbj0HVBztkgBmO1RY+UbKHI7CVOeprYr
ksgNKtqE6ni/te4r41ydNx0Tu5AJv3YzuBfNgkRGq3TAQA6m06spisnC1ewrq4+9
Y0WSCE9NJHZ/BBE121Nnif3hsJNNULMcD8U7bXn80HZNlwjJREzIdQLJxmxja5xj
Z6t6OD3vlrGrzrDK7e/+psSUSRo/ip2dWyTpJsgM3l3PUMFDsynrMNQcvzGju4+2
F6/cPIqnGpwgMecnWaXtMY4I4RxLU7oakDeaMpmK4Dm4zGjAVphC6xC1y5Gwvt0a
a3/CIrpQ1MJozVTfqqAiIk63BGOSt5CYxgRVET4UBDGrYJ36W02OaU9SIMHADxny
qns3nS95DsBvt3fdjosB4P4KHjoP5cyK13Eq2czrF8mniMKS89cj6zgBPA9MUDwP
uyQZWL3dnjpUiXqISlLw45b+XdiEMvk3GxotLntU8FRBcpXWrxT3t46SeNlm8wKL
WirxEhiazjJEiHJN29IWNAkHhsw7/FdNoJCDaRgnDiHDNymhjf73SUHnXFFAVbLA
tUWLrvAekdXjBDnxkGYIPAXt03IZVAfowcCugWNgwCBar2oN5Ksg6cBYJp9BB/0N
vsBQtxJQtabbUZjPqbQTXvTR064VeGxJoFJ1lQpuEZuIMwOYzZ81SEO8ngrOsDlP
ywO0czoWdS41sJ3YqOL2l7Dw2U1rQ9YORi0wpd5ZJFnXZYLu8Xf4RLSGh3ikZKpf
GrSF5oDcsM2tDZ2HZRh4aKyHVC8zMTHzrCscbj3WTUiFZenfaVg3l2AK3PHx7A9L
mJGM3YpV1q9sXGw474yD0gQkfHXrZMjiPEuVY4iklPhrvVlh1UnTzVR9Xa0Nvdkq
TewK5dx8/J68Cqb1gDsn0SYBbJX2ioWfvwKzcZxoSVXWu9RXyRDU6zcy/WlTMCiM
ueudfkLVT7AFeaeX0Ep3aCKMpIpmMYstLsSOlNm6dPBsnNWhUyCU9Ym4jBQEPqgB
hfxCEItF0A2RyyRhMS7BGpJmc7Xv33w5x12+8CoTF7MbCQ18ZVXNfMOaZeh/hvHL
YkKiT7RWwaB7Iia1N3n7UrOc5x0R6apQKZhcpg47oMVnvASO8juUT6meU+9xRojn
8j4D+4CuNgoC2fEiehEIKSjeZ2zZUZIRzSOR/magx3k2X7m3m/3hVFJhQlvnGsoi
1BUqtgOtnP55XSsIxmpH9nGRadKMqFNT3mG5Tvq/4MhD2o58OJmFwdegEevp7gLM
8Y1hQbVH4wM1mDClsyag5jYsS0F7HMIrl7MbSqZ8AB+nqMFTiYes3tymS/NttfGj
81xhtcu0wTvg/e56hkXBUMpJBuD0SPPGWAsjxCEVI+3kgB/2fuZRvgH78f2xqDXS
lkDkXy7eExRaUpYElOiSPGkUdx1Us7NxtNTKILr1b3k3fpukWRXoOkyH1ZFtNs9n
DZJPE5dNy1zt3TAbwxaFyZ0oTwty2pq5Hu0q06tSW5YQcmajHJx9H3ekhyQ3K4i/
cCAPOJ9JMseZHoz4n8HQvUhxm9yBrz/eCQY7Pmwzf3U22iN7F2Ky0oIZhsAFiDbN
7iX8J8oEi70M4/3T3P/RamMrhabumyv6MzaHhSP3WkICu/RQcj8TYlyVxLM+tXAe
vYPCC5bwj7B5qKWd531W/de8ORR3vxGdpo6trBHCVhRrKq5l57cXVmcoM3DTPXV0
zE7K//4R6pgPuewo5/Ha4bbluwAUvPaOzwv+0dVJNxelJr3cpLnOlbCoBxKamdlt
4N9vzJglPOgipE2DI+uEQ4AoLVUMc0EW9jQw1ZeypOipPPAuGOihUgR/nSVkByWJ
qmjUgkTd7wo65C0myJvVp4jFEYwZp34jqHicTmSWZFUuND+5xx66gT0RA350LGST
db7qhLr9xYe9i/AL5qVTfe8MZ77r6rrugneb8Ss5OE+zGMKMQcE3HGuI0vTIFctm
cKlarV4uKqn4PnkVIK+S0x/8WThQkXf9vMmIln7GGlmfwjZ28FjF7vA/e/PSxYLo
LQ5zQC5r/v3NK5b78qe69Y978q+ixmlqYRKs1f27vjoC+Rml/jFcKOEYhKtTQHl4
p1J0KcaZ4rfehS9t2JSCpF3qAO6B9YWZTkJy+xieboHKFk6wOAJxnOG3ZWmUqP76
93WG4CNRF+AvYOlZ4BokE7/c1oq8xxc7UWwy6ptp3Sq/+ZYqP0f4p7hIGG7afE+/
OwZcWYH088HfPvkXzorHcb4tooNh5sOdJIY+bcO4pCfK4lhiV7peHQWzyuxj3XmB
19mvr6s9xmfW3r7M8Oxiy23yFQnrD0TgmritF1Z5CWLVzFN8gGa7LxOUXutafs+0
tnI2YHoYbPcPafMBLxFR5sxUQiFk5mI4QrMrK1tUj1kGGyc57gBHCgANvr5GBxKh
ViYk7+wea1vNAjtUj4AmgI5pKhZ/F8mV0FpiLMOsIcFvKStWokkaN2PggXBSxMV9
kcAxS9K+jsedJrHOB6VhLoB8L84MmsARDyuKEZ3d4xfQqdDAOpS6Ax5sIUeToqP/
Zg/Y2SggXztGVNHXokFR4axyUH55YKZ6PZQMuOUTKopptXiV7CnqcozzzTLBgJlz
GSq0iVFLJaLwO7RsfikeSvW1CFOzmtn4NbmWXQHBrXYlEYzuLTYtHulJwoftXANm
t3PGDX61DOvCQMyUNQYnWpOrsnSFPPf3j+sBit8dNuMJ2txuNdMGMTJMx3ellEDl
G3sP2wiC2acb36TaDKWVdURXxIL63yAVQ/sZwAZT6BiInPoaiyb6VsBQH6Cklrp+
+f/Ip5EA3Ro9Px3wlRdHg460zWJh3EIk3XpBXUXk/6OHaytRDRrRWyheqSkOEgSb
YF4+R8Sd3VxBj0dxnl/4dlgR2tSWHxLG1jwIHCx42b9hX+qFy287Yfy/9ZWjI8Jq
As6+zIG7rdYdBM1piwltPTtm4jt1no2xFHuAj5xSQED6/qtFHrMa3J3r//JlaRt1
HE6tiX3cnfnn9PL1prUj+pVsR7ZnCAaliIY+Iqcs0ri3/yuw9FbhuFFx+G4hks4+
nkQaWQK13rELNIIQnvHmmIBQDpkj5zdRYHidsj6v9g9THIK5two+BmBLOqn6Liu5
sKsPXIMlOXCL/WtOUw7MQK8+dHk2034jaYAfj6p4ljQ6pOSxPxSPhvhr+WCEfYiP
rVyDqZPddwZfG7UzpRuW8pzins3iyWYhXzEiZq3U6hC+l36dMEyxfEvhKcqerKMl
AJfGqwjAZWq+pyhHYMxoktk/G7o0IcYUNERL81E6FfNPQ//NzsvavdcNzax2GTBQ
18QNC0HPYhAJhwL6AmW4zZtDO7takgeYMh/hrqPJlnkHUYpWgaK59h4i+VtDTON0
OZHo/WRIBjKxhiXJCKn3KeNqB+twn7Fc0KS8eRrh56zblYp8noJ30cKqIS40cW2v
vsE2Fju15uT1Yx6bTfiasNfsdjbFun4T+R21T5g65jdZZARIZFvnd6IchTbFOA8o
yoflF3DpyLEClNchoWhomozl26XsaAQwM9WSKWM6Pc87dn2EqNAUt5ECQa1Z1ejs
EYrI3FhjgZgfLM3EwwrCZItj2IMb9EJPK/gChmSiKAo63ywJBtyKP1xdH6QPDtPC
CfIeC+P1VTS8xvZoQMn+ur0Lw527Z7sOCFsLDNbrpvW3HN/jAKr++fJTotMXuU/v
2O6AlDZQvJ1QYBVnIPlM4pF/VO8XIDFqnmZWamH913un0PJ1RAp+yG1tdIhGtIO8
9PQ77/T92wNn4K4e65fWryumr+hK6ELlLISf9sBtuJ00keVZHYGrZozmho44Myxc
gRGdIHiotY3xIPXLIgrBwd1Rk1T7mzFgeqAm3LsFMWh5ybF9aPtlFE4uK/mrXIfL
3xj4NZCyQdLHVCb6P1n0h1MbO/q3vPwsXjeZTd7Z8Px3Om2haclR33nBcQKYKy5y
SLrxy3z+uK8nRK2sF/PeElUJ9aV99Kdd1w3qXMV5jJsn7ZrN8mouUwK+g1yVh9JL
JOJcFjc6rnFb3mZIILSwDAE7R38vUjC1akOrDkE7zmIeTex/Ba2l9LXI/aDMk7mA
yzfc2drQmn5krR6+DlgD9uFqjCczMjKsA2lbntDmCFXkZHLHdmUH5yguYTOFNeik
04Etzr1UbENKFHQzZByNGojoe163c+YmAFtvhJYzanJtV6iF8/dODVIBvosEoaQt
ioqOQ8Y/9lxTXchMcINgMZy7HDA9oMl9wHVqnnWrtzj9VHs2ZmS87IT4b/1ljSvu
OnLftLs+YgTRdtDkm2VjAYUJ2Gh09D0mmWVNZvI3vdfTsfYFGIWXw39PuOIkwKv6
CSf0rHSRHVvRPN0BUA7yDi2g0lvWke5y+STRqE1VKZlrMLbYZjpkh+dmanzuQuLM
133BQuZ72UD+hqa4gfzfZmQVFqg7F2yWmYgsuGXO9QorGZ2dotIUg4D9mTTltXWF
vAb1skETgflXoWKwvWN59yC2uJK2K111kiqUR63PdvkUR+SHOLZra4fsP4IW9wS1
nwK1O707IohYkMi7X+zcwT/WQPxR4AukQirJmpN2OeeeAyDi9fhTDPD8fXXs4IEe
78FChw/W4mXITNnPxQ0GrvJLDLD0difC/vhc/C0xy2TT91xvUNhNe1/49hkxD4eS
ysWmfx50JKSuQ0ahgW1QceZVm1xSMJfSoT/zHQAjafaX3QrDB9ctPsBGCWzpC9Di
PX5BBQrq/Zk+lcTJhLS6jfKogHvxB1a89ktyr+Mp9nu4EwwX3ISJOsm34jZaznll
JJWEFc2Eh8zzGM6jAxw74QYgy/BE1uZTd++f2+yUeJoOF+fu9KeNxvcdUWtFtiSw
wgKTxH0MtXc6j+N+hG0vpaX3omP05eiDGvxRGW4SchaW15sb4I3sTHE7f+YYbhUM
gqxEHVBvOCCd6WBTBPYCjgJzOf6JZIleHvlfZUzKI3bD/Pu8PY4in4O97YggtaSt
3eEceEQ2E6bsqOJaosQo74kineQhwUb1x8kanGqrirO6MnhR0YuBcWx3a3yVgnYh
GA4UA7CbKhsMd6ITjbR2487AUfLSQjuILvMrqlMBQqAs19EhEhLQiy92MpI7i1y8
m8rstsQAOJf1hHlregXbitlT/Gz+wPMBUnrttT5wTwwYNV0+oFBKBQzw/vuUdbCd
5pObOYArCnuEkYLkSsv693E0bRomb0jylFmTbRSw19W7cfLSykAfIa5hiWnjyIDs
sV3y+W8NYA1yJSPk6+IkVn2IQQs6HuqCF3qXG5F82jPm02Ock/wQB62uB9cXNaOu
DNzClLxLccmTK8m/fJC9S0TJCYQR9MRnKMqUuhsMkK98o9RwseiWwXDmDok0wW+R
divGS/0P0Z+ZBWkS9BkiF47xmXlH0CmYJ6R4XBxlOk/07R2Ysh4mqytI4FjNOHE/
th+jVbA9Q3GAyVs4zP1vxw7PMGJ9DRlIE3BkoagmHyM1R4/1ciMAI0HRQGuJon7z
B7//FidP7xZYpIBUUZODqqIVk+otri6syEm5WN2hU0GCv0aJ/kSGU/V4WAoB/oVO
LKE/YwdAcK/B/uxHjHal7RWX4P0LXjwMx7hN4aZQjBHfUhD8jX2IUqgck2poyAKq
IenJKF+fj6RS0LyVtUNGMriLMZvALZZlP9th6SPdQreyoc6kYgUeukigSWVFwrnG
tTiAE5Rh17gPrddkFJJ29neBtmazx6YObp7LzfcuBTIcFALkqrX/SgukluK5KA+Z
1XbGI0215HRQ/53+Sy1eW0lm1Cdk6p/+bdaUgWRvdvCWYy45zn0OJt3e7i3UnF3f
OdbWT1ItHbtJSHbU7k37PxYH2U4d8rO5YXVl6AfVmxA0zxyn2vwX2giGdNbaPNyz
oQU+WVSD7RkFmZaB++Cq9Uh4kg+rLF6dVU90srxWQj6cAndVvP+98F2oyMAf5SNN
IiRM7WQxPKTEXyNVOl9yV+Wshfd7udrR92J7fe9tVIHcHH2s9aGxTTixBVF9ni9R
Ddl/DFLJSHP8HWqygH74+JyrdwuD/v1KoX+H2DEAFNRcmzbNQWrQj9CiZtX1G8gv
H9bsG0Z7Qnw2zmOAszy4pdEoFCzuqNLeN7cGlYFC5DUBkly9ul8xkahVRIr7vtfi
C6TwIspiiD2Id1D1I8vCRr1hnG5qIrrFUcj6KxmLA2aMQisPtHv4YUcRQ5wThhtf
mY5kO+A3CnFmu0WnfPXialUfx7s1fIJKBBjrY0tkjQbA/j5yxpAHoPojF4hfH9Ni
wIS4I8QXubhQ0e0Yoh6ODMv0a/QqCku4PRQl8MhnM2x+6Fh8ISmQQ3P6IEQKXy5G
SBC6VE8wa5+Y+f0SCu+YxJj6EvfeiCSgIL1Q/MIpsy3JOx1+pJDzrra8RiEiB4ht
BtlIhMrT7yCDhQvIafwb7XMdO1JJNlNDjZsrKrcUK7iJYYyghcsi9Qvbmfp12Yn6
RHoMTruVAmerJ+qzVhpMElxOFwKIy6zZ1yrBHc6aAseskyQC5TAlwHoTOMCeUKgi
4MpZt88li3RABPmLZZxiSJBCQSKv2qgmRn01cUQxNxj6UPGMdpm05TOWS3iByHWi
zvzFb4udrWFeXyfUIeomWQqi6Ne4Upu4O0Lp10Idu1egdbv3qjnZy2foiLTuwUHQ
oPZDPOXPgNaBunXQxQ2FDRrqrQWaYVg7hVW8Cgi1ajEdM+L3Ngn4XcOHo67NlppW
hawd8IVod20Pr8hKTaL2E8tr5XuCfsVBFuMKbls6WWcjOOIkCRNagW5t2Vmeihzv
d0kxk0IgeI7yUVuS+30ijXCSR/+fEDgJcxz30OAiFvNqVjNi5I0q9oKKGMf2q2es
HwQ/DQC0VpthYULdTG676we4m2ZfWtIxMZUtRr70YrT1jnx7n8/trOln0UDuKgpC
YKu6zQJVyzhM4d8YPfPUc+mBVKM5yfhasTprkcn3rueA65peMpe6bujrhKksL+Ff
waox+tOdG9qQRz5UhW2cJrHyPQDbQ19YvHJlkmuOJIcm4P86JpL/Jvdi8vVE6nFa
81baR+9E4gb/V/QkkgOUp74kFODUSLfe+Tj7HBI/tBDf6WgW+rXF+URIT6GHDpxb
q7KdqMELPDkG4i5REgaaiNDUOTj6a2yMhrCFMqyLqAEeyKM7HjRrZs/T30EMQCBU
ENATYx1ZPUr4OqrsW2bP6SddajtmZzYfklI3zIdHqpTFxvmjdzEaCHoe3nLyrXuK
ov0jhgFjgZxItopSEXa6sI0vGT+oZPJqWUD74twO3/B2SKeFiJx2bc16xnES2VMg
cRrOK6GPVdDj+mFl/0EcMCkqjX1XtWPcL/r+tyjEsJZ5lSpwaH2PpDHD1tI3BjX3
XtjYH49y9FxJUuqQHtglLnXrgnBqEqSYMK+ugn+PDaMyXlDOv94B+4bFZ4Mp2iIN
U/fJanFd45ColqggPKob5FFuPHZ/SgGsxIguuupIq+Re3Sr8IYLSYS8yzqE42IDI
TkMm9uUx9zQnJqxjxq7Tu25sdEcwUa5T1W9ZryF3SRlrBiO9a2YqEpJx40uWwpFE
MeiumSayd041SSl0GpZ5YxCow9anu8I7IIX577EEvUQT+qtwUQe6b5qHnnygJbOU
2M5W4eGKl6FIHipa99xCHlQ3n7g0rE+py1cYZQBPHMYVAnCgly9ChSRwfQo+gJfd
NTnTECd5d1hGczWV59P4DzxF4qWZseAYf8OJH+avw1wltMfitR4cPKbC0cti6906
TdcPPKMpeapQK5mMNcGc4rUsehSVqgoRRAtVsaqKnyS1ka3FD4j20HsyPy1iv5Hw
8VsQLBPAhU4Bxzdw+9ZBtKutJXIDJwtpS/CWvq7EexOsuwRtqv1J8DwfAGzMYrdJ
0ijG05e6NgfjLrPohfyeSZERyJtTXQZP+bbVhjQ3MiGgKLul9byd5+V3fMnWjKl4
upPpqNcpdS4a3rwq1bwSvr8qms2WjdyJBblrPhmjNrELbZHJVOZz2mMZT4yJwYEs
stncjldZ+LK6kU1BLw3zHRsUHjYeqZz6rsWf4JjNfe8yBZ5z970yPftLoTTr5yGJ
p2yZmNWCEfYfYoVUB6IX+KhpNdCcGOpV3FnpAEfGLNm3ZntrTvfXKwQYnle8HNG8
0pCTPZSdUG2UTQ84Tn0WZQT6HzlVm3wWj56kJyQGT1NFJBwScxHYWywWcFlfTVdD
nM40Hf8msRqP2Y2OJ7m0uifyltMbYpi7j3l3aLuiCwkR2GFoLO8YkTnZREQ6+6iU
WbgGsBUS2A6RfJ2a2aUUwO8U4CwYxSHrz2/YWtdHnFPM7bwfyuwhtx6J9ENp+c8V
ld28/rREvrKAzvvQtr+gzWhCgAZjhDSmYpyMayX6PMaLZibEqmjtqzYKXWesZa0p
JADyYq2orYbw3f+xLWMHAGH27VUqfXmN3xjxH+20yLj/4jtkbZJmhRM4pAJpPZJm
8M8VNjDG1peqkYr2yfiMBlTAd+y+x+NXfKDc6d4beennAxyAe+tbAcLPmzDGpk+g
pt+jCOPeo1Wk6SjWIGdMKgMch7y8OWfOYo6RmgQlhx6uJftjWSYiCY9WwlNebgIP
QNg+T3MZfmlDtYDOg+gX/F2wd/+F8mzBn9KhUeNDcB4c1YbAFpi6V6elt/j6woxt
CZxfY3lW8KRk+b9ZQ5rzLbQmn6oNcAY7nWuzFCErk9ZxNqdTX/IyO6NjZOOyAQa2
MvaqcAMKl3tj6CvLBYUh/SbDcUHfy/J26boA0GdPJFHdnSOdsO0cOF90/0Hu2w8/
TLvBZyxYhIL5n8QlhPs5yTGrdP+/ZyDl6P2C2DCRStPQ+G2HVNGlDJdtpHKzj+7R
bOf8gCl8c2vbnUggPbp3iav3ox2w02KrLK96cUTu42Yz6XN8THu0prK8zumVd58i
leRS54LDj7htF6Pdr4aNu4rUxsyrjXc1AmMq0ScU3FKYBa7DQQ+cISoWeMZbsu5T
P/vRv5r/inTbXk0Hw85fqC0jGhL/P0SnVvKvRilWhEUpESv/NCsUrz5/nLm9kGR4
XVo4oCrb3ZWwVHTuGYMH3tyfWdFwS+5XnakPfg6Wr7MWLMUkskCCh4FZRDHYA+6r
ODZQh/IjCuxd4mWMGCB7tVoJ/6kBBKEko6uWTa0W8s+AadKZm3EpWQpX0eK1s1iM
an6bkPiLDhIrj3t8f/76JknvDv9vyyxxeMotF6Dz5CJeCZMYkDxWHcwRAfQhHV6O
TOUqgpv/gwHyhirFoWrYnYsholS7CCw7Y/inBEZWw6s+OShA4CdbfojeAXxw8ncH
`pragma protect end_protected
