// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.0std
// ALTERA_TIMESTAMP:Wed Apr 26 13:33:37 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Em5avxCBLL8I4twdNuqmiZx7UWP05Z4imOWx5n67B0QvA2eORa0Q5L/ui+DEH7Yg
TUg53sOBqe5m8f3RFX/KMBIoSiTzN5Wu/m9kl/msuDKTrpwHbiuYgbLqO61p6NlN
vrcSkzCRUJmRUtrtLD5Z/Iz55NwhQZvx5IE1uLwUQOM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 30832)
i1URI6RKBAjWg/dyl6HYO58vIjvAJdPCy/UpVx2jWrcNZwTELUAvOcEafJ41ETQ/
bPD9Z/S055p6Boc8jgvtoxJQmbl58pr2bOeXL5TW5eZLpWm12E5cLAW5cIum3z0x
w2JAVSrvf+zwfE1YFVknqxxxR2LmHsscXyiHpvjqCqp/b8DtFMzrOrPQpIwA34cF
j+95ZFudzhZ6LywGioHw0q0a+VfT3ruuwrXjX8qizEpGYN1M3oPR7IQIYnOZjhFo
S7wgcCgje3cgmH/H5yuIPPrHy5tLr83hF0+FP5Ry0w9Ba0otaL4AKm6M2Kgk1GYN
skjsmaAA2RAYciqGvUDZlDSRQSqoGEKwOEYQzJjEafSUUG7Z6ZHOnRFonqQoi4kD
iafWDAITMro5d4V6iZd+Y7v6aEzaQqwUSyRenfqNAWEtuUipmiGTiS/IOvaDyYi8
DfFz05U4tDmB124sjwkYym03kTRWr/DHxsZn1iE9C2fg18IiUMgtbVxdNk6ZxJEA
pQmBmjfrbcFi50uFWOIvC4/IRyAXhF3YriFHHFHDluQh0tQmJFd0XTjs5WdI8Ivy
kRufs5xradUaILUsIU2HauEH3+g9axQ5ThmDqYiDnSkHQiYfCwafST0JfueAsUkH
OfYE9QM4zou9onwpksCI2T0WGQp4aOBPhP/v4/+fLwKH6RyLdE+ox7z1HsXYmIHk
8HHOmlfk53bM8arAKxPRTAUW2XTooA655LHUbS3vAJx8n/2UBimA+EIuPS59zhpg
S9cDDCrzuMjkxw8JywMxFiZaPvDj3u/4EWlSo+kpZmWYyEy1AHPdMzx4EbeeeIz3
g57xvKEUkt76DWWq/ezicgw6AuVvinLplVI0lXg9EPV2p7WcCNJJpiyZWWsSEXMn
Yqt94nnEXQYNHt4Zp+XE2t0EFE7ZBXQmwPCTkmhwWHsbmp3D6/STSID7hIYEiEKB
FVUtyxrEhGhFdQCR/eYappWe0cXW6r8yIc4BL+P8mnSiguYdNcG16n7R655DF7GF
1DmPpTVyb76wKN6gV2olNqbPKcqjHWS43/HRxYrFDY3uA2fxczWYwXdGurwIoI5H
YKi0deTbGYObJERZrg/Rr5yVCYDChVDB05kyEl+l30pgSzaigKiJqpdRaUacs4RU
EnsyzNeSryQvSWLu07U9VTcFUg8iMwxiz0/Cb02CwC0Pt5cGvhBT/1Y24LUUs7Py
6KfnIboqAYriB1xByvEtjWMv+56fJCA/AXRU/Ht/dvih9tmP+v4SVWVAoOQnyt5O
0o0UvTEp7p3Gfis64+NpLr/KUaf6gKDuk9dBl60Z/804qMk2J5pboHj9YcjpKHks
CnTCz3VamloeAqRIvVcD24K2quZglyveB81AKeAlGJXBxSyqr1Y9cmcmfVnzVuZ1
+SplA51K3bhz+xDn3od9Za7ohIL53Itd9QkR4x1L7u31IvcFTiCCTlDQJFRe+GVu
VYanFteLSgMSQZKihtK2lkXlCAOTPrvPGIkzH6N7Q14X9H/CSz69Xcn7fbw9r5+r
stkIeDa1ZImbeeR2TGv41KdL342EH4mFQK7Wwfzkem2btztTJTNCN/Xs6ZPzwPVF
sMmEcaLTxwb3jnaxnc5+z8wJ+fwr6VmxE+Q1IrpnL9nWn5iAsCnrhe4EKHMGzYoW
3o78pBWQmL8vU4tmssmMSPFwmKCP0OUhH8J5L5w3hZGfKSNOzZh8MaLu/4Lpz1JM
iwytHbdikd99YpYncXCA22Pob3aX78NRLhWY0XEamMSUQpBaAPHzVC7Bn/845YNj
vxPUPeQZUv55If96oUQgBQDIaUksSgm0eMD5P927/vwaWxba9OZzEttkDFx4R8gQ
voQXifeO3XhHxWC7ujf6j34qIpD6XdhAlqlX+hqR9sET7hmCsonaV7JgOYThRUfW
IZaaVdSN/r2xNgXgplaOyxU7lMaq+TSkWPabrOVhW6jLaUHaZRnxxf8PHNwo40XM
GQ3rgAYyix206ckbufzVSg+732ookNsdfnHl/ADMyNfT+LM/PeFFWJ1I8k54NfdE
1d3MlhiG95Oo71GNYFX7gYnbXCjRcHp3187t1UtLT1ov/irkctwYaplDVMniopvq
hT6fNtC6kWx24xnoxuWb6kurbqoXiNc/zIVWrpRHJ9MpXR/zun+wAXWXcG1EzZsL
8IvSIMqYqSNcsjWI4anqbKgw8ovlrlnsfvkcInPG8dfxCXEg0A7aypdlLYWItQ6y
+E0Rlc0HYwn2BjL545PfVJ1k5Ees5qQAcbt22kr6/F4jJ4E0tEG55zlEz+zNhoVC
wIzXzQ/ov+LzozOyLirHkAFVlC6hbrsz6Wq1rbvwC4lrxYvC+otBDV7yGU4zeiRE
aNZ46vK33LoVWC24x1u6bu23tVoTTMvRJ8KESyJ9BEsGFXpTQb5zst/biY4cOr6+
EgRrpiCThxQ3tnQPtla6ZL4Erp2v9HYlbPo/MP+5F0BwV6QYIvVv9VtwK9bBTWxA
kndBq04F23iNs3LliqgAEMkvm+dEexJSi1yGTX+vhhYHiU0N6/MD2zQubudlGpK9
zztbfVgt4BJJYvvx391S1TRHrwb5iYmf+fueja98Q8wF1PBC0Wap5lGingoyMZ15
U2cES9WFjkLFS1Or0hkc6pFWlFar51RyYJuC2ruizgNmzlj6w1wXkuuDcEkMCD//
Tc1/N7iGwko39WbW1ygM3fUb9UOHwEtuGg8QphfPnnuO4C6T837tXxnozgGAtP2A
CgXpGi9Mk8UTrZZI81n7d/IxYkRuDSWHxvEW4y7ObAHR+U/NvONRINWTLo0LCF6v
72tOLuiDNtU4MjeDYsbMBuMLX0NJtAbxVKWN1O/HcH4dQCbxp3wJddBbdG7i2Y5S
m9o82Y/DusXlb9PT2p/uP7/+lzmUO8yCyoXQKkFd/RW1TtmmYr58cACKDHLDdH5n
3zk3oDG7RA2ahxxdOl9oZCfsH3LaFFEOiXwYSBEH4kCHHaYEtKjRhrgdfkYa8HYu
6NMv1soM45G9lt2dJHcQCqfHp0RPtTWMIFEvSJMuDwj7LPiEjhm2kWiPI5ArdARJ
WWPeEXxYZj9pc/XQQ2ObLyJBpotOovw8HqthTN/EeHNdX1Zh8iX5zCXeDImZDeDM
I3hNXxhTX+sXj+TpXE3W195s86mnlhSYmc37e5jy6Z2GbENz4nXi6EdDSlmTd34Y
ePk4AJkWbxaiV9QaAQKTznT0XkvP22r6Bo+PuEXWPcLKMxRRE72Sni5j2W+WG8TL
CwS99v5usc2eVWJ9dr6YrJHR1T35gjh7wum7AcyVVYxe06zDpdL2F9qVJi4RgyyC
J7sqET4L3H6WkrGO9SDiiiB+VyLS/JIBLvyJ24O5x0K0YInV7j+8828KkhzMkxem
u6rvpcaTqC8Cr+ajrWd+ZyUQNvH2l3FmMtnF3NMv1J4sKyQa1Aw30Cn8WHQXF2ff
u6HGZ+HMmSVJXOXc6cmZEh/vFcKe5umy4FfGQWM2WnxmqaxaMNsjKuQVRF3VWwGw
rR7ucFyn+d/pwCmCgeWAlWIaIwudjvlbt4HQcRSjisLTcD/Alu/y3Ej4NyRwfQWy
L+vjVWxtZ11i3rVubKjm0bKXRYmrJq04VRT1on5PK4c9toqE9XcudaCfFSdOzpev
lBW2W9CMVKU30wkD8mHvYja2BmPaE3O6Wtf8H58D9eRGS7YXCq26+ArY/upfxAx4
7pucqu2OTXFRU6w0/uh/M+vA8nZTMjir3LQOfVeBgbeEPJItQ32MQKqv+9h4zHtp
xGfk6paSYIhZ/bnM2zaW3JqrW1fIni4M76PsDiuHW1D4ChlxOM78LzGly+0MfGVW
2OX8SQf+rzTeY1RdTtc1lEUXWDq1FjBD1qb7zz5OJuYJX3JdFF5NYmZKros52IlF
f4yKBMwWml7u3GVptJt2K6AZfB1j+361qgAMkiBzP7P9dNUWA0IOatFecXi73HR+
rPtCY+ePr6BF8s5PKwsUZO1Y5UrdIvwva3BJUZ2kwJ6g0M0UFRVeqLJ6y9Uup5Sq
4w5SDlb+u5tjjU9MsFWu+1XPTGEqDwkF0ryrTHphPKeO5nnrzf8KFTZRehKBPj9z
cv53/hJIsRkkmZN4+4WKDmCwe5MP4FjMZYGEG67sJQy9wJRpIxAug4J5TVFav7HX
hVv3tjyw2leNs9yDhccGjvnEjB5+Hwf47a1c7xYHESLYtlBZcoQmIRAc9K6IYgl7
qjTZmZ5WCx9JrPZyb0lvY02bXUuyWcotl+p8WYRfPKFzVKluo7+c335EsYISbqBp
lvS3/n9DGlQ0CYWUPTp9EXPp+3PgMwqBlLAPm/Vhlzv8PdgHyKRSp/AI7vGUaBtM
mjcOJVn5pnBhIW86+3RyKdAbpWnhGVWJgiBVRYuCt/CvmYVJAWam4CtV8+WdsP7P
8n5qIv38/ekHGhW+1DP2aa+8sATS+XRAKBAebw8WQlLIfZCslqJ8Pe6QkQ/+e+Q/
k7iapeqWUP8qO4J2r2+hFVEwqIcfS65HeyIwgbCKIT6KnbFjZmkrfaG2KBlNgXmi
/kJlmHbxbHY9xjGqCFSWg9bUWB93Z6N+wVifEsNrATq1YJTltvSnt+nHEOzKnXUa
stYyjvIlUzdQIQqVcpFxTcjaEBkRj3/otyLVJu4rZF5Ycm3nUdmd2+QvisgapQMC
m+GoJ7mxMQd42wcq/F+FSU4EKx9mbXbWUPuslHGGcDdPUgoVYv/xJ8Bt3hEgibOi
j+sPO7umepYO3+Q3tBO1atKSyHMfMH0/vfsg8m1+wuoEU6Za3U4oY2+EcT+0dCy9
GYLbHYa5vQGXtbxcj8csihTNw9IlRWFZavDFybbwqIJ8W0IWH+H7smydyl/PXrp6
rdIVxY6bUOPicX4Nbh6QjmSt7vdyli/v0xHukFH0nx4uDHv79TBwy2Q6CFw4X9ZW
e5I2dTkTykodGYkPBfPjDyT+yUgOp/xVEgB7K8/blHktYrKO3eqOjPqd+akA1r5U
/yq2rEjfDKH/ecFJJ6v7bAAt6y4VmsO/iCmjr8CATNtJfRRrbyFbpy7A/W4M2cle
ST3CHQulRGE1m5IalvqpWB/bvEQohUHhzzs2NPGBEHcqkZAUzZMbH6FcGiNKQ3DP
3ftbMhrnEOUrHOabxIRy6VCma9sg7cQVD/pIHrCnDhKg3NPV+vNBYoKTOUKL3DQH
2nP/ttKwEiaxgE921vMy2/KVyV2YyPqqW5GcyfR6oWdn0lN35tJyBpt8eUDMz9H+
zvfZZaJdyQNtWz4vATktjRq1oyFTSei2fAgEhBl2mzKaEWqBocsTlYb/TQS3fti8
inzReB/R1pJ0V//Bxgyy9CVavWYb5lA8+TKo2W9VjpxVlD3rPGqjBKgM5WVsfP/U
ELU0QawknXtxEokMO6W7qG9t4ZX8o50MV4jAD1q3UBEsXrQt1ZFt1681gHOvl1vK
wKT+tLe0hkfLq29ILL+Pzw9x5gC/csIC0+/nwzgJ0QYtMrpgjhavIk3MLhVPUP0N
JusOGiKFw3e4T9uk716SWQ6FYXdcFAWx+g8vNJ8DxxcPEZj9dTz+r+jYyyq0jVxU
l2efn2nTI3w9qF9ZoOJJR+XYgF9JhRADAKwK9Ka8oRG0VgqQJA2/cYj6S6tg1iwe
5WZUnQ7cSupafpBkuac1B+/JsyVHcuQNdtQiNdLyh0y3vv41uh3re9WfRiUC++al
BBG7KTHmyrnTo6sMwH4DUBaCkpmG3KnS11XDAVKdgZBDBvzKje83tnexEuvlobNK
fAFU9yU6SvbFUKu/Yj/9CBYjXqPNXqqcSArEFJijiVrkqQ46AfPASYWtc6ybrInU
fV/RKe54N5dKFOox2Mqa2pS/h6HVcoVa2op/LJ1k3cOJ4wTNczPaVEpofKkn2lnX
lfJnhUB67xpu9Duq23cSEPXPmfjbT8moiRyk4HD2lgGJuhn7uUIcVZKgTR7VqfTA
0Jx7slk0ZJSN62ReUW9Z2AeCdpuKbwyb6ZQjkiziyqtiJS+WNqDv0CJR9jZNDx7B
ON2VgZg4JWjVl9jkx/0hZ126x26ZjpakfRU14fxapqedbiFPKpvR17WuFgZK41dE
OetNgui/n7cV+uBY0FnePLT4bprak/bLj0xSkTus1liOylCEWsTirZ+dZZf9Ircc
CUTx7TsgCHCE+dB4DJQ0QfD4aBe9iAXKVjSP2uU5zjB1s22oWW4VtVePrl4LwnBT
NVuBETv4fDrAs+gCevKYe9aDgEsQXt0zc8ESsWkesQnc7yk2FELkqBE+GpIVoOno
Tc187RvbY4TuzuooICIWV8/S5CIPRXOeix07CI+m0f2vscbNWJIpryRwhQRj68W9
hN1aMqu3qI5/Dwv36YoYGmjTuZsNUpwViLeUeAHVIMcXFQR0IYyx0iHw5r2k3gJ6
LjLVEhiJdI/S6PPFzCQmlTWhoXeoaYESCpNsojWkLrPLyiSP4hs3586jd/RlNckc
ZU4OeLOd7ocFwNP0YXoKUk4Q//BGa1r9ubMZEz05CZz9gYX8fuHxRyMqAMPh/IUf
e1PdkSjNS2vDA/jKNgpo44JJPyxumrBAXyC+mGnKtwMF2K4crt6s0k54OZu58tl0
0USoVTGVWN9V49hwwPbpL+ysAStNgJ1DnIZlXahQqDM4FoPmr9dLJtxX3UXXD0JN
sEplAUu51KKpwyxMRNMPeJlFqyKKun+5xUwEYql6cKKlHO5MUbzUtqOcKoska186
zs/IDA8GHFXmP8igjB7Z91K4IIxW3MNUhctbkrdSwyF0sd++JxphO1UZYuxmanUr
HPmq/L1z/gRylexRpUtzCn+swzZdoaqY+TQtTDCOZM3RQDSZJAAwfHQNmgcpMFCe
jJmO9ZQh8Gfas44YR7N7/TwndJBjKtlSaPF8dM+YElLK6YoYDYb6tdyPtt1/7KHk
Q/O2yzRLkzQf1AwsQ2isGkMli1vJ+wezpFWaTGeHD3CKRgPiAtJSljwLW+Nqtkgl
7CFcqpUnvb9HYET+L0WeuVnGdMoCbMMzgFQSRXtdg6Wqb+VRsw57p1a3L1M0BIF0
YjeIGCmmCc90pkF1kPlj2ZsTY3cvavE84T/JWhlniCQExICBrF+s72MvO4L/SEpL
+9ZXYa3eumoDOeHiyQAD/3px5Grbpdb+XdhztvfYLAcpbpwnxGvHe8Csait3yV+3
p1clu8qt9ZoSAho0xi13BHtYbqDM0hW2W3uNy1IFtzAsenBAq5y+V3J23mW7RWlm
beOdfItB10oqLs2tGaGa2IPOZTjHRZNVw2gB6y30sv81DV91NaiIGWTgFkovqZ2G
Lor271OoFIqyJJebBp3nPAnNIfeFroDk9F8VJfleKCAXkE28AHrNY9y6JZ3Rbq8D
I1q8seHXaGNMzE/QcFOlt3zOlkv7OjEzttOkt/bkJfBSgdEhW8HsTCWOOwW8ePGT
9ZrM5xYyv86K3xpyzgrf+7rByWXWrCsaPEctloVlCpKsI0az2qI561iU7DIoHSsD
CN64xIdJXQBd39WIiL6aSQPdmNN3b2k0NY+3iIQsY+TGNKwnLSTMRRaDT+oqcjdR
ei7QZD7Dq17KeIhlUvI5Bfl6+c57JdLAWXxJbrzKqW6RXHwVn9pFycVZlD9mEiOC
ydCvySOXejUBC8Bt+Kc1n+uS2pFJOGE5neyytYRIBRfI5JBN4N2CYUs/BD3gB40H
SSDjYBRcf9CYe9e9f7pmRuXyffyBVleUVzzcXMjmQ1UqxiGt+6L3HuS4xU5PjuBg
oO0qNuOXHmgY/yqfIcGQ7/JvcTFzpX/ugKvmPkgvU3uIsTY97cQpEO9WJQVXP1vJ
4SNMe3ErEsVjAEv9ldxLpfkrm7UHyNd3mTS9K9aJvlaLH2B3aA8BtmtVqTuvgASu
3zUL2lOAmxpjmTcc2j8H2pvTB9Sy1rNeqHZVAFZVZC8kvHL+KVIKsIbtEq5yjtIv
WmDX1qcgsGcJ7GhxXyySBat/L7kcznaF4/3DrVxt40tu5VfzONpv2tq5ITP6qE7/
E3CFe3XUGcWNyecoB1lZnOCMwGQwLY370mFL6L6Gs+fnhSNUVT5xo3e9vw3jWP89
JsVbMbWO76+9r5GNohAz/FgHzU/XIoiDNo8vWD/2KjyJBPdKdsSUmQ3qQQaInHU2
4zzyVveSEdgv0r1Jnedp06Hq8xUGixnF4/prGgzTau1nD9Hrjv8Z2v/kjLEliAP4
1Jd5Wo78o7Ov+T/2cyDj4lAnxg6K+3EaGpfg4hTRuonuWFE3ZHBrYgIhOulbUUem
GcfYyruqITH7hGg9rm57dOHVRGKKPTPbgYXrX/f1EsToSGDrRH4vS6//5rmgnVEq
QE1/AJF6sgA6HvWhJJNB8bUd6+LreWpYQl+LnDSFM/RSr8EjDMjmqhOpESX+lkPy
m0I9JEbfJsWxKCh6dx2UClLUwma6IItrokxwEt1WiHpv4aml8aFv9nG07hV6vODE
g7NrmY+kBvf4RcREu0SWxJ0bnmwH7oMZXWANFtgqJNsO+LG5T6xFPp3P301Lj6eu
ILcKFsqs7/yPg2fRit1VgtLYuUG0RmGl9zXNkhXpXoID8qlzt2dJ+BiuXcwJoTYG
aGeGkzpiK+RNZtrQRuTKSKWi4HHLW+eSBFinI+HnANX+yY5dxBqes0aWwteY/Iby
nxtOKsBfDfPJTC46H1+uVKucKLWQYoAJgsp3vAEAFLC36mLOYAwOfbsZMY5MqF30
8vpz0Ng0yqCEBImAhJPJDIBx8iGTiEmxg9L4800pn0DZYfGyxz3z78kkxAAwP5ta
HX1n7gb2SdVbhOgrVNUcI4tu2gD74eP2LlWfgHIEptStcknmGpghsMOoQwvEckOD
YvCHAE2br/EijjdOKilJBgzZUN0Mk1BPJVnRaZhbuy3b/ZwZLA9c5Es2fZIjgf/r
suOy9Wp7gOc6YTtKd09WQ/slIZEWJYhvwTDH4H5/b4o9Rku+hYEIpPZOPxqlyuss
t3THPc9G6KaRwmAD7GipjvkXaY37RaKfFTZWuUf0klpnU9jJczri118k71hUi+E3
HLt2Gx0mRDHx0239rAyODe4nk/35+3eIUSRuWJSVXCdXnx8/ktloiOss6A0c6vYs
TYIxZKo3lKYyQc2PjaZ6uxY6d5RvADxgb4OCx3p1MLnoUOwn+JssAyZIMpIIxSNi
mw44uL4ZFHpO3JKEB9F1xhNI6hUylzZXKnV7Cbq31iXsaBfi7wABZB1/LtFXgamJ
sCsaCvUl0262VTDWobWWmrm5Pks42HIKeOBAwjySmqesm7bbQ/4GY3WCgLNyu9Ec
Mxufe+yXzp1GHNfprfg/8B44F8Buqmz6FATkl+7tUTx8l5aJod6sQq4lRlKh1/Qt
jpkW4roEm96UoaDochcOIIie7MRvEcqLFkWdyD2dGaqZ8Zukegnqwz/w6s9ty4il
AyDxoijii9bVozInfEKKiMaSsjYLl0PZeyUAPXfh0vTWxPhINvsNX4aIT1jTzBXG
JOuTMjPbYtWIyu/8EcZj3DpJ787J7NoyG1OJN4fIcBThJPHl0IOEqIRviJvN6vil
ZS3teLE36SZ3ZXLDUZr3/3nAbdPvsl8JsvWP0BGgPLF2XxJ+R45bIHfvpyy2jdUF
+9epcdmQVzFDPKAOnFUIUjKQMPXpuC45nEtNFXc6O46qRDXeSQQzRjaifgjQIgXA
n/HuNqBFZAK+ssCOGxA37wgre6Kxw8QHhTnOIOp4P2WtF4Te4YPisgrp5dH8fWuh
qTTRXatYGJsApCGXbM6BvbENnPQW1KhfuXBh+n+Nk4A32qEmx7li8kNYOmbgExXN
gRPFV0pUMsfZwvtrjOI2QAxxsMwMl6TuknBnzUxs4XXfOdd9yxHrcQySlQxWJVR0
2PS5b4mXCmNTcRvM84xrICrqvuaLRK20SVAfGdLQD+BB8JdZgV67bSBTrULQdpfb
K0BvuaOk3JZbg1libxxBxsJkwhfytAShBWtrQMXptd+huYyNzg17Sy2ML1r251Rm
Hn+2FzGso93M7iBOrJj33HxhFRMxg0PYCW9dPFD3q5Uba7FhRISgYUb5pFFqe9tp
84WOfcrlr71ZrH09tH9zhPi7ZBOZdyYRN1c9w4ZA313cWAp3XvBry1NG1zcfP9FM
LsY1JmOczSDWd71GwXSnoUUXmX4t4UkwhXk0cVx5cMvmNQLF9GpWFY6ERoHO9VOh
aj9Y0g/D/BTHFu6HQEem4kOhT5wtfw2MAV6HlhyXxp0u9/IU4Nv5S0glI4Y5z4bC
EqVI7UGQVSIwXwE29kc02IVFf0LyJrb2vsEXhi5K+arGhBraCUBL74pQZ4emtZId
8K+QgwL0W698LgvOxZ6glCrzy7+t5tSub9yzX24a1wxcH7pWo0mCLVhuB4gPfVOC
dGb97LXDsK+ohe9qJiFS2BnuIfUY8E/gxyAxtgDkFsI5U8J4/lLIk+i0QM7goKHW
nazYVcKkg25IfG4BkqStgUkR1LGKwNMYql+q4v2+B4dgE2qsCeOw4pulyRwoo1s7
F3bvleOFWVeNPWWzFbD8+9GhFuamniEOHNWwFi/dzjnysAbJGatl51njRiDmd8yj
Vqt25HquMOqSevxJX0alylMS0pTEyRSEuXTl9uXycITZg9J6wlhLzOGZA0StWtb1
MdPzWoEEjRLCwM7CphkjxmIQUu2AXNhBh8DNnEPL7eIKuMWVJ0cmiig+7xpCXTr4
UR5Sx8OPS30ToiukZMoscLaUWCldY11Gn4N+c2fUN1rawbCNJN2wwiEkSxnfCt/F
SRSRbDItReH0zGJdupxoIu3/EjSjIcWyIiTDZbFv4XHOc4NSvi1PsKwCvit9l9yY
DLUG/WE0z1qfztPdb36+UW6Y2l32kQkP/hX6feztAfat5mJytwchLOZq9nGwHDoP
ULiXfCPtdxZbQ/Xid1R7xYWtWxoDdpu5IZgGdHh+AUdkg4AQeBEpsEXGSLHK0i4/
hjHFoBMi1hYW1fNpRkJRJ0iQWpTSVG2qF2HNbhFgseWUvnLgOQywkBm9yNR2oTfK
SPQ88JR2zek0OHiCD1aB+78+20YVTgQdek4cUvg5cYolE9Pd17SlxHlajB5zuT5J
lYx+Ofgr8F/avwVoZYEsP/FAoOg/khFQfjqG67eaoxY9a7T7gYpedd3Lea7qW+fW
JvFcfGPA9lIpUjhzK4VREciy3CR/Tz/xnwkjX6gt3qPQS/2n1WJxx0ca5RKBsu3H
WjXELaySG0k17OUh1eL2D8T2EL53LI8kT3tnC1oD9n/BiC0BR2yBX+yrO3mf3Ham
p2xlCtUPKEliruN0olCbN7bPjv/5H2/e+VfnsAKUDm9/ToU7MKw/r+f5uO2yDNgs
vtTUw29s3LuF9tj/EBVyeBSOyik82W8FjxYNS3exWP38rvSaH89lkmoqBoDqHvMK
bv9zVXugMWeANG/A0vYHMOgzlVBcdUJ2fGWCZCj6CSoImUOwSLPkS0kCiJODs2yl
zdfQBHzUbxt15BoFqU1EDkG5xWSJSjV21gK2K6Rrq1BD1IqbRbOJzIDoBma6zhAY
NvpY5nILTv6XoQ3Md1KxqbIq8loJdiDQepgf25xkZdJ8PzuT9qspF2vlQZ8QwSy7
kZHT1NJZu0fN/kyGbyH8+1chO1DTa60hLPtykqEljropw9WuLhqQehvHE42DK1gC
w4PEThzKAYhsc7d8E4jcdXj94d3vnOWzH+8cnDbddZF/TEATbklzMedJ8rS/5lPq
xowA4IPaO0IMsdTXrOt2Ei58jK2nKf3PzDR18KXdsf1Q4IPTSBF6EwroPGtDH/mi
i1kxqgBTIJgSsb0fvC6kUXdR4DvPLt6VkM/bo7yI1jOuVrfS213yDn1jI+g2bLBC
el+i9OSqSjoV3x0ofYkqojlOHkAnsdfMhpBZaW1ww+xHYvU7XSi2h/iOm2xYI3Kd
ascmHgiEfypdbK8isQNkONo54B9LUOfSf0HvOP3zH/EvluXAOpmtmqwhmvI89U3u
vLxw/dleNSuUuuYojU4AHxyPxQX/crPA1KvkpKrScN8etPfZyS2OiH5Fr+fQh6tX
y+XSCwikTFrbtQLDA5ToIGTSdXLa4D97ZmL1q6uv3o029KxzLOClUgSHUpmodi2g
AGLS0ZnUZ1WCqyozVUEXKD+nrBBhzpqPGOet1UFjLtj3aYklFLFrr9W/5Ecvq+o5
98uskWm3TN4fjwC297XeDgISHskKyvnhb5X9kZgDijvU7L5+CdA7BPot1vxdp4bV
G5bY40jWgKIjCKPxZNxfxPhiIcpP4urZuXkzxvtNtcAwYEQIyQ7kbEDXg/ihSS9c
8h52HizryjvZB5IIhvjVH7YcgwF7nhxrCuYb1GtQZWUwtGs1+Ug1t9pWatFrH0Nr
NgWGCXU4SdMO4WQter46liTtq+2iEEVjgVNScZCWhcjkDJtwStDdz6wofU0fal6w
H8AdKU2EWiuYo4Bb/b7PUvtjeSXZHxqwIgMYDO6hWPe68apajXONvN1OP7xBH7sg
Jp/6G7a4MmINknk/dmbTqBvGDIewpZsJYNfSrM+B2UlvjF2zTqKkodJV0VcyIWrK
+Do8EDgCAUczRVp8FtJvOML9lyot20zwblMr9r5gwUwe365rUyfCT3Tr8sD2GOat
wppXt0gbFM+WMACfZxi8QUlImnGBvKcjUQbjG1qzT5LfsnnaUxYfAfcq3DUxnepN
CR+OzBzlOctBQHBuppwykUnlSZJ0mVaehBtf/m1KhrDQlaaOm+Z1RqoKcZAoMefk
OKZieF8e2/CxBgJAfvcd6uV3hqocN0RPiE5aGBUOrgK0l8DQVmlT3HRCC7CMrN82
aTh5mhPAc5sND4qk2Pk/BQ0+/vnGeAPfrr3TBCnMpoq6gwqDFIL7eoEcMEj+W9M2
XyZ5JARv5XecMA8UEpdyNlbUTQoGpSmRkqpVr4mUBbzLsb5IBmf1W6Vj4+HckmQ2
f2QQdqXi0usl+plL28IOFiZqk/49uDSjYVxCgT268g+0h3kFK1mPm+ZnsH8z1kH2
Th6xhGlWctI9cKOzFcWCCT5UADYX9DZmpJlSzXrRma3znssUa919zXaAO/72EDz7
IkBC9cQ3fVONsRu4CbvuKwIODau1L9hxbpmmeYb2q1O+ElnRVYQcKqq12GCHZhnM
04ycENFeuZRp/eWYEv435spYZEbBEzkosBhVOls72+4W565SuPzbHHtgPPiu9iG6
t2l+hHAXGxEsVTS+Hsj+wG9U6NdRfqE99azapkpWvnU+UWtdUlKZyFC2Zbhj4eH+
cYoF7jw+GUjq6FQLrrK6utjDlWsrOjhzH/L1yX3q20jCzHLcG3T/tm8WUovQPwq8
U91jDMkCcVgbyOGIacCn7n2Ik8ll5J+2dzDvL1MuYAPri+WIxb1to7Xbi4rGI9yz
LJU1HNpWgfyyzokRF0C4LzdiX2MzZIHHbUcY+CJrRfy2VMjy6RqDJf7MUQmgGYZN
JbcnPgVeTUEmZK70r55/i8ygulW1GYaYEUYHZb7fIF30OFD6JjTiJ93ahg9NHEEa
lyUM8A/A49Ve7ui7veaq4ODuY1mjyhPOXiUWvsWZMlDDeuZ+KE3or3fnkaMGta9r
Bp4auPdb0e5qyi+11HsQllf+bz98k+Mh9+MPV9xRE2YUZ6RTtJKlKcc7dtMjtR/U
phvb9rw2lZgQC1bISsgVBnn8aGDgGpWFSNAOV/L+YmKMGoPV3Y9cCRpQf5PTaBrB
ozqlVpYE38Lr4nLIC6ZH0nd81TK0GR96Cf1SfvZicma0HIQrs6mRCNKrBp2ANybY
0wIe36CM+wlmzmi0jifLvVgVX2XdUkcm95nDLq4v3d05EBrtmR4co54xv9f7Mxt5
HjFu7sj03mbJPKxS45Vh1/x6gqV6H3+Mhfl4NxO1lWg+DpG488fA5z3ROjE5pa/P
oOp+Cwz52PrmF3Tq/gwLCSsfN06MtiUKFqbwi9lx8e57uUVX6A8GZi8Vbd7pMWXY
hHHU6bCdYR9poKZ2F2zRE/9iy8monCbqsYQj0GTPz8A+ZsAzi4jN5pTy6RTnkEn0
g/4fUdfRHhligyI7StRZfZv2PT6P+d7sPBGz9lvcAeH8QiIN4G+Q9239+GCwvrso
XIAxkto353t/HNiQB+yHfRIXKFYAGX+JQ5lZJs9koFba69OpqcrL76t3OvAJsfaW
ny+kmtK/X5IRFeB7om6wC8OR1yfLeExbqGtAnWIYbdOLmaySLNKozF9EYPoV0BZ9
ROh5QN8VtLXjfly1n5uf5lMtB+WIXMo2xDh9lfkuKkWikllUZGgs1UQpqChMnjWB
NdBWSHBxditlcLXeEtFidVGK1/cjo49f44UluMArlw6emS62RKvHWW/m9Es4HcjO
Std2xTKYn7DpPyg6y/FHGlBDYrq5L/rddUOE9fgqbYhbM+51av7ETFIysoO4/lU4
kJeEw7kCyQbLhhMRrd+JPMkMGZ3/ogPCMyXTT+ZAInssbdVQrvPzNUaSrKOrAcAR
LE01yjPMIeGNVCg/JhbEVBAjOAnxglQTJLg7KnMCIwJ7mAwU8xYec9+BeBur2KNR
kFaaJ7W+TG+Zh9GVZggjVCCSzJdVZT7vh2kl3VMSod6z5W8LtERTA9GUBfCCzqz2
AeCTrIaad/haAFx0onAnt0X43MJZik/rA6KFOoIt4Fsy1tK5GOZ9d81k9i5qnBpB
kbEq5fIMgjXCfo7jEd67zylH9cwax5OVBe2YLnQGXbVJTAJK4azUrGhLGFyksdXs
/3sDujQn1mvzjpKUfGauD7Q27z/BLxHqy1MBzw+pEzLnlVBgCjY8q/sqiZCxSNha
lHMpPVlFRlpwbd935ydOFEhFRurmebuKXHAlEQFwFALW4vw9DecvYHULhqnvEQIT
tw0wy2Ig1wsatIIGjvGgZSmXjLK412Hm1CfD733vCSANWYAHMDDh4tr56DCAI44J
+E9SKQb46dJmE/9eSZ2Sk2THIX0fL0PfkoxCb1LwdYNGZeaaDx6unxIaA/PIQfKq
y2nSY8akZQv8vQnF2+aB96WU9PDEPZPt6A11CAWkzQ5wNRac+br3TtedFWDqC0MN
XeTPFockVAKliUhAq9x/Fn+7lFVGlkxMlq29yKHEOMDeGRKUOgVEFzvKE5oA/9uV
XibD7DhSaHcLaZCiTb9LdHrN4M6KOF3V/Urpt6lgP3utaZXkLiJXLQTYH3L+FI8/
fVLCfLmXSpIq6GOpDwMNXYv9QCqB3DaAUgXb/PFCa97esdaBd53YANBmApe3jFx+
4TMRjnVf0YQBHwLDneZpRsK/vRlFhDl8KJ32XP6LZURq9h4B1/khA64xeZKHWpo5
Ngi+46UK9nYmz9roynySrWAwE2lXdNdpk7JuvXVSEKDkeh4ME1l6mHRlN4cDIKBV
Trf5qRUTgyFPA5bYPOsgHXa0e8FtFESwQLi43XPsBtfQhXXe6c0lm/XXX4mlWEPW
+aopnVa212LqW4eOhnrvxkFy2BauouAtkPCZKb5wEH9GzNqoapP5Iu216W+lnGws
Etj8noxvq2FQ1aHIvIfc3jndh4Jg2jRQ2V8pzcKr9aZAZiB0Mby0tNH9KRgeFT8m
ZFI2i12LwzKJU56gNwDW+7DMop3g5hIyClmabiwifWSwzbKD+LiCCoxFW3VThm3F
oKlsBIoeNZg6p/Zzp/Ykt+E/PWMPitGyRqBGzuUeqe9XEAUmuXVM2WOL/PE65Dox
VLzLD0vnaKEnyu4wqqDZAiaAuwvfRsGJ/IWR+74SvAgk1DXbiLXWbfjzxpXywIFt
0P08VuQs0uBjeEUA8n3MKyajAQR+WLyk3evqg5OYTzMjRcQ8BwrgwX7eouZE0cDs
9rMHjn6rClGRht4gyQLKgFL1jqV1SXn4bWldJCRgEAgsFAbsd1gGecojCqzApT/F
5ANsaBaa1e2sxMj1RVdmWb+eAOrKF/dx64P8H3EtVCvcd4WbslkY/aYptSCfL1cF
FzN6aPh9DeXPpxwqfF1AzuZWM7XJTkSo/mjgOGEDvoNjuIE1WeVgYQRf9oMXXlVs
WU3J7E/X2ZhzbsZq+dnvX9luNIa/OAsyt3rSaew8wHUuvYRslhbO2o50g032O1iC
3hC632Ih5ogcMRF312Nl+glDr0AojquuoIPtTjRTTsLBZI+vS97WsITma+qjA6Ys
EcsF8B4kdhK8jQty3yl+YVyXJKNxC5gq8zDzRdhCaFD3REAsdztcBjrGlTutiaf7
UuObfL643kO+UNRyzAy1wpL2r+qVUdVn2+TRF843fIfqNdP9qVXsalEGOLMvKrKT
EmZ0g6Gun6b+3SoonK7kCGMs4R/tfLLkzu8fEe6AeZrFEucMsJLiyY0+ixOyioUD
I9vw463aOStBfSfiQtiSJOU5nj8IsIfOB5cAfzlr/+e3iw9qGFIlMcDB0Q4QoK89
doSVet3HdILCRUxsdWxl8HPEbQ9OATk+N5Xx0M2Jb7ZnZ2mXJUpw2gKbgPebLj2k
94ZFhkKxAeQ0eFElFBYQ3t2OZl2ooXgzuSN0kxZsj+FsmFn/Zp7u1to6L4rLIk5M
UFHMx3Em9iqtGFe7sNN/ENbzh8GzQs5EkJjwZdK01a0jv1+tWCUNxoD+gbr6rGaS
OS/4Ym2wEEYHbsrigh8TP9tlBNCjlbXMdxJSB30+8/5p7CRcICDrPYoHC0E52YRB
pNDnI5fTtGFsKxRgf+gVsPk2vFLD4ab1MULNAx6fnJMy8ZaHfZI/hZ5wOZzAEXaa
vC23VmBtNJb0N0538dZ3dcjHmTarSczLSxijDGmMvh0mQIHt8N1l7U1TXc4maEr8
g/kYpnMR3q/5fRsGCh96J2zSbKx00hP097Aotp2FArE4kFi6cwpveAta7cBBCW+k
jdLtP4AFCqvgs0KyWWf9pIZG4qxHyEsAYqj23FRU+NC0i4H45H76zZ7TjRjWp5LD
kzOg8G6RnrPX4WRl6+1F0Jw74ztUFbHHqhsvJXyqeSRtu+w5Q1JePon+6QkI+Mi7
jF3hKJPyjE/2h8xySYEiNBRTz5VNg9Qx2gUTdSEywLQAecFNiJ2REFikzZc/mEQJ
7fkfug01eShyPTKz5YGngLL0qbUCVuJUl/bCnojYIz36ppL8NjSfR/gy6qN0eHow
sWekPS9IGF5UbUPhd7WPjU7KnPQE+x98MJcYsVzORpqMd3BcmuQezyK0Oy2JaJaA
SV6ykz6gl6rN9KkNIrFCmWP+e8HLQ5NNKqAGBt2oMeROpD70IWj/gEordiKtAo1g
qihiiCkdmdppMcQvsj228pt0/D6GBjTNP4B7ey0SWRSj2cqD9fhheWYs4aTwRDyp
CNY/sFoSEsUx43N+nSuuogJ0dgcEx17x6UkxR4sJH+V7+UEeHhtlYfEL6gFxkN3p
1wb2yg1m7DuLVw7LMC+kdT6UHfM2FffXLG6yc7mp6BwMWKD3ZrX55v9ftSVRjhy3
xRSURtYu1jM6ne/kjNmOwmCHWv8BRsD2W0GeCzdpufxEVsqi55mPp2wX/1oQi/s1
hqyyjmsnqrRFsqyXximjGv/iu06UeRNgtPJ12ob+kmu/PdqAdRF4Efn566FSvlbx
rDrk4HMBJ+fKKUO9oX5UjkTn8PjLF0x7gQ2h7ErP2JhUFCqVi94JISEAvEAv6cA+
AoikzeE/VetCFN1/em/El0rzCsqm9MGVnx6HVMJO/ArwQkKSgvNU30S6UqSDUQiO
CxhmlFAb1Ub6a6buK0fxEe2wlWYtTMalpjjqPfQr1Bt/4hkOC2cEGEoiDO8eeV3o
h2HNeeU6orIyVbXkGvpQB22JzbcwgZddcxdUsG0wmW+UfvXtMek/UslOldouRuTT
NZ+xl4GR6SBHSt59TXIiT/LQ8Q9TjGRDEtKKOkLPZxMRbB6+jNYdVq2FPJYCvCxP
qbqiTQlddZq0WEIc5kxNe6iu3iUDs3LWf5eOXYWpfEZSWoGEukrlVYXuXXudxQ9f
YmiOtMXkoGgQu436NgI+lwRY2KhapXb752jKkD1K8t6bbyZhL/pTvbVn7j8qNu/a
V+6pOthuD0ux02ql0dThnAD/lMvcdKZHev0nA36p6yWCqglEKNTvPPDI1z5OuXqo
PN7tLqWlBCAH/u8HsTH0R7cQXdyqBDzFc4vAiM2rxD8tLbIGhvJWd76i3YL53Vf7
idZJbQebaG9+JACxVnPAegj7gYxNauQiPLwNFpuknwqp1KCZpgpxpkplNcYJcftI
w1yAeLXKsmf1pGwTCEyR4Izdommn2k+Ev7a5qNtXYTGrzhJUcldgfUnr9f5EaThH
mT9QaRkNUzdydgYC78vQc6J40aOhX24xxaowhzMc4K+DObOQOCfk5gzl3P+hF6Pd
Sd9mPsZcJ35EfYxdFPPhadCHj1LK/PZqcbuhSU6qzfS0CPCLMVbUzhoo26kZS3rF
dwAVx2i8QS6BZYSjaGUaAu/JA7t5C03PmSaF+6QcIRJb5NzKkPlTCB9+xfCpgf7L
pNWaBHWtyCFWgunH4pfSUhAiqeyYE9vR4bKYQIu3/rZkX+JWU1lbT5lF4I2UC/+O
OY8qW1hHczEHiWOY4TuzAQdcx9ydlS1jtiLs/puiqp9Sg06FKOgTv73t43Od14mg
CFxQqFynh06uoPiIxY3uvvYMQcQCRBnRXWLbpb9NZ7mI/IU6jXWStTaYjQliBVXv
bj40cio2agN2AUBDjX2oYeRECCN4AD6csoXx6XKy+SDP2qqYZu5/SPaVbz/07e5/
4Ze9CXuuLMdO4T8dis2xxil2GVHlRbzXDwcE2tXU96SuSAQwuyR7fPPToLixX7Ze
JSPKST0mw0t7KIe3+g6DNzbk7xgxOWYER+/zIyfBvejjgimAQvstbf7ExENhVVf/
zky/Md2NVgZbsGv/LgaRoogz7ipMXRrw0GisPjscCg0XIoG6efN3axEnFjYAo+z/
im16xptjr5UHCNVKBpr+inLTQ0IFmZSRjQKQHHCbzFx2LsVQdaHiNr5YrB66hWZq
SYi3StkUxVpgNCh601bIMojGSRVQTomzNgHwMbV/68Z5g/6Od/OWNZuTUN9nfeUh
bSgrs54a/toc43pSxpjXhcYB6Mj6crCHzZnkxZY404eiuu3d6MUkyJ5Xw1qGe1bZ
Ld54x1nhJ/92cZs9czB7v9ii3pCX8MBspsXscGTW8p7+YkGO6NOF2lLSkxoj1HL9
qx95VLRoCYO23hwcrDOCI+0FDlLN0b9aL4f3vk01ZoI8oAKcQpT1XSHecxJ2/FVN
YAsFCkP0V4XqxoiM+F+FI9aTkk13ZZTyaARJs+/qT7BQiHXRYI8WMopvmxyyHYcz
4o2t2lTFEOzZIlK2ZsZzUEZKT7zp2I6pYiUvHQ8dw45sLc/+btyOgVb1fSOF8/X5
S54vNFdbx88q02QbhzJo3dh4gIypfo1tHYyDZ86qkQ3DsLFhD45uFh3lxF89cLPV
Z2Zk/d+glS1D/S92SxJBaItrZEnPZNP/RU/+oetnuBexDx5uhDJ5KbQxzHfQkTDD
3cJp5mVU2sFZlfQzFbYBwKAsecPo7m3OlhCnhTJrrcgjBWhoWHOwNWBSkrPxu4UE
iQblbxdaiGw/DiejAKhD+vMBbwU+jDqxTPa0Ys2O3isMYBM7tamBq/A0tA6h8xyU
DZcuuUOr9hMn6OdOhEhW64kKM32/FN9+FlUv5xsMDpo80VIzFxTYXMh3DaoCODVm
9weqLGmawq7nQIymXxtOY8IFdWAZ0C/BhWGh+gG20R7AdrTKG1gP/gu695RhbH9p
2jXOaKMlOYIQFLW8Z9WABzYm1QFucFE5NM1o3cHsbtcQb6utkZ5/gAcHpO93NVSc
jz2tSkrTQIJ69uhegrgGcw2WsFyQxXgsizPsEkhjeY/F9KJmCtxf14rV7W1O2USj
3pfT7MVZjPH9qZTBZM3p2tWO2+aXzUTDTGJLXZF7D/ohDmSf55cO++Owi5q1LMAQ
nAuYWi0BSz4yRQ8B1OXWeeY/0aI656blzhse86V88BKbsZcYZZIFIOamZ0t5m6Tm
s7N0f3H4jAT0sKz9drWN0ODWwBHvmSLQBw5n+A5bG+E411Pnqjj7KIUiNdIbDmfJ
8zLMq0L6pcjDW7q34T0Z64E92euf20YqwbHPoyzVhosYS54FMcVS5W0hFK5WBImj
YY0Yxh341weZQNttyF5qXg9tiLGVAGtgqRAHium9dOZxdXAcq7lS1E9nW0zJL6c4
qxtC8LCmu7ROCw0bl76kI9+EHrmgqLazjLRn/KuyxmXeePTTHD+uZS5oBDLgGvZS
RXJgeZpEUAo1UPm0B6FKKSBiO685K+6cL6RKpBcx0wwWQ9/C0uGZh99ku4YWnOcg
rUb/qR9szE25N5qiGbGpHYZTJNAUMHwSnitwyR06ObTn+OVLfd2GPhSnq31jKlMM
sGZnpSDZK1l4x69fK2BEoh46pUv3ekCIosLKH/BXVYQWTZnA0cdgRZp9wJjTWKGg
4tih4WIcpxBo4Qk/+uYScBmZIC/+Z/KIum4xPQc9CiBdxLPtZisvZX7qUi5LwRuB
KR5sEVIl+V6NytaZGpM5IwwioDROYqvFGJyMqBNTUjd1ithQzgZMFC0PkjC7+ICd
EjJq3Pq53nWY1pICLZ42j2AEUuNXpJhN5fNf0myivydteKYycfj3pZcTJYxjOrvY
banY2XeNEUxb0aJ+OCgEAZP+QaHkr6uvUByWHFo5rwW4XdqabirIBUVPGes9ZhYa
eylrJ90rmkBkfhAQ1/Gfo9A0AMai9+rUgt6e2HNo6iCRVMGOpmyA8Ezde9+DS+RS
rNwUguDtAoxSFDAUDcmoJGKYLcVroRPVamy+OwtLkMd4shtstHC4YAFDEfUVBrWx
KEcKYLvKcX/k4ZmKUkkidjC3xxB15pcdcUbDBblAyES907cG6Kdw9sGKyhng5zqH
DA1XVykuPNhVPPi88YBxw+oIEOuQVsARacB7INkRQvm3RRS122w8+8WvzXB0dGWg
ZAeaoLgRDiUIo6qFdxPpxImlGnLFtIpmG5t2JX/gXjk76jO59SpXke7U/fWeomHs
j4sipX3Fe0s+loamj6uN37dHTh79i9oqEFPBg60W7yBLqP7YTeKIb/yOfMz7i8GL
D0lLiwBBRz/jrXz323/6/SOu8CRniZCDF1rjbWbRlWlEiVRynZhrlzxJXMle1LPd
m0Jwdq33dNNj+pe2IckFgQLIWGIHhGwTkyDCbL1KeRRo3j2Adr6paGajc4ENHMSj
O+mVSMvwcjVUb8cTCzwUQwj1cjTcS0ULV6ja6HqczgmTMVIL3ULl0faMty7o9WuW
QwCwUUSzav5oFqdzd0lk4uiuQFCbdkJ3y1orX7o7AR+A8pVjeZ41qTO6V1u0QeQ/
a+Woq/uw9UpEyZzF2TwzYr8tZqYZM/FGrQ5X/r0kSK+Keiau9RPviE5qiv5QsRsm
I83HzdJJ+Cu6/enwM3tWbnRBoeflN+WO6Y4Bd/cqYC4/VI0H5cP7y0RLsaXwmL2Q
GbmYgOs/2Pw5SXaU8EbZTIIvZLqzBzwtfPtvYKc0VjR4jYDbEeGngYAXsTdVjWWd
AcLEPIXJWktOOOfQQSwMeni9UO4osJsZ6xOyzNt1aR3dZdgwf1nGmuMDBtXjysLP
Rqsh1u2WfK2w9XxumkHw8udM2zw2v2z98lP2ttYU/CGSGEMp0Hi0ul0ge1SnCqKK
5CCkuYteG37lzGqQGEtwX5YyY1ydpWq9jI5Xvlx5K9rimEuYbMVZ0bcSpaeS6r6s
DJR74J0uJeHDCPaGnnyxmYGOYRZRfohD1J+tOEaewNwCtuM0i1FudiP1lNubI3/S
DQZ+XyBfMVSk1+/tfzI4ZFIUtaWJlnAY8Hqtg8FL3dD8BlJ2oZoiVrUHaZzeUuFg
dyCBWJFiifghzJzTzDAMF9hFUBMTPdkzodBGyzC2EvKXcIq77FO5I4yEtQc62LDL
ueeJMET1s83tJf5UH215EBRAIdiFn2byBUgfL/cl5UazZCXoZKlZ1vXJirlRnjdY
CY9KCt9sSQdGn7TdOmHI+nIbPmAPcxfn1ZRisxs+crk8cWeIm37dOie+vNINSxdZ
5sUDDFVbo8JoMZoItgh1bIWOkxzPWYiDqMUmjAH0TXS5hO2mOufAE8Jn7BtGFz4N
lhG02EpBzB2brguVhu0bsnaXHY9IcTuXxWkjs2lUFT2rfHHGo4E7Qvsdq8mytehx
eGUzGqrh8gDaNrMGVloQQwSeIz8Zx7mi1rVCySzXggeOtLU3aAqlUZpGLC/jK68C
j1aa0/tM+yrSyDULQoDSjoFUI145shSAAVgxX4S4rJ1vSAH0dQY48GiM2Gjc0N6/
vJa38p4FApKTOhouD7WQMjhk6ERvI3+oBMYWueEVKQ1jsUR6YbbFNZTSo8u5zTvl
cqwC0ka475yMvaKS4pYisPSuL+m5qaHW+I5WjcJC/KJx3ukZO0sHbPD02AbhCSNN
RqyUgsCU8223qCjPbeoWjQI5IUQm2RpasOxp0U8UntrZE24C27ltYxhQzXfz0ygG
FMkUtZSCi6tsvwRVc1hQGJqATW4r11ITOPWf5Jd7h4J41W1Srr9dlGxZRPcH2Raf
ATxK2ucUHOH2AmIiqnQ/nScC8CDtaq289T7pjKDxscLk1VKOkjwV9tJ6BGd/eNo0
PSMfT5z/i6GVKsYF8HlZDaJDP7HePLyB2V6ZdcbChYUoYhCiVZ73WgoMKv4Uup0+
vZKc5QctdAgzGsAhFHsIrHnsWkLhOkfBq3BUrkGPHa+FETn91mb4OrILshbF0lUH
N0BuCwNe3tuTNP8xlG8TJhMFKtwljsy/683qONy1+3MKIR9kczgkPV+afgW11L2K
1s48kkrBO/Dhkjp/tHK5l/Rn3dJuxWFKa9j7KeJ0xW02hiBmqy71xf5Pbbr2+kuP
AhiFo6UMQBHh4QZbwGjT6PuqqqDp2pj1sK2j+/dczbOysklPUVJrgXxoDU3llO/x
nL5kwFnkli3N2h0Zjh6Eza+K0HZWsyZj4l04dP5ipXrOtBt5s5yyl5zqRusIVDIA
in0FFyRhBUjUXmC8wO+uBH1AG925u98FCGzNIsoGEDDfPSgFWyp/lNO/xH1+wJ4q
uw6nBgiQTUIncrJhz2eiAEN24rc38KBtP23VlCiqtWjEe+4O8hNZfWRRZM0xrG35
cIepXzzF2KhWDGWtyJCr3VYhtERXb2IxzM5OP33AyNMZTJIpdgIV7YOSJGg+944t
4MuJ5EVUPuX15euXDneqfrdhdhKN67ko2zd2bRuNGzcjbWSec7LZI1vFSEc14Q/L
uq3G+Fc+36nk3E597WT9IHpCmjzESgWQKjMr2h+UGahPea6Gd/UQJK8jWbJCXkq8
RrbCGw6I+CIOoDatsyq2jJsUMV4ftzpnjsJfidXmQ4sBvq4GtcY+wmSKIkwO4AfE
5TmKy+1HA/7IC6Ex+WKus2eTjlfzo7tPyBb8LGs2ULCuxg23O9DANP2EO+0xkBmF
iD8ip4IK2KgiDqRJjUheFRgsdvQvm0zw3CXLK9Y2s6RIeTlwKpbgsV8SCIW5PFxn
KgBF+1tOFDiVZat+eWHpu7PEq3UzurKhZ5GCct1pTCiQWrA6Z3Ozjo7r3q9baiN9
CyVwOIBL3l9gvpXQKpiEWE57vha/3/Yu2iijd04QZfjJR/gcZXsnGdZdErUPvt94
uT5dONj50ySzrf2pGPBx0tLE4BZ33/I8SBE4WgR9aCeTjS6bELDSq1MqiIIt6goc
a9AaWh0M5Msx7qBy3y5kMgIUNsWTUhK22nkNasn+1AWMuf5S0Pdl3RXYDZsDVdCG
A2hEo3psurLCYbTpqauhtbRLUzTbvu+ALBgdO6BkLVd6929ScZ3IrFAAS5EYWde/
xDHRBHDrp308ZnZayytFyE8/K/+HtqWIVmYzg3qBvkqIVCZKKrZHM9sg59wPhTBz
3cXTsXLYdn8W7REWaKuntB/+oP01ciOUMXTNVc4Ho8s/Tn51901hJCq/00vtX3ac
D+XT0LtgjuWrgFqiMwwNkWjkSSFWhq4mSYBedXaGfUx6RseA1cQB9tWc6vc4iFvO
/7tBN1uANObTHOoWR4wKyCegi7Z22LrZWm/srugm4wjrBMTxm/1LT71+XLYBmN5U
23qlKcwAU+mjLyHZxpv/cGFcBCywZ5tcrM8hCgMfIBHHJXRwHoT1HUuwck6yGWta
YozuF4jeFQVeBnjWDSjZxMOfyAlpnWR0Zg4fAr78/nIGBtdX/LU+rOTPgKoabgdz
ZNh37Md2yT0Ein1P58/PBYvxusUbEoT3Kb3O2tldwbzrSKckMM4mwO0KZbrEw6u6
yI9Tq5QURLpgHUNLQq4KKwh3XOLLd374fQ1T12YoDHEIHSLHrqAwKewuJuUORDeC
XOvhVG/Cf/MOrVT4dGwM9rDhweVMpAiENnwFIht3N/xKuAVLhsd1fEnfNaRUBfER
JQabHhZhueXjMWz+mbyOPoSr2EYKRlYdpKzmifV4ibTHxoG+zN3qE8VYIJsiaKBr
xx83i0XhAkTg524olrRM04LgitRS7T2yLIQR3/j+Qboy7OllfGC1irlh9zDR9GQ9
b44LxNikB9UDuyrwusZ4RWnDQ/uWLb209ov/ZdSM/ji2I4oCYCX/DFEZBq7tpTZj
551u2B8WScMx/R6Dpcn2Sm7sKqke3mjOyS9f9w8eXsCG19YdZykUw5BLR0qvQD3n
b4uX3UqdQKqbN0KsT7kRNgFsKsLFZ/PzGNEFbdZDM4IiqXvwyHFiyIl6vDk0fAUP
XB++p4Y6rpf5Jwt2gv9jz7WN4q6moT+/JczzU9Qp5PqLeCPZQRzWHy7kRQobJ7DB
P+zQVtNchOupsy23fmR/RcSIni4wAfFvHRnh9vN09XCIm2+VPqbPAzZBHEZBEuMd
z1YOs9DLq/YVKrfm5m9gmu4TDBNi1iGSkqtes2DXJgOVaXAzaHiwE3M//4yKUdop
Ueh6d2UDwjKOv5KtBHaeimFhNzRGGARxYtqy/4TaOT2KA/UaypKuOn+e9sMI161l
GndW4Wi4TlrBtUkdxjuBHicEohyyZe1tD/cUTM8uTS2oXgcHzj3DedxIpEzGN7ez
Q3+r+FHgRo+ZY7zKTfMGGgAn59+67I8rlyH4+Muz4uPPaIek6t3f4CqvwnpPQYpQ
7zJzkJ7JtG5ofhLgrkoasSAH5jN12R6GP14WwTADWATePFoCsGssUjJwSzmhZQzB
+noO6b8lZn8TYG4KGA65AZIQTPlS52y79GGZVKnpavd33dJGtSLC1qGFCQZw3Zp5
2DGUxKYwHnir0oq3Ppa7NdJcEEk9++TeqlRAI/IjMcu4Ksp5rI0dsOoKujqu08/r
qHPkhFw9mha6PmZU0D+8jePeZ5dMA3NcHmi7/QQNtESvXPOJyUJxeYBKeP7et4nf
d1DiHN/Ubj+IzoDphha/M6mNdIIpeW/67x9WPuvBX8lLBJCgHCDElYduBs4UIjD/
S2ELtPb5J5fzBOHul8W2XdRwNhFESSti/emh6lYQ0yNR+E+HF2J6D1abyeloka4i
r3nt2uTSVVY9AiIEhFt9yZqMAin9DMtndnJc1EJEbMrc/4BN1Mi0dlQ4e0cX6fbA
Rrp3ulPFlg5MFs6BY4tSs2TwGthVFdjEQI99GtdetjSC76/mIMOjmSLt9YI+7WiI
oMNxwFRQPWJ3pYriW5hvtBG0/hUncUO410EQuGyW6EJ04NVd1PH0ERWEGFz4tldQ
FEkHzqSTtdjhtqkgK3ZvkyJklnmQSYwtoGsXbYe6EBF7x35UYI44TPfpxgACQ83x
TSBF0VEujFowB6Txs6oFjlINOGsfHevgMsgYXyDLAmGJNHQeteb/Nj7xZD1A2On7
GObqyeNB3WhTTOHbvVMUzvlhREkTXHiN/ATE+3/ymRxQ5J+nPImNv0eN9yPWcZx6
o9fQtQBS0QfjgvoRpRyQQs3ZoGGETTdz27UBoAYZTHdA/trjWHA9UoVOkH245YDY
tQWStLA8PJH8Bd/VpvdNllIFe+tuwFBFZfqX/rhdb4KTyiw8erHAHhvRAREJp22h
9fjVqBSXp6+N7MJ1U1sZZjPhPaou9QqzjXgl8+yvh4YhkADXgEkgYonY9wd4uDhV
Qhmn9AWmR/JcAapp4LaLOhaopLb4MWMpdQHW0Y3bEaMLrKFU4XikNkLBPpIwvRCy
KibYyNXXkWhHX9OUnTugn8sjv0oBnHK8jtC7VXLsrq/XVfjGkgx2UOoHezv5xd9/
LLKAFd4O0gtwDl9+vSD+sBzVXKFFLVAIAP9hBsGXLysBWH09GUwQBbIej7YqznWT
2hdcVBh/wF2olwsLY8OV2DP2rVhFr1YjSfaMiqBgkhFJV5P+a17GptK5Qe2SHCRD
8Ch/Bc2YwRNL/yYFq1qLqVjY/oDSGkW8KEtJFTtBUVZtikZJDCB0wWs6/i93gz1N
cDGDZvnb5RNZs2xDJKq9Fyh7FfWeqebVqvRylf8g2eBfZcpXAZjSMqodN2hNXWqV
Sr83saP8N1dk1TRRlcEgQBOW7m1vJZ84lCjx1A4Q7Gmn8ko9Z9SVMftqSpcCX4/D
GP3x1OneS6nJn4VuxScMxsi+wQYmRkiAWBYCy28eD74Nowr4ueZKl1di9KOvWUjy
9hPmH0Px+WcIoSWBhgxKYRvGlcFgWLm6Fz8WpeV3lmevS/sUNTiRX70mCa8M5q7D
YHXzl9gGdKSx1b2ksj2O/OrJa6Sd1S4hvk3rBf51EiEn2m0nzA9GLrzyHiT99P8S
gpxuyVSbu5Np7KD8DyQrYXN/trjbd3BdIQtNufQEC3b9yffUKSB3J/G4PeDPw4DE
scBn2bX9NDrckT+vAGITc799AorTqt8OfTEt1tUXyaXW8OGsH8qtihTB4dpyDIVQ
Su74YcM3myLFxzi/dej73BLuGNSqavw3q3vKs2D8yZGdRWDhv+IIzhPErejMjiOn
th0eTSZRV9R8zNEhuaPvoelXt4HvhqOxI+eYVFf3PLMzQ9Vvah9jFkBaTimijzzv
NoXVQbmSHFh/J+m0y32Ep8DySK6HKDvBA+DQDqcAm/4WYQv/OOJ0eZyaQQrG4LvA
xaM4He0iGa20lB59Ji3Kq3PxMAsaSITlspv6fXw9cZ9NA86EcWdeW3HjxVQVaIeJ
8X/LQJWSL8yLce/LhEDrJE6+k79/QFupvCKTJ20Q3sRr+CgWUB563hA3NR2jvazs
fPnXl1RiRh8C/V39po2Mf7gfb4cruGBOSJ6x858MfkzTqF9KXH5Wntzs77hteNRj
nRHSt28xn3OyMc+x5lf4r45HzkFLg3qmXvacNALP6BfH+iNYkuTcK3PBFeM7VOUM
Ua2o1crohRga+UIDni3Qh+UPcLTdMAaViSKWqTy5T1uD52tvsJIAIeSeqMnG/UYz
V8dGbdA5aqY3d5xjcNvmZtCpylRz0QhDoxCgrcUvSd7XJge7/o+GlwI7eoEN8p4Y
3ny8ThUYKSEGTa7JtnYDNRrmstbeVzortV6ECc62MS08+VXIZTCmj6xahVuZVDJ/
DhAsNeeekQLY0ix6gm9QUszEv684bLzJWuqsAdNThR3VBhcMy87RqgWvhkDa5jin
Oi2j5/qsnzUMQSgAEqDVNe2MpvuFWqCJZZJa7t/MVM+mh0+BzW+WsATIZ2HDrEG7
GuqcmYXRgqmq5cPOs2r+LLZEWiluVzB8acrMHHie2wp/iOkMRWO1j97LNpuiwiJV
OmbXx6Mgnv8XrDf1n+pWpXZihKsYHCz+EeOOx/1tsLzXFZMdhPYXghrd9h+37ba7
1sMz6W1Et0xDZMdzdJGlibqTFm2AObhrLZQrHrYrkWyCE9Q+GCjoGA2AC/acdJ5S
sql2LJvX3Y1J8/fmQLkMh0JSgeTAWC2p68bGcfW/A6b1EuDh2sWtUjFJBXJlQTD+
DYe+SSd6cgLQ+QQA46mOVO13JGvrEloJ3U0zrqzrRpOUS+jckTWCbp9VC16/zIZv
yUE8jx04Cf0WLX3Gtn+2C5mnJqCBfVuOuzxCagCadZS7wAP0UksKy/QdPAE2XsQr
Bh9FQhY7M2vJSthCnlGtlEcRuylzaue90MfHuF0dlKIfQJJsyj9QtbLReXPOyOkU
A6n87gTqtwqUqpfVWFgvT0B504BPqUIJOxlEfaT2ai27SUYHL9xtb7G9F0p7+GaJ
VmHNGYebZsTT7U+XK/RavSSUYgu+jpiMNBAq+7WwxaAEqte05YyF3mHgEeqismls
RoLLeU4MpyPLaeRTE3MZ0heZ8zdsUWXKhpKvoskmuWBVApjqe6w+yJrdtFud7QBt
mI3whytLOUdNs+d6WB6xxftHGKZWYOWI8SpaTwHzi0dcxqeIzI4LC+4dlq6sB1HS
IFc2quMGjRo7DmYdgb+pWeeBY+Y9+TRrHgVoF5Rk5ut6JWYCXaMiZyG22WB05oXx
GKuOEhBmFdz4T94nn7KEH5VJ1W7xdFUbXrgtErOs1ICgr1cM5KGEoFP9Qu1svIvv
8+R9UKcSXCnmvtNNvBFrsEeKRQzwc1CfCt3RiHtJwQXNrsOAEsRQpzPsjKJpSnRH
X5MMM6a5rq4aMciF7/Ex8qGvgdYi/Y08b4Ux1TBY/utahZEnzC84Qk/I4qAT/mbV
TGasAfHEE90TUQASvJZwD2P+fDrwtjl/pxwCNioOyA1jyLSAR1JYqUw/I6lazbmk
5bTpMGRtUBCzsvCFc0dEj58nReYHqARVE137Mh0l+z9ktJigclEHIlWvIs6Pv+g4
h5JHZmsM0nSREZcEeQTm+TCSQ5Ec1VccwoUt3cmi88mjbqzZpfjyOe6HCSwRmxgC
tAGO50JiqHdpx9jfrTa4u3xF4yYjV14ln2PdZd19FGOHKl/XFJ/idFNoKOqz+x8z
fzSJPcSdCr9CX7E/3TNreBOcZ1W3+RJEkv/0NJ7Hoxuarp600AI+yXhslbX4Hvtl
pyvFRKmLIcEFpx1OHO+kBT0dix0F5DCNN+s1++BRqguYQ1oCSIkPHG/WkrlNM4fo
P1qIv8BK+3mCqfh4MXO/l0vHK3nGXJrSdhlwFvKgxg1qg7Hzd7ygssQSR2EZH1v6
pB1iURlpxNrQp3wLK4ZDgc/pQn9vu9TECL1y4p3RUiXSH1AFfBrHMMVeuHC+AHBd
zIcmdLYTGnN8xcH2vO5v3Adnydto0pUQqZSlw/k7ZFA/zuG8KSYre4y9fyJa84dA
gG5wXkw53oRWms2WkGhgAem6ylw0hWk+ZgzHeGsQIKrjAjR44ofJSIPs4EKcetYL
5ZIcLG4EHg9r2bijDXS6yOiw4XmX7eDeTpcW4s2pQRV1egq5rcLjdTZ9coyL/xZK
+QoWdStgrcihZ7GjfSr5Bfi5r08APRmPiTv7E35CEItlGQQJ7KvXQNecsZRryEzX
wocx3I92KI3DVlMgaQddTpT2GMdVbR/Wd4j2HGuJW0g1UTwolRF+8alYleVIreOS
rXeqpGpo/e1vEgPa9dMskKKoNj9Ev7Adh7GYCsXjaSU+GEkJsNfzDuHMZ9L8bpfI
KnLAH3t5OPjAHYwS3XumTXuMG/g383fn19yHSCRu9doVdepjYxqTCTxfqWpVVV7Y
A9qi2wxPVI+D1yGySxuQ8wwEEi+ztcaolwLR2CGaGfezia9AZNVZXDWRXn8sDJqM
VMG061+lCIO4xMonr7O89jaeM9rj76IRedtOVJFEsrqxSRK/QGxO9Ujtuyde8uYI
1tfD/Tat0U/kRMaWWxrQEvN2fzf1Te/vOcnMWIiWpvPP6D9vojB9zj4q3cA7IIKT
Cx1ygqppMlIqK8ryjc8bNbqu9AxRAbir2S7WUWtA4A09j2kTqXLrpXmt7VIBx9UV
7PbI7NAJ+3J2JbaDjUtagIydgZ2Y9KKgDyGSvgRi1dAWYHzHew69IpKSk9dg5hSb
cKmVKuDPGlDzWmTtLOahp8tWmQElfn6yeqLnEa89p66sRgunR6Z5IceoNZoFknF/
Qwb2vKRz91K1tzU/lmVZguFYBv2YQ5oThJzG76MBwS+e/ZhAh+DksEXUTQHITpiK
0matISGS6SafhHH0r9snLQuwHc7bobm+/WqjfSckflx07jxRdksqC7faM/yRGotC
rEDXSbL0tfsfXXxBEPPkku4zmBrgyh09JAv1W1iaNekBlGGEzbndKXCfbAmX0erl
2ej9GWSncE1fsLXvhAoi746D9vjilXmfsLlY/6FmMMLboKnpvUK07SdNxIYUg3AL
xluWoyInOeH4hglJteK3rAbKZRzjp/MR+n6uX9AnQm50PGGUlYno5KjUu8rHl9Y8
YsqXX/2oZnFhv5Tvs0NPk2MgDGwn1WKDFgGalaYJryC7Ul7Y5B8hGa1i4x62r72R
DMPRzD7MWe4P2TcOgWW+AxslcBsuR+5m/1OmJ5ZS9c5BFyQdMSfKpIfrUnQ4udiC
mmpSiXMyOI53aZxKx50W09Whnepmxgwu+O28dmWB4JzDFJuXjzLGCxIXOlXmhZ/G
8S6Hd97HO2au4iHByR7pHcuqDKex7I9/n36C1VVFaH7hWmnR5QawkKuuS9QPcLOx
3vZgKfmLV43qcRcS/hqUAYAfFpmnVDPLM5zkUEQc+n6Eq2+J8pLkqYTsxi8Dam1D
UonzinPBfaw+TZrUcEQr7Ysh9VqGuSk11Qe+aollm5bE7dJrHk/kcgaQW/dTBBn2
7RAPM9JLB2qjy3fn+OCrjlX/1Znu+ZkRQcOtz9JmSwXntqmg9sOkpHtsJcCvA3TM
bUSQkvY1JOpaTtUvUwx7pZYovjya285zZ6eZeHcLUDTYaIXyPAlKiPhQ5K4A1AJ+
9ge4a5WCcHl1hCjONkwetB1IBLw2xqagHu5cvw3oFmk8H2Vr9agmqNDAMqADjceB
jk54maMDX5IJk5KwzgcXSWgOSHyNwziWUKi19wODY2wpGJRxn1o4yFekpXfvrSDN
XEs646H3Gg/VSDcAqtzW0s2e/4of0tgqpBWqakDGI2zi6ryEKMmzfkJfmFWVswBc
M7i+Im2bmCNJ7GAgZUyKDbH0HtPYPOsUhkfudDYCsJFF6KGE8HSyTLKCcpAQvyUH
Ee+N+6qkQgceLFb0PNA/E1XlAVFKvyKq3MHQOZajPWXf5e1Sa9aqb57zLRHHxlYM
uv5il/ekeOaLfx8tVkVuX5JbXmXo7mwgm8t0S1N8iyh/9ifCMzbLB4QS0Xxqzemv
eAZol6ZzxjvjdCFxbppedfaHS++11Ww+kBnY0uDAdP5kYsbx8+/1rLQKZxJSBK3s
ISWZ6JFzhJn7Jh1ipZ7+f8cEcNlzlu6wAeo8Cfg8NmQVOwdb7BjRgLCh9ksuaW2B
Ykkncj7XcQPwrn1woDNeBHNMJ3c77vMHDC7Gc6BXi7aiZh4Ol8bNffHRIWH97HCn
fSzL+ST6XgOvJl4QFfCiNubRWDYJBKSt/d+EJtsSxeMkGfylF5PzHt/WW0QQ0qSk
c9PZpdNXK0/XnXqSgSwo7qCt3P5RT9EUhjozszdltygAUBPQcBMcbAGMgXDtMHH7
wmW9XLzhnIkxk8m4HnNEH4Ec7J5ouFJphqHU0dNOnmnEqPX33vuvrNC3twCtdYsz
7wZOG7j5Epm+8hF10MJVwFbEkh+MX9xcdfeLaehbJL6NddnGmpBpDaWBlKixiEND
+J/oh95VDcOEdYZsd7YOa4u107ztZZNjBkJpboYCn16lth6MR/UGQpF7FmuIruWl
JOE3wg7cr2BWfWxJboQseSM6xMsB+MABdCKn5DJaA4dqCZO2IRAbwHSZHRhhpftM
DOrGbFcDGBq+ZsYToqUUkGHiZ5mO5pdKhq/QKN4gFSHARZip5dZGZEh3vJ/DPC7H
rvbUkc3ROuponyx2SwT6yvjHVLiUe7Q+QRo4wvi6Yd5LyIBpITDfF+nBeUSIii2n
PCVG8UHWZsu1IGcZu8T4RJ7NSI+eUvJ6JP63GSb2uhOF8gQsIuBwSDJUQUOP4blE
5DWMgwE9AFguJKF9xxtu1oa985a0aTbraO+6cW/+eKneloHa3emfZSGlDv6PnWl1
Mp03kXVhOPJq2TU4m/4KqwImaGmYh2ZWs0bcwCKXBcxLMCMba07NOQN54yczoI5s
UkUPvreP2ZcNjXtKGiobbgDnss4PxcQSoQTx7+9AMezkjb11JQRgCugbS3+KqXuA
7iH3xdp6ixZIu7vtJEOAC7cqKJwKe+DCf9hByrfyAgeCyX9VXhv/1BKYikg8+KE+
50DJxElTOfwlwtuUf5X3+H3A05SlrjMNL+JloyHtg9smP89PlGT214tOWIJ3gccS
C4beBIchNogcIHQnefDg7OO1TbWRq1FdRCEgE/WSEAghQHopklx6XahmYZ7lhx6M
NaWCuEJzhw+Ptljd0vCOP1iFdUAGM9YihfbyMrIh6rSU1HfMTeL6htDRuIh5Eqm0
y3Ciqw66oLa2AzG8g5bFI5qLDVXDLACNtuHqhOU8bqgR4AWY0JU/6GzjIdZBLop0
VMUpdsw7xMlqjHODM5UHgRcg4k0gT2AX5bA9IE+N4FAtSdMHKFDrQDWOwVrSUbZD
iQNqS8p8oqiHdQAqY2//uGi9fNwsybb09QcWsrXUrgmtDttijRjIYAbPYel2o0D8
qlN6mOPJAfPp5YdBGIQpygHu+v2DpJk6H6Qnz2Dhxodzfe7rUHlWSRnb5MObFDpx
5imbWRlVH/O4gmPcA7xls1py+2rTzO9Xaf6d+cQZvZDGZqZYuRjPN1QpKx0nPQBc
TOupwIVTJFg1PtTdwY6JdRZu/XWURRsrkGPjJ/aib0MVTnZwEk5wBssegwotjDOh
vUMKMI91THxFIYz56et2Ma7yB/p/5GSKf1ZEC6xrocYOFmipUFRXv5gBmznIcR+r
urU83oUUpwUDiaLoZdH2vLUnnYB9nrKU6RySIwx1wIMUog5knyUXDFbkq42kV1JB
EkulD0NnBpm3OwRww+5Z4eebGwBj+VdN0epE7WdFHXOS1vBil3cup2KcGYvYIoCE
8wOiorlhd+p5qbF37rk4CYdrx0vuL4nQUgX0s7uSkbBxMQ21S5bVwdgclNv4eA16
J/67zyIa4oz8EzxobDXfSsmC+CCmG7ijHLk+CMHQu7l7AdSGzE/VYlTu0e0VYShz
hi81TIr8f3nXkpUU+cle9wJMJhq04Uzq18UYOE0sw1+WQTOU7kSDit4WQD8MlfAb
52dy228yi9l2YWI40pZEnWG/X2fB1BpSxJB0LUsrBVacNtR/9D4J6pABllIe1dp5
29gkql+OHIAGkbpQG7C8f6XKhQeFmSaAWaDwHTkt+waUl+bJlnPWE+Qjax10GSqv
pXky/py6n1RQ+mJ59wKYBj2ylEAk2fT0dsytZhhmiuD0wuE560s8ffn7sgNlbE9u
7IP2XuIu5IvZZsHJ4ntdNF8z7DVRgX9KFX6i93+b2Sy+JIhsSk5aQznDqMdzkf5l
1MvX+BNJVupCBw9OouoYXbzC79sraopkMJAt0EW/Wq5BKbr9O4AICWmHZ0eGbByO
qPjKA3d8ZNQSIZgdmyib0Dry8B8h14bQ6zuCy23d7uPgtOODYwYljMTiTs15HDIa
jV9Wt3929Yk7ukK06Me1x7kPll+JAJfYbROW9jRMfygjl/0jCvjn7uVDhDKczK4A
8B4Bz6gnnW2ulCqS4v5JM2PwTbqQ8Z22daoPfMlETgEaCnewyn5LznFeW7gp+LBE
UJnD2zeflAMmuScwdbTD+xOFz8L+0Z6UOjyT90L5+mSCCnLzOHV0ebm6E+xZf91N
a/hGaRQvwDitmf8xV3Itil5/vQ2ZeYp2CdRSPMG+G1KwwCnitg+Ht3iSSyrYLXpW
SV9phfHNQFM7f4uLD83V+H+bvZWl+CrScGWFguLBIp0w9KRbttfXn7Cl9ehwQfau
Bp33dr+y+VYxCzJXAW3qMtaYqxVKauLj+FCMVDZhrbol8pt+dQoKfTgU3zjq4vw5
hsqmmbm/e+u0cuctcxpHKabVyaJlCXdSbz+sETQYIordVDyip99wQacbKPcPLvGE
VJrQmZZbrXtNWqJR5WySVtao1xV060EHxpX8BoJaCPcf9AblV7mltXr5uVNe+XfN
OYs3vLZ0Vd3bEjK9q3Q7niZyobfDmR0tMcsH5uWf566VCp9SGCxWuD+B4l9XLD/Y
cjg6Q/RHGhCVLoT1KEV/wHtDdUvt5wCL9vHcDnGkmmC79MSL+2lKHfMkp615yi+O
pXTpf04Og/yR/w/grpDcGYH3C/GleTgT7bT96v2NuC5m/8dEpCiNsk0ZL5riGXUW
Py40wQEcnvOg3heEVfN7DnXJPiTp4QZN+2uPj38BcfNn/by81O9hLN9BXgkTCa3e
+1rDW9pFMTjquuqxYR5LdBNLrr5GSTctuy1zNDH7ibyjB6DATUbEpPdYEG98Oq3w
ayPPvbZJBm0N/hgPEnha39Pd01v7YI1qpLHyffIdZRoG0i2H2AlQDDb3gZnI2zJz
Xrnxl+AhUKUU3qddk7DVvgq1aN1qcowB46XgjO4VwmCmg7kmypmcY107lpE0FoGa
0Tby8gTzuv+M9DQRLF35mPE9+KElgXWazjA8cErHHADmipYdY/DyprwR1k0sBluF
JrQoxaF8YRuXC7XPD7IA/zIVV27TcroOz64QOoOI6acVZeG8lORDhbQph9zx5r9t
rZLe+2oXIkShwB+FshB4ljqN6xCinFqX7UCUyCsSVcIFhaGXhHkFbp7yDB9XF4S+
jR+Tg5mR1xOZo/17AgHzcreEWxJULo9qBvQsgQ8EV/5nly2qos+HGtu0BI31jrl6
HnYiy3uzXqeOvoDhHcxEQfwwXqUPbgDeIelpn1StmKUYx6Me5nb7eR9EE5X8LKAL
HB24RyZVpCZYvutqrvaQKgMuQ8SfGpSKCO3NTgSPUtYkAF6+jBi1c9/NJOjBiIWC
3HcAuKDAN0QMkxYZYFp9i7nZaclmAg4MjY85CDStozZ+J4rfU8x9S1NMfl8rI0CK
oVh3snBEkg/9xaweidgX5f+kdxY4065jGko+vAReVZp/yTsM7yUKWS1pN9DgMUKm
rSlzSn3z0o/WaQX4xeOgjTrdj2s0u22CMzR8c6uvpn2Ka9gpGhJgkiQssU7yRot0
koa/DaOtJrUUuiG8fRk+WG+o3tiJgRJI0DxCOHKGJDO3e18BOxu5rXwjEdW0wFtf
r6dnXIX9ufDyCCk/a05eWTbb3X0CwyWwANmYBKwki9ch5tvmquJmtIPi/gD1XwO1
Eq/JFWxNcS92oROObMyn0jArydiQZeI0wqTBCB7cXGybhALIvFckPsOrXpu6tegu
a/zdbY+HYiph7IHqi8SxQLb/t1KB8mrDsCaJdGPajD03MXHbHbmJP3yqJT8E4Jsb
P3KWRFy9FUQHFM5ByQyYIe9SQcCZ01Wnps/6muQUFq/TR0N56dBAp/cy7cXkJlVM
8eru5SQj8/Wp0mBlzoG9tBf8shRMA2HbPKOI0QnTRlltCAG9tQCz9faCLfv1jFNh
8EBSHmdEnfCrJbyi/uS3Qr5ie3n6OHjvMIMFJ0KyTzjvxVpm92DeMOg8PXm2DyIi
ug9c3UkGQE9JIEJ5AZ/+P8DoR9WVmY863Rk+JChiqxrQ+bL2kGCOytHo0Hojpaiu
+vJVChzFAprVwShMj/KyFTOZwzuoRMWbj3c5r6/skzCMeP5KhxTSFrAS4O5I8bAb
QLuEsbJlasbroodQyB9t3e7LeuKFlQzoyfcbb3S775v8xuwK/99jzYT6OEIVJrXn
pJc/Ofn8HmBiepAaX7qSPugSMV4EN38x4GWVqWkIjEoCZQ6MtLHzpuL61M2nnTCR
6yNsKG2p7nKgMybQRauakYJ93tKf5i3h4FVvGyflPKy4UYkZ9nwIzN2rkQAEYsdk
yYWotD60FZf+y3KY6vev7IKNBDAsVvSNjZCWwVEu7+Cd98w0qR9zEiprRgkGvYr9
3U9SM/DGEylPVeDk2MrTSxawkDUWz+e0SuxQqFiW+ZbDLFGa39usvLAuInbltddS
mKOpWrIUDe906e/kISpE6cn8uNkAJRIpkG4Zjp3+TZWX6nOGW5xWK4+d7oLpbG71
4IxX9RZY4JV5XD8goQbAQUVcGIBbWc3KWCiPc8W1ktrvE1tA2xWYOBYy3bNQ36k3
2fVQaoXBO60WcyzHKH3dRwGt6sVEDn0NnGK/ujIwLYPtRJSVYkJmqhi0Lolxg2HD
eW8YH7k+pQzWHYFx8i2yqKuWuXXkVKaEVpsKOZPiw1jk/UyVqLCa360ocwU8XNyA
kAczyK2O1nSr8Ra2AtWUiQzVrQCHPJNJ6SqULyH4a7kwxioBoaZ24V5ypnBC6Y1k
g3523Mx39pxUlIyD7B7KVQ+GtgZ895ft8IFlcP4czgDhNjEPVYNTg36t6+E8gP9u
lbZ+08jDC71MVED0jdcaL0P612inaXQttjPTu7QOUTLWbEIfUovG6A2LnT3CpCYg
wQK4M19Xf4JlQFsA3LbtgPQw68WbSpAoEJDi/L7/ltWiOH4663fMYWYuEdRX3Yhm
7TL2utB16FJ6zr5pazbF+BTwXoAF4kIVIbTrDSdtfMsIwq/5h+bvCCsqAPbghpZb
Kujbey+Ldh98CS/aeLB7kPa2Lj1KhNdTmYXXum+WG3398Bv6i4OyZr76IkAlR81T
W2JBn7KIlJu74FehRXr8u60bC3TQM+VvugkNa0WPQWBdReihx7Ncum0VGL2KLdcv
+98Xq7KO21Kd3+KWC1RPIOGa8LiTT5KTVOTqFRwV22W0MeK4Pin8vqcWbPuUuJXh
1rIekoTyj9Oecd8dSeIJwa8/AUA19odkCAN1B0wbxsP5WrdcTQubSNh4isw8TBld
7UQHT0hBwewy2eAmVZrFSvLqw3slhwOLj6+EUtfPR3COA2492365Jhd/wmXc1H7A
GjMQGzHvt83FNbHbNNF6L2Mig23WNWwRkRC98a1EwyFaPxMLp1vj9tn/Y2gcdlsp
gwb1gbVEM84xcLRwgPEBu29iJorTUex2eEDgjUKKgtUJj+nU/sg0aYpAvFqNVrjS
tgeAgBKkEY6I0nfCaJ+mbABZAAtK5EWLaL5KxYGuRQiMHxVCjfByQNxj1IPcr8J5
q3X6kl0FT8jgqbs4umf1tYiSNQahJMtIbD49os676F0i974Yt8WfU86BZi4LNl8T
XSHir/QNLTvGUzmBLMm577IRTBFDn5gCINNpbb7Dyg283smox0uYhPS5CmaLFGAy
lHgNmbjdQEMdF3CNxwSLWBodjJyAXjGW1CJrlpnBX0Wmum7W0NBu4Rz4hiu39TrW
qRUMXXxilXd3b1YpWHq0SpgRnt5g2Bjk9FrT4ubpUCX95FTNZhBz6/8KoGTMUVkT
LYNBEvE4fyBrpMQ8wB3WmxenGZFZmWBif/H5DJvLEc1aTGIB0lbaQgcHK1W+RVzW
VZ6NIU9GREZ+C6HRnlw4jOr4D6ab4hoLg2ZFepiLYRr+u4ckSaQ6dNumbA4IC89i
kMuuTHgfsbLiN76ZjXEtPEBGiLMNspYYng+4wrdpniu+9yKk4oKi+KNeKnvpii//
2FaNAQMbXagLkDe3P5nazPhE5+cdKPdUgcbCO6vRFIavJc1lpNDVkAm9ZXz0PjqL
uo0tt2BKrwh69dEHq4fnzOAmtwbtcjdfMPEsdy8WwhWkCPsNEcD7j3UZb4qQJrW9
Kc3U3YDjZ87At6wlGmnFAG1UvQwt2NvPMcO0o3DTtAy1qMltlxD4xKdXp/m4mLrn
B3Ol3gdC6r5q9JSQt3T8H1xlN6hX1fSq1snsfaEgQn/X9sQ1tHubiQpY07xZUE1K
olmyZ5QTUIvCN2Uo9yJc6kx7uDx1pL9sNAi744//At4HISLs/VMNjwfgMsmUSWem
pZn+LlECuRLt8iMSflsVwfUVW1f19HJBjCoESLMATvPqVxgNc7HhDBSQSIDaWvSy
63Z7Sr+rybQ08Qz5ZijyOFuwibdkHWvjGJ/cv+nVD1+26FW5aXKnCluC5QSHFtG5
EAKK9eSxrvTKxkN//4mYg46RlI3IASy638QqWNVKwyLX1zNzV8rtFxhcwD4/yXNa
QWAVNVnigXXj/BuicGswMoJaK+0wKuAuvGOjJ8W3FYZ9JBmSua+zY42WhTl0alDw
W+UGATcsKGyLlu5qjSAV0LMML0gLwBFCgFH9MzUKSq3jidpv6iuRpoceg05V0vSW
kLcIzHqXqT+njaZrl4ou3/pJrrbNgShWi2HojfZ68HyYxIdJ5GqpX6H027b2ecCi
DDII/PeLm/tMHh8VFzmHP6ndHf7CL9VouesM74xm1zpA2AJjCiEhdd8xnB9w+65G
P8S+88tAtbXwIFrNo4AmQMHUoVxas9UaqjXW/c/XAJkyCUH3847UPYjIqaDQTylU
CxbE86bJsVvuWUu1e9lmi2i2oSMD4iqVF5OgwQy2b5qbJi8z9oj2MNmjBiGVNHQV
IIYXkjO03SsRTdlpONylTBLyStaRmKnileBOpjZS5l5+6rNBtL4LGkpsrz94C+KM
W2/2lifxpd/QSPXlgPUnDPHTPkAd+T+SXNuzOMTGuDEXwo52a7ksvcCng6LC/dQD
VphvUf8Qjx26do1eCGCKY9jpHf1EVo5cDq1dqLPDMJhSikohxr0hdToytkUMPAQ8
qq5ryunNwZgs4SC01kgu52CpC5B1ehuHaj0B+zm3N2QpMeRPzFemizI0VoqP24WX
FqKhDS9ZZKi0tl0cgDGybO0+qqC/f95TN/6DKRAz8sKg4WKp4CfAmZNCBAQUkD6Q
0edGTT5C4DMLDE/4i/GBqMc7ARNM4tlUG9FOJJxXuppi0dTHoppDXCozpJwsGqdA
7kH5zgtQsFUCJAPim5FwxoA0yxlpDl0bi0p940BPnW7HmiUN3Ewi3ZycYT0mrsyx
vMIjslXTbc3ai3NAMls6C6OsalT0s92ERTZ/o2Z6Ez3Qh41A2K7/kOxf2zPElHhG
s2fcQoSVhOzdFad1VkCC4RprFsJGm5/bR9QwN1XYhW+ZPoZu0igKFCEVqmNQxlXM
OGQhaMI0As0CTscDKL4ImFOnUfJmco7sWwqqbN9IYftXjKxMIyG6TV0O49oXqn+r
uRp9xnNYt+byU92a2ACjDRkHgaUubeKGJ3LV/SkzVwwS6iQL6o2AmUf4dAYNbqbb
3kVkYoob388yeZsKLh0SXPQLCZUDt92k0oJgO9Sn9chhszoeF2jg3JcLe/OqVjyM
XiJTFr9ldeVR2vhIj5IICTBn74Yn6mK8d0ZWEwV21mcSpbiUG67+CLPWJ1ES8Pr2
o5ZsUpoSppkvoD5BY5rzkW5NuxXArMja1r3XUhvtSgeVCza3FihSPZzGchybB3tl
fTAdSdvWLOe0cECXd1GrctKSPINSw4RCmAR/OEvu4TTvhhhL//UXN98qdQlZ0+BH
zaoBMexIv1gkBZraY+MzFuK9BA+1WI8sZU/wl5DYueAb/z1hncV9HbvccOSAmkCt
+jbHIE+RMZcHwfqfgwidKyAU8gvwcHW12G723O07TTPQlog7hndPCq1k+4T0svKE
xG3pZOp0DBYjV6LxRhe+nzvlh57oAkh7B10Sk7J5HQ+wChurajgDKN64E/Q3/zxH
pC5jh0i4jcKgXaEqOJnpvzH8ZcFSESg4k3ejSfiUBx5iSneNkFLg3yYKXPShpNXF
41KvnLq1EjS4LMSuMOBk/SJlSJl+2aSw3GnEb3xp8PKbpJCrPuy/6Be6pXJg9wlR
kDB5QarsQuzqYYqGteh1ziDQN0GwA2pubRDO/fh2Z7Mf8WnBoJDQ/Em1XJRuEdxf
z0YNpkYdecZpQbNUvOqp4t5nEOJaMbwtDR91RBgLx7/L5MF3jZuU7uuzoOpFlQEy
avN28Gtc6yfj4FY3oTzUZIXhTyZkn5jD+U07DayHxKbO36GeJfSvJtbp9Nu6WzH4
gRKjXcqJR37fWD6xL0Fm1IWSWK/yir6BzZHfzNyfNgI2/wjfhL3fmYefJbwT0eNP
NtZ9vH+dIsdmp5w3sGcxIe3J7tbtfHEbXmAyJ1exzlDylDb7EqZILgGjYmXGVC6b
bO6Ne8GTbkoynt68DpTWkIhwxRVyrR7MigJL1slQpsN9o5QuUSayV0KrhVTB8HCp
2VuQ7C7Nhef5k+5FiFYj9VSDLRgMmes6CB7QUVp+us9LzCfswGr/7HseyagxLmuB
lBVnHIccBxOudSoHFguAZtLY1An+BxXDSv7O/kzRUCuuQgNnMOFiwO/aA+dOT9Xr
QpKC1PsP6YRt2q4IgVDmiuyHpRbfzZj7XFdKzdFb9yssSOoRb7pC1t1CMjpRaZcA
VrHDT5tvUXfpMLNrDyuFKH6HlLT6d5v6fTAREZEyZgUCYrlZYH0rto/9MZt1mgMe
/yJjTEHnqW71LC2tYXUbcVIhvq+DJEujVpXpq/GZUw3uAiXPpHQ6tMLnK5u6fYWT
jYktr2Fhagn0wlpoyg6TrbCKdJkyp08rSfC4yxnP0YNI7YBHodXqObp22dYtA02h
PMBFo8F7ve+GsjgD1XPLAadeKbhbkdoXnCw4aicSy339YlHZfeUTBzQTp+eBFfur
4Eq4zhxNC2gDP0u5hx5S6y+Aw/2GKJsxiuAPWARJr0LCqTHKgWgxJP2RxHqVDXc/
n5uOX7V4dhBaUHrZv7zky1Gkd3DnIe7kD0DLKfB1GRsLGt7DskSpJRVOvhzC2Vui
8Ne8jZthBJOGKSUfUajD77oX3g64Q2PqKkHSh0SjHsw7/0OFq5GIiiVnuiVzEiEw
1vhXdTBYd1BC0WlFVWQU+dxGdCloE8FcfopnCCBPQBM6LwfwaEuTkfrlp4RjLyh7
JsdJeASUQ8Fw2t/0ZgLTjBasF0Bi/+6BaUEdK2kA9vwMciAdo+x99Uyr5hUXPneM
p7Af06BA6HcYBPKPdt/IEggRkEImFJbSPXy+5Pbw23JANT7llSlAcoTM6mVI7loT
p99XvltzInl5PPIiJUBtJFI08dssAbmPFt9G37H2WU8bJxESj3g40K1qjTEOChSw
JiHlYL+nbV3uBo2ENjgHUBiSZiA7qT8YWSKtQVrurIJd2gKjhrn7IcKLgxN8+7FD
nb2fUMEQ9ie8uUVpgOBLcUgEyVcPFpTZD7tpVvf8C/Syn5USOHy7Dc0Nqsp7A6XR
66p1yITxwBN95N2bjtnSkMaOrt2M3+aus64k/daKR7NgtGKposlxBXoOzz2jk05i
UqaD73K014+BTlNmffJb+Q==
`pragma protect end_protected
