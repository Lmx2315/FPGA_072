// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:32:32 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
UbLcCubzQKynlTVm3ipecvjqPfXnSEmFw7NgNqqB9wPRK3gEOWfRQjPVYIepLi1U
9Vxs/Ddw6WqXhGRUgQkL4U7hKUXW5JETzymZpgXLySb6lTAzDzJGdZMX+ZEJ8rgc
8LVlbmcXoJGB24Y7yn0qxFgGwSU1WG4J1e/sw3jMrio=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 22480)
65GuL15pc9tr/dtaH8yeNUHI6Y1TT4DixCVPrApzag5IYuEgcN0/uaK+/0sGj6E4
EATx1iyATZiOZ0gKLKtK9mQi6uKedcgZWNq8V6xgpZD0xFug0X1xGIO/cg3PpsXz
1AiaG42KlB9QjxJTxkzeYb6K4dHRaIGZmAqxZrGMjChjl0YVR+tPO4dpuPBoCsk8
u4/Bg+EWFvT2LZz2TrSbhpNIAgTYUdJtM1Odu5d8adj/Cyuy+vUki9LE4aU96zQJ
rxHmUTO2e/4gS6mbgZbpKC+P7yKjU4MTPEqLBl8d3BYuSEtJLX3W/Wbgiqp+es6x
kmU/0tizYa7plzOFcMkUDkOmMq+bkt+SKgkblAlhiik0+vwmuxxQl+ADODC5C56H
ukWTLAQnXJoqPoFHuTW5wObnYjArbyZP/FkjAuzN6Cftpqo/L7lLhGwY3i3ETA/r
8C8LmUNnsUAzC2RWo5HSZMYfGAp6IwBDgPqD4j9tjVpqjS2T2NQrtIY9AX+VIDjY
mZT/2hT2TYuZJSsNeoLgOW4xmSoLr1aqHEUIzoI+NnE4saCkSxjazUS6t5WHFsx7
UK6kfjeKpniy3DrS3IXN7gdqhKwtYrRWIRwl6HVDWcitknoedHcDRF1Y9knH5jIG
jtthbORxmUlKVnqq5EFFwS7DbWWbhO7aWC85om+moKk5XaZgR2yuxu2yYQB0D1xB
Xz5iOc/2GyDKVUCCnjNDEiOYHNL6Hmpnl/NSV+CTocLDspD1lR4HWnnpT/CRY8Eu
9juanOBNxIA0n8GDsT83N4vTN3aJboAyQhgCXRAInbuMPF4MSjbLq5BJ0WqsrMDi
H8d77iKw0Hk1hl3CK4wMj2I8fRThBS9QeT+XY929CGrtvHJ+sJWmCEJ+FkGi5DIZ
P99ilQzTk8FsGqK49B7R2UZHgbKdIeeqH2JGpqT48+uLeb61P9RWT1Cwm7vZU/2R
i6NRczcPI217/MAjrYtcyoFjgA6eeSaIznSIvoW+SIZTpZZKpcKNuaGvrlfguLb8
VmISRzuJynkbkS9EVO3IcJS6X+O9z8T0Z6Tqq6kUR0/Z8e6Gs04kaoCmRTM97OkS
LtJexQnac0n86PK4geyf5A8U1fXrc7J1nghfjl4QVXpwcCXXwxatg0hUdxYD1Bcz
i7EQUyeqI7AeCIEX4ffWLYp/n2y7Eytx188H+veYClNH/LHOHJM4hMWHk6921MYE
56kfT0RoaJ1A7yII9WWufAI5HKPaYW/QKSWzGPfMdQbI5Rl3vlLPcwybauxI3Tg7
+eLubcpPxjIrxV+zTkbRCH5RwgNPsS9WEEMzTivI4geYSAIPeldkwu5byxymipzN
DChQulBu+vPJtg0hBUwxcut8n+f45s1qLj1mfB5DyLBNWv2hCfT9N1/EmtUmClmX
bdJP+fjuNY7Kn/9DB5sLznVOsnIXC4IVLZdWhV7C+RqmQv5+cqg4b+5K7aUA6vqP
lNVP0skr1HmEevcTbtI6X7qvoerIVk7WPs4qcwOgYlh4YHrpI46scyjCkQWqtJBW
4FvXbivHq2+lSbNb9+yVimOcq7k6TsmGt4IglGheYizPogDE01Hqrh7QDsyJNJXT
58sTWTLX9Lf/VnOQxv4RrzIPyW2xALUhpAkDmSZ8ntxR4QVSpWNQCbUpM+YXagWD
4+xJLS55+YMq+VwqkvQGwMMJ/kTbugW8ExNDQDh/JTG1s5t4BLo4hnNK1lx0BlL3
vramDhw3nNK4LZYSEEabR8NBERf8Ht5KLOFqEGdSKwaT+lRUi6jerY1zJgMWT2mu
u3inixM+TZ4iIswVArOVhTMsdUsjT8lnYKulAo9kbmd6w7y8LMPIUmFSmnurAsxC
lA4iQ9bWH8oegIZif+ISDa14qAj6GfRHEMrjSSGiIQuJssetN+c1OHuRm8FuCIwa
xeaeTT8gU8MaiVWvQWObo5LhCJKDCRAUbd0oqfbyJx5/JDQh4DHuDssFojm7YnJM
905lPYkNvIyVzsOn5EC4BgMfXZlkMlEzVMrrlun/KiJUCVWDCfqzNlbGRXSg3N3R
VHJ4HzAxQlFuQ/+ZMlWJuxcHdcQMZ6I+YjA2E4CWh7nIo0itoBkkgu6SXDX4z3+R
zWz9J2njafaWA/6sig0UYW4knSoXZOUkuOVJ9lkroJ7TRsNdA8DcXLjPtPtxeJM/
Ac+Sn82guJwDckwBnuAGL41f8czpvvzdOfqAapISfYxCnz8yGxg0kypbVdPBu1lv
ZXmT6rut857IE9UEEFVKU5iUT38IOsOLBTAdT7wZde+ztecd7Z8E3Fx79apyEdzw
PABArZLpna4c4+2ENb5e9blqnOdwnABydm36VHBMRcGS97w3In+yAhczXw/qiAcy
71X6JvnbxBsWoxPgBvGXT5xjRmxttdPHHGcVFssVGSvaIWlXMSxgKY045qT90XV6
SJODL9rfT8pVmqqwPWE14L9m7mxStA7ciEcMiFUwKPdlYwzP9fg72cU4ROfZWpQT
Qlq/kD2mgV/mFcYgUjmvS3gI1Kgm527IXdnwBMMsFNIYIXnEXufa4DFKFHFKmrMX
mhGsrwszhkuMAyfaU+TLULkEvOhXt2G36PMk3vXkhslMYkxkqr5Wbu7ObklEvWXe
aUIUMJJgqVHJBiS2NlC+/YVKJDHD8AUS6EBvbFU6faH4DwI4/l0zUy2hze975RIx
CTgihzaf90gsSkHyrC8P8r1KEKJT/GPcak1BUhzWFC3nQ7YciUctGMeTdXwGmGIm
QqgWNAlsbR/3RCddturXJCVQ/82TPwwRhjDjfHokFp2D/CZNIbg9+0NSM8kbi/Dx
M3YPsp11bqRWiHT46FSzRHoLBUHaDC8tD/DLk9rM29+MBh6nnDvsqozbniVR7l63
df5Pq9xRbiTwEQMsktrRxdMAm3BVgCz0nzo+j4GXcUgrA6rvSuo6enA4Wf69Y376
2exMFWasRTihL3pE0eObSVDaqmpDfsLyvFp1Xp53PeBugX/XlTqn5wnN82paSfy9
0tZmT1g81BtgBTo4StGYZdm9JGIgIJwJeq3PafFUI1gTc2+NTI5CZgg/f5YMzzd8
8HqVvfmMjlpEmULcXHSawTbvz3njmUDOvLhOHlDkNdDR5NXTGJO7dsbUFkEXmWaf
F+EIK8moxEcGm5CgjyDHeUdY4ObkJlwphwi63Bq0iJuD9m7CnTTrtSHR1LMc821B
/eH0tbpDET2nOx7HBSJQygyHl409nHdyH6bpFx0ej2ecVsv+kunRTsiHgos3uNNt
O8IAk0fI503S87KS3bcnkDBhDad5VsNIZvXoartl91QP1kI8ktRAi1I49mESgkyC
1uptv4F8Q6OdZIyMMo6/Wlj4y0Jmu6tqZz5D/nm81doVeQykgDWUB2iZNGD5AfME
mMgjkCfjT1Pb2arb5Nnmq5aYJl8K4ykHhZZIOZ1meR/PbLyHCvi3A6xVyxTHZtNe
xx2cffqfj6a1uMRO2QytQWyle/eDCnM20QthuFQctEdd8Ftec6CZuA77zGa7Zbtx
3LN2MbnsZhIBKd9ASCYtl/0lBE36/j2ob3XCrNiCJJlQEG0viewKfQ1/zWMGYLVI
kYxR0u2PEK8I7iKaW2g4I3LL8bZbD2KIIS7na0qJbMU7p+6iJNa4mLVh4Gyj/+6Q
OutnNLA7N7C9cEjOUIfQPAWSXKM5D/fEqL9ESkL8ETHOfvUWY2725Bp34eND8eJ8
TN6o0eGv0zPeV0PNIGlTd94otRWmoc5GEGucQzf++OupFPCounhU76X6zUL1ihWl
FQbGB14JOs3o4Rhzy5kyxA+IjSsVWKz54I9WqwnNzJjTe//gctCM2c+pfrT3PGik
GJnT70UU/rwkHs4sTDv9d6w7kPPyCFhMRqMg1cdJivNpzXio2mQhZJCFA1RUHjZ3
ivSgUBcGctes9oJmbVRy0V0VEhNY5E6/TKd1slbM2Ih+lITYqvW2Ipc8kVgLy7uW
yU7jcRK9/sJVhQyoRBNMtcDmYeW1Lc3prGouCxzwSybwMc2qszLG5jY1C6KISa4m
ZP7HFX9d3aUU97kQDTWTX/NJLy197AWqQgRzXgrACKegFoyAq+oNiAPuSVwyepWd
eG78Vz0i+akHwEAA7jtbkh7Z9NChxmPjUVYO93PhJlGtjxoZtd8RQQGHVNqGYLlu
AF2YzAfobskyl+KHlSMPSBIAr4t3mxYYoO/ZRyLdt5q6eFSSJ+gQeQC2RpmFZy4R
XtH3vN1NSw7kMDyHIGd/4K1edXBwBaoOJBy3OFgH+IYvDB4HGVqHeg5NObZefmaw
K4WjTbeUEZuW98IOOaEB4klsFtofhnlD5y8aGQZjYEUMdxst6NuNHD35E1e0JF5j
tOjOYJ3aG8muSgEsSl45sqVGpWzHoEklivxSDnZYmjln8o7kwurtwEqzGWwoqZwg
qBlkPF3L3ckayrm6VQeFfwlQcl8dUrs//ZwjZUH+/F2SaQrdlWsqVNcBxeuTWOon
5nHTZNFRieASjCfxIb+yFVYsf26+0ZTS+aRkrZCkOA1ck1MoQGLSAYstampSDrxF
HHaKSdZNrPdChJl0jpzXBar96ayOhE18/h95WvIjhY7d1h4Zap/nBBCilg/mn4BQ
7OWoyMMeFH8YJP2Qw9qvaP+P0JRl8VGtYf1xhVOFLImaKBPK3IBienQXFXlBL7/B
c6mrJiw+PDLwyHlBxeIoUFQXiLwQMsVgLYATQAj72qeXbSDyEvXhkoDRthhmU1j3
mCngzY97TvIHc5kyFrsiuSNr2pqE5QPPONllFMGNE5go2xssYkkl2aAK3c39+5pa
jXcXGoAUNfknytV+LjtpaNNtBBuJsKHtrWplegYW/LXBtblxuZOQABEk4o28VjpC
CQETmZeSMfBEB7AEoJ/mn4Oj+1OA/jEJUA12SRFHby7Gd544RDkFLQn/hOzkRX9e
4DnENnM8rmMp7Uhh5RaptfswlkAFZNYcZwNoHWqCYi06hmFKJ0aEx3PRbJUPwhr2
pgGQcRF4XG3uVtgiTfVrllph4xpTIxgWGLN9MZNtPmbZ2OWK8dfsJSJjFgGPpJa9
GE7RG3vAVDg4EQ+GdYBgYE/nIb3f7P/DKDadqeeGmkE0yU9lmDUVLtlZOf78ZPkc
ZTXQtWGverzltBy27RzQA3V/0STbwt3oWPSzCx4KfS5CCjV9U/9fouPpmRZoyKvr
f6zy+j0d7VG3Bd2HReB729+nK3ybPVbjtd5bdtncBwOSeo+Y6B3OqTU4aHMiQ3jC
9gmGRSfNPFi7U9NZxRWCPUk+hnd8NJW8Ub9/Y7sKDxI+z8q9moNzMOVqrQ27AeOc
0fI85HNWDZdPNwZ+GNb1w5h1UW2c/a8XwlVsZB6UILePMZliWhHPNnpFwU7uRZsy
E5ko0HcwyjpJGp7cM8S5GPFow2vfTo/UcSfBMcKqDhLAHqoFNVYCyH0Koxlg5BlT
Ur7EvTXLomTiUo3/sD5ejGUDWrB1T/6c6oBMCvKDsS4ygIDEp8Dvim9okHTDW3ia
zhMj6uN6FYCuRfciWT58O2rU6P/uflkI+Vw9zNjVp4WWhL/10QHgafeazBhqLVM5
WMrOW4eke97EZYkRINppx8hOoxpCqZrK1TK9pow92tpcd9dB5wqsYnmdtMvk7NT6
X6/ucsKsr9OwDDYqxNJ/ynXV1WL+OV3aO2QwgJuHjxk0puKRIRcY74kW1dEw5RbX
jaa5sXnijlEhgrxVJk/mw1lig7b1zjDWjMHxK19M+85i7SW5wa3ckLZxlRltJEsf
VqtiHH8XnXi6jaNFt8MCkpPxbhAkxC1/C8SZ1t8Th3KcM3JNs+KKYoh9QqN1hLRO
LehxH2XMJX614BMmRt4igpi1c1c7R+7l5HSFw/GR2FdgGfB00DaLoiyH/usGbJJn
gFjR9mxfoPzjbZlju9G/22GK2GxtJbyy4Vu9kCsQVAJde7AZKkg/m/67tzt8PeJx
4SAhEhHbaLckNVydZNVkAF/l2CY8AE7UWx44YV7IxOPnSQOqDmJvTB+a3XfWhOdD
OYGigqIgbwl3k6sVL6hHq8za+GJqg0dDQqCdkUdRPnG5jEQxmkWRnbBfSZLytE2V
D/7XeMwjnxQ1yKYA0Bgh85ifGjqi3arcPkplm2C6MK9q2B42yHAsJxuPX8H9fRJd
Nu7sYuYh+PAY3ZNyI8pDD7ZX9Ne2GE0YhOQuYSnARu6/qoWHEc0SYaA3BB6WEpFj
Zc7iHIWzhzC/COIvVc1v+QUBttDaiOc1S6SpwZuNo28CLKY6rPQWTXcUgFftXmtG
LP4+zHF9wPradb1RmgM/TpGz3//ML+Ag9WKCvOW3zdJZ91jqkezqMTVoAazI3WgL
G+w3myWRb/TUnfK4FVzO/S7I+BbRwJLKPF/UsfKMZRPBJRjBeYkIaZ1a/JhpQC/b
P6XZ7aeIZSc1E0ZwzN4s9XuoGJNH2lhqrgRTG2UuCQLA7bTZjzVasbuIQcBllnZ2
GpLWeUx4Qwy7IO0/nhQ3dPh4YL0bZhmqI28w1tH9L51jzQl+fG6g4Roi16jW2Gfa
mANyyhPzzv1t1O6K4fb9tb6V1ZheHF2Yes0lMPvklfTr+bvGWK3z42ZxxAroBwT5
3/JnLjs5rr8ldiWA8/96yS7ll4a29gTRgUD1FFyKjzv9HIPqWT6Nrhur6srjfQNd
/DMu21LOolYiXihRa2wy6Evf47QuMia0OZbEdsRE5B0wOfDdz5X3USFy1CPmL2YR
yfRpTIXtRGhtiS/4amxkFm2vKL2/iMuL7OKGDbMuunySQHrzgjDIScsTkP0N+Sbz
63efH0HKlTQRReby03Lc6dqe/B8t/xFXMOkWuwieFzr9HCJ1/uPJhO1MrOH3S8L+
v+qk/4qnP16MLNkaQ5Hk1u2TGVMEuZOmLTekYEIVTHQVeCWI0T5KenzU8h3aTSnp
1rTTxlZjFPD2vRm9kWL7yYfnPEfqTiYlu/rxjAXj2QyY4w81H2lchu7eVpqG3dqn
6HFjf9oeHF3FlKf6XwolO18sbuExIAZOOWDM8bJnubwlYc8YNzuJ1h3bvBqHgpTL
mYQ9d78D9Z38GZ0u2AJ/4N0a4KQZwjl/1ZWQLVUw8GRKNmUU+JwjjRDRetL3b6nl
fyx89CMVJcSihKuJkOpixmdhvNm9g5H8TeRCyPNf3Z7DhN2w57Cyj59nxJbNmxTZ
h9u6+wqexvaM24cvRuQDbdrlp/ffVbrTeyvLoyGDLwtzOD0Ld37oWMtzQU8zybMs
dJp50e79NRdNrnGnjTocJzPsVDslFrbbvlMF/xF6Fa7VWAXmsznM4Kpq9RvADKNd
VWif1ii9jjzmFN/LnyEMCHRyqQElxFAWqafbMCuqTIyDVJnzcayPWyzeByJfsdJ0
lm3vZAl3gszmyfKGKqTybcrvYljjGzHW9s4/aISJQ5sNt+qaWAGfE1PfU10iVqPD
Z/HopKPHjukvm8SrkUuAifLjKJkJKq250DLG4sKVQt45JNNDs3Rakxio2jqVGKbb
YqgLHw6WE6dZOy1KjfLjlx3ED7Rav9y2fYI+//N5bDCT/qMyBdR39Q8KufAKbFx2
KcSabWz9piy8WbM1/wia+epDT+qBNKRL2Y3OuK7gGiuWFU2K0Q7WGyhfKC34OU3Y
0x26ENND5oXxxUkeSfx1/I+KIA0dwgFpnui9B2/Fswyc0vghp/6FE6GA2rMboahk
pH2RjleQm+f/0NOTCc9FBcDjS7Bxnq7pRycSP8cswNBrKTILI2VzDcuLLAf1fh9n
trUeMUbDT/26wEdl44iTQATQwjgg63WLe5Ho9PkCrg9R0MfNriVfnEBRWaacFCxG
LLUSjmHbu4Rf2oATjY2B9bgDbLfPbwqUme8z6Q01/C8NmiBI4oYLupnGDayKP8vv
dBxJbYIzklcj7iuhagwmBog+F5WJiE/0mn80RbOybPq8lCf3+m+v6Hdc98qH9ydt
Cyvjl4eNs4m6dvutNh7HdscQF5h9jtVw1C9CO0HscJ6IMnYmosbLOipjnFiBIDyn
wrLYxOr0ZDekyfKDPlal6I55YCS6aaitQz2YJxymEHQ/RsqQf1PpEAorTMokLK9q
dq4RJHr1BRAyWVwm6E+33nfVKb3zKvdquw81ub+xChYYpOjPKy9RohcQU9ynYWBS
auPg+IHurpbkX4TWrrdJAghNybo3CT9MACXZdb//kyXCLHkAd2wBRwE3l8g3GP3L
lO32lDxXigHsjUEoJa+zkexU2WP/osvKypbR1N9wMwa/xfPiXVKeStpi3hfzXTFa
Eqchrtq58rkTG8ckop1HoQgmisOQRvVVyuxtEkAStkwrbvJwLH2Rq7ZoXfVO+h4c
Y+3vdx7C9SGITe3/EBz8AflZ+QG0F4EI4azaIMcSQfB3KtaAVT2wjzaLI275A4IB
1OX8q25M8ZAZ9ux3Ny6k4KRy5f7mXS+WnqCJj+bK+EmEiP8c0VyLgs3bqLwc0uM7
qHA64Bc9zNtx1xlwA1FnV3kiSQ2cBUunFZhLMKhXnzLuha5d9UMGaySJQ45O0BMP
NlRoNcrWg/icS60GKdPvC6BZn8Amhn/jy7gHlJr97PlY9xRqPcVyTztgUCpdl7oO
YuuuULky2fl3PyuqBOQEiFmSY9r6ylzGRnZPPZVL8IfO6+bOyjjbL5FSujHWvbmr
gCcGPFgMq1YTkB6/PWtrwUvq6KsHYFrkICc2AziQDk2bArSCSTEIeLP4UTcZNF8R
Fxl6MyyaRHPxqMi1G4F3LoC2a2rmjK0Fp3ZfzXEcLOALuBEL069ftGMZg6STwboL
yD2xbeDHcNjYXZ6J1BNj/o3ud0/tUT8ohAuYLUraRgJiEi9Lnl7gVgD2ceyBtWIb
IlHGQ/kweYMK6rkIy9LhRUZLGli6UoT1zKwTS0LsB2/8ueQUKXB1Q0NINiR1cxd/
MpB0zi/TLWQ23oisDCRD6SplRA6PadSXisvHeBPurTUfHwoFGMH0rJcP5qs/zgzH
uwGXQr9cAcuDZTFa/IojEKR035SC4+LOEYF+oLTtGogzWJTvnjocIlZvZb23Lz0c
ZYfTtMWmXbm/ODJ8gX+tuJb2WjPHtlo7Bd1XrkzkV3mlEN4l8qUNR27gqIMXmbt3
9rPr0efff7sCAUSfTanb5kW0bx/b5n+61N1xTw83MnbYsiL7Sv1c9f5CVr7WA3X1
2GXL0rux+rI/dub9RRgKDvdxHTVmqMSNw0tRke5w07m4Lh7n3MFZDE2VHGyz9xIS
5MmZLKWfV+f3qjdlM6xMpDHxBIV9ZzrlhmjuzqQaxZKB1OIbB14aom1wFIGBPgl6
1U1cwYb7zJR1prFaOwbxWoNC0RJBbd85vBkMOqa6SDD73lhO63yAOGEk2lENS/+H
38ccbkNuWy6bejbfVWh+dzZ+NrBA4xvoLLQ9lrqTVz+ynmHbMBaLG0H6u2iEzcm/
f4FEjyn+85iQ4GOSZhTeXbEh+bBwuj22PD53CoUWwHlKEhMkcP7ZnRJ3BAt/tX6A
QbnAgeiQlJXTs5v/aCsetDuf5PYcqxCGpXMg6PQ/q95vJB0rULmlHt3pfyhdFM2B
3FL6hM5euMDrCxM/Swr/4HW6ZCFDOyB+WelvTEtPbJ0VW77m1otM8FHaFX94InBo
RYSqUnVY0puVfvtXfPE7qxBv4fwypDROCJ/SROzY3eNf6IWNU3zPFXsl0plqw+WM
nGcLpK4IJLyLR9AyzatdDR1/yUvPFkVbAYps3gNFLDEvOTzy5uIhLqfKGIbeVu3W
5QUwYOHz2bE0SNSBJexBESEoe0OWWoJSF+4y2t9bEWVNNAuWZuYVhpT4k+hZ6pDp
E5pLNwz9sT+KiUCXZDzrDDvYCBznOLsV2cjdPCaVai/Qn9q/7psh5EB77gVcfugJ
E4kkfQGqcYYyKFbF2DfSqUNxacH5mTgj/YwqJFtzDZEDwk6NOz8T7sd1vexurfWp
YqVvYEapziADn284xolbzBap/KRldr8MzTuiVpMwXjESdZYG63Nkystj5311Ruh9
VFueBBncXBiu+qh57gIV7w0wu9jZBnoGdyKok/i+MSUO47NzUobSrOz1UpUY1ak7
B/ZRMiHuJWxpv+LbaOBASNaDyacmEUFZ3T8AcCLUKuA+wbomBX/yl1/u7diwvfFb
MGjHmYy+MAW+T2lwXpPkIOmgkfF342Mg/IMkxCH5r6zx3WqiebilG7ORHFtf7erR
y9LXvZ2LeqIF4JiRpXdFUbShAliUK/QDU8nfjeOnm7oe9Z7OGY0MQ9QtsEBC8G7Q
Loqm8f+vt5yBg3IWFYclzuhgmxlPKur3ZnZrDBGcurwnpFSqZinzshD0qQMBUXVC
qauOykChXIh6qa6bP2D95wMkG4+U9sI9pxQGFBcJAyO5iE4+azPX0Ivm5sw6HTeC
hxnIj48yU9/sWmAo+15u4K0saNfZXCZzYxEVPRNsh5mxT4wPrsKDV7e9C7djGUnF
QuApKgP8LHf8T7SAxfIuEljaPTwneHx5dveR6bMw5Vi2SfyTLIu2uH3WlpmYkKaO
uvhQaWvQkquVxAKxRnS4W98lxB64KLcXzNjeXl4Ph/6SdfVtkouP+BRv9d7ywOTm
qGZXygoVNw9vTgq9iSKAqCoqHkVNfsa1bgsZ4lmfUdm93h8rI3PDgpZ+XDEkf4ZF
rqIf6VcUbZwEvmuMhccmqfJ3w4GnVG0JyqoP+GWTJ33+Vugr9o+9wLhxtXFQG7jk
7Na/yjv1D7QjkBZxEcsVYxBthekgleiMkpBMFkvwgTKb7cMdJpLkjYYsl20Pd/fW
VcOzFnZV+1vgvJ9wEFBs8SC36YJ8nrRzatyREcZfweEC3j/GMiaCL2sS6YJYcye7
pokqTw29Se+RnUxt5yXTpuvqdeyF6sR53zc1fAN4+AhExJ9BBJhQ1VKsw5ikqv+O
b8MDfskndx5SocXlZiD0bj8IwLaQz35jD/A11FyJs/o1Er99Q9bx3TrMWX/mOge1
ruqSNW5eVEVKt/Y+NXnBS/0RSGBv85jUlhWy3USG2jNk7Hz3Sdca7tCZjfqBUq2h
HE0e+5gExEdVVWRPnZ9c8djLJrkt/0s/ahWiIeMSZyIQEUX7MxS7UclGMIT8OvoX
4REilJmhh/B/jvOJrG3RIcue2IPWDzTjfnLxmDfGTeh8pswaNOfNezd6aiAb0Voo
jqvvAskTS61H1RZ+8Oe7fDMoxmt3d8sp+aLmIhURydLI4xvtGaO7ahkwQP7VccFB
kHUhzr5/i4MBHG68GTj29WH4PUYR+2w54fEStgAQlkYHuSRZLBrAKgye+eLUldMW
peELaPb9SmGIi09TUa7rlKM3w0NdUjueCJRwtlxWmB2QLeonqefSrVzVzXhv55Ec
CrnwdXdqCR8YUBXOeZU0RtzTTdyEAK4jqOowEccTOwJ2yqRogtkM80OBALGdxxY9
X2oWfV5a00mhJYZRND28ciCQHu62reFiVdngPe3CsDRNMQxmKM27k+z7PoNZRypG
JD/JU8qpblkv6vnha1VR6Ku1EyQEMXh0qzdCdASHdyOB/N2Y6113ANn9iKUKYNHW
91FN/kGmpfWD4030V7vzq0GvkfLzAke+C9fAZE6D0opG18DYeCj8dQyGrVNzy+9B
+AtPBm6qTk2efRuCa9cbewXg1YplgexyZw1881FVljt/SGakYLmfoKDYpJlY5fHZ
Tyo1K4ibvg2sYXQFReksBnUT+jO1h02baM7jL7ix3GAZEAY8tkuzyc7HM2QEm8mv
zwV9Syq/l/7by8pX3xnhVTM/6KnUvIOPZ2XbsO9fk48Jrjb64v+plFhkEu0S6h9V
oT7JNvVDPhGen4QHiQQbRCgvxCghXICaoAQYcVV/wkNiKzIdQ/h98JT41ZWFlOpY
ry788QJdDxMXsfZ0ICbAQSY8qMShvlnEq6OSvLhPCfYe2onKA9e8t4tXCeLOUYZ9
FvjCtJYzauT7aP5NCzrtQFv0k4TPQBjwfjnKKn4AqCtaTBJg+H0ElGuecSj5N679
gUglZtqR/pP28gqXZ4wN+59g18NgibskYShr4jaGasP7pD4ag3BA1Hb3ThiRJHN1
vKEvdfDULNwGz4Di8G+ED13kqdUj895NxRvzz5mm+uqgnqmEMsAGlMlVzg/F9RGn
oE8bzJak7b6HI+WgRfJuRLkoSK16knavBWHjYqJsa5rFxlrfaAWwUdSOzVuctcxI
j/f4gLY3z8WJmFOsdsLG55++UevJHnhJ1U4ILzcHoRmmYnQ2XnXRuMoqyRCujlFr
zjSIEC6k7gcBiEFOeKQ6nV/UI0SeW41z13L3wWvLP+U5ClsCdFVJZrw1EaHio/jO
/ERTVQeKNFpwUkTviFdhYnlSX9xmXsrlwNCGPetnKtSV2eGdQZefMoME3pjiA0LJ
CvO2wpxymu8QiFu7k6eiwsLoLILKyOmxherkzDScSGh5mQy7PZ2Ha+fsvEV6DaGD
fmC/Ke4LN/V4s7CUitSPNKczremgU2N7DqY2o7jRbLFWntTnc1SDnvsWV46m1Ldb
no0jv8C4zMQ1YjvPSJASsf0vByMKBLzAoa7+QD9WWja1ieI2PDDa9XQWfHyiLUj/
rotuIzPgR0HwTteUhSzOkD5osOhtmuGWn9zOSwHLp6BZaZ/TiWKOJm4vbOIhI2G8
25RSwRA+LWRKygG3KfdkJuKzjXLpUARD7bGs+m3boIpfovr7Js09Od9SBiOpb36l
OVZQfRoQEQfjZRm0hH3RWURAHQkaYc2u7zVyAK6i7gQHxpVOR6JqK9k6XUZk13Ot
CIBQkPoCjSpGsn11OBgIR1yN89Et3QOkE7qSucLNDz9touRwMatoblvym3qU2+nc
LqtFEIurx1foB6WrrQ/k1zEcUzmt06YRrLRPJFSysBLLquMGkg852oQyV4pZHTk7
jOProsESMA+e13DKcFJWglEoEsbYfvMbrf/k6kekRitqtxxLm8xJPJmcksaGBj5W
e7kf4OjaN0e9elA6rJGX6k0wPsRguP7Z8EzmcFY04U8yRk2NGPlWZq7pGz5UvXc/
WQRdvETxyB96XY43aLN54oqdLRu/bRTFS4IOLQyW2ErBj/HgU4Gkf9tp/itRCKZN
rojLSGemKEBzuNN6lTwcZ4RbQN3yB64J93QVrxzHiGT+6FV8ij5l2ALBmbf2afFh
3rcKycu2ZypyN3aIYq9Qxr8Q3OwoWhh/63Y76FsZkEttFwYvC05m1vTk6khcUvyH
UnEBv2S5GshCemq5apsS72Yh3jID3xX6VwXQk9/5nZtTV88lTzvSPipPO7w+cdwT
h+CCLDzvkQmWDjbZxXZarM+VgQ38NatZvfcVzPFixzY6a6+/jO4typHR60Ec0t7c
mFeRCRb6eXSHuAX+N9tJpIZ4adVZ6fbUrVndSkaa9uvcYlGbAPLK20wG/pGN7rL5
+9b9gQvw11xeJVuXam/wVYjIOoV8FGfWpqLe6Xz8Nsr9Q6JSF8cDhB7Ky2N9CUl+
lOVqTl/uh4f9T1Hc9koCwjOWipdl+YYczgsTulmHiMdpeKI6oFkkiToS5Cy2afEh
E8mSahSq597abjriaDZb3zOqN46f150150moXkQBm6glHGVY+T7uz0kbwtrunhUP
Ibt/QKg6oMpTdl5C1ll31wo/asvmIY5lxhm5HR4IIb1D8voPN7blNnd/E1f/y0zd
H2b7KtrDVRprSg/z0gZupsTnSYRxgRfK5G1f8MgtRWXHfdrpqbPv/WN4mfms33uk
72LcqY34NSIk/5+0pyf3R2/CnPDDuHJxkSccvvwgo0c+193ObSiROaHZSEeRCbXn
MnSEEHjSLNgmswLcxLU5EHh/D6gS6vSVShXOcJiri+QCdBWbDBa3Ghqda/TkXa+D
6N4wsN6YEK8NoUYI0bDK7N+5A5hWQhETpnUSov9KbcxDvg1jmD7a3X/yMk9vdT/3
Wc9FV0lyM6+RkvXn/nVuaOVvDjKwl81bbIex32D+TtbzXJG33XiWIWY2XfUAT+7o
TUX3O1g30GuNe97q0KqzAWf2533x8ICIyjTkxOVzgfQAXwU5WLmjvEbkuv+fIfOz
Cqlg+BLdczZYUddVvmpcGTS1hRKfYqcT8vqpsS+G5x50+Dbq/uzEBANlsayMpA+A
iJd+iUn/Xhneo3zshlarlf0hVEpiIRlIwK4xsC7ozlEbDEEg1lzNiUAl06fwwo78
cJfdseRUmSIq8oUTSYytGjO34T89tAdqbQHw4sFbu3aryaWqjUZtao0SBJSM7tGk
fs3VOO2lt/HYPhjBIQwyC5yHzCRBSy+BtQRyd/71l5ts2ZAoa89ZUGhDnmZWNwjp
Xo6ioF9iJuRbKN4uiVUCu26+4bBEo2bGcWCIIWDneR8I9aeiyViFJp2FiL2BhWGE
95NrZPoAHLmmtDBmkJDl3Qe5lEsaMPWeMrc8/vpUbhCsZrL7nu4Oavw9ffgTz0KU
TP91o979BFw3IigTXiw65731lJUVY7t7hXwBDdbB69xojlj9PU1W2xBl+W6UV37B
GfET4jx6CJSkK3H76ECiTWIBJI/TqnFvk+4z52QPay/iT7NOSYTTGS7XIXkIpB1A
qKvbIhU336Z1Mis1quL0cW28DXICXAbyVmBtB+Ina/XxZlyRzxHtst9Kazt3oesR
TfuWaBz9s06IBdZQ4F6Ugd5xhtQBIa04b1ohVMWym6xcNVB4NpkZgNfKHAOAResM
GLDztRTBeqPUl5oeHquP7fxSnrwkr9OdAhozOrcN5lO1t+Kwruat6P/sgjgvidUq
vRGUH1wb0ZdD8akqFkTYNnZZhAmkAUSXzx+lhK1kYqvSmEn//oi0Xjv8X9UjdIHf
4pGXqDAJ3BUQKcDAp3UwOYJDYGIKxd9f+3d6q/49RHrQqqfu8aiYwybRxCmdRScx
y0n0XNv2iMTMpMj0TaSwigLDaMSItQ60ZIwWhhctYU2ty0vZU75lCQl/rOIBKyH7
VKWen+02+Bpj96Pr90UXsu73909O3c78OPKXYpL08v6auWJpqfWkP8UNZFfCxVEZ
AUUwo6myq4lJm3Q43F76fNCG5C377CztKtjosFfVQRw26pr8VRFRJgPvaT2iT8iE
C7ryy4ll7FoI4ngIvp3nCin8mlMcf1TGxGg2lTFt7JvbObbdgA55R2u9P2/8h3FT
Ykg7A+IOohtqztK1joPvbP23F4S+6xDhecYRYgbuE6BNpxKcxNwSWArB624nVBB/
cxVkFavDO5Bq1vELBZ0Ogr2KEPAJnqdxyIlOUkiEbYbIF7iuDgFmqXugSCkHKBzT
FF/ZpKRyzDdwIFASybonFUOH09G0vR7qY7QK+9Ra2mplJeMP3KTO35zPV0Jr8xN6
BP93X7N4aSBRqpfdc8qDxqusQekzBn0ecU/TAPDVUX8fAI9U/U7HelQ3VEGCkLE8
mMXUP5M8yMnEYnl7EQSvqEgVLGCcZphhQajO5hIJWQdY/7XcJLQdS6upq/oWGgSM
luWtB2SUtbnlGb42wWdZswRrhHgS5bviBYov9gqKi1ybrXhu/vnQUCBCvIAtxBgJ
NBi5xb7yhi7PHAC+hofpdd9nkYjWBbhvjzp/BjOnevyIngYZyoppZguQ9iZTd7dL
dUUiE40KUsnZnvp3Y1U2cFGzeEZLqHO7nTLurFGqL8uqThOslHjF+CfH288gVj5N
cyyRU4bfAChbKWY5er6MoSiq0157mH+62rurI3zPE+vfx+82KFhDil7zvAqkFWVP
7GgjJR3g5bZuF59zPVB4x8aFDSyxBffroFaQr5N1GxizK91BK8Y9KS0VC7w6vU5N
hrFiIxIbUb6yOGC1HLiU/uSf6uDEBzrkzgNcSGE+QcB2wQT+gL2fUgCnU6mgAXsi
QJ/TU5uZQz4ZLOrL2yABqs6+NC4VUKaKwK9zhwIBipGjE/2LLHb4ag8c0wfA8fDy
D9PnR4fBcVSEOlAKLwjE4H9P7Mmbfo98O4VJbiH8np1+IXnbWL7T99V5mf5vfmtG
QrGsq+2K4DFhzTpnp07HCc4LumfbTe3bOYjxvG/gmKC/MvI84rRKIyDnCC1s7RmL
tBjtAtDjcv6i3lwbr9PaUXDFz8Cdea5n+r47mZp0EJbo591gyZG51M1Q042Wf0wy
X1oY66g1usO5rHbSvktN/oicYx+Vj1rin3G1T8FqgmiR9bnxc2OHmB6Zuv1GcNB1
92pZVCdWuWvKrSZEsq1X0bbtmqOSsiPbNPW7QpxY2WjoERPgUT+TaSMizOMtL/oi
bX23VpoQAqi/B0l3ZSDLRYH6RLTp6j2IYdoBVdkIT35yBZ2aWsd37d7fSmkCE+s7
BPKjWyR8Z4F39rqWKoelhxtWSUV+XnPXSORNd7hCg4z5+M+xBy+0E/1/uNRU2WU5
NxPCqsBtnS+1YH00Dm6Um92JgubmM4hRDmKnqqPvhjvhv9RjJG15N0y/mkm/YX2+
hID0w06bZkdWKTQzrsJUrTCYWBxEXnRNOH2nD4QHP/geU2m+JD/R/VmhRZ/K+X85
c9eY/tebS6GjEZ4BifNtS+ZnfNOBAPzBxfSwoYIt1KOI2pzE4doupKbaBdBN5L5F
3x4JcSM+5FpBIBrCz2YkE+K2pBKI9Z0ghSFeNHnMSnGEJ4b9mHffzDTmrEpKq7BJ
+qBEnmJSXn1pyh+xPSrUwJhwYiXIS6gqiBNez3fDKG0EgBtXgA/m4dB2jDSOhZ9N
LUQHkP+Keg5gDN8MYpB1ww0fz5NI7VwuecdS3yuPX1LaVnPzGin7uJcj7PBd8moP
e/owXeFQA4W7xsQE9hmxNvMalCgqYgr8RPfZcGu+1Tb0765shzc28sCgvy11bmrQ
pURJBMXyc+x1AkUG9m7EqvfW+8ObPyEOQ47sSDF6H/uVNKVM2hl7RlpnOl3tNE50
rDf7xWKItqkGXgq8n9LoXAWMWHpwTAkFVEDT+pPMderNywlQpKmaUexx3MCejRTE
PMB/HLB7igzk9MraA2A7iBy3g/ZUvPN8Vs3TcS1pFIIAvVxiRsv12cEoFlLfNgst
8q1nbnJcp2thxYi1GEv3ZwnwgewFEQxjGas4E7cztqM74NcRjZm/H1sBNqDBTqpC
pPtx/PAB9qkFLJsvAVeg7p7kulruu+xZOZHsu0AkON4uila4qbGY/ycT1FxI7uv4
BBP7G5zRH9202Hl65ZdoXe4wmyhTcPXY6ej7+la1y1Ke/V4t2V8W4LmktJPpU2Yf
LdO2mRef9K2n4pD/ScRFP1/MXWLr85uD8Hf8f/i38OOVrfBwOASDgg3sXSZDHNTQ
raTw8zCgwP53zgu3GUmGZWsymm4GWKkFdJ2gsd8qkoEfFWBnbtRkRJ+aA2vRcuar
egBhJ4zrsVwVdcrx7AZyGjgnZO/FEjAi18xe+f3Wi5T+mAq6Ty0AhhNGe6PqIk8f
VG9DKu6rpfJKfgufpPyQRmVyeEo2kPnYMpe+aTg6/cfy9RMZu2RAMGke6pC1+uHp
o0sw+LV3U233ZaqVqkLAdUMnwIQJpKDDc6DvxfJQFgo4/o70TMSknpdZExa3lvrp
qb96s2v6p5p3YpcKJUWcKbNjb3ALUX3+6FNDw3FWkNRQnuDS/bMtW3ooERuL/rDz
J+ixlrStubCdP96wS/b5e7KiqvQBiGyR5lxrFP9BqM+0JuVUQRfwyw2Gl8Iw8pBf
doh0ENyrsKNHy3WdRq8+LGgOvDAa03K+MMKxZEVodzAPSwPvHS164RNstcJbHz1y
5aGxLtAHH9VQREc6TRFtePCuaGd8+B9So0GQthwmt5MCZjPqOJ2D+l7n/t4RhTB3
Zuj4mna/rGCrCVsNs4sEUniLVgw/G4s84hg25rQgGSAwDWDMtovk2KR21FTimmbA
6XvvPIj/XjL9TjUCDAEglY+94xfRxU4+23Fx0z0ruTpBd/u5Oe5iKftG0KM3p6Hk
UrvM1I/Hk3djdAsfzM24Q6hUqC8KowtRMHOioFyD3TqxXAcp1oA7M2Y5ittOKdvS
dMpu3QZ2LHfIJI8Or77MpZPntyeSZ/7hbyMN2QfaQE6AXPpVoxR3Mrgypt7LhLkf
CqZ3bal2l0ipVPJq59pUcVEjgC+eVxCDatwqwYh5joCGyqsbiaxPlNVV+gv1VlyX
fU9496IKY/+5JAQBkcf8q3s+GzAOTw658zCmXCUg7tqS3dUpJXBs9R+iNCogWn8C
WCMzgPfUvlCgquuPxyA+aKPGDHHcEQBlgdwK031VWy3AgbYzVsRUnV/Q/SFU5g1A
fD4m7iijOkjW0pwAXRzMLrlr2WyrWh3hPL9hyHevv9Em9Rhp61WPjNhK12D45PU/
rHkbwE77H2XsNSdadTA9mUgvMx3bRjCIz2VMU+35xgWUeni0zH5anJvqcPaVsHgy
IGh9ACC591rdf5+BSH6SKvbwzatfLEWDz8Xe9Ql4nh0pa1DEHgmP0/aHrwQyNWtL
r8Kvmqdf7ibtsfIyXPof1c/iINIrMMlrpnn4/zWSPu1Q3qGRjdJ5UN2O4A08vHVu
xHDJe9XdBIHk5sTX6ZmSIos/cSgUFeLwY5WfpqSWxpRFNHdxO6pD2o6JySzPsATN
ItSPzKPQlZFlZnj1NX+3g8LroSwAqa5UDoNkq3dbE8zBh/7MAuS0d31U8ZS1TtXC
9F0z4DLr4zdpCfJ/mCf8IpIORnum/6zt1+v9Jh4+lDyHzzpy7Lz+s3Ow8pDNMQvB
ErxBZ2A3/LbbfuuEo2uBxKRUTuy+rj8rb1z+iR/FkCHPfa4liSO6n+qqhL3ui6XE
ZPzR5rz/ye2ATh9xKUlJTNkF+0vvmpDn6h5mzK2HZcMJtmojl7KTGNWla2eS2N4C
LoiRfUmCr77Cv/HlUHS0Hx5wfP6zGQj5t02n0cpSCbQ+05sWsTVadARho8OKwKxs
1JDOX9tKpNVrhjDGjBayNImqu86yiysx0iRIsskK/3G9s/Sdj5O++LkXrl+QYLZX
GXMdxJ7Fy6qdhXOhHLNYf3AaJ+n/VETjp33gsWjCgpl/TV71VHgulS+d403voro8
0WpGMdbjS6waM/Si6unzAfhZQbGlR2MzvGqWZga801JQwt+LT2Ar1l7FX50HRxGR
cwybC4klpYLVTa4lXFMdTgvE318DlqCseqcj7S/YmXQy8NcC3y+hEODBbju/rXUO
M7slrilC9vhCxNl6Q7ldqft1GBHSbXKArkZLPY+nApNUlnUWXzQJ707uVv5KDLC+
9g6PegEHSJ3ayp+tEO+aOdbu+7SIG0yDqx+/jfmiZWp9NYxIOCnY5kX8NjJuw54A
6cRr75SrjmTDB8TB1yAYaf1fXIIiWKsOrfjedCpmvXPiJtfE1HCw4b66HHODNby2
N0DvI3QrsG0xYs5G6n0rHDbzl/aSwOg5r1HRWX0NXpk0OTffJnzOlEjQ48AoJrQb
xauqVVnvj7GjEA2wjkrHBAjr3OsP8gpYUuc2JBASxOFGBS8xqZ/hJgbVy1TLdtt8
s5ZyYr6tZWa1rtcwXRY23YffkZEzxRMSAWE8ptfAxhbrFzzvxTJFyz7vzWffOcI+
WDkucdNBcea3FyIFwUx+sGaIosBAqKDIWxdKxhFkGwnzh5gIUMpY/7E8Z4Zq+N9l
ejzT/L1SKbvqSzAtNB6pJYrvWPcAo7FOJGks873k0KvWhSCQ3GVMA2M9BqFbIsO1
XvSnbq/zj1nDUHhKCIjZJ8LtAOhPxAhbFJ29CeQYZX97DfOawEmf80tLkRu2Xo3i
alRs8O6w7rrqVyBXgyGUaSnwIx9FsoPXMFv78P5XEaZzrcLGPNZcprgOu92tDLXv
89PPQ0RNXhhk/ytqCQ0GDOY0p8MJQt/37B0JO+NivoXFyUFv+dFdNHn7H2xpHMR+
kgfeFyN8Cw5JlweeTShnRUUT922qyA1HrCUBi6XGEU5qTUYl2enK7o4tgOGJ50Cp
whz1jgoVn7Mfk9G2Si1/HmWHHsDdqJGvLUPjjTZBKVET0vBsveaSZAeHMOv08sg0
je84wjEUX+IsrhpD9N710501POS0FSthYNas0tsIvI1BKoDZPI+n+69cwvYyV0ye
dGUEnBdwO4r0+WN2MG169bVWFPykf5d50BIwgJmSlpZz50axRrfZROW0qxsfz4Uo
vmyBhir4kjk4ps7j/IQuqHpVdC3FyBwXcgDv319xjv7Euiz3KSdgQ/HNe7E2tkFU
DHO8Mtc1OIcMpWMPRAsQZfqNEWwmdtlZDkQ76Y5SRe7m5sxAZDN9A56nzT9heW8m
zhcxLtUJtpIasZBkz2CB3xx2Uhp4YNFWz5fgJEMrtoiDLLsIUneFQLNkjAZKX+H5
JWCKjkz6wKu3jKyRLtPCFezR1o+EH88M0sD73X+up1+3/715Op6ciL0NfA8qUBCV
NgCG5bgzRQR8++WuZoWwmpqRrTROjoVyW8hu8pAKFCAsIMZQmv8n2liCIoJyDxMi
20z6zDumxjaKDa5fRbSJ48urFICER416XB/E3qLr5mhT3Tvhc13/dsGcTt72ph/n
YTQDZQmL7dGdXCBKPT3XoVa9L8yeTpGLGZqRzNECKau9tQiuypvDLWhD+Kaz0tRW
yMT+/qeO0joKQWjUKT3D8cUHe4ISwmzhmKpBCMAYhnXu9G9lpbSZiSA4wRkTuXjU
rJw9f3EYJkPSDFtf1prj6BmyDgDzV7viKV4Grl7+sqfL1FG4chXgmzmqp6K9Rlxy
qqc6ynoZKLV+5PeW4Y/ljSWQQla4TZhM07A+R6L0axTr2s6u7sMS1Xn8IXdDgvGL
7f2tTdbTYCatjf7hFtOuwjf+NsGzKoAB42MJXrvIwUiVSG9qnJLRNkiMriQH1TG9
DMQPD8tfpYb8gyo7Vd47wQCk0x/gAp36SE5yPI9GMIe4lu0G7tGcdYtVcZqyXMK6
xpiPvhBohmT184KVHUHwtVtHrvoLH06y5NsvctBLHXWvJwu1CqHLL0HhIlU60x7M
QDAWF5M27k7JmGC/8qkfLuoyyV6fj2x6QUJqg9Gdrc3k7fdRwF113P7oJ8qB9zkb
VB2aIQKISIcngE/mRffNHPsU4pIt+CXVWCehmVRFv6yO6XunJ3qzm+XhSf7HyqZ7
OddIm9ixgnBsyhRybZX7Hv+p31tIjakyQ6VREKZ73bQm7y7ydpXIl0xg0fnr+AQH
zhVuRvN3+0nvATEeXrSOY03iafWz4xOEdwb6Yi/U5kxEy+vcGEY7iApbMY4+EYy5
c4LMLrszaMvCo0UEranMGRRUXcBZZuFXfuipx6FP0MloP7B8PEH+h4rU9Tt92Pcg
bnXSdt52bF+27b9pJuJ7mh2w0DyZfcnUBFQJhpW63zL/nH2r8M2Ap5wjopNYLZ24
lyoJ4JaTfiQJmRocFJhLg5RoY5Kw8Q+e/i7NfO7kK3FGNeucK4Bxje4EB3L/Hf7N
RtxVGCZSuEIn0U9dXKNGxQ7v7bnXXiubUv70vPsm68nvN4dneHEk0zkJeq4SB46+
blJCqEAcUVhWja7Yjz9WwYx9U2gqCKS/hspkIEd6RX05KSS/835L4sdVlyBe2CrR
2rxij1Tf3UvHgUAFf3Hf+DTJ7ZQlYlJA6U8azFZgBIELX7mQoCzjj+FE4xuLjkxP
5yoUwvWzn3ArHHguJNjCcZ2YyZ0NRs+G/yKXS6tY0v69uXax3iFN5lLLXrsKFwIq
k+fX3VN7V2Mj8yMvj4VUnPH2xt2mUmCDjZxAz83qmGS1xIv7rPL10SiGrpSi5o7s
wM+MCI9z0QmgiIMT9/q48tQ5/WZhvpBFzOrtbm8kMQPLDU7AahOZtZXgp2csUwVv
Dh7cnh4+4dskjWVCRz8a3CNBShZHY7x9X4XoSEblCY0P+J+Vqql5Ji6Ieoqmb2CZ
BmTejl0N4lt/9eXclVPWkHxilsKI6WVyl0pIlXHmmh7IUYegKso459mKSrpDGvwh
n074tnGSepi9A++9/pRxZz5fX2TEV6fgHsu80xfVX9i+rM1b0M/ZS+gxEhudH+1u
9RYMidPxr93xp46CszSALBDJr6z2p2JUekRJ+KYr7/3oJ5eHGKf/bvrbMssROAUu
xMTeDztgkHosD/VcoMDb+2bj6FdHp1pHcRF2u2JLmO+sX3DbpkNSDznUmqSuQY1P
/2KPKLp2w7efpn6he+yORjbmkYvKjKi3BdG8zDoWvXRyHpJ2gGq5WYcxd1rbeKwN
nqSPpizw15/lzdZKflOUqe2sPlxiIK85p/TwymAB0gL+cqP26w0AAFdl6V/tjdPa
YrgMw6vs70jt3rWBkIGGjkxSQWI0oOUeipXWm3iRCU9b9SBUVWxaEGif3Rklf8wF
Rlkrp5LO0ftaZ4qOtSaFNcnXSeZi56c8eQNHTSsCyGiQ1TU9iWqijjaBAATuD8m4
csQryxc8At+sksTItKZDySLeW0/E2rRP5xbUjAf4+zTzzOStqk5bcd/a9sBeB9On
bOKdtMCnIj5NfVJ//qv5UaoYxyA6Qcgq5kbGd/iBf5VZ9F1d912wcgj6tKXurGk8
KcW+1nEAe4a4jt7Qos6GYzZuySOPE/IdSR+KtgX3sKPas2dbMLXLOSEzCrduWV9s
USLkyfZnEFUm/WgokKQJmEjMYKUhw2j8tzpXbHwGkFNFD/5I7UKziETyRDwgzNPh
HgXuQk+0i2/I/mARSGg0oMRnfXOA8ANlVbb/0CUTfPp5uMUrMTXnreU88LlmJ9U2
YQxmQpYZTwLIBbDZtJBdrH071Esferr7UQ1gksQTcJ9pVCu8NhIMC+ya8qmqeY8b
E9rDat9vU8fL8o1sQBHOgtJgLW0O2kYrm2O8OzmMgHTfdd+3hXk2LpSKqOYeebmV
LJ0blxaz2DIrS3dM4XRURTahVJjIcqSo/3HF6cITnsgfC6G1B8Mkix+/k+CxdRoG
YWHCtHLua66rqslERWw0hba+mAiH06UshrVy4mN3zNoDmm9kjJ9RnfUaGrsjKRBs
t7w1okvP6GkqzRcO2CNfnIz7Uzm9JW+ijBZj+4c41DiCjbdXvOtiRPCSLDyIQSTX
1aiwnhyPaaTi5H2h8oduDDl0Np2IBWnMfNrqYDe2On0qVF7HFwo1QsAOhOW26Bca
BGDx3K2N6cJf54gXJvdig2lT5+9lFQ+XHTWMS0VUCZLeW5yUPa7O8XCK/8wABjHa
b2SMrtx+5s9rj3actjcbu/y/QbjNpPig18T6V55g5maAcrRcKYxVa/9K0CkwrWK6
gGZ3tNu68RDhUdcvB20sDR90LirYo4lI2EjtWPrmy8QOguwFu/6bxuk3zPnkEYNp
FbjRnn5b2LZgMUiNxroMXCK4flaLZTnvVr5a+L+Q6/kyJOBATldzrFc1B0e1I8rG
IL2ortkxUeEQcYgUds6vdc8+EXH/FkfOxCLdl/1tsaHe1o4N7guhAoIqK3ST5pJp
JOpqltX5B0rrxJdts+fv0kocgwkUc3TUB7S0z+YFuSka17ql+4fVgOZef0JnHt1M
DwM3g6KdHEBrJwErMKV+ApQHpbE/FTQHh56rf7pi9YaJ0yOy+/vjX7ertv4Sty/S
MX/Mdq+t1lRdsgp8cIAEBabAJdHomS/2nzEar9GKU5AB6A4194lYbhM2c8DsWNhD
uUqdXg4+66/UOo/QyNmNDAvKPYd8pwdpS5lBCKQWPMufzsqF3pw3wX27Hez613DU
+dksaK50WiJ3L5pi37uLzImdR6GXglij2tzNrQRpR4KpuH0lsZsuNlCzHBI8ncf+
63/M10bSLzyOrcFS5WA+JUxA0FSxNsuS536SIezAcH2uQ4i2H/diHLsEI8bnHzX3
8FdVHWNh8s6yuxFVarnIaUxL/EpCbKUsA6xBIbohiW0fN6Tp6zbwcEKSFETXoYZn
pz5ZG2+AbHpjKPdmPdOBTl301TvlcjUuhCLzyTTtm/oyvlvfWsL6Rx/BKruWUZst
O9N/u56I6FL9MHxX8N5N62/09/QN6Oox5ALyfHwToistbG3APV2iZjmhtEaFdjer
PZZI/1hXmgBLdD28ROGfBdE3u+y+bCO+EYB+FXwVUA6RGdWz9RLNLEkLiUx8a76N
WeYVw9sx0z4f5LuA/ZmqCc9pV8w33xRqAWlan3/XYxuJUGvE12vcYh1QjfM1Q4kv
YhFSvN9eyijq7HoztayWnEI2/wXUg8/bXKfdZXAId/HeDusKbEb6qR4I+EPgcFNV
wTiRMVj60QDvx9paCtWtFXfUVCTbfrPsDfMXwcFo5g8IvNcEgKIpfB77bQX4zMl7
0x4cdiT5zfBzvjlrrR+vlO720A88Fp/+k63QXQBk/e6BkZIAKAx/VuUoq9dZvdpc
8sFTLjtjfH57nIzIVu2gABWJpphETveuA7N+kJpysl4baPWppI59s/jtg26pPzz8
yKvot0k+/biD7yKWVcELd5fwHydbMW/383Uszu5502cHO5UnWhHsXsfTNvhyn95C
rzNwAk7wHidiYZhCiQ7SP0H8mYnGVTOj/fYX2XzhOa8bniWvJ6xJ3IRMhPNiF4Ws
028RwSceQxNW5gGv9v76RVudI276yZF5LMN83AmpfNv0K6UJwODGdA2zFKRBuGP7
LBnru5bFquaHkfZYIdjInGR2NTf3ns61gXuk1DIlTzZ3+J4gECOVmhjfAaXz27dv
NG0hZ3Yyr+BoxwdHdYemXsGEG/2hwN8xdDofM4yS+OflOs5S1AVqPcb9eOS4RpM+
vtPpGKsUz4hEHtsDrr4y7udk1oULTAKZUOLISvRhKYNCfSY5fBhLQGx6/x3eTgpP
jv+4kQOPgTOAnFrI5EQvp3+Xd2C31pNJz0G2LYplKl/YVsAZ6eFLtiNDdXOtmV+7
h/Aat48z0gsg3vxkA03pNfLsfR6LR5LXE7XWKaRouhJJqOv6tAFpHzbIppRe79xz
yUR20TksxclezXgEb9yQGed1hhX+NXGUTbLEHd7YrY8KYUKzozeeL7tFHZj8Xt7Y
1IHM70FH3XA5t3LrU9DN5GIaLvb0OHMFlmENBB2zZZAIIN9/lz0gPFxDT/NWdhnZ
YuinTu9B8tW8FqSkaoAUwtR/U8MOm/kVekrhCkuN6hRN5STI/HtkVeUnNkPRVXTK
LhxwPqLplBhA2hiB3uh6z5uU2tE3lJUq6DZW4WjB3baFBFPF9oC/5uRvESA4ycT0
qCcJCCAdsEXQxyWdIuGnf2734cmfQkGDbDoP5Pw/7bRJ41fkMy2F1OKPWQR3N3iW
YVG0An/G9JL/qOLi/uRS9+JWSSxIWx+7yNO8sRP7i0+bi9dlzzaG++0EhQWQQgEq
3Cwk4saTgA8awRJruoafjPW+UgfvYS7NUpFODCArdEzn7ZwIyzTaqp6XIQpmRQp0
9y048/gnm+MmT6X07zYfN142+EyGQ8igkotiJeNa5EnBvsPura0BA4tUucXCLIBl
li187rf20Xhon2aLrOETxHWkcxFE/7uldowNY0NcV3gRainalsOHEhg2xcwy6Dry
rRVyKjuqdBSlUBcbiORSHr7pNxSG5oD9KbkhQzVgVK3EESC3CC826DY8ZgSXMVDe
92pP9dSPznIGpggDKQMQiN8NR1UHTUEg+GifDtdCltCjD4GOdCcs3d+n43PiSvR9
9WRJs8ehx4FOCeAIkIWyCRLXm6S4sN2nmNp/zVco96kwwyDgwRJGQCvT2QkIgxHe
H14sJRoHRTv3GJmAaffpgDO0/0FG2xrwxw15xkMqNNefh4CT7ZMHBBacRYquZRtN
hU+9MU5d5r+qCMfyoicrMSBzBvaiHrzDFaLB5+LqZ8ZhszmG/faGPHsfGVuoYztw
hDk6sOS9/RErJ5TFt8CH6a0KIHEZ5qKYAggnzxIjaDuUkBdrvAjgSuyTP1Jde6XF
PineBdwMH/+WUqYTYxftYPNBzOOzssnVGWwSqQOX9gUebQsVq9K6IEpeXf5TPFqj
RunYuBNXxiglkh9B9V81f3Jc9FKv/AHgc1ZAufB0M8c10oYcVW8yUBJX9UKJflaN
zH4IiHuuDnjdjfm/l1YLSn9W3YKOh1yPSLaqu1azJjrDScsl8CnNiqsKk7zvlt2p
06d2wOf+cOLw0L93lYvQpIOUVpQxVBkxuvYPZU2IWiJUKt++PlsnE4hXfijPEF3U
QbDlfAyiCKJH4Z0ILyDFOh1qNiHzHVg19VfOlT9/R3pFDff7LP7cXxd1kCELdztC
p9Gz8cb1iH+Y5vYtjKE7bCS5UwhXeYVZHAdM3CaXF4fVolmEzQmeI4yFbi06e1xT
ug2Fpre67shH7DqScL4xFgcVKx7nzUgIf5GkPs00hMue7jI+V98EgLCqoL7GWub0
jhR4UiT79JAAGzh+iM3z6rXXoE7g+v76eCpxGar05dvG5vhlO1Qmn6ZElCWRz+a3
VxrtqXDJqMCgGtwmh+XpWEnm1x/qmYzVgpqsSkWoMh7tt0Q255v17/yZS4VfJfsY
THMUM8xArjVXr0miAYLIcY4/WvQ7I7Kyxeh4jf59KjsJOBfjGrN/cyP/uKoDpod6
6dm69gSiayBRZZIXJAN8R4n5peQvF7kGZcVEe+hRPM5A5xcZNhQx1BhkmRDiH6eg
YaA9fWv7M87UGTQbn0gHdU5nICkDziLgDs4TjXaMkWP/g+nGJDkiGuC1Y2HX7rQc
jQXLVHA7S83ME49sKs9cJUz5fT4A+g7n4LGJGvV3kzk0qepPpYgr/WP2WXq+5Dvt
dk1XYWAQ6xanSCh5tNouCBF6yJxu/GNUuuQ9eP3IIsAINTKtSaoYdR/+Gsn94+qM
QFc+MPqidMFXaKTMpi2k9fhRRw0dDx5rdopTxJAkIpG4+ZOH2wCYRt9xaDq95ZfT
vYwolOmwV0HMMXTxGbwzyNLxDRX0Hs+RSbN7BtyE6vEiYtGtoJ4F5gJ0DpctLxFk
iVv2M6o924d+x9DDC/GI80vq+1L8w0BxThzXcmz99sioho4Dx+3PrnS368+U6ChW
hSzSblINEfLRK/lVeK34t42lU2QRp6JDqFPdMa84TCnIATR8Tei3T0UMoazadU07
l3lq5b7+AZEmSUMIVPp3+ZHIHhH3sPG4Yp3Fv8Rn2FS05inYFGjo8I0qQy+VOwK1
MRIsOibp+dDjHxYAWTPKgdy2GmBfAfdahTm+H0di/pUnLVpzVUGs6+6kACSVf7py
3htwfP9q9zXok5DNjFNCZzxmrvsLFUKeIU2EzQhvEf9yK3ljAwRQfNG0fBa/MvSJ
4nrnv6CzET6E+IKuW410J5OYBjhmGwQ/8GGCGtrfJNQ6DBeFlp0+LwR1H+RVZJ/o
ZYnkKWd9bvP1lS7MBeKv6biw2yyOqEZnsHF5Xjv2rdXHRQQ7UQS14kEjlOmcFYl8
kcPbqtyJZuylk5sI1ZAzr4RLIOdyVF7IaMzUa5irIx4SOlDxeiaKvHLl90r8qA4H
qLaO4JI3zwfzJ+bxOpAEA8+za6idH4qN/hwCs2n27/Fp3i15Eczo3X1QM3ZlSoxx
bhTJvK26to6T5cBAOlu2zmZX9y7yD4dNNCNZFvXPNiYZQs+JtJtoQ4FRKojRW7Lp
gE3EWcIh+ZsBcysMbC1BRhJABChk1PL8ex+CzVDq0J3fwEu+Qh6L5Zl8tg5/eTVg
lcxGw8xrHcKiP8ect9ulZFyr1cvJVKGlLxmz3rFhA9YMhtP12PPmDMVytUryji03
sOwx5djU7jLuKIdxeK06F//FaJrzvXnB0JUw4IKMaPnO7PuPQjOCxWsspNKUyGbI
PAryJ60ZF/aHqd2kbtRSwmWGJxRwcVnD0K4uVa0e5B4ZhY4wTnlVUhV88c9sF/ZI
bPGGkoPSNSneJnhRDapB4gkgFjNCbtlEuZjtlbjk1/LOr8bxVgGZmJ8NzVqQ7AV+
gTyoIg/Qf7Rt0HwkDoclC2Es/lCqYUjWENS5iOlhaDjvAIwxGWRiT9yb3wgO9J6W
Q+kRM1I7GJVAvxXtuLGb6P0y/qyBNRueBQDGnqeWxCyOXu3Vu9StngqKB80DH1V+
1NLbbGMN0oTFcIR8Ry7v6M1BU0DF7P1mCW2VPqtRn9gNBRcDXNGQprEBbLgXMjnM
ZmjmouQ2xa9vGazn1+LApiIg31Go04IigydALKpX6ds7c9Z8dH1z8f1+fhV6gFsQ
3NruP3h7hKwuAHm0uDKnHCA7Ot2KmRWnwTikoe4AnFmp9YX1fDucqJ42y3OavNfy
xjX/RzWs1aphQiqU1MeXbtslWirqSp1Car7wts9P1Spc6YeVt/rr94xKB1s6BjxW
XlT3eJd+U74onHtolOcAZHcaYHxEErl+tsePGIJCJP4kj2mRnocnISZZ5pDPCpf2
GjHIYZIPu1v+9LDllf0Oj+2IxwLwITcdK3mQhKL/ItzOTP+oiZ4XnDHd463w504j
mI0mVIRA5tH6YVv+RrO3ZauzbO0JC4HCtoUQ+vfOKdsAN/4TRkFBaeNLnlj4axaK
YK7M3OBB5/Y4u8GKKgoGXK5Wd4c8p2jWEUdQbXKi//Bip/Q+G5Q6Hnwi9S8JwvHb
VXewqlxxy5pnBATif/vuNdakNsL0TESlFranhplFZlqirOiK3WjWqkif/xRgElCe
3355d8GNoxWpfINySd39fEdzPWDxtY8L0wnngibEk+sr6H7YOpQEnF0zmhN1meVi
VdU4wdKErTq5q44OmkNiVQRTGA8uNAY/ev68afgax0owsiifMsRB6JT9OBeNWLw3
xsh6Pqyxuuoxk/VFEsgqwGawc+4BlqA0whFj8C3r2rHBySdS62LNXzt8DUTH8BQK
3y41SmdZnsGLDvBy/deXNmsL171Yv9dxhQvWy6XcoDQDlu8Uu8fDBAxprW03p7DC
/LRVhuNXTwWKt3uYe8zB415I3T5TmV83oQ7u6F7Z7ePiY/M7q5gY3sMr8j9tPicq
MTt61HEo3Rbk9TL/Q8MgbRtK+HO4Aj+fi4YQZ9BOwsLFQo4wxiV2VEdFfrP2qPEv
6bDyd0XwrVS9NAl68O3F/IeVN7kyV5+5IDgmqK2hquAiHed8PwI+0/ksPe8P78GZ
TzuSqLwJIAIy3YZmmpi9khsMMzEmHr0FFDUGpHPk6XrsKdcI1w7NBd1btZvnhK5V
hXCVtELW38zFENMafo1RD8bEsUPDME9va7aEbtrRORv6VWiOuPSGzjw7ySiTMmFD
yoLZu6TLFq7SxD74b/9kYZT0fhE5J/HIWm1XbqkbT5Big/MgJqe9LdawQLNgDSAZ
HVMymx8729bqMFNR2U+JL4410Z+kC8AZUurzs93xHQwpoGZfI13/izWDs3ZYr/l4
Wjmcdd6q8YD6fNChaV+p4ux0EAKA1TJvQ2RmJI+4cQ+SbxakNu56Y7fsvFbvyOiP
9iu1jeI8ybC/bMxqEPFcQpxOYpCWOd2ms1X+gK2LvXuNofIU58FQPwup6ouUuo5J
YlCOQHbtc+1TWWnh4nM1FMz6MsZ5yHQpVCqul9Qrj7xxYgC3jCEDGXnoU+RRrrbw
6c8WMuPrHrUYa+T8hKVx/zuD4O5vP1IYb1HAkOcIR3XBJbyXLA/vZqGZub8C6cCa
dT+w+8V8UdXlaR2b3PRVejoirVRcfPefJAojSGMNm/+Z4YUCAHWnpeSiZOd5wUFS
65d3++x6FQXmVbaFEQFWk3o6uJWifS7qJk9o5Ix27fM+67tmwx3zYERE1d3TF6Ee
D43Vu68jjj6pP4cTEJ+Zg7k8S57tID//qBjA3iiMzcnONHCKJqfD2LlQ3uYJLmOW
PDiSohrx2zO+THya2PoDF2WNKxIX1O6wFLNwzSnE4cv9+M2JbqvcKRxkgYfa40YH
B6vf2NdjWabX16XiwG7G7AxP4rKOTAFrKJtti67ThjL4Vof8ukVEWsP+ZfDbSeTS
qB7eYXPAJs8+2SN0OUEX4Tm8ALu7EmnLovA4AO+6dTtErPquRYuMkpKE4TxchpFd
skh+TH3Z/eW5hBkEkiTQ7cEmK/0sPu0b7gkuePlVnuhF0hAjS7FzeByaqdHbnBXe
AJdDnWpTHBH3ZY8AN3eHIDnmGjOZRTE68K2v8OIX8VY8CdCGknrF0vYF3hg2A1w0
aUVjC8FO6/LKRt2PE7IkYxAkd8eJvDIhJ2niNu1HLFlLM10jJ9ZbRZl3kAXfogpZ
JpBqsuFrFO/g1XebVlThDQ==
`pragma protect end_protected
