// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:36:59 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ZM6LIju/GvAqDMKRHbfZRSDAoK4wNbSE5OVc5mem1p/lGRemZLcDo2SZK4GIqiSi
a50d/eicSk854Fuc43lOzUDF/zqG5InaND2g66poIvKe0I0Ai7oWRMEDGZ/Ijhw5
9SvE1D0xWK2w1vzpxqZhX4RianC52Tw9QoJCFJcrr/4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8304)
C/57jBKkY//+GyzsbNdw71zl8N3MGwbJP0tcmvIsBRegNQF+Z/3B3B7Ze+ARv/2Z
aeLESweEBSMzeLccPBuebtm4Jd8QIZ63S56FertE1jyfFAg5SGJIegW3eTxgU/WQ
+Lm3muVbDO8nOjRTJxHn7c8IhAYeSX6HlxtdutS88fkorB7j9zaRwWvu3VZQXTC1
hro6hAmPOpk3TF2jm1EF0baMgIoVf+a4/1Hlg2qH6Rjtr/UJAPa2lVICZdijRv66
h0lEtpADEcseNUmoR+d1Q/LXBtWMyHSmIMXj/SSjmbU8IC0dFKk9MacTbjXgLLmL
BrpZw5ejqk1G54HcWgdNS4gPqnR8qb/rIUPslB77fBr1X1aLSqkhA1kbss0Q9OqQ
+2ytoajhC81Al608UrQxIIzJ8DUM5z1u9zV4z1J8ZrCjIj/obonFjjuCKB0QXAla
zNhldyPL4oIwtup71S7Ek2/SYBHcUR6QOdV03jj9edj3aNSEM+kLu3xKsatfqKsy
+sxjkO6u9M5rlYXa1o0xtmcEupo/BNE/SmS7U3z/Vxchz2Nade4AOG3QbOL2L4Bb
5jYSZrMNYQpsPjisICIZ3yIj2VGAtFZFbu/yEXcGCJI1+ERaK/OUuN50Ckk9bhFP
1wjjuvpYwaCSlqDNwK446NFjXfZJ3VjeOr5KlTGHmJc9EsCHHDb+BcfkFKaLuAIN
AhkNEvh+CeFn1c7/G2W2jVAQ5BtL+JvPPFA8KGZkAooQVGKAa7sbwYIKB2CFOpTD
8I6glzhlZUCgdr2O14xGWxcxh0oDj15pP1gLEKhkwue0xdd6KIOzMJva/oJ/JemJ
FbUoubrlkYcb8woTIiwiOY9neUvvWgY+eGkqy4vtbnvjM1Wy/AVdUOb4OA644UpQ
tpOgjmGsSjUIUQA1JwgpXNYIkKgCYIWN5Ml6yAW7Bzi87W30Mxvg5taifkMP1kmI
Kyh9uElCsMQnoBGQwgzOmFGyXABvZe8dpiqEIWimas4yIkkpyfBAEcHYoqkagYmK
H1BAI2XQ90VBTGoJiFtsbs8/9cSreUz62tbvK5IqdK+P8Sdw/rj4zkFYViH+cCAX
bYmAyg8cwFVWbFWTSgxzelAC6NJx8Wq2c9jaD0yf1kt/k9VuQ9RydVGGDN3dM3MX
B3BTvs61jrbd/SQjFdyrwWemISPxFHIFRHIuN9flLOJb1rFb0A42oF5LlMCPJk3Q
nRhsRwB9IPFib8iwDBQTC5B8iI+5R5AtPLR8MslpiyYRmfmY3gX4RoowyhA5sh6s
AR2AC3UUs6XrxD3MkudZSNYapz6ZoUTfmfenre/ais7Sc6K//GnK3NHYJfbYKMfS
KcJbmkUIN2HvjnLWMrZ44CfrLctaR5tL7/HDzKTb9ya93RL9L/SyyR08PfE8I01g
mnCaiqXE5t/XjJghD0kc/N7Z9URw8u/nmxgujdyX1Wx1RdPVJodPNyfImbfPXSqt
LmOetTZchs9EMkyzA3hWDp5otULkF+NFxjinlYYNJURXW7y+bTNgZWfGanjz9yu+
y/3TB5p1xeSiBRzbxywG+xcUFuNG6iWDhYqXv69Ug2NFVR8kxKGgxxkt8pmPF3ij
I51Ks0BQo6PPEtaIkKe0ryyINZtV6um8ADkEXKOvY4Ejt9YtZCNRtl86ZT37j+iw
wMTNP5Ot2WG59/zd7dLOkw8pkCTV/wKCyZ+UR5CwiQ7Gm6tYdxfuX8l4rQQ594aM
ncLTrf9lfhIQL78007DMg+6gbvJcdfPTeMWeSHj7M5quvllc+puTLt2zdsP9ukVt
ILmKcJNN7k7O98HzDEN3s/XGFaBJzNbttPnHIXZotsrUhzwrcAKpRb9Gwk3NL2NP
h4mStowrFvQp89qwUHGB0FySYlODo6Vzq1sto5q7856abRPfTQbj6NGWogFBBmS1
MvxCiW4ZdhBAarSHJZrJIKxoJjc+QO2/zHSy8cRVDjRuDCSx+R5VNwCoto3kYKa/
I39+gS/vv7Nn1m01CO7VMZiPaRyZh8XSKPnJ+94EMJQLpN+RHPcijDtFfowAHHEu
V/0qfcmOG7yx65++punh/M+AcWxcW1HyJbQmQrSLQu+DkXjTXDRCQCAhfmwMDp8+
5QVO6FoRCCsCCmAIku75mCn6Ote3c+aF5r2zu1dxT4adddHFeDtb8vY6ETD1cbXy
+OxvH4jli0rEgGNr94O/L+vrjnHayTbTfijZAM5JiDmdtc3vtiDGYLvJOcq0pN3N
mJUbOEi2eZ9smnW5hAVf836Ws5cTj+32wHjUX1bDGWuMLh+vMbpajPiC8kznAZdf
gsnwJIQ0jmOAjQHYvyUDrpSNabHnXdl7tQfJDUHaQmqkWQTPEOwQuSLj64bWp8NS
tNTCq2XFWibYVzn1Moa/TW4w0fRDX5HdqDKVQfP7TWnOajQWXAocjjUNXCzz73Am
xf5eGp6Gjm9Cw1C4p4OviXXZ2P5M6xhr1EQhdRf1XPuM3c9vOXGDhQnLtHVNVRBo
FyvMM35r05B4ZC9m4x/XprhowpM6lGhv8QhiNKtGvu5/C5z76fVMD2PBSbSpGw7p
I0lr9QwFgCMl1pbQMaPusvv5IvfA5AYQ6y1O1nzN22VOqafGGIcPARYZSe47AQ4T
6FTSvQfEJ+C+258vJ8WFcew7nPgRkF9FF955JKDPNzqQRFHi6jiCE302flwe3Aee
deqHnvRolYPF47bMREASniSzlX0wXfQNPezbAC5z935Hcq37wbqVwcJQtOOQ0sEx
hB8P7ymY6Dmj6hh0lrASOMC0HidRGEVymTbqri5vQXdKKnrhElyOm22fb0wrba7S
f3l5H22FqDuRCkqBJhRUDc9Y1+UKE3ayR8IXO5RcA2ixPage1MD6IGb17v7sQjlO
jb3KKYxQdLROcKEKW9/qeJpYUGjmgLV4/5n6eF0Jh9ObINZQWNw9xBoqU9XOD6mk
wY1NArEXw8iooaaOp+nFzOqVQ0z75Got+ezBOAnQu/ntsd29SIXafQ8VC5UPnNpB
uklROfaWcXRwwBvJM4Vb0T2EISy9Fm2knOLZ00zibw+N5UmZtQt6EawVyPd5tRgg
qFveHm5+Y1e8uBzHQHoPPdismw7eJSB/gnTU1XPA5NHwhCH/zEfL+ywN7FlOkRu5
mmOmVm8MWTwkCuApMOUCoC3quDiDKgpdo9iH8OEGZu6jJDCSlso4goNqdZkug/9N
D/ClZuNuMCl17kOrsKBgSSRnpwQqC8NkMIvtzr+VRo3CeBSbBqFYAfFptZfSarPz
mpNCh8Y9EIgqO92hxstc8ktnI47lyL+GDC2kdpZZf0iT/DCbzBEU1Z00iW+Ugb+8
Yt5aGXHi6mM8bhRuEP2jz0jYfAxOcotoopE2cdSTk5CbQv7ZwY9Y4SOnmW1A3auE
E0VBPFYWEfRHGqI0ydQmD0+RAhanP9ejAbFhdJwleZ09d13lkd2VWUYFStiuysU/
K3mwsHyAeeFXi9aJYuwHsAQtpQYAVZDRbeqVXRkduEZW5ScAuCkhiCWDWV5tqpOS
1LSWZId5taVy6LYjlXVp1rI0i9u9Cyzx72l2uBk96oJOVC71rPah72arEdlcJ7lM
dmeONMojrZchHyN4JCKnCY+fLErCf4TtVyiX2y+x7QTwini2rIe9298HL5zaERj2
Uh+zevf2uav63DX2ovZgeYVOCvigAKc04JlAPA85zi8/htU7XTJTCSg05/XjLQs/
mi26M8QttISRYpIspe627IaKTW0fjmOj1toRsdjEhqIlW6qI8GbE/hnole+BHFX9
fj5/G2xoqmSjJH0wJIyL3qoXEXNHOqnUP72sZ6HQCmxYlutWO22Lt0cGvAvByk92
GivttphSzsNNZmL++FUwOWRfTXKu+GiKpM44zL7BCEwDWLWxxkuYSY/LuHez6mms
N0PKax8klncAkBLazyIilrZgLWZurBJPpaq450yvkNl6El2VZb6773wZ9xr6jHJX
bZ0H9DURtD9iNaK7hRVhI11dOOeNsYQaLM3E7qiT+v+RMiCM+B4V5vpC5QWgLf7P
YcdDO7B8wKWRSJCDYDCY65ydC8mqfN+aohCYB/Y2y2KvszNZ+ygrOg+47CeuyTdI
+BzlmFKu5mYsk7CJvYwW+qWSyslGbTcShKdySuQn6ESgSG+/cKlZx/B9R0GECdUV
pl3F9VUg+E2QTv5dgqDhbB1YrIYzluv1fIk5Y4QeRGFhK4r3YBak1RGC4L10CTWa
Bg0/yvnICE9wN/yvyHb8cFMeWSjAURxus2lTF/wLpL5jJph1VI/d7ZD7/z3/rTyB
DYH6H9VJAG4tqlVbQgLWf9hNZVoN+KHE5udTCewOTFoloiWGvLzrkB7PQFbhYsJ2
uyB8b6xiDbpKofQqYwWC123l5p6jntv4RL0m/ElDhbeuxuM7wkb9vwiM+MGsV0BF
BxPdqEgPPgeK5oOWMAFxsm2OUeipyOmZiHJgA2v8lnNBtW5tAPTq3sdHVTDP/279
79mMj4/gepU0eIZoOXTSWhYucKV7jDrgoyfKIg3JBOu1tLlne/FzVWG/f9MZV3At
xVUq7FQDt2ockrWDeMwEbRlRIJ0mM1vlHjAhyFz4GZbHmCttCOoQWRZgYocp3xtx
44GKdyfdefX2jZMgPWK4Iwg5JBfK6Cb/OfXpHZVYhhWbocn1Rzr+R79dRjaZ/L1O
Ruqqk7KVKMrbHDM91uCimJqFDTW9n+boDcPmcgqgYvVzW5cF3+G4nVaJx9C4/HLN
8GriIqo08I6pwlKnPcAIVrhmGSWlniQ+zgcjkC1i3M/9ytXGNTDc2OsbOzm9BmeS
ffUVygB4weRYfRsMHpipUFPEG/kmwvzs97EulYaIXFcmKO+4M1Av6hHmRKch3Hmn
Ly1z2C4Dek4IAvVUTKi1vSUktNwVKAplk6UTNZTfxkFmLAWozVXZ9W9RhuNrM0/P
jxdaPekhTWIV3OAGzAvPCoExhoxRPYi4qXLkdcGg9HaMsC9mc0UJUlKU798VoBeM
b40LmkiWASX28rvdf3BV1SxqG7tHtnJB/yEzS4iXoojPHiypFtbloST4XY8Z3z7x
IDGqj4KsZc2JiwLzO8ZLoAA10wV+1yMmjgZfhFIdtDXd4+9Xne3ypWmbc/VpOC8/
jjiDP3sk3fW6BQm/pJtqFPKtmHSxJXPK2HLJ3MnWUe8zd400urQiWX+A9YToEdxP
XtDRXg87DKVbGai+tkvk5pqPtV3/MbTytywRFa6dZyavfgSfY+bXpHQvsOP1r1wg
s2qw91ZhAqK9/AOno8qeOWxgwLSR7Lk6Bn4SxbFY2ncCkoXeVwSGI3flZad4lqUK
1dFeMwSDevnLEE62a5e0p17o/BG/FoVHLo09YEzrS+Z9G6uBLvipTMrUAO6GF4Lt
9XtAVdmxBoqAENggzj7wqr7lL+rq0t8VjoSzWmkAkHB9ycam9hUhwCu0Cn4oTa7O
5B2h38xgwECutWbq199+O/Kq7gHbSB/cew2qLX2+DKaRFORj+mnFS2OTKECP0oF/
i2mwwKqQDDWy5SQZm3hGEzSnMGdrRBCkFGeMRpmXJT9RtJlx+/ptAvnUY7uP9ZG4
kq6AMrrrsfwCZl6eyd1sX+OTm4P5gEhotDiQI9JT6EnVrCtXIyT3n74QenEaLjEE
n42rFVM5JFejGsouPslqcyORITD/xe/3+65u3INRuCXe6tvjTqYsDbmbvNFli8/a
gjw42B3u/dK3XZtlWlqPKp27XUWGu9K2Hkyztxnofnl6QSFwIp8H3mf+sFwcGAJ2
oFakSp5hoRMBAmYqjliYQQQnU5I9s53/UmEAZZ8QcrLy5Z3mjbxZQlAgGVsccBlG
OQyzjL7SkyWPMNaDp7ct5t9WND9ZRx6xiZtQ2wEJvVM+QeDhlcw5uUA5HT4rrzLp
XXUTJt8YL/u++PPMY8ZFx1YpZN938wAVDJdHJVWnKgwW3JVUEtGd0hd0GTfOj/qy
cJpZ3R1IwFngwhQ0vx+jrrA/a3TgMYoPQI3+v6/EI4b4hkhbbVmQFo9tj6yshTil
cZu066BJlscfvesTkvVuB1PJQCvS467wTFOwjkqcbRKz5v3YJLaq7F4LAe+AHYAt
W9Tl+vARIHNiBdMQ4JGbmJSw7XPTH4t9GRupbX5gM7D3XgIi7Eu1K69ol6zNXmyh
fivAvdqGp6+bxO4ADu8+P0JdyF8qsdj+mhCqglD2I6B7cqW6GPNma9fYB36+CGKd
J9JNUFhPDbTUofwZJ5KcN/F9pxzNNcjfG30ERelFOGa7LV0sCpkYkgaSNOR+OVKv
hkmwXWxWUPE4v6DlTKDlI9kEw3RwaLczW8rCPcZYGtLz2dtDD5paLDz5dMaNIPhF
kyhgqZk2zpNB7deUzRJ3rU/3uC4meaK0WzygI22sEwgZvKJWbKs0v9BhZCxRKaT4
U/Kotzd8afUGj2zUGu++OsBVsq5oqRd5QVNe/rvS18kd+sx/iujwfjXBKNFPkttk
ujTvOEzQooQNOk9YK0Vm4z+wy9B69IUDc2XBaRMS/aZQ0o1NCr3GNQNiIW84jJ+W
KO7rLIsnm143e+bAtPTasB2jKkmyQ3yIbE/40qdT5Xjn//WBekt1WL2WNgPk8Htn
67XIMZiDjw+Z/LVSYM8P4IPzrOilPOHT1sTOgQztOL2bzPT1787uouMLmoHyZM1a
UaiuvUpyvvz8AzETvxuEQIiqLNuB+1eI5IGedgvzIMZeKBCmy7bYKuEnpKCZhnt/
ioDqflVC5tzm5GH/Z4Yy7Ns89kRodCI3r5/w4KXIM9/AwLSbO/PUKsszv3xIxyIQ
slk0fED3GaT1P3BkoDf9fUgvjM79rM8LY7MrV7ecZ7QLtVB3163ieNJ1Awq5UJj5
bXm4RgVvKhJ30TV6MkGxd10duRR7fIqSM2f57S9r3dodOoNHTD8ezQBPG+SvYIm1
oe8Fb38/G/Qh1Rc+Sq8odPcWBqMpGPQKVAp+Ij5vjFca/l2V4DKIy9ZbZnA6oLKf
IyQAGAxBPa4AxwbGRIM3PSMRncHhAhmKg/wOSIeTddr1EGIxTweZ+Qcp6QhkDzWg
I8yUZBgeR3oiewYj/Z6JVhcmHqkRN3yoHXVO4mtpsfb9K0eWD0SYPj1oOXlgjjYB
gNn6XHEDG2NViu9zbKTP2BgVZb0ya89JgFOndWp3IGicqDT9brkT4RaAWx7LYgFl
TriH/k+LQkf8obPGARALuFKo9HGXFJ8DUEaR5NV6XObG35LXUeGQ8sEDUMwOJgVs
OxkLKQoerfLJN6v8ZxbJgv2C8jY2YYY48q/6WC0yz11bS+9fra8GJIrjhNRFAHbK
8F7V/u4i7AsBeVlPh75TbuQ/qYlaX6MHgUwcWl1JuhBA2t8f6lcXp0jOPrY9DE06
/NdvarqPn1hb7UTnt6R+HOwV44KDlDz+S9zHMiF16ujWm4vVxx1mVCZodENBH8le
kIzJtHr1rN8b4E6/OFnUrsxR7OTTPwDfNWs7t1Y0eQNZRo1QHOQWfrwKVcBQB//i
uZilwynfDkfNrDwVLy4MXIysQruLmly2+2NVAlj2/cmI+yVjb4nRSsClRY7P1Ae0
K9GqRlDLwRjYY4goUC324ZasGyq4nlmGdp0Mso1Iuy7XFwRtIMJKgIDZ9RMU66uM
TS6iYW5xsYUNKVwxhmdBov4fjyqw+rHeSLhyT2G4adZaeJEX2zjCLeGB7KfEzr3R
xj6F5JDrej203rtZOp4pn3jCCKXb9oAO4YkAT2cvGy62HPn8vVrOSv9V05exlpdx
0RNXNHvIHAX975pDf48Ra4NiznrChbZQ1sfmOaOAE1/3rU97L039MskRDA+ftjqK
x7FKNi7oQkngt3gvT4UyjdZlG64l9kEUoJmE5smdPVtfMwyZToNOtD7B9XrwexPM
cly5rvoOAd8hXZKYowBoMl73bbfFiXnCAtEoYSXyl9MOqlqrXTlv7xPhe0aiJnC8
T458X6o4oebT1PTh+/XUVWLEtFpFyPoVXIr1UTO0ssOZJLiQFe08DWAiwnBEofPS
9UVI8EZnE8/8m2+gxEupPZQ/KtHXb4x3FTiK/mSuMzHiLJ2Up38WWs4YkWcIgNXA
jt+Dv1iyFM4jGZkh0xtYIq3RKjvK6ZO2bDNOMU8ZpPn31PuPzOqg4L8MerqoUmdd
zqV+N3SfHgA40Ym05LhjQMStGfQBuvhMxdDMmfZQfl7yhJyMTFUAjH3B0OWo+6wX
lX2mTv2NEk1vk7GF3c2QlEJ+R8K0keWUZV/zdOXiPXcg2GasY1APsgsg0ez8AN3i
sv5bOUAwb1MfedImc0keUoCqclaCLlwwZRuaHws5a6fGiCRsgNgYpDla94b5jNI4
jS7UDh06FbbKytPaXdx2WsCL//3233Lr3lNhqxSN3NXnOkVoHF/qIeiJydXl93ag
aow5ieYeI3WgNahmlPwHCBgdgTx/9p6dq1SM5RQWrxh76uaV4czjdtF9d6vkmacb
z7MS49pa5yVMAoLbeJL/QmDKWxx4b742Xtt7OqioyH5m9WeBTWPOfav2M6ScfD6f
3AV1pwiNhW3Uuxohy7PIjaRfCYK2YzIq7PmfDuipXqJHeX6snRGz+zVx5KoLHgRp
K0XY5CxgIbQOHtl2vXfOa0wJTL70cmZFolaGSFepNi+TcEgX7zEPFMl4NwYpdhcq
U2hXiQIgNPygPUCzfiUyYqRv2JZHr4XI0epCr1KE3jI+UCO6LIsv3NZ/uvZM+mi/
U6YTk6JmJRs2UWMRCA1pxQTv3Lm6bNLzDVs8/iMSpqg7+tu3WmxmkvlwAxOwXCdb
i1qma87i8ydK4OfbJOAyKuhDl9MIAaXSVPh/SS4SbnKX/PrF8Lp/jT0JGF9g4rc9
OY1Y4zvXLy31fe3WyUU7YP++Uk6c9sr9OIB3SxF3Mxfrq3qxjHpaqc3ZVB+NUH4O
AToI1BdCKky9TnnpTr4BzfUQGJfh4tcYhfsZEltwf5/6jJ8D2d71QvtobQukP/Md
n0q/QmLhImYsKQxWFKJu81/MW0KQGrTxQUDpIUrTzKSMZPm2H0fe3Zd5x9TvARer
Jh5y4Jj9ho1DkUw+LOya1dVN7zVu+uQYiR72VLNq340IBvaGZTim/lInn2Fw4l3k
d3l7RTqN4k4d7XMMU763CXh/B+UCkjgchxJ9xrp4WmMI4hmoFXw9QL/cHMBpNpcv
PmPqpveSzP2ldqHgd796pwxatJB+cl0cZeBjz2zHci2eYTniyt1Dqjp231XXJBID
fY3ckW9l+P34gNRkluIavY5mJUfb3pb/ItmkaHRW7S+nW6kqHgGQp2IOX3bmucSs
Qv1KbR7e4EOwWxlmbUE7j/kTkiwWrMWT7x87BSJFq7bYsuU3dYO8xzMt6NxiOrkZ
D+ClTjjbLk/Hw1PcfHSeZ49zNLaGSLcvzu4C5pa80qLyjEwX+aCuMdSlycBYcf7t
xF1K3sKNI7hvYlvtczLn3ebA1v+CNc/9loum/n6m38vD9UaP4Y1SMTwJAB9rPTJ0
Nes+HT8u3x9CrIK9MKubAzGFM5xtZIUC0mWLJ2Twcje1zj6Cm42qKn2f0kyMOF2c
pChEI2Boxe6mu7BWR/XSXfrKXhF30FYaxUjypE8hqMpUEb5k5DIubfAqf5s0PtrU
Y9SqRSZXWQMZCKNj+HfnRDsM3ukTwV6ddj81kU9R7OZlJmVb3Knq9W+DUuiINsBQ
WqGvpzm6W46sHUHO3nBJrphPmFHK7qKSmNThV0OaTuuXr/sd/kHCkcmoLPURpPXh
vRQb6oD7Xu+nmveASQOuqpnqhEV4JXSqsxR3BAVbWShCgmNlTdpMmjJou9zdgzEZ
Rz0SbPOb1QWzHo3TBRRXKsbfcOwLUsYrZsUNOn5JOjE8GDfsfdv0+Iz+PKnHtUoY
mOOgGHPpUreanQbroWvhoOVhN2lXrDptVrOkO1x54NdE9hJrVMGKQ1GZ1DV5fefz
UKUZ5HOrhYh/xXNncD/Og6da5/CAAe51faDCa6QNmfOU2u64yWqcN8fZlQgc/6lu
7XG3uSM8k3CCEBSphjpW/JfzbsmVpA9hvNJc3GRCSd0/WB1dm607l9HMoOw/VPCT
WFZj6dWM76fykOgu2MkrCMcLsH0WwY7kgQuYh6msaoAJpgM5jFWg5lTQBRDRJqvR
0ymG0BDgs0QnSzqxOsRA0Z5eHplmIjoaGdAEDD+SAbhuufhsoZvo7m4e3o1ym4ZW
ulmmgXuIOTM4idFiT+yVn1ckfnSy/AiqOUqlSJts6UQf9grdVELQfAXHCrOxbDrH
d5jJ7h7Vkp2H4bw3nDpGthD36VJk9jmYa2jx4f0sYG5bmx0sV7Fqo/kn7BZ3xUbu
3j4h7D6CZuoWUa0on/LJ/nfhpWtmusKEvqZ/pCt4tWQY8U5d7ZpBObz7cY459yfi
m5VrGJBe2bw/apXh7gC2qDHyQUQEaaDIKeJiKnPSHz0tJdu6BYkPF2pjvlNX9m8l
xjF3jKDQ3j2VITjN6CijV3viFXxWTdtufpr2UwgyKq5XtX6CZKJVyUYjnsu5UAa6
+PCxVDtIOBavURqLIixXMrqM/n8IcQJ2Sqlp/bW/eoSbOKWKtZtJ4B1augp+frZ2
LbTjOjRVAX6gNR+NA2SWygJ7FxRIg6Bl9b9UyOfGbPqyf3C6hGIYCwowN02eZDyX
mzdfN0i0sl/mkYFygJQpAQonu1PyEh0NS8WNOfCeHrJNuFQ2RtNpNr8HxqI+m6e+
8cMASzMyMjuBn90A1RrFL/zAnNwXDgb8Lax/RnqW43i8aDpC7mJxUaytHozkWypt
nhpx6PP/as89mtZrnxrZE+6a1iInlNryd5MXE4fWiDjhuI27MYawZZF0PzAgmNAR
gLJ8D3iAFyBWP3pwPfrCyPdxfqrwg/9pP8n+aV+GlqVVSI7W4yD45GfIkVL4lh4m
sEBcyY6XrYA1uy1kuegjHIwaYXmQolHxWVvBxGxmkB8SJlj28sNDCBlYvk4UXvxh
8Iksz/8/pjORd21fCBWXVzvwva7of3C7shWJTLRyPiC3HeTWiOT14orm2kw2bTOW
ljyyIppuHQhBG2oKtX2IEs5125gZJ++P6z8Z3CWPIb6QfIgYv82aHoa6382cGjBX
`pragma protect end_protected
