// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:37:01 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
HBdQUQl8lmGq8O/X/5XpR1NUJOOMjyZaisZEA1N+hgkvh565sglj1btf0gdG1Vod
B74ie7mBWELJOPbSlZbSa9ydCI4pd0v9hR9hnShq9Z4TDSfty48oEGAFsu6zxZ+P
MkekrMFCqpMKfcfV4mrB5fhdAU2Llq4uAWUYhfDg+mw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 22448)
xj0jQHIuGNXr6SsMse8WJtClDsrxd3eluOGLdpnEjfKhnj5vi5LA8y3rgqF4DZ0g
Ma2uMv7wDqBCkAkPbee2Ko1SChG195qP61ChfVAEGdwc7Qvrvj2nYyJ0Bur73tDV
JfCQ55rTZRrjb889jR27X1z1j1+EMXLTYf0lMspzc/0d0/Okf18aFL7rDISC6btw
k8x3lBNIkypIcVDjUBDrAxwmLWI9znaKW2HfgleegXNNwZoIoxwySVs7TmTA4AKT
L30Se15rX5jLSE0M0GKENOWUK22WLbh8cLZiGzxQ3gGXQ60jaToNexTbr43NQYu+
8L2MR68x93cOGb9texepcKG4ykZBXYwCY4Qg15ZFm8YNb02EdIHaA+szxoo5MNUn
3Q5UjYBOAwbEwcXHUL0TIWeZGJLT8DVDk4RA+H/bTDLQFJBYmNK6V4a6NFRvh3Pn
ISFZqgRByD6skkEobcASFwqN7iieyFf8+vOU2EOlZr1oKbaT0LUHFYKQ+0nHqUfT
pLh7Ay1ySBlO1Gcpw3zrypzPueShlgqAjHcq5yfdkjS1jiCyq4RiAyR3Nc/sw2y3
q9BfP+6g2EZl5jSNvmdlGXjgtL0fQgNQH6ozeKp3JVFZC0D+sIGAV1QgCsebZT6r
/KeJWjZgyUTAjc67jM9fBzl8i7Ui0owWUFNcMrl3IPx8EjpZRSzcTPIavCUoshJC
Gpie2IwOKRS2XyaDctgngjOSmYFRZ4MNG5uYVJ8tGa3mbbU09oYlFdKk7MXtjZ7q
vHxp84LeTI44PJWsZvKODz5vS9UKw152XQsb+laT3gWmrL+cDRGgUXIQsvfI9USs
BUAA3ffFomD4jUyyXb0SmZu/THvPLKxVveOjol5T/HjG4hAllIy0jZsmiqSnCf2N
gPXoZDjHtB5D6iyhMNHnnMBlrnYuMHaAb/TGDJDVpT/5ozG6smypsa4nEA0jWqQi
W5moPJq8q7y7d1VlZHh7OMmx5q/iOCIyzMXZUF6FIkADSfswZlKiXbn/3hZHQ678
xoDQx12jICAwjAIBVvTki1rxXm0QsnX4O9uGrg73LqugkEzWtTVfQC29Zbt5q1d2
MpJa6Xs9+tlhWVFKmCVQPxwYqVmhhUc1WYZIet29yvE3sZuEZVSDEAIuaMPeivuz
aNeKIW6H55CU7Kaeu94SIjukgBBBnABYNQs1FlJWntNvfza8rsVLXul1PqiZmRpr
MO2i2arVd3zKcHEwNDCa3QgWS//6l9sQ2grevq7bFOx6ODWCNj2dKoGTyjeZzEEl
oloUijwPJNLimmz1sLoLEoaanc9TAz3+oc0DLgpt6GYCOrPT5MoWzfknB1vgFoVs
lIGXBdoVtyMBlIWAqc5tYXTGu4YG5128+kpYZI3sBe7UWm/rKzeUdgVkAe8o9JQI
kTMhTq68V/Ox13VwphLy3mf72YDBUqKx/eHk5bj3XJuzU7gP4BucSaNAIXRNlWEs
zOrT14uCcbpTq9DjDcyujA+ZMarUmaHh3Rz9Q293prwc60lKwIhr3jVabryfRHF2
iZxY9d+6Oli+yLDZlT+n8Tz9r1akHIgkbaWPw4oIFImPsSmR/JBU4ZnwY6b5vOnc
M1pjR8Iom1/JxdoXS+U8zCwio0A/kOD4CIi92IXxpWatvBYMkxWTp7lWfiqmVPkz
Q9POzqStivYMBBj9hGrdXzdUFgDFqvdLOBFlVE4O2UlYmmMYTbIr91VAga3KuRIs
gvgtu4F40O2tVBJ2eemgqXMtEPYPRvTccLD+l+3VQdlOkG3P2qGaEw7ux9f3RWb/
kbFWesAqJ7MgUql7uOxsB5623a5BlmCzT1eG10vO2WJlZt0vh3/r5CgiJ+WS04vu
9B9Ye0s4hQw6xAkuBz+rx95wSc4A/PLhTgrqlqBgGLYET1v4HqV5nxddpFDccx12
PbGAQ/D87mHOqRYQNCDHHCiKOKfVeE5EiqfO+4tJ1R9Ae67r6Ia8jtW/Mk1xo3SH
mjc4pwNpLl0l6w7pnOm96jq8BBNbMbbyRWC7npthVt8S9mbSImfxedMLPoOpD3HR
A7Fif3/+NddH9jhXXJO9tPF13UkPfx29kT0FSSm1f0++nEk8+lc+p0m2PvERgxXA
WmSbb9v82VEvra3LzNfRjZZe7JdDVHRaO8dI0PYYqo5e5+I5q6FZ0yF2BbyK9lAR
a5vbIz7MDfqkz1uAoldpH/Ek/BnT5UFVqIjONOppXdoQPGSXJAM/xvF/Rz444c89
+Pa0UjVECM+CTRAsTEt8K/jSUQKqyqbBFuLzrXMyGaAQGrqGOOi3q5hG0Tg+kywD
NOJ4mTcjktfLd3OZ6EVU+nClGvHHPNbfzXnjs0xrl6APB0+XG7gGEaxZYbh8iWqQ
grScLg4dDFyk75tHsYqBEVeRhtWYPVJheF3p74U1OrH72GoNaocV4n7PZW9eeHzh
WC9oC0sKaDKmFp9t7iDb752q9Oe5cGJIXb4wAYjD97KGUroYLaIQ8PAyXRMA5Ddu
mGqaqptIDkWbhuwf+rAnigHzeRdc/DqaF7xwFPRArnz8Ldm3cKDmV0mbo8K+kIxn
b1MEq/9Vjrfcyg7koTdcXe3w1eSPSzehQbIiuE0cUcPRK5wDUEaSSTOf47Fcd2F4
XMWgfCU6JU62uIDXRtQWmWYuaPuhAm9qDSaAdgx038c1ZobpHoX7e4jX8zp8Dwnm
hMqURDYPKdROWL76se8WNoIcm/OJ0ZN0hdnE6Ht3S7lj7wPUXsJFCUINPUuRTjj4
iP2Nmyj9QAgny7IFkFUdDn9hXrsnAtrRYy0O8l3zups77gFMgyHG8v5GNNtiR2jL
Lthm98ZanVocksjcRHNOFp8RW1p3nc96fhrQ8WW9kod7k/HcbYrppwyl0wY6KfQZ
clk3LhDH5CsfRi8OjI7MQgE0aQZFLSavpj0ze8IIX8B+zelMsewYE1v0570I6EWo
bTW6nmHGDETsFjO24/uC0Zgpg00VnGSnDaUxnMpnXDsWVrbv1/Yx6Su5kMtgehFf
zwEB19c95oMFGU+jvXhN12PLIQ49QzS+JwKp0M3QfK1IYCB0gMVrSGXfX+gBELel
5zJ83DpI3w3xZxzaQkK/e6Nu863xqoLPe/1RpVpStTB0xptjyrOxqkJHc6Jt9NjC
jljKNZCsACFq2+B7Adowwglog66yzoz/vZvExjhNS/8YEhU22KGVE7Yxf9Fv2sv7
BjBBhLN5lVlcNtQMRdFTwlg4f4IJnDTGvp0tqv+ZrmO2TyPXgWUA1rVQh+i9Vc2i
J4G8rfKPn8PCVxP8QVoo7X4/aK+yYrxFhO8s+XexgFFza9qG698RN4wXZf6tbomf
su9Q2IwmGo8Wr84A21VoqoF/VNKobmx1EQgn/dy+4rG9pUAEF+J2sFgbTiTGnxv6
Gns75QclAQi6Lk/KgRPJX7y+J76V91qLkIIxLfFiRg56xApTVlgiqLYu2k9M9UYN
VRepx3u4yEEmOyBd9VDTELunbp4W9WQov/bFXcWiPAo1dELtVopVEixMEIR4lL02
Ni7CJfWJTJimBXHJLmyyvVt1BJZU70HkzyqNRhKLKpaNvK6bip2vbg0HOw8k+Ovh
aUlpMX+BFAcsPQ7HrfZlvyec7lBAef2v3jaLlU6p5HIfWY805c2TClY8mMXZ4W6j
Y4P03YTUf4TrFkH+Su7DGEWdx89TG+3P1AZXvawhS9wlQYc8UxMDSf4RFLbizsjA
+YsSD8FjXfAzhs75BBwbf09mW3O1WRJFSQNIWAxc8cJAKqrgC5hNJ20EXuPHEro1
2w1Aj/fACd8hb/NrsBhLM+luHxMiY3N8f8wAb6tN/s/4pKSkquLA/2Fur5qat+bc
jqXVzRo5IDpMQ4EFO5+S5MG4k8ImAdFp8AkAr8D7UemNjqWGnKLoxWx0/HFOJhKL
6DtrsaukoLQqlJFsW6q+I/GOAX4/F1HUd6yCxKmmvFCV8gwFWKVgrUsdaSbDyPtq
Su1CDLpZN9ck2b3v7zmyDNv6EEB/ZTDnbSBdr/Nb8PWTpmZI2hFereT0k3LaqPSQ
i3ncD77Cip/2qfzK+mm8e4kEF9Jq3L8MlixPY1YhIJetziQvCQuYpVUY2XvR3EQ+
EueV/43kvJoV4l62Tgs2yn04jqynOEnPz1mY1oWqNb2DKvl7387ZTE8f2arqGQtW
/zTEmjN80n/XCNKPw2fpXeFa9orHucuZ4ZB74C/sxdBvTL+9aqu7wOrvvL8m7HcW
JWuxS8jZV0vPSWeI56UbfHTOGkWAVKJeME/JKNw+o6fLyZ4iwNQhYuu29A4bM3Zf
PkNKtCjiKd5+7BT7A9wFLitoXYpIDo/+8NQtz2CwqvF2ZAyMu1CbhZ5tJycpJFmA
+VWGHc15zbFthhaeLx8FlOT++U7IT5OWZqvGaDrMOBZob/5WMHL0CkAszkMvefKv
z61gF7SLIvelgo1Y+hnIicvivRe9z/eWeAPBK2QC2clEIFh6gptGiCOa66nPOqKD
lcORQxPwhhpalYLSMbNMH4WFuFuOpdI7SvJujzPOL1DuQwOcPIdPjAk15IsWptcI
Xcd4GVfUb8cnPcfhsZ0z/uydCZY57v6aic6qAMaaf1fzxV9ed9Ttu0SgDtXARVv1
eToyUidp/duUKP9bI4g64GzsnhnCqYhqoXN8QweY2NaLjbtdwPtKEt7yLC9eTeNB
hbVsYL2U+xVv8yo8PgIwR5lqy/I9LuuDWYc3mpHokHsqdUjpVRqoFFEKE7kUmWe8
i5OO+sjExlM+nL1FoNvcyEvjekTTrGQwVVl3Nyfi0+SDwpi3+ZwvqWBEqWipMnPY
Pc/01txxox/mnMacnbD5MuPsnhFXtAnrZ9XozFl1LUfj3DX5RdBh4gQXb1SyQ92q
uKDPJ3c9pTs9ARa8qi6G2V2ywQp+Wy6Vp993hohh8f71yw3w900BXKDexY8sdXKM
vuouA2KOUzyMDisqwEgY/e/fgEfW5RhkbxZAq+n4gweP9/UsEffQpb1LDdhmsBIB
mlvi2HdElgu1uyEgC1rIgj+0DHCYbA6f4rxjAMHdLkLgYfTi0VTTIpDj7OD9txdL
HgI5KvVuIPm8N8FHjzALVH4tvCZNOROJZeBJC9LK2NHL0x9sX+6oudusFFDLWJxT
sfKv+4kZEuHRmwEVNJxQ62Ctuhmp4NQs5YuxeoX+Z9/gJLB+5dpwC/nWgp5TyOhA
Wi84wG4TyLmdz/2IN2S3mYT2B1XCez5ZPzCltqTR8SQYgm19xDvyCONj9A0jHISg
cp7z8Y6Q1Ia4rDR62fmKUxMl9peU8MJK/vcdVc4Rk1dJmPoJCw0t7LLIGIRXfrTn
YX9Pe64MYbfIMgJkyzgI89NwRTsfO2ViFEZ4xNDr7SvTFcry6p3XNtApFomD3ABW
L4FqTctfTZjwA4YElnqNKJcUNq9bJOp8xq0zkxAstjWVuvBB+pNVf6+fnjEUqch1
AUmFCmd6yULYoGnYzbNklrAy1BHSWAcn7dEaAz05nDNPHkuHQuvRuXVo2VZeRpdm
FWNCbfg5Bsr9epD5oYvci5bEDxg7sSr2Fnmlakmiz7sG7lU7YPgEzGDd0zVLapnZ
y+9ylUOYI+jjT8Gbx9vHjzCpnuNx1Xrzonn0Czz94w3O+mCNfC9qTraVARTPFCHr
T4X6RpkBbxzsXT6zDuPdLlf2H0GgY1D5a8PgVNNbz//Ju9cjLGXpSdgY06suiekT
S2G5G09NlbypIho7tb2jL3loJi+4WDlXSzwD13tH9Ej1tqo4OTgcHJ5vGoAwLVr6
SDLzmmdWzbE+1onv066rXHFXhcX4jLnZzyc3NcMFc0PMP2bOtr6H1ucGjRCiotru
inNfavYg3B4jzbZqEcOsArU+l4IE97GhfM38FbLVcpVRXR954kC4bapkLgaetFSc
pGGa9KQ19o0iVNjJG+HGzD8tou+35Mw4cDS8JfT3ULVbMsAu1WLJ7jCiLStHclmf
53dnzEMV1aapOI2ZZkdJoun4gliPAg+lLYPBZiBty7yjAycCjVxFFFmij7qdefXO
jpfcHdZ7T+vZoRH2l43wBuDOpNzEQQB8JFB6Qdi1eZRcrmJ/1hd4wrplB4MvDX7b
5H2ZrtlH7OWj5bsi0uw4YWZF65IVwjc8TZ4Dfv2E22vd3fg3J5vL3iqtLM/l0O8W
ebXaPABrUwP4G3Jhvs8A4Uy00+7SoSHCRmSuEwNAq5Re06IxSeOhb7H3wphPSulw
BlOElGxUOsQWdMeAY/EF+REsoFvXDYLNYZG9My/WpmjpSKIhArSGeOOMrng7woLC
5hVB7w/t+gOg20EjuWjgTLdNbNaTjlwL5ytKHNA1/5aNdTHrVwn54Xemdjz1YvPM
egEVGP3w+ySnj/y18TM6C1h5wvieMOZEug8/uiCvpDpNeN2xVTrYpgGus44gq4zq
rlMFVfaJKXGrLpWyvvimk40Oq4Ofw51mvKLMOVW16sWJ/tIIn8IonWkf42youPX0
at6JsKC2ZIUrwcDEU9ZEU794rCI5vR7q4193p7pgeQCTN3zDnBcqRYfWmluCet68
fWrgohhynnuXdSnfPgUzIgpjK/6V2A7kXx2ZHGPSAd+hwjuUjO5In9tPC1ZlK4Bk
O+js8SzHhD70AOb0eMO/Wb3+qkzLvBVTPLOcxveTh2o5eY/HouBqvWhT1CGNeUte
hH3nueZ/rPtlR2uKoMX5e0nPW05T0oycN829TstQ2zPc75p9cvaR2nZfnj8/tKMf
vn7+/w9ErrhNUiQCxI8c9fBBH1ZZvsU9dbkRX7sN5sJtIhEJPqMPacltExKXZA3B
X/toXrY0gDCVLpgJRziPvq+//EqseLBpcqdugM1yvaVyGz/EPAYVARvpcIfwDZVm
hQqjm+WhBic9w9BUhdQuYaPufa456B9VC7v+Khmkh0TKVMOm31irFnuqNqbamnPn
FajFC1pTj3yNr7M2IKpdEXMSB3alRUFUJm091J6ZqvGnaiMHBqoqe8CTyy3bSSZg
1wOUWnZJUZjcbjwwSFXgJJlZS68aAI8Xb1MO+YneZNr6qVJn263o0/k1UyMl7Ftj
vV3BxmlAZL3yMZOD/crP6C2J+GL2zKw7bvNmgvhu7vEpcuu3X4gxqoI3ohUsqGB5
wFgDV3jSNZCeHYrTAuO4BHuL/yCFGQNqIL/c0O7HFzCD/8llp1djhC1SkVQmyifA
/Fch0LLltuu90PigYLuYKu0N33gIE+qOkUF3TG6HYrrgULLtBE/xa9x/+HQTNVAA
WME6bLg3thrmEyvUQR6IwbkQQX8j+340mrstU0G+oN2nv/fdEVKjwM1vA1i/jmhc
Zg/WdBFLpZfHvDcF++clqLFMwKZe0BuQGpy3R2zhNv8XsHEvIiXn7hXVFJjJXfZk
YOll0PEaIseNNHG3WfkKbJUX66VNk3GP1i8avYJENXA58vIvRzhQ/m7oVHbumR4p
J8+jSKyTJSpUfjamhwnlukf52tRDpQEttJb6yMaYde/wx9BLMkZG93/wjAQckwVt
X0H3ev1SXSAATa/aJ3G75t/Mu9CeYs7an8EeNn940JAzhB/pDFuGBVIa//7xP48j
NNFXaH77ELVmaDu/wl1RCGKfVdE8p8uVndAi57JKWkp10rDpF5zgYolrxN4s8ksL
HgzCgl12m4U1SXvH0+MDgt2df4EQZKsZqttgtPPN/SE1HSq7Qqtr2mypc8VxtfIF
13XfcfcyQEIQ3dEihN7NthcbbKxFKZyHlpiHGqtPv5N1PHehH9Fgdx0w8xyhU+aH
eLTqvFAfhViPmgVkY2YlQmt15yPeXktFA9PC+z3JtSpupr5BEfKI2s9vqCGZ+lLi
EfRGwnAMHLlQd8cbufDBfOIRUnGzXEnDMyQMM3qttQLyViYjxn0R0sdTmPDjreR/
kf2KEZ8PrDqcAJNdXJeY5gCC9IicXFopM4P23rhMqdCIFUu9ugm9q0PmBlDwTlsu
L6t1C8dX28tbYWeXxR81NAG38Y6eTrP/Wg+kzk3bY1v4ggxWFJAJEZnz1XJ2qThz
jBa7JBVyQV8VUjtGerx/CBXWbK1u+gWNJkb6c7AX2oEXCNQcCd3emAGBkmqd0VEK
4c5HdsjYZ1Lo6x0cf5rcqDtjCnN4jKf4RU3jnvaGa8PvSvm2YWf18N4qa9lcZgML
+Jv/GRa+P3zFemb3tyE2FuC4HkOT1c8wc8NV1cbVp1DoZB+NEL2yGZcgNmHBwMAP
IRVod1QKGafx+uK0kx6I0cIKglNK58hqpvcNuqabJrvbcFL7T8sUEkRYhdp4Oa9v
fhSiOpalMnHpGGLBdlmErFaQuXqzIcrYP0ZknPLN1c4yVw7ktIy49DUFCqtCdnOo
RSS1WmPiUbX+j3H9QG5OETtLJy5OYlm+f23HwzSZi7PianT3E3VWHCB9+7I7pp8+
Z2JEUHxuajtD5dQtCGydLHfIrEsO5vtvm1QyYqH6k5hoXuVFPC1RRbVHKyaoE/2S
FtQAK8/z5Pzadpbvpcv4AydVqYITalunlzw4qh6iCod1Y8kxKsw5pEfygSYQC4gt
SA9uqyQYAZJvb7WLdiD/ybgprUtW4Rfph+1MhoLKpi99hX+/phbhokDlanssO7LW
uK8d8ywXtxkxSJuUkRRNg66RL4RvPU0tzbDxelD+dkVjAjGSvCjDh84NxRroPwCB
iFSC8yhcEA592XvymntNUxn3Hz3aRJOlH23ffWNOsigDwxFSVlBd6n9N//gwL2/f
dsAPvhW2kUhEWWHO10zxdZiOvecNXEhv5NC5xi782dYmosmLY5lC24Qn38ATJ4uy
jd7fdR59be7KMk414bUBTYDY96IcatPuNrWZMspJ1w7xtuZxzYVHsphGFL+S3gzU
6ByIWdj7qyFCZZXuHuro26NtuzVbtzw8lHyWf0ASzCTzjO2pQhbOlksbsOt5Isl/
GcBsoeAdOAoV5HBLn+m5r5gIxBeb9H3bfzVACSascVSBFH7jxseMYcP8IPNCo+QN
o5VXs1BOfDLhxZXBZfaCfMbv7itVvDRPQ9KPVxV/HmHf6CX+QDXuKB3jk/s/CjSO
VUEcD7Uh9KekjjEaDyL/3UWqCOlUnJe6MLlsGZWrUic+65277a5t87HQxuBX7c6N
V5Dk/16gyv9pKjohqFxwibn0xrR51/g4evhpJLn6cEdTbAFgX9IYrPyFESfHnU1/
hODFBC2VKhW8suRXBZbG9yhufvTSjPVF2JnjXHkQ6ujPtSAaDQmqgoYE1R25Le8M
8SUWGDnHOekNZiRlkQqKp0GBuu/qkup0J5W8OOePlaI6PsNfGUIQCuzJpW7jgBSX
3P7slZksgaFoU0/a9zrldBRZNvX4tZeJNW+bz4pHFiBiPTBDJiocCZGy8HivdmDe
w2L2pdWKV5upN08xLaXKe+iI/1wWTnvztCRVHoPVC5ZqI8oU51pg+kPh56s0eMJR
DFozPUOZ+4vHEJC8I4VE8oCineEPwZ17iJMp1NCyq4YJlfrkx3Iwu9HL2qRW/LfM
ivNcZpxC0tqF1mAPns9E6pAvTCDBmTuh7KD77gp8RPymkEQiBQspNh2FGvskcajv
ssOfnYcg/1NsHMtTPJ3/eWRddYyIqqx2tQkx+Klzx7m1wO1xYpdXzoe4wvg5QmTu
SKzRRCn85jqaOtME9c3rMEAd89/l9uz5leazT7mgJkF5l7Tv4IjlF3w7pdWpC4Bl
Ov5ziTtETmcbUBymevFrIzViQU9JJWRb+NCd8cDcXTjFJ7L8ceNIWRkA9o01XSNf
004dIPO9eWn7vp8Th6fCD5mVOvVbQGCsk+C8AnTDvr+eR6wZlo/K5i56J9H6ARU1
zr5hZR1RwmQE3+9QqojGW6INdiz4v4vDc2HMzpV9twuC2VT7JN5tZOazqBELCyWW
8jZZeljYu3berPOahu3jR+lSZ25PphIyF8jEQ/XovvPWrWko+U5w5gkDOrtQZtgE
cSb5THbLydhXFS4JMV+U/fMVAklie5CZmBFnOeihT7Rovy1RUWj2nL6mQwmaoevz
WB40zCNgXyHxLXAKQgVpolHt5RRJGvIervjOyE8cNNzF7ShAG4E9QSFOGhWFh0Cn
GFmKub1h27BH4Qm9JXZgsl1tqFBBVLpLzsz03cp8DSkkiyskGvaPQ2n2IPM2nW5n
ogiczbPtwLKAtOit1eOstUe4W5NRq5fFsRXYofUhoMnEMiv0QHvL2lnYZWfLEQu6
Ao4gVlJ837CuHawmWAeX3kXsg+jU2LarEgF/p9yGWsGV/RNBIlI87glUYpJ8ND8U
8OT3XA+S85M0hIXTy8v/j7peeLi7lfH85UpXi6F9lYcJoVGMEZbBiwmOO983Yh1q
GcmJ3KqW2ZkOQNdKfO9zeJsDqsVTnPmBGg6/zKQaQINum1mFFwhJoJr8ABpfya8N
ulnlub0tgvq3VfYrXxQ7bqUOYM9jDMJ4wPkph882pmtNOB3hBKaypfiogDAsCuzW
gSPt9UBUFYI3tgNnSbz4v+4OZfcgIV/tBTakzblo5CJKtEqGroRNAdptmcceOvZG
zyujAv+dTd2whqlg+HytuBRTfBP26AWWGCiI56kUAAbpQLow7ALAIyOYHi1M65Yu
4D55yNerAm00d9+O8jjD5m64k3/LlhZ/QgQbdi4f8F5BFR5zVrf7ndBW0skrvI0D
EhYdIHIqsYLF6atwJiZJfbjpfFJkWGOVK2qkI37hKlV6m94NkL5YNLdZ/s51ttnq
zLNe+oJWitM+sALvlpPmFV1rJYWu7a5clHhltfGmlrs4OrQK0GM3U2lzfeaN3oKG
3iEhUYVegEsOKa4ery3losEBElU0KFRkoRbGgqxH5PdoBVWTbfDpG/V7DJb/yxoU
8DJw6aFbIjS+1fl9z0n3I8Qx15uufMxQFqEUYJkXrFDv+uxOC2626CkxiOzR+r6r
HqhHfUb8lhtcQSnGpGKZTufYoij/BdscEYR8wMRz6EooWCFYJh45p3h5jp0EPTbu
hnSK3rPcNSLByh29Zc3HWx2e4k6AlMi+lMPLsHJNJDxiDFjahp56TUR2R5+s9LyH
pKp05HBfLAQoxsKnqMujk6KIP7gY+PtZu+heFo9I5X3dHjLYEF71lqsyScLITc0p
GJYa2eonr1pUlTd91/1Sf0STyEB5/EEaHGkaYK4eFGr4oTuCer27OYOS+FAGG+XI
VMFdbncfDLwL100bvBm2EWevtaoO05h+RcFmw175klwpERvXIYDQ0uleOGchB6g0
sUpssdg1Nr27Gxxe1r867AR0SBjsb8XCOXj2VkiIOk66yp9xdnLn4NklVdMilknW
5AJKi46AAv9Bw8AlKI0IxeZA++sPKm7Ijji1Udeu9TD5z8UqQr94QPiqDk7iX6Wj
ypEYODNHkz6mOfvKnOmVdo4XeN9tW7k0+ZKdq+WUY0h3WFN6HkW/nimzPwsURN9R
1N3CYPpCqsyzGK5jPakRBsKQVvtC2N9dJqE9dMY82jfn256OclJ9+ahDa6w5po2P
GHSfKOt4RXw4fsqCxcDb+kq8YQEWwUNaV0dA+xnaRwDgbtXs2um6Tehy9W72pGPG
btoNCVKaX4uHSa2jnb1hjfFzi05yTs5rAD+m3BMwsHi8pwAUSmRe845OHSHxAYi5
ZT31nCx75rAgIDERMU/yiPNdc8JYt7Unet51FBaeiC8bzaTQmc3j9acIl1l4PTeE
b34nOIklmlcJ7Xul+w1xyYv9k+iYklT6+u0aDPQkUAoZmp2E3plGw1nMEmd11cpR
cvvtiK1ERGuKslxWnJVlhr3BhM6aRv7+refHXqb3E0UDa892mJAa+Sncnflbr9Rb
aqq3DRqlx+rriUcZNgR9qMdR5YM+aocXEtSMVrQfwFtP7rM1FYowNTn+f5gscFmW
uPmumb7Zak+xo74tMvs5oqK0yBuZDS8EXwTFXmh2lUN9dod8kqop5Gfwr8Ud5n5J
IG3lcLZX1NtleODlyte0T+6WHWJ1ugO6e2m0edufxATB7YTIF4Ac+fYH78kmQJqv
+EPXkZb/1IgbV2BH//BuYNHGEG8XS92icjD7JsOuY7c2btfv6QRWfpaA2p/5T+GE
cvv6rqLW0n7X2u7GQHEPAOyynQxCofk1U2CedN6zvYiT3qniI5vHNAk1T+0BcTS8
0j6KncNs2BUKTBixvYzx6HV3PE+xZZhem8h4YgEnkqR41o5hqOJMRFYQb3z+g2kG
vJjHCz70Y0IavHz0i8pd0fozArM2cYZ3QGfNHsW4xYTwIEWs7ADxYSwSaxCj+wQ3
A7DS60bBXYLxxwbw+OGzgYfujf44enAxMbyugnSnLHnVTLf/Crj5Fvnh0MJKhs4i
bgpvk22H6iY+wIE1PUAfUTnFJLP7xlr6M84Gn1owkM5Rjxqwu6+/y7qfXVnP97Uo
fWznz92XqCo7G5zz011GmZLynx81wEvtEJn4nwoXJp5LmDTmTaAYVhqRZiOo48IP
Pan91r/pKKXm2f5TskWNy6lraLPqZHoZRrOf64PAltkbqeInu08gD4OuMTEYqn/4
8Y4Lz135V0HWCVIHytsk0x6yTDPG9sHi6cGoXQaadzNY+OeXndxssOv8kqk83zyr
pKEoCmoWMhVLiw8t//OXr/DyU/BWwVJNqynVdMGquxcQ+DnKMi0A2edj0+690ec+
2GyJC4jIdobgLTjO8av95+Qyybq8AKDwOgRNzAhtulX4nrO4RbF36BTx5gVTfoT7
MLaEaEQDs44BgeTr0TKCAoVFfU4FyBrVXirKa4YPwPNMCpzYAM/ztWHqa5+38bwb
O47XDx79GP4VKHlH5PhNMReDZx8a8kGw2FrNJwKM52I775fNHcqnUlh/HIL+W1to
1QAR/jtOYk8aEgbrqS7B6jh45lJBxyF7WwsNdRLHwQGzz+m8fuJVUvL+xH3UE1V8
Ao9NqGS2H+cGlfU8A5gvE6ePf0/VGFn80hpbtMYmpHgacJePCVDgCyfCPq3sf3Ub
9ot0IebtI+DS1ZvG3cOP32MXjjhs4pKl1TOYzi7l5TRPkVdRgxFJAj/x3VW+EeSl
4lk/WCZARRRbTewJ4uJPjwY5QggVvk5R2SDP7YqR0H9X3lq8tVTTnwPJYEQm2RYs
uUMmdmQ23jzqxoN4jtzR0XZL72e7LaOkSkiBqq/iIzjTCqre67S6RmIpc1licq09
zwF0kbjtO/IqXywVtF4QxUBlpfsKvsAAwgWjUG/JwWbkz2mr59335XzBsq9/uB+o
IEHquaP7S/X+2hZhirOgLqWXuC9q1EtsKy+cZpwL3AjxK8VglsKOSAroHeFhZRhr
czTFWcg0CmTzIjL/DoHbojfpz6x7EC5wJC2pnHogOB7Phm+hxsusfH8let5kCIeb
FmsSbcTq2owys/z7bKMd1gYJn5SswnjkBlTeinzeNSJg5vwupER91GEOUIz9DMd9
nyB2ARNRK/fa+tdHRKo+ugk8Wq/91fRIBwJjqbJOkB9kobo2xd8dujw0irBfTWp0
odr4YxGI//rimPOkGvE4Mz3SjBzapsPWZTpSGoPvFcQDyCOU/Ffp1Q5g9qN8Hcv5
LCR8O69cPk3QAom15tokdva3uGTyGLVbCqVwgmix8v4gVSqqJhlO/+RGjrlDudoc
WaIr9QDzu0X3f2+i2KNam4iu0o1RycuHeOqy2rE6c/RoPhT/a8XxUNURoDeHj+pf
y7D/xM1Wmj5lBnyryOIWNBf7giNsncMPL0uGwpBjSOUVXFVwfKtljRoaqZYtYm3u
zcQ4ixerXS5C6Z14jOEanpeIhOYSy5i81qfeSnx2BOd/aap+SDYl9ixtisiOBmRZ
XBe+GKuWg368jS11YMbezKVwxzJTDXrnst4K5hi7EbvixjW5XQni4DapBJgRxjFi
b+TLsSDLbSOtMGgPaF0zuRB2n1bNOcXseABronMy1frlgkJ09CNAIDbRjdZNOMwR
tnCHaPgXitjf8IEkR9onZWE6GtNJtjBSFQg8t8xLnfqQ5rQa+lFPjdcd+iL4rD+z
2aSkmSfZaF9iQm3ZnwO4cteHUcTUCmDeRtkdiwZPGyGZykD8VqGvxFomtVuW17hI
ef6VDESz95fSraeLIgZnr+15y1lo4C3pMohDDdzaA3JPOWLWYJS2x8pXZ2DmC42H
S2CFI8lMfnb9CYFwhnKU9lHR7x7WZ/hmtUqjfg8WWNNSuWWKr2PuqJ3kAi7ne8GZ
yM0xOEk++CZ+3zQhxWV0IlXMTiWA8c2GQQqhBWLyZY3QKF4PJur952wVWVS3F5kz
La5WLteJlaWrJ1w8ydUIg/gaqRNcZ2mn3aQyXdgit9aA7jX1eMEveSbOuK8y+ISE
rlXWpOhd+auqleGXA2k0eDeszIwHGFQ2aSMSDceNqjr2Chj7xguuwn6uKQzhAHiI
+rkL6iyzDyf+bVT68whlavTcCbVfhmaArCZLs+oo/vFZBHDYvKCNugMQEFm1qetf
g4twXSCgnVVXHR2cRQhiokEG02wfNhXCFjhhxclIFnwuY8AqpK7SFYFOrWfCuKK2
xR3ix9On/kF7Ef4WqCcuXyJcyU3169i7Rt0MSbENBGN22ODqr2kaYnP57OTKgP13
fhsF0r6pEyTJyYlVVrdwIgV2fXejy7B77GNAhi2pKOxe0yh/eBT0u03w1soveuUV
4K872IfHuPRrSraOC5EDfjYn+8nhK8z3GAJZkyrhjHZTZamlxAkNN9DbLXBgs6QC
E8ez2kvPwbHk3jsDO1Yj2+6gli0FatwpeMYVAT3wS95c3N49WDj2Zoq49CmaBHu1
Uw10dQfaugrUd+DBcQL/Ew3X00MzSxV/cvSRmy8nAzfwoWmw2JtDDWQMciJ9nviy
bAE3fElJSA5e0XjtdyRlJPrjbJjdBBZ9QwnYMHq6+5QsZBIFVr9o97nu4unPnt2J
hLlaUf9ycEv/b5FKOxtARlLpS+uCepLTcmyWeJ+cg0lQdcw0FECQ9AQuLIdt1AcM
ihxiPg2OeTr4rqXvYJrJQM41IGpUwlVESLpc0zMO58MIANGg+enwhInJzGFLQYBw
uY9mY4fX2HtWXw6cZwuNFTXjxzf5J7WcC84poJxyZPVwwET0hbxsTLly46pDqIry
MKMqh24Z7VaEMm1+avs3BbNpKjLSCWgpGiLw2TBmHtWTchuhDiFC1Ntcrg9otDqD
ZSqxgXgpIGXzrWoH+HckCI/IW8gQug29FD+PhoS5w6aESP9pAOCbMmI6aaJadkRZ
tDBHnizlCgKOzLOSmWJ57Z8iXj5QT0wsMKxGDJ/r+JggSxuRkJVJ/7bGICLVFD0i
ol1O8bQjQgV8kI9EOTIj2pHb+BcFCxT7/IYilYBbPcpKonPeOor7i1N5Y6cnDt0w
++lnDV0apZL07RICgyP+wB8bwbtxsf54AnWbXSiCAD98fgp9ykR77gNBgglH08eH
lye6y6inHqsVDiVSJIpLraukbjpujh6SWcOoT+i4696FWCmiBX9IjA4nsrdfk0GB
41faomGn3M23cj6QBQRMUh2SLbaqKBcQTkPVVknjkddh8VWETVCjo2N5f4AfFj1f
zCqNmBnIS0z6SaLZE0tN9F93ISx9BGRBxcjWK/L8tosYJib8m+bwLsOOjGKQOQd0
G0kQdvld84iEl4rTnr8veEcpMtyHymWsoGWdUo2rmM/wg2Byu2pfmEWvqfczTWmA
McDJA0oKYNmO+khtBcHiOrLYhHBfEkLnND1bEhr4RM+3WHZWFG+C1Cf2bpREeORJ
K7hjNfRNAarYFnH12S5hdI2qvtmSrzr/w4GYt6L3cBTd79B1anD4CV5b0Bt8HxCH
zM97ccHdRsMrVZkMgcZLmnDo2lwTmaYrnslxT99a+kXkeyuiIowq2Jk/hSGCFpuL
+RpZyJRKG8klZzbfMs4IXVTp5xacoeKF2iy2WFmdyIKyrPj3SVbVL4MrtA+IRAU6
+HnR/p8ukdrsHvy2rsNRHqYWhu4PtisJbEY+t9yyW9Y0OQw0UBNsvOhxZ2eogZiu
nW+50mVaEypdQo8GAvDWLnSGJMS2lWCvhDXxOolZoR6wsDtKDZs23yqkuBJKcD7q
85riNeUZ1SX7A7JsCanXeRGYTJti/Vbpvi+mbSY1TQiETRzFoORO7KB8Ljme27nd
vYQIGry9h1dMmr4tVdcEdTOKr+wPf/mL0qEBjUzyToo8SBPDZ9MkZau0+pwyy0Og
3osZvBhin/NJxboMQUX95+zotm8+Fz5xJ/BNsWB9oUYEJG4neDEZsuq1K8YKRoCh
ViyjeAIGvjckXXylHhYZdPhnpA5u+lLNudClJ0g/0qF7Esvp6CBRtIJS+9PSHMqh
bYHJdVZeD227ARdLb2e2jojRBYwjW2ocsZYs1ZMyAk0OfVAqHD2qEYmhvLsTMEj7
bDva/JuYpub/CJUaajV1YCNOFuPy+siODYgSx7060enlYwljN6io+1Aj024Kf8RN
pMNnRehTnNjUUSvWWx/UHyECN73ycRXBXabnxbtmVKgz9uLbDKHEUiGrWdrtYvkq
x5Jm6VulfCYDlSTxvX0tpHwhtzB6N7yGWUBqnA1YazynZuLoX/gGhYHE6OqjeNve
Prz78XfeYfu+t+eCuR/ERCIkMAHimaZM3j6ot4zP4yrmTth8Xm5GUv+WTEidJY3x
0Ui30pPC+L7IC3l/67Pef09gNO4DyDplv8hlC8I643Qtq7yRAOBhZfzP6bpOAEGj
4jc07y5CC2mZGRgreDphHHEem6aZPvvqWzEqom0ntwM3DMaNTJDQ1455aA0zHYFt
JH2Gjws7+PeK9/PjngrGcq1RptVhs3y+t1PkvGilYH2FfUXfxH8cZKkuItIylF5+
fd3V0vwwtcUB9LBsvU1owxKAWWT9nYhRkJoA0p67gq8MB4W4r8kFPfpr/CRW/auU
FfUusP3Bs8gSmV907hXPrVgTwW0GMbR548U4/Nuxk9288DA4vPSAaGxrLFqgqsa8
gMgbyvQt/Vn+TERC0FuJZ4mwyHZiB6lMWPDqQLTsEpsbz7c804M1CAfF5L6BP1RI
I4Mx7F6KljU1hRpTAKd6wuZSr9h93XsO6MCqLemi6kgoRrxdswZWgHRriLFQmx3D
NdYPgGj3GyzowAReJ641OKpPSwbad9ThhRmEphZs29ewFNZvL/UpAtd0Ctac1FG0
PfAXN7k9QJUK/6tOP70uF+26DQjpNigZodhkpyKmlM7w2LNgkqjWL2yOprvhdbjl
vW8urbSnIiFoFZytxnY86Jc93kddcfa4S5l4imSqkXOhvHum+130PewFi8UalKId
6jMK8NaLsMaBUssFy0Fi7Z2eyryGO4mVgi0kjV96nQXBKxiQs7d5wPJk2qQBathF
OFOqzeDfLtnmc+l0O235fD9Abzi1zH/XKhNuqmmoN+5jMHvBfH0pO1qf1iMlUnw9
+b98NwBKCaYs1exOYNiGWHP2SVBqRfUWe9Tt4/LMHw7XfOb0zei47l3BQV3tzAUR
qAg7EvWbRkZ2qbv5GIiBkuO4H0nJDGnavuCoYZO1FN9QYdXq6DHIGPs5Qb9BEcPq
cjh4qvO4IIgOQLACzpDbAQLzbZbJZ+jK/v8UnKvx+alfRlHk2nZA+0LJsy3X+ZPf
uYd0H7+sdFJGBrxfq6+rDAGYcazJpYMxpyIOwwHfITMlM3tNPgm5DXLXFyPIyCL+
hl7JHf0bS1WDkvm6+IL6wHA7abHvZc20NtUKVZOBIbmT8YO0Puuf0kkoegLAOF6z
CcBEA24VTtuynMrqCf3t38uVm44om9uUyTFx/pRQjd8a7i9SP9LSp3OMd/siUZRR
gIU0seniMfMjfQxUtH2psVbWCtnQ4cb4j5+Z0QkLLVqAtzM53qj4ZqaDlUaSQOQY
NND5OmGZWCweDr2J/u0DuuLlIjkq1RwZDh+mlglMPZ0TfCjn6LmsWAzjTlOzbjYj
VKBf2Z1pAxWG0cvTiuzf8g54d8PXq5zqsPNoOpuk9dOt9718RTbB5AcdPUmG2GBb
0XWRMEsGnGu2NF0YF8McRA+iH5u8WWSObKqT+oq4D5pJrWSgZdiszRXo4uir2/f6
pYA4YQ89NjZWZg6HQfs9L/oKo73ZS83BnZIvFqk5FB9irV8d/nUeiyf7EAlKrKxs
852Mk6i1ocXk6IEmrhDB3Mbw4MP9meUV9R9sT7FXCpWz2yDpVqyCuzchqTeqa1ey
3DyAR2YQFng7VIVAsdPwYXYqEHRCtFFeq9x6u7E7Y8NG+LRmWAZeG2LzXQbGCpQZ
trJwcxuqeaw2iMqswFeu0way2SlisXRVIBf9MOP5E34Y5Fksntb9qNrq5ChiSJah
ex0EGc7xIOP/dXXOAcuc76nO7YqyxYwuoA5t5P0VIl5DQ12aZZiePs/6MFwu7HhC
C09Sq0051S6rM7s5fr//wV3kCmqwJ9RmOaBZFSHuTh2aHOeLKemKfcfrutjIwVVn
iI4nrW5xwriAeoKkPNJXvnk0t23dW+q0EFId0P6A92EyFzA0+HkI/rNQqgBGW1We
tlxK0DBe0002eJ2kSkD/nPvRFoI0WsJxiYN78vqn1tyenwE62E2OXryXDxVQTUG3
c6NjYaHnI/w+YhOIT8FybuNFfYmfpgO/wc3sfG441Yt4yqnFZDmbDvCS0u6WM8kQ
rDusInafD5ZExOGE/vDqaGxP7o/VpPXcPty5ITmVXaxSnVA929lQjlIzCA5XGbst
wKRGO0E4yWalCpi35NibZ9Cb5nPwA9Y4uOthXDvQ95BG8e7IJ8YaRHofJiI6LZx7
s4r3e5zlcmQpHi0ECZJtKbaW6Eq4s6YkgnKRq8KRfpHfQIM/koF7rJg2mH5MZ2Pj
WcC9bJ4vdlHqgmoHBJnbZ8Wmqg6Lg6ww2dhNZJ5er9YFuCK9s4aHBQgp2BEyYK8c
HxaLoyrDnDEYuxOw/IZ2ZucovcAiSzBuq13HNYEtY2l83BoFkTxIR2hPpZKRVf50
67kQhHjIXlfMuH4TPvmqmWJ+M8f7qJv6Ybnpk7+lgrwPjuKBKYRmH89RrlhFTGOS
daT1Z6FAPGpnX+ITnFDG7VGC+X1oMGlKwmSPNe0wOZyEoCNV7+xfVYCs2Jlszwpb
MLKU3/bmrzTR0I3UTI0fHRTGq/qnZmgyX03FpWhVNm3sOspMe00xxl22QCAEPkrm
KL/1e+n6b+P+IIrULJO2YWtNMKWnC7lXlna5sR2al+H5SuEVh5/RRmhfAZ7jhzQB
EOGeLGb5FFwsvbDNOY+/ZF6q4BF6upLmRKN97+8msMB9mpiIu7IPth9bmfZjKp72
d2yg6D8joMX1SEfKkMXWzrexylvg4+Y8A5pe7B7HLebKlfGPf2MQQQ77v0i9jDpj
clwzKrYv6w+sl9Thy+HnYCKzbVgcUgiCyUxScnhxKcdMWnSuYKRzwuE64Y5GBtDv
G9MZ5iwD0JNoDZDVr6Xkabn5AjmaQXVlbqCa4tS5K7cm8nRefWJ2ghaDbDU9LEyy
5IeO/4SKtgU9SwkXQhCTp42aFmxSmcTA9OWWgtVE1K5KOmLIgHyGo7202eIPlRQI
hxlVxVtwZFY8rL3V2z+12WKCIzCKtGq3L2hO2v5wZimzxVHrbAiyOA3wst8dKzeR
l7HNgvAN7SIp8IM3d10Kbq6EhAnlei4IaDN+0AVo48fXVvxBmnzAHb5VDkp/3TLd
/Llvefwxg2vNFrMDCp7GNNfsae+OGyDIzwUIRv8rq2NY/EuPFlidERRadz200SVE
gI4iMSDcly9ZyNA84fu/7oagVb/A0qPu+m8bBJR+3okGb5Oc3wWvJzSczDtSw2nL
o8A8aK04vRJ0ZNZPuvCf+uvLmIr/8LTc358s5eFj5qalZRoWUmIBPvj2DwsoBCYW
+8FztG5xCCCAx50bCHWmAalN71RWIydkveFSMLIq5BrqMwRzSS00QWJlN+/d7HJv
YTJH5Fvqq2IZCpsnT6/srlztn5ZO8aTdHLemgvtWyNd6kURyCkhCKSk6AUxRUMsu
Y/7KnmNl4oCb5YTWU2KzHBuyqE9LtluB1n7WmHKm4wnVdPKIPRZhSMbqq2kQuBV3
a8Dcoa3tB31/P4rqYJ4cDE+6HGzlHtvAXgsQ5ulba2vLtJLmkr+wHl5QE62kvVv2
p8ZaHAgD69MkhveElb8d6SAiYlZL1TjsLPIrgoGjZJRYlFb3c7J055FqvF6+Vtd9
UlGXtsCSPlHw5O/146Md2htQsCD+E/UEQqFcnf4oMMNu8435Zbodp5EuVlZidZ+j
0hAap7l+BREU+CAJ5wPCzIGzMkzSM2E74bDRDd5KN+SYDvq96pxn2RaPU5Xgvp3s
C8X0+nOjm7KfpGsk1vCQ2ROjYZ8bINVfsGdFHffFJ+7VrMD0X4uowGtMSh8/txBo
jKRXkDi8LR6b97Cvl+MxGQM7YJ8Mk7RzYid+4kKBE952IUd8ZXEconneh4aHg0QI
wSr/+a+W3CaTMXDtwkWI37ib4Sj/xK/Z6VReRCxInCI3nqRJsptx/L3PPrL1Cb3c
Net2zK+B1U7RL0fmbucuZisumSIaH0Q5fIVbUfZ85n00WkgXYxb7LctAKI9F/igt
+sZHEAvZ5VL80tj1qlW9VdLep5FZ7wMFKFLgv/hyHvXY1bHWvjoLhL/jzTzoLTet
201TmX7SrTTbWg7aTKiJD9QKHGIHM1elt4mbbZIYCGhvzT3ZR9Em4x2ut+4UWwoX
40gCxDGUtgaJbDCeA5Z4U00bWVF4rDUEVxzjvGp+Qp8Dg0UuQvvYbg75lOzIagGJ
w2UeL5pvud2BqAjIxEYh33/NIGUr/NTI7atCrWaKqCz4jQ+jU6ftjEqH+R++FoQM
rQ1gI/wQwQJFC/f+w0vy3HP1tbMAzWNSCUm8sIiHCdfizLe3qrgMq0wxDyz7pPjJ
mo+ZYnyKicifoC8H74sXZ12se0lta0pk6nlXMZVGwFdrZCp7dbRUs+S5IUtK0nvE
BMxuceXnR+Ehf2zOSisvT0bw+PPdzEEwOX3fki7skePKvf8mWSkq6k6d4sWNQHNi
saa2mKiV08lI+jTTD8lQJjuYUqJAnhfHwUEqPgwut92y3gxgcAE50vqUxHU9KGmt
Yw5l7rHtOmr4tAzOA1yb1rlKxuOSVRdDbX162C4yCj2uiu7AOiCPL6an6UVsVtqB
k1IZznZdyBIMcu1V5eFjYQzlb2cV4HKXiBPsohffhEU5zeFUR02+mFbUbaH9LiiY
dQFdtvNtdB/Q0Ue/IFSBnFvMsjkINpX+r+4gp4TZOvJmj/K4ylIVnpHNF91aW9FH
Jg7LGK3keGDeHTvqwN4MdtElpaViOimQjYFodOPx18qPIoAsH6CCVDBFh95CCVTe
l70J+WXU4vfDTk1zdF4WY0KHiortQ6COOnQnJBbunutTwNJjpa1tj2ypI2c4XDrv
Ba7VxXdaFeNkMqCjeTwsQ8HoTxgPyiP65+OclI/jbUDECl8ptaYX2BR88i7blQ1L
NekQaiAh8pX4U5IqDRPyauKbkDGQxC3rADGdaL8A4Ey2lq52PbPt0p8Apj9V0Rp3
v3vDKT4mdJ4XtPjRSDG5Er4Q8iD5oVcNkbAPzPGH9kq0YD+oJ30+uH+24SQtHzYB
gD2PywHGQdUyw4G8uE7noJ+ZCN9hQD1BVzABUhQJclwlNl9kW5i3waZ4N4k9Zp/w
v+BWVpeJH5SWwn9t6Xj7/doGcqN/zUxTnpfpwwph5q9JRRKqFgg/AtyUz6LUYp+I
ohAIqtILBnI3e+56ueaXj7Zbw9YVOjzKf8zM4jompYt/dSrkLovmeLdMxGpOg4lm
CxlpVpDmqlH7tc0EeGvk7q3NDh3x3HHfcG2zoTFO2tmRnRtMLphG8uWk2Q+PXE9H
zFXhh5QG4jnNb6t4GRjZ43NuhRNIbCW8Auo93bMCFG7yEPJjOGEtg16WLGFSLMxy
9J21GShEMR0eYWIgI/w2xLJnEFKW+K0Hv/ZESgqTHtibyKbvAD652LN6eASm3lfu
tekY3KGpO7Y7o0sIJH2bL9/oAL0ocR0YLdebn2R1HGEQ40dxe9NxuiY0CRTdkTXp
f2b+CoeOO2D7URPlESPKhwWASDcw6t6OHWGrySlJ+09D9rM+3vlbbgeSsSfsTuvJ
KTGLo49F0GIHopmHkwbi5N9YzCa7mFGTbs0Q65JKwJlkRzf7tPztRs6OA3oi6G8R
PrN9rzP7ZRy7I0U03uYDc9wOUSsaxXfifXR9Fbwb0Pyiji/Nhlec/sDqNMm/3yag
2G6GIUZKoqweBltX4n8U5ceecuwLPLRuOHIWMYxQt5QTGVcIP2TY4XdHLif3p33o
BIngjZvI2wAts7uRwGy50lImqDrw+ykHd89FzrNm0AjK5XQmueQlIshPdRQqOIIM
ibEvg1U12ptug70kvXitiJvm40OYmkikP0Hu5QO+mDtCFM4pivTf/XrO0NsDYiVK
1wYfu8W8YpzRFm+7iXi1evvhDg4XL931layOpyWjk9njjGphdnxDIR4i4OpCbs4o
slyArg2NFxErkcSyFCre53mQCedtKqPZ2iW5NcjAnuGyOC5XBrvHBKIjy99OHQfY
/lZP0sRpMkoBLzXSAznShT4edpTtmj6xagNSX4g+TCkoxLGxlR3IYLOELwA34nWm
FxhSkKjdJzUL70NOKh0L0SpEocKDagmx8olqXIMTJn9xMHMigdokAdfYfC2Ao33j
PpUvHQyQx/3TO2vB1xBSNv4Gf3/kgtuj0ICpcYZxiiDwS5ei5MH9tQN9wHXUQSsk
5CioMEEwGTLwtCSPIvfRSLXvq9fno+Gkq8l675Vdh0viKys+7uI1+o4NFHtxdBNf
b7m6ui1kcw36mX1aC6WaUXAtl+wW2zTdTw8tJJYC2c5hby4pkITR+Ou0ri58F9gx
32LUkAJNZ9APq3s6kzb33IxzxM2/nxzEJ/WXsqUuqdrtr+h1CzB9SIQCg7mKcqeD
cjUBnslKL77LjGHv2b3dF9HrFzWLqeqauSxMVGBoRRez1UAaPcQriOpwq8SniLBH
QcP9SNheFcMaz5bK70x/sL3HB/ieWzgUcCJtAjJZchPC1W6QG7yo5MfU/+JIKthh
tEpItpypbMik8FpOxlvkmTTqfoNbczBoP55gZocecIukFkz8pTQUicpAbE53eI+K
ZvRqGluGYh27jX7FcM65lMhzcQHfYyCz5xXx0rgG/5he/hL/ehHpZE6qTf5NpqoH
RtfgnjFJWpGdl0GVSiWv1hQemeR0xwgi1hDiVaKVVkVKCf512MX+OiuZ2W5NaSwk
gvUvq14UJBC30pajj1WuO5VqEgYrnvLk9WXjyXL5WY2Jxf8F5W5a1YEPzSPFSDNz
Ww5Be1/KDE7d5B1RIPiUXXvNRaD8FhD5JAYAU3R2NQ9KIGhIEgs4DknKDP50Hswf
uBG0L1yz8NhDSTexZDU9QFF/CYpcc5dmukEOPkCjTVKaEGZXv5TwUyR94hcFRLVI
uzHpb9VZVff729Z3xaW3DrVHsAIwUQc+gzK6jx30AW/pWzDU+4Xx0dFgbUxWJ4nT
3TbaAatS5vH9tPoUeyTrMRKgLSR3pzv1f6yb0qCn4+w07kY0nP6Kkugdx9eIaKa/
MvKKJlKlUM4XATcMQqbfe9YCQ0liuapgI2p7grSTkrnBfbuT5bMSWGI5zPCh8O4o
m/zHDQNCSHfCgISaYGqOI8fkWXY/VRUGoWYu+fV+5B0cM8xW2ltQ5kXEMc3dbQlR
JMtofWnaA1RNG+1wqigCyfGO7trKMJKTGTgCiYtbYnFhKL8JMIqY8WgL49MkL+wV
7w2AF5ltuKAq6S24qc9czJjVNGw4AFH0rlprUlBp6EnsZpMLFhjzmLxzQwVS34m9
TFRcIM1N8NTt+lY5uKfXa6lm1UvMKCscT7AC/Ay35SdLo4S6dUG0zltWpj0kGyOJ
h1o3aREliQ9Kmwh9T5nhBeY7jCcbKofWV5TSx4YtdLwfsMFBzr0YDgfDme3yRUii
Ej9yEy91cBJ9I/oQ59MsXcpVKz1PxGFdOIFjsTGKGF1YcBMOoLKt1eRkyrAXZGyg
oeN/VyqXilB9fH41m2o6D/JM8qwzoaA/DzATTZAzFnXSK/jU9Vo1vfll/fBW/xi/
jAD0Ou3hWolyxk1tMPvupqqxI12Jfujp6INnx2tisONIuUP3Il606v1tYE4ORw6P
q1AAjHhI7nNzduENm16bffH+6oAKFqn6jMkFqarOD8J0z672oEGKELvr0HFprcr+
DNwA9NuxjKaKExgR6uPpozfaRQyepxDaUmHLBd9sBtbjRSTqGB5irGF/8OC6ZcFI
Bi12fse6uFravvVI+rz6pP8tK/7qL1zAFsl13Ytge7Ah2izn649oZNKuMKsOCpVB
uRYYz1f02XX223OuVQE2zrovZB6lGzZns1uNHuT1+KrLyWjm3A98jOKe27DsK3rw
wQPrJbR65O6UsN10SCyI85NJKpusSB8fZZMkrc/SFAPv2VWHqogvY4u2roCNepNg
42w/eDiQEoQHqSHVvNktDJbUBq3bjsyhC/tPCFoeHYorL1YH+6rl+jyzr/gnRiij
0ALAyAh57SOcdoO4F5fYBhqPOQIxM0DOXBvM6oT7ybmUNQhHAl86dOxief+yNCpO
IvBkmcP0unKXG43MLPJoWGCA7i+4k7Y3/H97Rcih/+qYNESMLGWKhKKi0PYkOyaY
NqeHwKQPYC+dYJcoUGsRBnNQQkGCD/OqZ4wn3fcsBLUy1/5GFhqYHBNJZ2NKI2cG
jdZHHHMsN1mQs9NBmZ96IeGwGxio2anVbM53MGVNWXhHnFk3o695gUV4/oQsO4oy
tpU6PkMEIQ5Xl2aPxsynkMYnmUf62iYFQZbfz7XHocxvlH5wbIwuwut7s1qQ5UyG
0o2Ck4+uwsq68I4sYU8sYA8ZCFudPRCT3SR67uyny5Ch4vRlE9MbH+DAoZNVe4VJ
yedu4rSV23KYjyfRdN+hUnn3P00EPeBa9uxBwOd6s0RnF2uZSJliS8ZkEJOy49SF
TIyuRd63tnmneBW0AQgqtEzoH7BTZmfis79pZ8HFc1a1ujcQ0vWsoQOhq/CrdLee
FNehB7fV6/N0ndsWdXg/g6JVolxmwOJQOqErVJEc8+FTAzmWuZis/4Coj9B1Sadf
CvDsXidV7DjmQB59QI8iieKNmg6mUjTdKGC9KhJ0KKG3kc+adBLOboVTvvW6vnfC
hcZbdDUmdqnMNArATiJra0rhbSYLBnCnm6YBQ86M5JtYQsN0Euz9WtII4tJRfuxW
XRtb9h3Qc/Vyz8baCHkeW6usraZbKYHDjKUsB9IBMdI/rvWuLJ41A31LqPI3Af1e
4zvuyZpK88LkXP5Q6PXt53qizL73d+shkSJ0ZBbW/DGn+SGYHBA+gLcDIHgGoIRy
hu6bDLAEcS6l8q6l/Zr1SIUuApUcW8xpVlKv/+a6LUEOsxeieqZZq0iHVwiZ75NL
KJFydgaOqcpS3l8nLPrFnoE/g6FSOdky/KF0tTKiCOKF2rgclWFSrwNZf8mVYAO1
ovD5UNx3b/QLWH4h5h/+az78P2fUzTUQzPA7i+T+Mcbw33igvAUb01TnfG9zOR4W
p+O37Hl3g2AAOHCNK+32n+6dVgWP6UTKCiizWkdfSF3uVtNy54cUCs5FPuQX9x9W
Wh8voQ49PlDoFq7Q1jQz10waajQkejN+GjA7Qkosxj7OLdxmd273fMPdc0uRyuLk
7Qa7pTiyPZ6X9DPyERj1haip0goIXT7JeuKfqiHmguPiQGn7F+E2/Q0+OB3IbW88
GPSLfl/2jI5VZy3TTtXFIz18Eo5mAvAWnlTWhJhUOcCtz+HD6mKX4QpqCtL8OakY
EStPsQBcfzswXAbkPeeqXkg/IR3jnsct+tV/PA7q41UZN51c2jpW9O1LCGsZx6mE
iCDxcxiHms3BUqpgCNw8Z4Gknl4nhg3gFRPPq1xaLswRAk9UjCg/AQoZm39PLAXx
o87mfYhg2Exe7v48DakkUUzqVWiAT0ZVwp9cKaMrXauESv7IPghCyns7f1YpAO1Q
/komdze+Mal61Kz7fsn3OvFNp3bkHJFrCmlt4neK5cyWtxiHCvjPH6wFGrBFDji6
Q0xIKPfrwbaAp9BMoy9Ypb5Dvf+LjaLAMhlqZj2liwv3qBgg4elDYKH55iQptyJM
zUBy5wn2qTVugGJ8uAX+9iidRH0ZAAKXGx0qBfuP/WgdJkfWpnKFXjPnPNt++FBr
N4WgRGnsTs5knTsR6y/bDHwUzN0V3AiMdHjmQ+RhLaCybAvZ7EByX6UeaYXFhAuu
QHmP4yBckc8K4J6TGql2Q8t2mIM40ujxyjShrXz0WYHyyxRWSV+REpwobiJ67SLJ
2cHSNB5bfvjAiTGUq/7n46rtNYR1cZuKn/wGJ7P2Rm5XUyCGiQ3wdFAzeem4TUhy
uLk/menPqkvnS34JFJU36Qy07ycSpVWEVUhjpED9HK599farZxUkyPuUCJXzJ9Pc
YjZicC9NhhPwmlDCnVIkW9beiNtjtHP3FxnthbNvMxbT1gXYH96oRSseV0Rs4Pyg
MWYWZaG6OyNoD5/fA6yw5Ir/uk45csZkOscTdBxEaN47fIxtYIlxImdTD1KYsA4s
PesvPifgn3tIAYntw7sUASKtBrG7K0oNsZntQF/k4zVfhS65DrY29RgK8b8+109V
/THHiNY2kY9hlnLme2Ay6BQQ4zgG2kZRwjqEuntmkYcdz5UZtCc06maVXwkIFiF7
4MLn7xQqbd3M9hlLyuhrLX4cCFDpKt3aiCTdCfOaO1IIxyKNPQhGaXlY99C7DiZv
g421hiR8M1sApUvIFRQXOi054W23kj0FrEZ5PwAL+kH1UzDCNI8DqVA8YyOOL3py
HqfMJHGS8ZvjzwaCN6O1IL8RUCKs7bDZmP7qh0n5Hq1/nnhZoqSxQG0If3Sdr1e0
3QiPOZRtlTR/LAN4xaI9BGRW1ZLF8Z1NQWBknUArRh0XVHkoB78mDGgshyDdjD/4
X+I9F9frzAOxS7Eb9W1t7dlw8r7zuRYBhC+Nzh2hrSm2+UqyyeF+VmM21nCgcZfh
WmWoMOR1IWB6DnDINUHSzppRbpidcySQSZ07+QxdSoIuVkGXDY1x3cSwlj6/hVqg
Ms/hV5LYXu5EMLa1Sx+ty5Xii2GaI7mt6dRQ7Y6F/f8ZjGlVfNxK/CuUaAjflxxJ
UbgA+OMe7t092lL4wSQ/Kq3ppaZUO+NXC25suT5vR6ifoIrya30EysJ8BQmH1bBb
KEd7rKfseaSp3Cnhsre8hsLA8Nn/DuMEGg4YCknD4zgU0nX0+JHFTxshFc7mJqDN
+nuAd0e8GK0TZviZc/toWjwSBQ2qu9N18YUIDDYtuoqwNV5ybDJN7B75HsEE88JT
YGQuWhnFn2KJATRCvfZuvbjOhm+VqnRHpvx/0K/MajQvjA1+OUyEd0/MT70TYlLI
r9gGAdsWAmAc2dDOM+Hp/IUHKjlnY3ShXga3ue+lHB2fxlD6zmfa6tlt8iRUi5wB
jd/rNd9DU6CzTxzPsYb3xiGLq8dKXHqVmouDYbPpNn/32jbpQiRfAfs99JkjsEQa
4StJD0GrCu1rgNrEZqDBWO5jdw1Pc3oTjpeLKYHuy1Ehqic1WPO+k43OO+xy6aGO
Wmi05KfVAmjOgvKje8OMWZFtglHsTyD+DEeUoqHVo2gQFEKTWuF0CY2x4IBDu4Oq
Qxbpn/lbCGMpMhfsjVWrFtDL8M+96nz59s5P+4roY2CWXIITj7SN9/Urpn7MLmg4
zxOl54bP91eMalfVcR/FlQXN1tovSoOp/tcLX9q8grq06858CyDks5Crnw4/XpLx
+Vr51Rp//75reGs7gD+ci3nanGWPu5xe8cEaLxGX0mGcH9oOQR2H9eRD2aXp9b8s
VMUnkyd2J9u3CmMNYD27GplwA19FzMFSPMKdpOIQX75MJV8egaBwvJ4dzJIVjI2a
v27o3sISSR0rliAuasPkkkWnhEwfdxdoYCl/ZozuoqXT1gTZ9f+Ut0al6/LcstL3
ywGJ2XgogpLhjXcrG+Rvg0Y2/wxOkr3PHayzlnFdsDSl4SUB+Anv8XFXL0jIziDJ
yLQyqUJ2uH5iHgTj8JIO0WXKGCkHo8Yx52mb29JoihTj7ShR4eumFoIU+NCWwjdO
+R2Rs1L59qOM/q7UFxZ4nyLLWFkmJGCUVBvE8K71a7l1NOmjFgnMdXGbd64Cvy8f
cETV/b7LrieWrcPYtNqD/yRL36jADF67HlY2viN3tRNLfzXo1UpCwUYsavRjw2QY
lttgHxIuEds1Yk/PhRg4lOy6HnNMqBgb87y4FKJlLP1+sllbFQGS4JbDcvuQ8fub
j1SPJYx8IJ61KTxDn5RIIUj8Z9Qql8WbnXi99DEtWQASgraiuGcwzAQIVVR68SZR
vEO1/oXU/YpIvZo1YSotNxBybMFIStfzd34PjXpyPifUbVE8CA3EplaXfpjnhFhQ
vjv2PFtT97JtpitKm9l3ix66WNunmPk20Sxe3pWThOarEV9+up704jAhyaQ4Xz4n
MrGtUIJeHExgV/gU4JtY0rUYRNJg2CXWghH3Pfg+SfTPl5P/vCj11focKETdQ1HP
DZ+NpoUvnFfGLhdxrE/XHCDc06Tq/fWxY8LaVmsLFZM2bJPk+0Xt+Yptzyo7a+qV
Mqq9pKqLAvqrttcXBQN84InWI8I1actvTJ00WUhpTRH2CMq8vhTCaTELUleEJbqv
le6h5usZjEB2zVSR9HNqn9Sst1CTYA5ircH9iq4NLBTj5lM8fMQOdKERGXEnyY9a
cFxEcy9QUhFoMqHZPIu26iIPeHhTuzPffiFnZR0Nbs9LoQJVf9T3QfhHf4mzCzpB
BuUXe90D9Fw5/uGYYG4hnfdz1F/ouYw7q0Keq1LYyp1vdcZXl2Y8h+ofTLTFB7/C
8iMfZY9Ew+hTpb/LKjCggVR9CUYdEPtegU/BbGTbZbz76qYio9dF68N6d2ovTrif
i/hXHuyNJ8xLV490kDNY4B4kGvDpZHSz0mLP+RsMIhuvhCzmlk4qBxSsTHDp6Vyn
HrVQx96M691jjhwSMEtoV8XX1heYjemme5HMTxNq0exZXWsxTlXczKbY7mTu4Ojb
uNURr0zQ88+6nsr+vqKF/vz9X2TijkrTp+J6CBF6np87K4hdi/qiugpjVMD0zob+
m90ADROmm/wv8P3FSxhYLilAuA5jFsD7NwhDp2K30KJf+glvr/pKN2+VTLZNNX5g
oGFRLWPG5lmCgr282IuerDx+GcjtHrN1inq95j/zqHftUKiHIDFlGCcpQTo1UTui
Qjr284QQLDEsXfGuEKVnLdcbmggCyIB+ZmAWCpD9ShXdLJrspjefHE9Dokj3/Rmt
IkuJr49IEAWujsvlI3KwH3FyXZMPVhirYIzm8BYcp11YdNG69l8sXB44QegEHIdd
u0WzNR60Oc0aVXOUIZbU6Er0WZZtUjgEl8UN3bSK90EmdLYUI9O7ajKH9HoOlcrA
smXpwlN3P0KQoHNjyLdBd3EBfwsWnvSBDCQZajuj1TixhbANKC6afyyhV3Nj+/KS
Jys10QzwNMsACjWk0pBs1o3KnfgO9QdASAyf25ubkM4RjqmLXaOFSJDytqZ3BzI/
/LM/yllhbA4FhpJ3K6bk91IOrsJxCGtjOTJ3GZa6vO0ws4JX7ckoGH57d3IzKEGK
lgJoZ0dwhZCduqA1jYN/TBUXn7y2uktLk5eGe1ZE2VEAWVP5C51lgJSFgT2F+XWG
SLK5DCPl7adVpWSeuHYCicPN1dl6XnptlLoyUqxpgortuaNb4QyDaQ5YS6UgJHeI
kLq1LHXXO0C8a/UmVw25C39He6eoJ4uDIOHVseiZ7CrwdEWmSG42WtwNbTD4wfOj
nfbB/lnV3uEjCsPI2NFSlfnW4LzEgkgxhrNG91ew0ZU1d+9PlEnVYT33yRVCOTeI
FAhwynaqvqnlkfQ1WEIgpimJvmKwi0DKBLsPK1kRYLOu1HapwjyYIqkFXWP079V3
s0zXTOwvexSYrLOSiSavtpiyDqJ0TuxeoSjDFmu4xfA=
`pragma protect end_protected
