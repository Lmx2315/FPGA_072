// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:32:38 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
G2gLO8XcTEXb+pfNL6m/40mP/8mIWvfw3tbpVrYD6l2jHZzTzAKGB/UAs5Km/e4n
vBN0XE5h34BdufpGXHy7iCjXU3ZlGN0hZrsfeih9E0jv6d1WVK01YtP3FlED0/EX
wv4OcN4lHiGedq4sgO6Y+clTEzZVPzk6SeTWsCYO+OY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 104688)
B1CaPK+4X9EfAKEaFEnnG0F1GKvyJ0SgfhgBSGBiyeGQGiLLvafkfIgQQG141TUz
h/QQGUPlxl1ZBypzB/DgzscLz3z7jcl5urYVjsecIQC7V0y741at7jy9zhWcj3mj
OzSkM1+XhYlbUs/18bTs7Vn4ajtz/a1Z/VeeT0l9rJCDNRamboGWOu2zoLCtTZRQ
pnAiV6lRH+v6FwRSK+MC+BmxXmm6XIjGN70JHEEqT4Yvg0/R+ocuroKRsZ5D/TSl
4xr9vPnscnfMgA7QDqY8EcOJJvOcScgs8Dxc0Atj/z+9M+YKC/j4AXIk3lyCbBDd
SU5+xx2+MToK7dhVtiobOiv139nArBJD5FsA0BfHYPQAq2gN47HrgysM0h+VU6IU
s7fpYaw7Ki/Q7AYtFJKL590FBpXNRYzVxuEz/HBMl1YR4Pi+9Oz4EASeYuCAqscc
euwMS7gM7YlvZH7iZ3BUMCb1iP8SzujS40CB9WK8zcD4ueh9Tgm10hdibJgVrPft
IxgvK1jQdHIYAu5YPR7nEXcG1VuxQA8ucOmz96gvp330PPJHi1SYUsl1NwB6RwxT
txCR/yiJumDe+MylCMfIyyZhQ4zBWY5Bo1LLPkpiQWhS6t7Exj1POhALv6p2CblB
6N5Ye22ahsUY1zb9fcxm+OaJGfPHlj7grL1R2hTdabPSiLxYPPpOL0uEER0ntBJc
bkRvBs4E1BCFvkdT96zkER8jw2Wqyqc4XC/9xfJcSUlOR/lyFs83XEbsNHLyLNft
aUHZqKlU/dlxmrtEJx/UadnUQbnHT2+x3txJ5fQlyRs0U1Naut3NcnGo8zPko0fs
rtuzSTmACjGFRKSXN6CWu3SwBrLTRQ5dmXFWMGQv8wABwJRnk/ApaZ5DF7eYO+Kv
CfIViOs5wF5nZ5ftAnGJyErWN8RG/DxjEMTBPx4F3wCoC3bzqfZ7bTD+SFP8hwh5
dkVHtgozTsgrIhxrCuGkCOQnuAQg+8xOu5FZ36We6Q659y3UkxTWSTrSdOrK1xmp
94wWXpraDX+8sviz+VVJl5+OAGYA/jQmzZNVbXTs6xD2MMZN8QGKFqFhfM1RGHEz
FfJoXLx4z8d+oXkR2IVmJTAmWlJYwIDumcP/PgB0CZ8T8E/yt1mp62cBdfx62dqC
4nINfL9TEbR0B0vpEDXiv0CjNJY6xBcFn5gURUgzGK5/x4H1w33GEOl0RCvalMl5
HT01nsCQnvFyAwoB11PcSyGp3dIviodk9ij4HKD1Gh3I9wrNBOPMYhv5u5+21ptk
1rYwkDALoiQ/G4DmgzjXTuU8xBt1b1Pd1/uv34bo7QGkWLvcuopyr9deHwCewLD4
6Kiz/DVm0BtU2NQCg/G/ERvN5WHQLOGBHOvNfSiB8QGwlLMXu3rhjWheTEGq3IL7
PptNPe082MQj/Ge6ZW7wvf6HhEexo+Fchuhv14tgkbQFkKu/3wT+7MDAwGj/kjbX
cZNVFyULvmbuCHj/f86XP7RXK4owhOG12461Cvlxy+KXATzzGa9YtsApFdVouT1O
tvkX6lZ4DSSq2+Ruo1BhnW+G7nJ8Ms+ZRjxmhWkQeHe+nhnup72cBcFU7REJ75LX
gKsSK+yPjKpyMZpWg/c13XHWv7KnBJcaGUeLiGlXW3kF9rydkGRTeylfSn4o4vw4
logIgovw6tnP8D0+ezmxIICb2hXCmma7av5Unj8mG9H3goH75GpIKnTq5rgxZmky
AbGM1maNACogkGQzEMkL5YJqTnLRYq75ZokeXNjhb8znMXPhNeG4NNFR0MopMhwd
sd/H5pUhtaEey79ahHJdgxMA9bQYbAgMSjkyhZYjTRjwvSte24I91iO0bva61fSG
8r9Wt6yOdQxCC2rHkYqu1Gv0MTazfnTuFurwuLwLGQPaMbY0PwoaJtTP/1QWdISz
RF2NpEjLJb4ePC8I9Czv0kDtrKAaAbqj+DNrujhMmeFUebiqMKSrssLkBGDd/0Lq
xPUoRWkR1NLeISzzsq4EyTdn4ESrPF3KZdpmAWjeXYYtziqN6SWv0HBmfjTHIIwg
4XRaFb/JY40oUlcOQrt5LOtUK3UhAEvc+B8a6NLbr9OTi9dttLenco9DM17/4mKc
cQy4OfQWVbigF5wnMMc837/6G3cHdW4itlAr6EhG9KtEDgS7Uxw4gT4W+OHf+uXf
2QZJG0llIZpewzTHxOo8PyRmgECF0lpHryBPcEAw+OYNs2kUYH4afQXUzL4a6g3i
RKdYSTOnK+IdFL0j+bFJiSXy8nDpIVbkyjhXoJ8RZeErTBR5W4NOnZufz0A0Begq
BecVe0k1ZDA3svwmvBNL5Pk+tVi4powVeL+7mInOAsnpchp9x7nxQrt2RYsHXXdp
QlLEGs/BkA3k8wjGsFNY+3hPWuQs1WHZDYEbkAtGZeEgVfJ+JmnPn1hByqtRA0tt
G1qIj2S0MyP6J2AGk/XnZDbE/CTsKGSJyvyIacydYsx/XDeWWz3hJJoMXwME86ZS
GaBqq/vk6gVSwYWhUEOX5IToYZESsDP4lU/KXeCXT+4SDX06J60zkFJA23iaMY2c
0Xtojd4YMj/omZ96gZP+EupoNFl3aZgVEywY6Q7OO+21fE79/VkSbpl+qVdyaLi9
sonCPlLKohp6zODiHVUVx2lbEGPBYdUarJS5PlMkjCmTnwd1NLzf0uTmYQ0oSW7A
sR9ZCFUUcfNkp1KELPlyVx41dMoauYWO0d71FqC43CmS4v1RF+s0ATuXuZm5JkKw
q58fHU9zzwazLYAxo2WxxxaiaT4zrNW+MhQN1Hkjf7TK7ZTKvVaLBFc8WF91WJZN
Kw5ntHxHU/gDBS6qdxJLyy5wlMxK0eTo3MJiim75muhNIavFGfd7C0ps3oaQEKGy
QjRJQW/VfIiDz7Od2Yj5KkJPRks2jJJRqxCMwO4A/5v/BBlluYdbikxg4gZDz2aB
SmvGvPP/HSCVVu2P7mXC/wXTFKtQU//XBAEX0xl2hqQ5HUqedFiKsK1F6oilgFe2
voTzq0f2Lscg++9EB2xl0hhDK8r8jVE6ASdRQrlfuyajzoKJACl/eNXhkwUYa/PK
dHVnzlM097p6iq6N/vNYqKrTnthZYPCl+q8RXr27TjUwjkT8B+OQrC6NV4x4wK/T
5UuNPMUWg7uZ/q6saivPsqy9sGi16X8h6tqVQM32QY6TlatICZKxPoQZHmsCAIVM
/EvYMt8srLBTmtCNOHOMM1zAFPkEEdOLg9ZvSjCV9eqUdia/MlzJPjVUG4E67y6Q
v+xR/iRu5x9iejgLukffjbmH7jW1LEufj1Ni4HpEimMRV8imGvVvd3j8ISBoGrZX
zmvxys8AgEZ1wCqByHbpAJu/nNnk34KJ6FUq5JGEmbLqlsLYS88+TCnmmDCPUzyF
brE2Q2gdz7SQmu43bIqeZ7VetV4zgYps+V2rg3pSp5pKS6uHvHRd6+eAejdfOI8e
Mllb2uY5RH3o3q/m9wj2/c2p0eBayODwf5GVl9uDIeQXAlPNBHL7vlw7nzPRo0T0
CHSSGD7zr0wFU31Ub2Gx5mC1yCAcdeE0c+fElwh9r6MlTJ/mbnEY0KHB4jmb12iY
CA77Ti4K9x3VTc/ENVCroHSjWGaSJgLoMke70mHdMck60vGI2rX66EJL1TZCUxO+
VSt0wCZ0ErIatcVaF8e4eMR6n76qUylhJJW7sCqUfSpYT4X17xNqYXWKPphgs97p
y9zMRaaBqe43Dh/kdNcLHw9lEVCrfDXKazGRpOCIcMGjbJoIA52wmgGFKpOl6frP
WY5zRA/Wr4s4aAuy7UTPhN161JnejXYIQYv0tnVW1oyOdWzFsmqbyVvzmDWYAAwf
AHuZqkm3N35cJoGNFDzOGtrG94jYFhEzMz3ncRsPFw4njfidmEPshkwlfxa85cw8
fpxjlzJakJpgtqU50NaRLFYbT+MOi14ORQSKd7DnpRubwlzSlv0DGnRXiZ4P7Wuh
6i+5xKAYHsLfSIHOiViYHLmk8Y84qe0cLmB8x4CFS5Q9EMK5dWGksSxEI5SC/hsr
COgnC+kw5jHltQ2DH6ZFK6OVVi8qlAt6cIoO23O/g/tjdE8ckh/mCef9jZ7DglI6
QAotAFiIw+4dHxh3p4kiJDeUnCj7vgS7nNbFMQRpzqvjQC89Vo2MqcXH5pPJb9mC
cg9Z7+6oiUN/uXZA4RaeWuJrsz8mna+UmL0Gd+wlLfsswKJgmI6Z84iejMsaDl8e
/F/CvwYpYJ3UTW1CGVIZuM1fCoomzOJlG5WRgAuPOfA5uGibzIskWmoukzUL6Jv3
bBPrNB8bVMRSBmAZdx4y6393E0E0opxJMAiDEsQbRnKnja27omeNe9CAxZEGM9lX
WFhng9nKS89VtSv5yNSVL1C+rGa/fWUGWh14cIWllzglr64OCfhm1yfiyWg/y6D4
4D3DjrK8nQgGUBO55fCKsJcCIasEO+PYEXO9iFUOovF7uBaU1wC4p2u12tCOt6wg
/ctl2w71mwJDBo4tMlfznpLj4LQlXe6B4DTcjdSb1vqZAB0MQqACqxKu6r1IB+Or
sTGcMQb5Tu7bCyjmmlbLavsILNek7IZndH5JUUO1o2WdtmuGjPZvZTxSMbEHLMDn
pr2AaHBdT6Knmn+0qJmp1T4CDq9UmCqp9ZyKSc3XQwT97iKmfu9fMmBFE4zLTCsm
CJ49+PaxEvLbIDTEo3vPhLQZyKhaXt3xC8bPT640w7sy+7Oyi2RDPJOojCcG8dFj
J9081QsVghW0eFnssNjYlm/EMU/tHKgwN5j5xlWe9kjlmu05qE+Qk2HVlWWv2ipd
lHblcCwlkLYCg9V/FNOIFBfQDpfvSXLBOP1da09NHY/dAY9VU/z/rGvGzRj6MKRS
kcuMwvrhmAAx2V612kR/QS7ZiCXh84/sbQ6DQZ2NKq+5a0oWFGcOYG8rJHwG6W22
Of87aXp9ZtHX1PjW2fEe7K2mHp35ZXsVD6bW5Vza4iI0SwATLKKAqkiAhcv6qGYZ
eb+gVZHBp21ZjPcsVHF7U9ELRG5qZYhPdf4jqkOHLwrkaYs7Ot/c4jV02PFyZmgy
vp1aZUt1SaafKo0xBQuVq5Wi5GXPNVn+CqtMrfKlk6zMbeP3Vnl7R8KJRMcJi4U8
YWODcdG5tlqetj7U8U9GwxA3UOseuP8y2ZgXlr3esHVgkq9VWUfJzBKed7aEgouo
3SUcbibDL/w/s6ZNIxihvqNM0mj1tmBic06M4VU95cNLDiWl8pPnzVQOmkSZ3c9C
+iHR2GHVrvnSWDvg+rUoAme1fSlOc7rteG7MPUm+coxLAXVt017vKIXf9W/dEJY+
OBU2+TufhTjTm8HJFIMDUlMP+GDcbzKEWiOAWnSry021jpLJO9NVQB7kldE8ZuJR
uNW0Ew8187LSUYnyT580ffaUVPTjmpOrjDs1sE8CheRIBeKC3R5qRsmR7DVlBOZl
PxCvzdxjA0y27Jch0NOrZbY+rxFZofLzp49+3u5qC8Sjs4enT7y10D3nYlGAWhds
z20Fyc4MkYx03DAJ60b8pIQmWhnqBvDlz9joqB9V7c+xxTX6bKKcS7CiBP55gsdR
EpwgLASgSiIxU94b95vM445hUbc6cKC1pkdLbvngHOMkJSJ2MwQIze/v4f30f+D9
dEV08qwJR5V0vekHsb1/dxu+UTC5AFwVUcdMmetqAp12yRwX+IUtR6ZU+uZJ84AX
JNSK2Fn7JgO9g2gbrOjKuR64fCkteaY0thI7W6Iz7eZm0MRUSXcBfmqJiZ4+hjWz
Fa27g46LkjdGKYcdB4ZQmuGbz5Kcx56ZEpB6pkvZx/4gW0EXZmsHG5BScl8CbUMk
X5oFh2nf0BuDmXa8oL2VdQfMeHOmGVsme77pks0LE46rnHkgnU5BophdSP+tygFK
88MUaEjozHI/O3WB/e581a+nzd7o8kJ8Xk43BOkNB5l8vYPOnTA2hokTvJigRUu5
wjee3nG553Ath6FG0r2Ef5iCi+fsk+DRX+uWyWkMCd5xUeIPGTt4x4+QridrAj+p
sCaFeL4Z0HRQS1KxGo58ZG5mUGS3OhwoWO8xhqmS04Na6SJioAPxRTQc50xWtumI
jkgugnBeDQ8fA3FdIRJJ1U5+Fq36P5OYVmvnFoGAV+gce7DxiEenRdpXaVwV9Yye
PFfgHpnCCPrfIxko8spu2LPlr09IHlphN8G387SAc9hl7ZfOAkeCrHiwFIEOUouL
tcokUv1FN9J1pxw+uEFtSTWgdHYvPsGb40GB2XUagigxI17o9VwMnItFdUBoS/Q3
4y0/Ftxo3qPz1OH2D+BTw+cHHzjLfONVRft6Hbg3BdcjnbSkRbgyrdcSf7oCxPFc
nKpldmCqB/+b72SYkXCMm5Fuar5m+H8mqKgwX6wysx+8NCBgV1OV0NBaX8XJYdww
IidUSfBhX3L8gUTyP4SkO0BUHZaxYOvvzCtG1KLZS0fegV0y/QlLbpGljL9V3wsD
YX0FA7xcafeU7N6aKeQfeKMqUkjIyUXKyoqdgNRt6frtp1tbsyAUY/Puwat+6VWH
UsghmnITm7mBrOTL8QgpWZJ7C/JtOIbSH0odgTOBmlYIA9XPcjNkHOhbDQW/pFST
prbRxgvHoVnWIJjYV9tAXvz06EMcpoD4AINO5urbrLaaA5KFWuZBZHV0DJZB4asx
KjnmfEqqltWS/ktR1jNpnifucjQQHKJ6qF0/LTGHCaa2rIGqWbvXujm6WjJE86D4
PkzG8cGmJNC3yalGCvnlWsJbMuudI+EL+cQ4IxRfd+6El47Jelpk7NSdbrfZV1l+
ZWR1Pm/lADDPLfo2Z0ORBiSzt1BL38TMDVptZwhh7cs/C+cdWoyjM1ySyLC6jOQq
LJu0T2rR30GDySBthGG4ByZQWCtcHfWzpyyknIU8FbDe34EG/8mjD5s/EMtDWuyf
5foYfjfIQVBjHpcmkM/z6YLUgXNnkBJ7ZrcEnYZHRJTLb+trr3XEF5vye8wYp4wt
6pV3Zqxizvzgf3BiQ0KniQKE/O0Kt0d/6y4yh7cHM13k9mX7JgeU61oxSLOOykuI
iI9lFaq0A4O6LD1RUIYq3okAlpUgZfO4WV2uyR6F98/+12V6Rz8WSTehq7Vbgk7R
QkutVn1hI2+NzltS4rjTDYWP2YSryLBQY/dCCybi7TLadzjXxMX/ob3GUyBnnXSW
kGJvz4mdJOvvWbg4FnyG0fdcsLS3WS36jQuqdRTGps0NqKo6G7PK7y45v7lV7BoA
0ITL9fby+z/spnRU+6hUl93uZLKDBB+2eZ3WhNXZYrMDF8SWlmjaD3o9ek0//hGb
VESJV+SuIgieiLB+Uex8K/J2sHYjttLL41J10Zbe4HEFEnA2MSyqRc4hJsB0G4hb
8CztFYzM86NQ4wuv3maanUbuQZ0/u48j5fgJ88AvzN1y/Yelh89V7lIAd9LpI1Cj
iSPfq1ItM55lLg/gzsdEOGq5Gd5pdz8OREcrOKGwpEsRH+Z4KNtzKtkkIGIfwn1z
zsLoc5DLzpsV9VJBBjjg4lMcaGZkbFoOrK6mzTRcFo24xgAnYK3uBbbKe9VkGH6C
O83/OYRM9w4igZYvTtICX1rZ8LyUaQ5h7HWH5y6TVy4WP0mNnjf3Jbz+xP0nET/E
fLs3jslBDx1AORXL0NnHWlYLSvEJ2Uj7jHpqnABb6rzslW1KzcW+PdOvG2gZ8Y4s
jMhb00OjQ0idqi72LXGa6NAjakjwj+/GThpsm2zRw2sf6UL3JhhkTxlD0lZ1a05T
oNBJz2+7EjycB4rNvBpfJIVgacbWNwpsfouQ72igdKhApRvXgp/RRrmz/NEUIxJu
rJSCmgAXFyYASGKBHTQkDrXZ0m4dF4ocjhzZP9JLQzbdNAceVd26FL0QOv85U7Gt
1Gwh5oEcy61kGIpq36+7GwRvStFTzMlA/ulrzsGDMFX/Gz9KSQB92sDxt/6EAcRU
rTbdQe4muSEbMXuxk25EcDEln1zTCU4A5dK1aqF4As7PpUXfNSa5dlZyWu/ZRdbs
X0ktrjEPIDMOHt9ChXmrla4j5siAcbq9UYyTStaPgNW5JAGYCr52i/iQNEVsDIC4
8tnwGDlt9QXn85aOcbydInmVhNWZBUWrgiZ/YZrtRnyGFpwguk3Bz5EGJTDi7cF+
AQOzRmxxh5igzZf0T3+VepXIVOOOy2bpId6+HLa+15Jp4a8xCj5G/CqvSnQ9G9cf
dzGJ402SXfyAcy7TA79Qjjx5F+2QkWNcJgieYMIBTuiecXXNf4ZXzRdo4JZByzdf
/N5nkpLRyAM1d1LGzTkxM+IYYcjU4IiAwRTdMxudNdYhCi+bs/gujJ2SQFck0yAs
2mDFLEbhaJ7H4KRCorq41GLwG4diIggWg5p+KYGrMygx8cG7Tv0QdzG3BOdbHamx
odPeQWBoGQqb1rbM1lYA8PpT3Juo7uEQ390Y3IsPJkEvonXzXc+wo+65Twwrw1Ps
JErq9FO4xDBdLhR53YdEtdImQuQ1uCWYrGfxIBKyTmRO2jFpxn+WZP8U6C3s+NRj
8U1kFJjN2V2FHhrTNgNTSlE9/4B5eKVjOsdZ7P8KIg5OVdZBmjdLhnOcgTdzJ1jh
YmxuxKFcjOTOOQT0L4BE5Wxm6dVZbqzxL0VZM0mmcOAq6n6C5gMvzf0dl+9Fnkp3
BgxRz2yGjcGP0BneGifMmlkg3PG7ioN6nn9HpilS1XvrpzlC6raGYhly0KqE7e3b
bXEdaNckLqHahKH3PgGEXBKW0DtJtydEdxFv6A9oeSGMdK8BcpMAvKpJSBkvFUPw
FSxxwtIgZuPwXZnk/NeJgiMJeDCylHp4DawP2CH8ovgjoA2k0pHLnDOLjmrtkA5s
8nyGJvPoGdnBuF2DSTCXTV1GbsdURqjvAs5YsBdwscR1RJJXiCoO1gTsohNc9Ao+
74AkINT/gmTTJOY4YYbMeGfJWZi1gZuHebpTYXvjOvbBlMCysH3WxtZduyYqpfcS
muqrEqnLrHr5GZ/wgdVLNhlcPCxD5Zra0pAfBfungmOdIoUNd+XqqXzwm8dp8W2t
iPFBqvNXloo/PenSIpGzszPX+uKc65aG/1kfLp8OCpOlGB++bALeitNEFyez3mrn
W8ZCzlzrH90gljA3jzuJc8u9g8WXVQ5UhIu51XKejCFeprIJQy2l0LMUhG5RuHrq
w4SieAU7bb4xXqKN1XJv5jRJnHLm5WSba00FDcEvL/rS4nZia7Bi/KhUbRHq4K4J
/Y2ZuCvn2oWFlRXcbXutDs9QC7B0yBPV9r0D//q9b282QsaMcmM0toezwXG/DEhg
b+yeUK1yilhyfS5A+gBf7tkgk/1lewgyYOIKlxPGVnnlf7NL3Tr+yPVRNi/EQwuK
PPOV7y5+woAtYIbSH1QJSu7w3j78rLaODo+VLqszfeO7pf77jf5fn3+ZGxaGoC4/
KNhpmaN5CNWGxVmHvkfEBNZgWDF2Gl67USmZYNjO+6ECVexUAg95sPnJa8421u7O
2r04RZyUFjRT3LlvFMu3ileugTe+lP4Uo7pRuHa8Vu531B/WeNNBSREzaG1WApmF
21b0eiV2BR6BZLDxpsy/EmJlZHxpNA0aen9NysCg4vJn9GwOpU6As2e5VBBum2vL
1oL9NSw7LEsnCZPDpVgkJkv/PnaKGHD+bMU8kzc9ctM37Z20e3HDUJVv18WGWWwe
mEmkvhKJohrUN5Q1NUOyZiVm6vEf7T3eEmQVgHKCdvDl0PiSiNQfWIZSs6pUdq3e
ONAzMwN7xzDMyUZK0gDEvRLlYxWJ1lh1pgq63IMhTmMUYvsZeiOHYl4JdeZcKSd9
/eo4IZwqgDjJulJKlp4Jc+mXGe/oAtyXv2IV9ydwDDKHauYkhkAtT/hKxV90/SZB
OJ5/J41YYyy6JDR0W59PS5X9jHpqG2ejNpUh4aQXKHP7O9uNq77vXDzJt0ELtjHk
X8gh0c5v1a3bZzwL5LhJO8bPmA/ts+uaosBLpcfEPrFvlN3Bk/YFRujZo1CdYqQu
ug3WS1plclZCyVUVxyJylMaXTfInG/KFn264YR13YkU07CZGLzD0ywkk+IsPs7zZ
wUrMzBiI7sH8/LAGlaE8U16IfeGm1DcM+E5x8iO/DBO3Jwn0etqPo5IkUMR+8dTr
eeqbuNGCqgnT8cGG7P7ixBJyoh8EUG91ZpRsLAH8rJzCrurSKqoWrmOBVST8xFkc
jonpvC4C6eD/l7ClKiH7pG+PKzTvdbjPCtNpLiwAFfYZA8rdVsEafZm7k+9fZG7Z
1Lpte2EfML+tcEYJ8MaTtnWXXF4Z0Lz9GuCdxphdx+kjvLpzBKr3kaPOqBPDaDa0
iqn302eTNJnCl5rzmWWnV4QPy2fiiBJGSxo0QTTdlI9804PnT6ouD5HC9cMhS4C8
690sZIpNmtlGeBzQiWEbqsCAeqFfb1Uc/R5PwzQis6i22Z0ty2BHYdR/UFnEqahN
9kQWq6EKz4noLldyW4zx3BvC8ODso7jwIQuCzXMKZ3R2MSfNKRlRy7PfdfXRdFOU
crifo2KG5YfBVe2vY9VmiOnNapWdIv7JJhkkKFyWGGY6mpGctbSBHLdf1ilv43Qc
G8tML1ChdR3Gnqkl1T/jmWl7rIo0maFHAxhQhjfZchlMYWo5zsBw4Bm9ITqYR9XN
EaVSZeHMwFruRWhz5rDrkSLeYd42E9f5LFKtOXPW9k6AtFOb76wwfJpxxlP56IbV
bI+jBBUTdoTgYY4gk/oMdpCmYCpCpVAMCFrSD9SWPOvgoHOIY6evqh8TPAJVLy3o
i0DffIZGyU4a6pHIORFbrEsnK5G8d2oKJ/XggAoCYpRBNBvMHdL94KwXDDYKwc0Q
UFn+Fp8mFK3GIWnBJN3uGZ1J+Q/VJxymBcUb1ZoGkTAs/PyTiqeJktRUXCZn8Fiz
BIQd/QiPOvWfMuzBzWyWqOhMLAQnMTBEKmQ6oOQoXj5Oo6zoaxg/pMZMkNlIjQ4M
OduNuBZFPbTuKxB6YpCP1ScvjHf/7FtHz4kUyLCTrzt0A/kbm7PQZ2GLEwRdZ3uY
EemBNoYHA5v4wmFrmVUSAukHYKF+r212MYfz58BH0QBbpjOCIh/dAgno0cWgtCz+
0SOzKZ6W6tGjEj2fhNO8K41xbxvOYS89XxMVO1NORwqPEyCX96eUkyAa5F3nJS9o
SFgayFI5dxIO6VzeNfAJhXhxe8c34m4jmNbVEt5fkigENz6W6c7XTbpnZSfbTaqA
WdtpkgIY4of9YZ0H4X5/XF4pl/0GWYAs1JdkRFjBwaQ9KNpM0KpI7Lb+ycTldXiM
rv8RqpHTLvvGAzoD6tj/+NgdgI2CZ4OfKQ3NDJF1/k+QGUtJKyCbH/Mogv3S3k0t
u04Yvj1Os3dfxUR9xCTkQnVNtEumUGQ25r4X9IpBpBKuhq1Y5SUIvwUVCW69lsH6
Hyt1zqHJymntc8uMhoRssndGT4LINmJZEtfmJV9AG2oP1avtgVNMlyOarFLBTLq5
hsAZPY/MfmN7ISkJL/PJYSBsW09sGYHHiruGeEKq43e+jUFwAEJigihSRG2rBJ9f
RW1ENDYOEqAn0oLFk4JMBuEYSpLqdoC8cD1B7K8FAuCaLRCpezX/JuDCOyDtlMx7
bTnKfl0dScZ7qZZYTocczy3OWRezwysHQZDy2BlaEw8Lm1bgkgp+eKCeHRzKdIqb
Mpv/8yqEeln27BQSpWXLrfAJKxwZ1JNVpEgAqrJ7blT+lRaxV1RzOM7rBlVV/cdQ
J0/KFo3RcFIcXmmRDWfUQxyrXzQTnTpfPsfJPvtr6R5t3l7zUBPsVwL0viMa41b6
4fTtOX6o8DX9RUlDDllvrxWmaDzWpvIqLBgQBOY3l631jUNa+34UgMdtJ5APgiP8
nl+9RWTgF+L6QcY9vSe+gYUpQqkBOxuEnjb5ou/lLt6EFqVWGLif9tFg7RPkurS7
fFWvNGWXyZUk+9Vnek3laXSMgtrg8KhzrVx5AJ741/wFeDduvEquK8RlmVSC7n1u
3vMnwEUZlJrXl6k9mfyIWeWVfetx31YMPlWBQGV28pFULY+4c7EfYowvYk8Bm2Z2
WxUEe2bRrHH/puqI5lY8GM0Nsc0yc1aOWmkR7sG7fJkLUVR9tdQdPgj382YFqv7W
EPA2k384qVIwXTBsPMI4BfAOy47s9+7TLJm6wBiPJXqtlrlohnuhIOzEWIm0HE3s
IRiGWdK8zwL1xcAPqMIiutefKDtVvnT6xD6ji6flKiivJGPN6ITTzze2yjSPxkIu
IyQUgZW2XURi433wDSbVp1klDpNet/s7iWqdBbh3SBN0mnHg4hdkw23BC50Px+5D
6icL37B9a7dx2e9Ks/vvGt5Alfx7gfUOr7ZqJo0/VZFvFMIXEeNA+2BAKqhoa8ZD
1J5vJy+E+t7BtB1IiUU6xzpMO//WBnzkpeYibOp1TUsVM+fFOvhnAYJT/dYKCwFy
O6peN2Cnzr/APaMxKu57P1Fqgt+qZ5bmsJu9KwwvX36zEQ5B1ofz3URlj3u3qf12
ErkLdLUV+5TvmmSc5a2rlQLKlP0OFXuZcHF0Byr8VXkiBK8tmctMX2+phIWfiM6y
gO0x3c/QQ8eMvZrNs11Zw9kFS8onlPsrR1g+/c/mgCptgyEqKj8XZoXHiaY+xNLW
UtXWqy3tK0nKP0vhO4Ha9YnxY3A4MJ/EGcDVFwVDwA/FGhxB1QUiJD52a58TNMRT
B/s2KShHXU5sKMNYiT6OVVBsi+XKwJEWht7sVgmY+miun6VfkeWz0OVNZYKcFeT+
XJx0In0EXbL17DC1rThsd9g970257MEFJZWQ07GeOIG+fQfCJwDR8j+lWOtX786M
ELo9b9QIR2QXDdMF6rHpXOPUnibVr655mO48MjB61QclFvzY5klzyZVn9z9MY4RG
0pXOA9rauMAzx75RQXgc/9rz6UdPmYCSzvOY/WUAI62ZM2kwhmTUo4SyP+ZeRLh9
vpe5anFQ0AIpgNWSp2kBRoWNcDxmaD4klj05fSwScvv24kFqrsXfvCcNZ6rStSRs
j6VZCrHe3r1qRqAkR7d+w+vW91/zY7yIJ8KoxUtV2TOZQG54o97uDpkLaSlBTbBz
StlYBZZNQGgJO6h1LMOsynzcAw7AZG0Av4zy8+HKfo4vBkWSetnqA9qOso03HSlm
gmq+PrLlef/PXXUygORx8wP7NqLRQ5iqQqJOMIaQHs8gg+0DykcJR7a/si/U9BjU
B5n7T0gxlAqIhcVPu2x7f6BCM4sGcOJhg/UYftbolebjxrOhcCYjfos6iy1xMfG4
i0U9g5TDs8Q6879wDsMMcCRlAePLtHljhBj2zV83r97/sRejaekcvKH/5B17TZsF
mqg725939JCdn6mcqExFEdFGQIEzqoedDuJFi5nHvEfmv4+gn91ywlV2AXst4Hhq
bYSCklDsd2sK+BtG57BhceAvzgDLn9txLRAWpnLFVbNhssHQ0vvZI60hidDAmbWp
10SZDwkcl1NQ+5h9okYVzat1Z4MUBIUjins4aAhurTAKJftSFHzL3+l49rOrbcb6
CEXnImnSFBPjwfdsH1wCq10jmTuS+M9gLl1rJ+rZmdgdsBCV9b+QawxF2hFvEPlQ
7arOISlr18RTsJuL2A/zCSiylGU0gzM578xkcQC5jJ2VtJZTT7e/fBLgzmdlfaRQ
jjeRsVpCdjZVg/JTxLSfv72awk16Udm+jKTWyVlhQuMzrg4L7j1YQiaV6iuyJJ8n
klxvUVhKw0PGxEzT1sVKrk3I+cwCADDQZu4fG+iR6ovzQK8hAr32CJw7BtpckEo2
sSePn6Nj0JllYQEOsXgLnjtcT/XS5ZzAM3elUtEIpEofmQGXV6vK6asXdY3GtpLq
NO9TPsYusL0NVAP1NNVvIdt3xuRmcLDYEmKvupqyMy+95RxeglIKTKnV3eS+Gk99
rE80TFfO73VK4StoPb77WQmv+/UAm62xVnIABslAaTCcn3SkpXsUs1fue9uwCZN/
4qpsp5zoycOuXX1p+OJ5MfslroxfXk+gNVQ+c2wdYBfD915IPQlZn1mK9o3sNo9+
39xzP5hpNKiAgZ1yBthlliGqSUwWNvGv/skDZ+utp0Lrv9EFJwf3xCEu1z5soqEJ
QqdwvXwSJJODXFBCK4HiyNrt1B63igwnP2Pd0WPApsAc+1O4433uDRuSOJ1zh4yg
hLi/cMzmWWNnUyxPFCRN68W4ujuQYcjbfl9cjedIFswS+hLj1kZPgmfif8aLh8bs
lSx3dYxIvJgTTc9jZgWgB0TZLDzT+uvNGOoflSU3Krlc0m8twnTTPurHC9OvYE55
cFgsx0oEo5GQgp1RbN0uAD3fG9ymYH9JkuucbIq4eZ9JTFdQ++AZQlqXjJ82qebS
dJ7wVEN/FenMW6NYjeLJu1mtCn8kwgYtlBYRRn4U1NhtlRum+/gkEcaimttNFxvY
7XPd/+3PpSuY/YwT0mg2DOaX+hwFLJ/RNmDy3fFdnKlVIwklwMi/z/lpDkuKSJP2
ixAsh38i/Ehc/5j23Ku5UMtPHwanvhyDKMR21SugHjB79KUmC0EHG3sedMcCGWN9
Oqa5nAACDY6jVxsyKeAAcp4UWunl2n7uENl6Ue7JAVQ9C3mU/iXSQjH9PDsj6Tal
9jRLZnwak2pGwlmo3KDQceSRcV+c6NRAeV9N+1G9EvqmoO/yx6BBlgpQLAQa3DVI
wBFr9hn5O3ZdLKxKGmDyP/kk4+bLXZXTjxuygNqpJDh/ESWX2IW569mER92zOkVY
ebYgTOF//ciqCt+rLPEt7JQ/8VpamjstoDnsXZP8uCCJMEAcI6JaqtPbE7ZwDXOb
DleUXaJx7Vd3JN2R0C3dSiqPeyVBEE8szc8SDbuEzdQg8vLeog50efurQpxMTdOl
0bkqb+Nludu/VWpTQmUSmP2pSXfqnvEQdsV8IHwM3M8L8Dubh2C5DSX42ftUqEHu
Qekb5bLzAxsD3qwnzbD+/W1/etXXkBuyGtlMCc5jpYTa4C1MPJ5efx1ySCunIBaI
mZceNrEOe/gKt/mgCIXeCHFPTworiEogzBBSLUJlruRvCQBoqILGVfz9Q3w5S0Rm
KKiD3nYKVQ1SRC3yCPO3yqGsnCckzw3up5VkIrdPmqXss3+UqIQP+DF8J8TN0ACE
Wsg1vB7opsA2KV9eZMlcSP5n77UN8zwoVmKMvUFLVt7/cQ4XjImCePnSSJf2lJPe
+3DBcMhut2bnIugUAwKNKVMl9xgGAq8M4dTZqhEjZrTOUxJz/CsVvcu/hxhoZUxX
ueDlVaDb33uU9QKSNmBb32p39kPi+u2arC5/NWDL4cV0dSm0lH0apyipohLFPYaB
g6vk4zsOQUSwgIO8TvKp3pYfEEteld+CLIM6YTfiUKjZmS58UgRXsKzk1EhyL0Nf
DfAeSrcxp3azZp85cH/MR4uBXDB1R2nZ6PS9keMz7ZE0P/6HsdIw8dzRPy44k+wr
wJdJhzpojEHPIKkHg7xzCEdqSRCo/CaRrhP+9KYMuXyyxg9Rhc8Z42QLJK9wP7h0
a6e6J3kCu8qCKhyECbrU/3tnkSLU3ON9ONGjI+mAMvTZsWzlEuguTxHs3Hswe0F/
CZv0t+XioROm/IJ9uGY4Xic2HpiTiU84sbdOuF0xFGP8BhTam2DMSQ69IdS9m3eh
j35hJbKE0NpnYYfmilmNC+gHeFEBwuQ2SxG8/mTH+lO7wCpNAyUw9SecXzlbfZhR
XK2J42yGZ96/AKIc/7JUWKCtjvLkIb6aa3p/tfTe0YlkMr/cZY5LuUnNudlSYYrh
rFk9+6QFoB8QeH55jWAHOJpT25FOkU5LlPO7lKxE9LgI7RPMQUYQVUv+ChJhR7P+
CQof/jATrkgSvKCAbrWJAQHtYy45VT0KAJCRJYok2qBZRoZErlABpmc3/l4F2B/P
H4S3ll9he0+SRTVJvi4hwucLROCioR7BmS+4fgmyRRXNwIxBxcDsFkTDsEHDUOoB
gVAPErhZywJQDpfDhqtacv6uH6V0/TAQGbf7huIR6ECoqDMfFah3kUOrZ/6rpmA+
S++PUaTR7WUcqZRZlB9OSOUVJFMAZZKjOlTZQuhhgV7tioQfsIfMGDjidTztotPG
Sze284mORRaII7VGcLRRU4k48N+DgYWfPddk3EI7YsTNbLuWwHy9Ypj1aotiZPr0
k+D/oXoQ3hHL+OVmfDSAQEzcZ5whS29TtqTLrqGu8jPDOpCuMYH7th8jWmdwZJVn
IiPu2aWdsDzqlTuZHYIt5fxvp+mdLTFEbctEEstxOipBLhp/Qg8SNUgieohEi0Cs
+D2uCxD0YUhFmkKIgnrIW1M3wNqUiwLUI/YpO3DGecXES7DO3ipHtNtNVhdKp/u1
iHjIMgyw4GnSSv0ln71xbS9F32GXSXbPchHmNgkcI4mB2U6Vbq1ws3/v/i67FDjr
8SjFuSR/WCwcUdYHMgK8SmqEgxN4nT6VjIakYnffO2CgefCV+sHiZOLeDn1iuphi
U2DDrdERFzkKSl3cTz0FUywp4W06llXlqqr9U54GLXvpAn2T+EQbBOQjZwOrcoCK
4r51L6aQtU9nyZQR+hc7ysEjY3iOopdwLX8FcUEUSspgQSobsJpBzzSmNIncz6Cb
Zwa6ZJpG1PgWKMWW98YfniPmGvlkJMFQdmoQBWfBaWjoMyFG5Foq8KQwrpFoiCRL
SABG192+cdjFGkEL27Zbjglt8vevYvtZcg5vd7cSS7jMhtsFhNBHlmXMrjZz2IWh
cg4gJltUlqhvV4eCffNOHcSeawUu0sGkwegHxO/f3A3Rj+YnqCb2vLvSvWAJGBNV
ccjoLNxccAau+p6SBk3KJW0nFN8E+n/CbN/5BHhVv2xXq3isslZrwJYaJyfQ66gN
K77LmoixVvfpB3Ofml/PIfzpiGYL2GnzV8F/bb9sw9h4ZouvQX6nICZ3d4FggSBP
yKmFQ4fdGIoaIyEHt83Gk8PChwQW/UGVzz0xJGwmXssbzOMNzn/ZsWVL1x4gLDiS
9GevVhb69px52zpkoCQm6GWwQu5QS0zi1LUXVKUHF3n0P7GreY3pCwYZFyDKL98J
iPZr/cr6QfhA+KZWoJWnWPx1e6EZzblxY5bhZBeBBw0RPrLkOmH6tzvX4lD7MF9O
i+P9ULNstOWL0wxCfYcQeTFfyd1UxHA4GgJ/iqXoh5PgkOgI4VTenS4OObFdJz8+
MN76Dh/A06HbCejrGMQYO0YRC5Ce8VOoMunr8XI3O6XalVz6XH0LgbNmluf8gW7+
dfkCpp7owW3VRQIVrPrF9rH4RLXjSx/VojNdqFZ7F7m/eFakyQH6yTBc1WRCIkZx
nwzvluLuAZ2fvReDwsl0csAcDKIQ3eGj+lwqV1JWkWsCXL+R79qD0HlEjpbeUXhq
vIRa7DxjkGzMhXc8N+c7w4GFh32cV7DHWX321Xj6HsMKT14G042DL7jhdelQlLEP
5NwJ60zE+MaPsXqUqvzd2DuKCvsEV8wNP0Incb/OKPthXqGNTF+lA6r7rykqQI3X
HezK/xSKhQG/GQTeO66TiiDD0jk8hZ+KpWnVMR8A/3c00Hf4VthKtz/DlAbhiPyQ
JJNHmQZz+OIiwiqP618YfiElFMc8MgDK0BuIHtK0XM+rAeL+Bqc/fOuDH+tvmQ2A
P+ld59KWNmnFlCB+CPoquIFE1BU8ExRapXFjHWZtiPHjQQCQFWs1dbezFiaxGOB3
ODz5EQSJFTTsMZGEUC/Ancnmy7AY326TPs/0Qm6IZAZ2fNN+jJz1aO8GzVc01FCk
3Jfy1HrIcpr7GA/tVu3vkoOJHcSq/UHSzpksOWu6AfyN5HNNnszaCIUCV7Fnw9+A
g14Janysh+xIKJFXF7wgZZXxMifP/xMbjlzWn1OHJMPgiwIwB4mo9/x2dmg2r3WH
gqUsm26L9BkMuOmBUDq1V3+tPMSEaPA2z6UkRZZJlSUv7BMgyDAghJcB2atw158S
WQrDwQ+cLFEwUFPemxNdiKmqSdeXjIGwLNx8cjlKEFKt6ziSWwlUqwu0OCskU+an
W9+7wKVXym7tWHmgSghwuX+6+txYdEkotdrgkNM7Po7Va1oW5u5q6xDrBIAGKNXq
kOWJDPlBdvjWXuzfORkHpVUdaWp9BOv3wKSVB/n68Hlw/ArLtE/2/4EDZixMoWFa
uVQDO3xcje2PGwU/ywXiM1+ptULkPmtTyf337+tCfL5VAuBNp0+pcCBLej+R8Pas
4kBz2ocLuWgMFqahy3mTwhYWp+mXmiBS8AHvJJd/QI0XwyB71GfNYsXl80x9WNEG
Ie7Wf9gKCjZhvoFBPnVy8DmwAe3CFHDhV+M1Nazs9AXm1J62gLqSkpWdPsVaJ48e
FafysP8VU+CtbFpwp0pHpL/rJUANB2pTQvDd0TV8hggalJpfAdAYOs5GrG6oy+gG
yQonPpFAZXS1EcmC+Iss2pgqQxsZNI8U4wyXO/lpqqWts+4+Kc2ZOtQprS5kOsi2
kfTXl+3wV0K9oVl/1gO4oixAOCWVMn8iAnRs6zPAo0XcSVaP9TU0ac97yKKLAaD1
EyPpeE+KqquONXo7EB3Vg25xhbU597UnLF/WeEnX1bCQIWQTNIqRU5MN/uV9afIj
0u/dLrobJnzJs2p+OmIP2rHhy/V8sX+KgIu09MTuIA9khJG4n/D9k8d9WSoHsXBM
yB7TlIV6QU06SDYaT3Ogr+DPWKQW1bDrzOYW4WCGwRmZFLs6F/NQ/ttHjY2FeiFk
Q3eiBFGMCYWmCCxA6s9/yAwZ4vqts+uIWyIkDLcFsUsT8akHiXuP63qEQI6cj8Kj
V9mUEb/HlNLoYelcCMyQzn3EkxFgFKtrNmfkivaQfSnvFV7hmH944okXRfE1q8cD
bbc9HasyKlC0TZ9JYivEzjs0gtZ36cNcMX9cC3I2HayizYlPFGwMpvyoxevNckBl
PRXXNtv4KE6vp+Ahnr47FC/AnGqBgEqJG2JWvc4jNrsG+l+4actSzZWcJYLidMp0
wMwwX6d0VTIgoYwUIw6qVt61YKxpyqfDOtQt4a5mXU9QALQqXygzQEGyPpVKdw8m
pKNlKnaGnSgcboUdG/5T9aYJlmQIR5ydyiDHCtjDDreeyGaho2nQ14lh9MJroK7a
tiiZNrXdlrWvIy5Fmm1rxVKO8Vmn+EDnt2ZbtGDAnzMD7G9yP/2/FwspKnm0Ul+m
ovJMMcI84KFCNTO2PIqrPGcOTQnruLFKR8zieHytkNFn5YVXEdLoZGLB3r+sqshk
6vnp+BBDjFQ67spw7l97mn6QyxLRIHBB2wIIz2Ua2I/6YYqtzGN/b41DNu6Ak6NB
OPprv68zl3k8/YCbp0R5MzNfoPXPuFT5CTRtcQr0U1zXCxx/VeltomRlF5jKl5Lp
sAIIKvgCuDdglMMjnb//5Fxnc9guUVj0zu5CVcE5tSA/U+F9DnV6KrVD0ie5KV1v
L/Kf99Al0knCnZtty7QSkBD3+17s7ZXv2Etr/tVXJdOIafudqjXUJtuNw3yahndY
JsF2fMo52MUTtMzDmS7SJxYKW6jqGjaeaRNbrMDQBHUTetayzISHMZooF0pyEdVR
POYOVjOESwkTyqZf2c+TG6HsVpKm557EWJojZdlhw/AD8Aa2xz0oyOoyBkpmN8G8
Me8aZXgiCuWmlUF/dKFmKzL5sasGcNZYVDzk1qrBv6Q/tsle5lbSqFqpSYYiZofp
VRDmKukDisb8JIuAeyl/Y+lIFzUlS9tbskf4nrfCeM6Wffl9bB3PihtjNUDtLCSp
tt9b9b0/oCT5LP8svBVsblxfVwowoKpG+PS6jqlv3pc8CCYVOVpApslIO0nqrlTM
2gD5ddJckn2cZTGpyMbX/L0A1GspFkfwPJBdlU0Az2Ka9dlXAT3/Wse5FqxTU80o
ctq1XZXuqttGSMnrMfyZEvUSVAPoEh3iRROoiyV7RUagFjFSvpRyoM5m7jefMmC6
k3r2lSP9uNypGqelDgLjJPl6ibHaLpkJlkb/SxR2O77WRIICyxnEf/rzU1nSEedK
PSQXNZT096v6y3Grb+CVvKGlfepDXjditfi2BAsZW8MEqMc5bhwgafyawl4qs0Z/
+6pdKNU4m03m9GuEx/iBJzUYliNw8+Wb01LOt42D75EaSq5gMbckPj1coA2j1XYV
t7N54ac+fca+5w1DZHQJtu8A1EEy0/75cZCjP855eovyJO8Uw1cddCjqs+UaTU2b
lrJVZPoIgqcryezlf4XP07EXYXsFrGylYWspBqNx+DbYjTvdly7Fu/JLHcsmJWcj
QFkKv5t4Kzg3V84Aa/djsv0X31wmjMxC3Y5xQLjG3lluB6Yssplwc+rf3Lg3HzY9
k2iVygG09mSLEEhyq7GWcormIcWnq5gYHHZIRTf+FIGJ1FvuY6mWHcJ9Hc/ySgj7
Unh35gEFPL7EN3SFHNJLq4qyo73/U34VLytIBkMMGKZweCF+AgvLYit7rsugK5lZ
IzwtuoeK3bA26cyu6qaW+fqzL/NZAQaY8hZmlaT/SK9Oj7RuITNLrRaHvQmWUXxU
no+pGTby+4wpacerd3PgXnXcknvnuXaXVVZ8F3A7sYeUj8jfOAXx7j265PAlI+gZ
zz3ce8DDuy6Q33PAfiqH/HPOA0uH3HHg3c+KnGh2Phm3AiQxLugISBbNcJvAGIZT
U8EdaxDjBe4qxVfmSUvySZ3hvpgWm3SKEYhNI2YJtsvQjVRbdeQAEMvPU7qrsHZS
0pB3oRDjt7AQEqAKrLfeU7LD34O8JNRf6dZRuAePUbqbYmjtHRgwqIaEz8f3Af5v
45Tif/s83XgKFvp5psCcsvYcvT4PmCM/CJ0pd+dTstdfqaQBDslqpJPA75aQPH8U
pqtKfv8vj1kcMkE3JVmO+ngmJttS5IrjsXAURiGMNlK/41aaV65G5qyJtTkFlsSF
IjvAWfLZwY08nmNw8eD1QKUbKAmKjxBzw7B0FFLSiaPF6pTS0lku40X1m84eJuVX
ChWGblDtnO3EXdWsWRU+FBj/iqOtKn8YHQG7d6OMcl8CSt5maiIFzjc5le/EiPIH
59s3KSg/3awnYofrhx2dm3LEycO6hpX6j746noMQCDQlgffbzcjOrPM5d11phfOq
4UIlqufUdYYJ+91ooqNwq60YYJbXaw7WMQ5arWb+a4a1HaoHWj+kuAtgFkAOgUAN
pCPL1gbDQ1khOcaH7F4caBgPYExIyFuQrYf6SlIfrJP3W74f17ApPtS/v4h57ixF
UAQSr3ZyoCTX/Lt+fCjkJP6EI8BJeujZyWirLcUi0mAMWJ0x+D5Sa9DSrikNHOox
t27xWiQYFLctV0JTTP81MZKZwDJMq+F1uPSA+fvtEw5lqRTUgKu/Q/tK6p3yMnpD
A6nFdmAgKmVNkzU3flXSxa0c5BMEPlrz1ysEN64LNGE4pCM+E55qsi5B6CJe1Yvc
7IUBINOsIapqw1pi5pbDaVSl85EC/wC18fymM1cApAuZzktHU/ZpjhvNA4X8YQUv
k5AXNou4ExHedN45w7cfWr+pFBLzIVMIzSu8kFI+tT8tePogpAAqgcJA7B0aPvls
bRX/YPP6+pQGJNqAhbspOo8ZpwoXn3W2QkS7dQc+0UbLCu1qfot8YtWSJhMSBjlo
6SrMpdDgRuhOqgI5T/slcAnIr8o2aBaHsGOvyMKa3dq2v7qOp9FMDmMe6QtIds70
Bldb7Yoiy815t2q4Te66+OQRA/TeB9zb0fHX9azbKqMSrb9a29icW+e+hioB+0EX
YaB/1pc7uNcRu5naWttiyJhvCW0eTQ6nKuB1Y7aa8PzyVeMkKcgh7FFmSS+7SynY
zeR/QdoEe3ogdfU6Dn7Bn7W6RrTd9O/+uilj/ccpBwGlKRadKj9zzKUxj+e/5Zlr
ks5ezCftd9eWLEnIzZ2m1jVCxqcYO9QoeavstQSi1fScxqAEFs7SaDeX/cI+Yn9s
YHOYY6Kh2taltcwgIwFxU5bzRrEUV1v3gchmvtlOHfuj+Qv42eL85BkQp6q/LQZB
KnYMfLSN1d3NXzEkHL9EcRzCisRcH+qHPiElatDWzk5XRKgLI0lGBgEpo/cIeVBd
pNg421NL2rzH0BkYPyAfalNUGmncPW2WiAsEYGvrhSnxLL3w5AQYdbDMs9nPrrNo
BzLhc/h/eSiiCqnhakpv/C5BYIYOdOMm1L8c8sTeqRcnWGGG3y639jTCpB5BIcfo
hLIvGxG3ZXq/TJgKaOtZfb5vbzVzcSdZGG08KGkttYUB5F0EiD2OZizMK0HzTKDx
cT2bSP7YWIjU6Rv/M1fHhcV7XRznWyyWz0q3Zq8e3+ae0AM6e49WW039v97Mf/cm
czla1/7VRShODSgfCNPIomcW+nUxHCW/t6F9GI62MYenkWqnqCwfg/vJqElyGQ4n
zYpexqriDg4DiN77XOMkH2pG99j/RnloWTE7YIAa3WChB/JXUQIiJdai/JMFtwzF
EWoyfkdU8/VE2v0LO8dieIRniV8XMAVA2vWWrP+C3NcvSJu1lS/UwZd04ntbWfu4
VdqaCzbjQfyJrO6gjdVPR7o8zVLH4BUla05Mjp/3glmFwlBROd+MmUL4KvlpMWOD
e/Ts7vaAos/2zrbWnT+mzo0qnel8JSMXcUpVJjxhijYiW7pz/fq8HzwRE8fnLTsq
b3Q2gVviV9rOzvUBLTQoGV1I0U14vkmuGwCV0D5V1HlmxMt6P4oRWgJ/e+eJt3z3
Nft/8WoxrhlIR2/8+vP6kZjLkZWaxbMojUBjwurojURHt6z0SIibjmgcw2p9vDMP
MBM6MunpVtiKW81QxWx6/NuURIgYR6KYWiONCNAzSNG4kaYnhKKoKo3JZFHI59+k
AxXQaXW2JrfZD5iinX9Q4gZxkSDyMiQuu/NE0wOf5Z8Ux1dr9yDvO+mL1a8dtHK4
r4UFbrp8OmlHqOmmbixEbLV1Jw1YNYc6ggjZ4+gZ7V8UK0t9NHhxq0GAN3+4kn1l
l/IQe6LwIZklNSN6rGKJcoqqOBSyoj1ejvac0ZLDDf495LZAZ1R8e/F3LUyeKJhE
f9pIrHJ0ngsMEGeatdpbbTJmfPDJqUWMjuBMjlk3EpKOM/p/APlYZbS1vwwxR2MB
w/FL0ENwP7U3gA0DhwNGUegTrt5Gx3+BDabFd2d/1lSBOlhINQKwb6GfoFqeElNN
xAy9Q6ib/Jtv0+Ltn8vqbE3UA5aKcN9oUXRMMO5v6tr0BpDsYUVg6xiadOfPO08L
la6hIbjC5hwHyY/mRYCiUQ0ZAFaibKW5l8PCDT8okP5EzyS/9cPAtR5XGl8h4Ayp
Rev2uZUl4Nu6iz2Y9hImGCz2Di7SAXasRW928aOlPRuKvksIRbFx9soH7GoBawgT
k8j25gCnA2LVfDVjHDqstH3/Y8Ph120akowKH6GIHI7iw8nF+5AscrnHvChSEAZk
Xt2NEETc5JbcdMR0wIdbTIJOIhQODq7dar7qteiHejIkMh04i/rklF6T6sj80JQL
nsJ2ZwjOZtVK5C6g0tq/eeTeIBiLIa/fiprz7Wi0Rz2BZOBXkGQSUwO9SS9ubJ1X
frNLiLt5flbfWC2h9Zd6A5B3GVZPJ6gWrI+KWhGtU420uas8laE/9MPFFtC4Nagk
mVSfIungTIH8dtP/+CiESRCWKQha6hcVPN/uuU9pTBeGRCwSTQiyT4LbWTL9eFwR
41XR9eRdJqXaXtwG0RG72rTWDDmcmagDwvnBQS70Ya5YQu2tFguWQvsDSictk+7f
2jtDRhN1IC/BbNGO1lFGuUNDBsJUTEeWZCPAIT62TW25FgsE2cDXUlSim48c9qMg
FFHf7OGjRcPiEN7ggKcIxiGvw1B3edAlMhb0FoK8dZ88qK+g9BV9hlNuzgySto2O
6Qb+v2f1Vg9r0567AeBftkWejzt5x6AVvzoNUlApcUggFBeI+i1mEWyftpttej3Y
SVr2bNGZx1kQhZeYRTumD6nTIbOdnicqpO90bY1xKbazlaQv5zrul7w40J8Gcvz9
TdRe6FzBTDdhv1Vt3k/2XhH3D/+QTUzRdLci1mpktJnFy3K7v80eCdMHH0DuvzK9
oU7ZBnPK9m925LVosLqW8C/SFFtMEnJO8LY8MleEMRFc9hPO9cVFCdeY3wcbXkoU
DIOHDfRVnTMb937gxbQgrVxZFq/LsQLhvjQ4emBNVCwOgTBtu2HR+p8xcZrlKtLp
QqkaltYW9fZRbtJVzytvcRGehqDzzJoUtYwLtJT14nuJVRuYuz29+DA9r4JxpoAQ
M6l5yrAW6ZNMgHDM0CTViR0H3dFhfbDE28Tv/djh/7U98Kdi5/ZBuN68V4gnAkLP
Ux5HkykaJfspf7I93XTqjtzTAUiGgpV/txhaDlhXwtqZQbLdZkfjBKzo8gCAu3g+
lEo9UHZaRBl1dpTNRm9l5YnQtLN4dZi2hoKb19K8zv+EenfCH+7m0KKvqVaR9rXh
vj77qHshXfjnR7j3MmEP0dOWyJjamIA0CRcfuEtZlN4gW1lmhQ6EKIhTfwFVDL/v
i24ynJU73JtdWmMA5a+m3XahLYPIWK0Zq2eEagXOmBT2W3nV74rxt+vzhu2o0aEx
53q52xS2Tv2d2f9xLkvs1qHudO4bpa7NGP9nlMmpmGvqKpJjSxbZF4FG8IVXy5kl
xLGIHgkcmoGCtwILcxmFDfhEWvKMjURN7AQl257aEfVV8BoY0x2aGGhG2sEwOJju
16BrWx+LdEITWFF4uswZHHIQzHjYb/hxqWD/0530gJRDpJCQf8IIgIvEDonGisu7
VDBzEKA/wzjEES/oobyLsVruvkH+oD8dNF7gS+S1BHrSGVt+oi8+qMRm5c78UMuO
1PgPwCec2rJCL2IhOjY6G9L+zMAE77i8uI5DG3PsWpUlsLiimEMjg9UfmeDBIyX4
6lPDikn0VsJZoz1tHkJszGWKOjitaJOSkIN2XOMdaLxPO7wjadNR2vEe9nia/47r
/CB1IiLwJUgbH9XZTt02sxkiRYXty2asz79SUwHW12dx2Zf4PQuW8hhgUeckJXk9
0efkIR60IRgowJob9gjKTRgMeLDJOUnmKPkFpX7/A8J2NtCnV2k2QldsbCo1VL2M
gRTGbQKwTAbo4rCPJZaEG4Poj7YsLJUMyQzsJYM09SyXT3RwR4E5OocroJarzkjE
4tRmsJJfwlo7anjH/GIuf0nooJ1fEWBOK1zTGFADekSoCF8xIdeoHxy+eETNwt1n
UyXai/AUZqDSr8Xz0zLN8skCwz+CVgJdcFBcbUZ66oBM+8xJRLCkF/zRegrWp/GB
dSFXjtHToz3D396NFjkr2KNhnA7cswL5foBbQQcMUYMBaKHCXal+EzElqrCRlCY9
i8bs8saShQd5D6x5skfLAPy6f5B+xLJ8DwGQYqAY/tY7+sM9FfcLAhU9G1XexTiQ
jWLmfjD7M7woyu0fOjmLgDbqjCt0pqPTe8TOTrI4Kvqxwjrm3E90jWNTM3fUSmNr
86WeD5ds7zcrX8+mynS8YTUICgmRUIzDLtVSGFt78dk0gmg21iGnAojjAQP+/6Md
myvbT9kc7LItzoNt0mDVczXreumpECW8Gn2lFLJ0wIQDSfz9pHZ1+3zEhpUeOPHe
D2QScf8UTBgZCz4LLSzIDKvcZWNKzmt1OJjSCSwHCq+ky5S+iWnjuwrLxmKPmml2
a23hnGr8sFTtXU32xZjVq75FUkK6Fr6NOFEptQIXZGObhAPzYPp91eAzq01XMabH
d1P3nMF7X8Je5VPZheSSR5t3a+fUiht4qV20/qCmkp4cTn/roEjLsdoWn+QkSF0y
u+HtlTrgchxaI/x+KDc1rOa7pasLhjTRSVceLoJO/6IVVEtv7p2LomT7mrAgOByb
FCpVPIo91qCCEbZN/ZuLhyICWOeu6k3IFjjh35KZn6wksgsSsyxrnm5wbvWYThV6
3yFByz3Usb3L5iXqssxmYBZ0WfimuDfORQMq5j+Rirh9Wgf9qdMlOj6eOLq8aRwh
u7HUAkJnGJhJVzmGDujtvCO+NyplZjyAULIZ+2y/yRsmy9KT0wAjCJdmsxOuw5ld
W6RSB4lsmO1YzatUmlar2CEF5hSwwPlU8ThNuQm9hNGDnCDT5wkJjCQFtRy6ZzSf
aQU+d9QEEVnhmb+33MljZDNDpGld0e3ryCKlbJBgkqs+iMi2rnAluLNQhZP5cAsM
+kyS6w3mgfvf2teeC88MEP2H+kdEKhjT/5/gSdLNNpJc5RJlp57xE5M7ZwlPYWwy
+9IBxDIF6bFcCP5gUsfDdthr0TBhkFsfzInFoCpRh9aJ452AbunlyscZseGX+yQw
ZemI32PF/4eygruujC02QF9gZrK8uJf7w0ndu/EO+/23RHom3SFB6oUPYVQ2OR+a
c+/Sc/9f+EUV/y55Y21TF7ueRb+I02QGtc8hBKuLqAsA1tPc2j/sht8gw3McCzLR
xXZhp1MdWhQ08Fhfe7EcRJ9laPI1y1LTvbuuYBoMr3VuPdT7JbSnkmJ18q2H8LlG
DwgPSX0VxsMm70vwXEIoRcuCCuV7WLrNcw4DbjnxLjWUqb5TRPukdmdYBDDawi64
47D7dquFr/viLAF9S8xgn7ADnkOMNW+FulKYYb/4yHMqNbl/Y2zwwED0WA6pJcVk
QihZcUGXUFqE0SPHZcOvHVRCQM8klFe9CfKG2W3m1lrYly6v7qLZsCaNSsyEBuyt
a5IF1WynrXhi14A/Y1Vl8IQUD03/X3uw9iaUEVw2senfahnBlC6E5ESSsV3Z5LCZ
EbKgLYB92Hc4GvWdbJAKWJ3GOUua4mC6dfBI6076xYMh5cNBkf01DgtHO+NHzFnO
lb9StgD8x4ZP29bIcwpCFatQve+L811kNiBWxrTQcYJYtV3x9y7piZ2rIojYZs0b
4QnrLeKB0zrrBBRmvm561/yONZWKDYuJA1H8CQxz1cAwUB7Z2VyhS3s3CNUhzRNE
JcSjOpnrdzcQ7WXSv3tAg7OOv+8WmrjfqKr/QBDzaHZM/XTjU8KTYRDviWnCfKjQ
gFGfRp9C/bcZ8qjI/BRoS1q+Lx0VoiKuBIK2bV4O63oTQUA6o7PhCgjolYiuwjhy
lldxRx+GTHhBn4zBrQXmlFSCFvHH7JwXa6udVzwvzlT2IXru/fD0lh4iLNYaEd4I
O1RvnnZVW9GkxQqkAljtp1YVE4ECtQxNPXRP76Odmdl+QmZMX8/jBHy9kifspgSf
okRGZVrCL0MF69sYIpLm2RXRO2vB21HSo2z+yT625+6udxZl1nbJc6hN3Pa9ws0M
eDNPj4fHaqETuRpmXM0uUPKRI9yTa73CAatxznGg5CsxC+b9KdnAwGEBxRnrRf1i
1lGSN3ptm37QQRijIcdX/pnpolD5EfMpPirJN8pY5XTNr0kA0aHK0YlLxeBf+NlE
3TmNDFO+iybsWDZ+HS4TEIlLAwRvaZfpQ1ngmSnwBa/5ZbnEjqc8t6lvUGDiUOzW
GwaJQozoUSLA8pnAygTKiJBa3sHNjohKhxgoc4X3fnNtyTy23i+01HsIdp/GPOHO
wtLURuv2l97qmxd1qNtPVRSrH1v+DqSzTCINFaoqIt7IzsoosWcsDJtRdOyQv7dl
GgtxCmTVKvuYZUfrXcpWnwhlyxdSYd+OYDAho1mjiQ/4xtwfqAofxGRq35bI1MXS
1NLnVEpii5o0UsuoRDJowmQoFBBLdrtEI60ASNbSNTpU0v41Y/88IU9L+eIeWZGD
1FBmkXrVheo5vKeAZfjDNhLDomkeRhSubkzRy0xyTINHq8ooMePQsi5qGD0Q95Ql
ShCxfHz7bJ6NuzV21KHjBn3FK5QdHE9tK6EXf8aM/kgr6NIuX0UIJC/EsNRS8KS7
GKoHH3Y1H2hJAxyNvx1yZGPQBVYYlRIUY+QY0poFsY/DwVHf7EE4c2Pg5Zs7VGBT
goffgFOLgSjZz2Wm/aYjULCdeeqdYC0RAqAvOhtGEHy6vSbbLhQIVpNnOHB/spYO
8E8nwK/cK1JfDuPhvuyV75Qd1D9Qqdm6Jf5rmv4n7dErsQpMH3BBJ7Z2MC0nwmwH
jzrWs9py+LnpHjkaqKO37TmVpOV/kNRi2rt2VSk6gMo1Y3ahhmwphEdPex698CaD
H9ZNVL5+cPqXUuGHv4VTfqvoLEIJfqoAC3GwbTuBkgETt2uPRp5qlv05FVcspuY+
3cOTdR5f456GvtrDIp/DPNorgbg0GETQp3ToFKbvNRlvAWmWZI1nQmbQvD4+K0tL
CKxFRigctWxHT1eL+ZcsGvWzATdpYUOtV04/q3/G6YMFr42iZfeYoCxeXQxwKSF2
RNIV36i/kvaD5McT6uQQjvtRTC0QADtdcTfdrQqqZGoMLpLCrc0L8XZ9aAHMH+pb
/G5dGutW11h9Lz4wXl4B5IaokDZ/XOMQZvS7Edv13JWQ4lKt+hPuS/hC5lpKAH7B
bkKjZC+PMuIAfbqDPDG4c3bIxyKQ3bvQRF1mNWNKNJkPOveQ327KPnr++0YYnSFH
cOjJZ5usJcd/X9GZaVsrET4TvAjk9LPXs7CHL9fE56GiNp9VJ72XJPjbrikv3Gq1
kabCA12Tid2JdPtlq5za9GCrRCl/KY2labbZgAuVpDTNrsG0Wkn0mYHjRBmPYC/r
L1CYaKLFi2zHhpkLwGa8y6jCI+jPQvHB1Ym7HvZnlmC1gUKZmfJVWlxHwCxiLodp
LCehDV4nPsZuXQeUSdV0fjllLZQSgh3GasM9RURKUNBGAS8rtGmYJPHZ/C4+oQZD
U93P+5XlKpF3F8kpmST8aUszCrALzCK9Lh5/VxnPrzO516tqrI0a79OFZJPkNT1i
aA7nO57pFeaSSuvpTz4SN8MetmB/kYV6fwshZn7Y637DklgYtCe1GBM2x/c1Jwzw
K7/wdSSi3D/XDZEh6lEHYkmHQfoliyoKGcOSptP5G/QTgLj24+M0eb0T76/c1vbj
xl2I4M2dOk5xro6IthQXvPupjbrbPebQU3CR5o6f54ytEmyD/E8uG7FldNzevRd0
B9WZV3WZUcmMkwFIZpyMpJf0dBU3SGRh4fTpPX7JMHdVsO3mAedTBDMjJWDHNzPB
43Zq4Y5gKrjLkSgFeXby2xhYsdomzAJKqbd4a60Ocay+eYIG+U4lF9Rvsl7t9iKn
fYHezssK8gD/gT8I86fp7NjCilpv24MNuZAkm8vOHjoTGQFz1MAMtY0/19bqIwSo
vBr9UO9Bo8SRzHo+Qy6I/S3IKZYVjQjJxpLqw/m0MOHEdP1bV/7ZFZ4R6WU2tQdc
DSvoOLqeTNme2IjaluJvT1V7a2fxLWofyJSIZCKE+il/NersAmHFST/x17eAZhcI
GT9dHwasllPaJdOLzwjlXrJvpIb/jvsY27iU3/V/cRzHzFxWmQsbVNS7vbqxapnq
IeWn/l4Na7MYCiGnqlOv6g+LjMBOjWw00N4xJQVj1VkfhEXYcmpMiP/6lJNqAiJW
NfxPJ7gKTPVCb85CD+j0VSXoROYYPNFYkNx2oRKFCoX9aWgxAnbQYqg4Hq3J4Byk
pRe+HjW+kVo3Z+8Ptmsdu5KDzRnC7zRsoGKDJM44GO9WQ0V4XLAvgXjc0EudoSbX
AU6YaTXBwo4rqQ7ftDeOc0KDMVgsqYhVym720ExzpdrdhdsVyuiPV0WRrv/iGAEQ
e6VTWJRCCoBhLU7uZTOvjkN9nKmrXootbREYCH3MSOdA7HO/dtU+fafmz3cpEeFx
doww4JX2Xgd8zvWg5zTaOgw81VLJP/+gBGjbkWTHGaMsB1UfO7eXwq+Yw3CQl0rz
MmypRV+WyIC3xiEaxptv4gLVNdbDMfp8BtkwtgBOJvXCMEbPM7kril4AqMvUhLfa
LO3wsEXi2OiUwZXH69zTUNmbPsSNN7wBHX5umcagv93TgqHnIM2GwiGKXkhhqacu
/gCnjcI3emrGgtwY1ty0P/gkUovwaa8eFJq9IgDvNn+u1BnzDvVOt9vFupsDQz5U
KXN3DqaZAdYl7qAkSa0kT6Nms2abRkcJe1BUk41GcgMfALNxRRoF0NmtIW+W98BU
zw9A94ryAv4rUwSoAOkPcZRRa9qHP9yuraXwm/vB5LXBwlKa5KGe5Hd5yH+5R3FA
Ta6zQVipDIgTITztndpU3PHp/JvpwJud3TGqMOKGoJKtLYkEUUgrO8SBgAngx5Tz
YVcto2g3kpiYb5+fIOOdeYEU6xztCQEv4WzfdMOGnuH66r/OCXcIOjfdKnB3RQVN
FT9kUyh7GN163l5HMgLwJOXKEdGbz/MRqMwcl+mbDM7YhEvVISeRaVyY3bd9ADt0
CGj6Hyc1MHmEbqrU+21Oge18FF7xeUyh0jZglEpKFoEG3RsrhDzMpW3dGasJ12dP
aJCUIg8DN0ypmVpUNIgSIOZNtCw6TLqqkpewZtIyi0rD8jgVKNKLc2obln2xiNEh
NKxE3qfSqODoaAAeB2hjzvwq44g3DlsIyyC/fWffj+4ZJIIIWBqZOc6pGwKanP+J
NTyLBaO3pTGNVATOODs8Gf2XMw2PoZKk716MHpIlreV6/3RutWlQPWa4C72pJQYN
xcqqMGxHjkBEusmGXppkdJE8pvu1hV3BhkLfXqgBjtc5uPEeNxH1ZIfNMuWJ2pjB
M1gqZ+y8unIoRAWtcpcx1Ow1eQtG+A7ojhfVkMayFsTtYBPWXnwoYPjdtDcOEO9F
h6Sv6w5vQnxc/Vna51+P6tiR+opkRb8nETQ5/qZmyVXfPjT6PEglM6AMibGcbbPj
LN7f60TmBRxAD9weA+Tkt2lAu9vexNrIL84yeGGWSoj306YNm8JV67JVMBLiC5yH
FnSlK4d9Vn2VHiPerM+sGt1tOUdaX3rnDO3LBZizD//463ZxKCDml8khRwrBUQiZ
KZa7kH27y6Mxj+vX2UQh+eBSsviBXTgBUp2dGNEWXPypZizv1Osj35FACB08OEsV
KdrU3F3V/FmCLG5LTMD+1yzd91pYSNDqCGsf1a0TufGQJsJimkbayUNJ8Wu6P7Pb
nmKrVCJVbY9V3hrRYD+9OxGKuMsw7N/kRTfc2WWQdAo+B+bM2xZlGHZKrFdEEECS
6l9x/tsbaw009ldiXn5ZrwzfyX4HgUM564UA64lp4xESCP+mENeuTI7w38jzO71P
jUGtUaunsLevavlljmhI/Dalr9mKXFFF1/KAu7fT4GBtU21yTB0Vrq/vi5k8zMKO
B/C6NpcJZB5Q1cWn+jmXNmsdZM20Q3uXwfI7YKR85yUINkJzurg5zmMwnjI+tDNy
C80vhsRmQZ2AAacs5s3ogP5PLv43wHqMGwrNxCBsm7lx1G/5zHb6cdDhfl3Mrunr
3zUNz3Fvn2k8KF1T+TCz0CY51NNLTCr7QMdRh4wBkKIBeDM/+kcPHda9UnJNHga7
6yXzjlrsSX6nFUl59HLe6AYzGuLjaszvOPwFSsooU5I84C+5sIVe/5v713HaHTuf
NQj2dH/Ga6DavawUlHNCh9KJsXWxKUJ3hSsy18fiEun3ydbV6kSN2s7CnkivVqcY
5uDE9CYhYUg2qgg16wf9PLVmNwqjU+8gvqmDLx5WeUN+1hWGdL54Jo4SHRMQPms1
D+EJlpnvdOgdWe8El6812eGLaJdKLX2vxZSdByy5x3Ufyd8jl/7VoM937C2mmx5o
l9pbKJaSKZx42ApYuikvqgUbNHVRp76OvoQ2YvwCi55/Y1Xp0+g2iVsp9uo4ZnpB
FniCZbFFm4egG6U8hFPdTj6mqokWdvXOycQjBI9rXgrVbmns4QAonnk+Ggj+ga7j
jb0/oNbPffS2DT1dqHaW+mH88KYuk7IcuZvdnAt3jSt8FzHZaSnjlUxlH946A55l
rcPpYVbYPzNNq9qUzQ6oskl+tKjn7rStLLZiWQnvxKZIejVf1ZwjlW9RbrcoiuTM
T6cOWcPv3PrSYSVunrOoBLw74o2ZM9r1+q38APGFkTjc07VUZdW3pdVIrfK5wjeG
CVTTGozJ6hMgz/ZsOEJA7/xdHC3dzn/VSLuchXFM0lrXunBiAAiOJz4xp0qdKbKO
1mveO71YpmGUqcqbsdgcqwkHZdf3HSEY0H2650nimDj2PKinkWfBiytnsfY7/jT2
GbRsxK6zLYntuMZZqyvvaBMgJGsJodd49aIDLZ1AkRh5JnwHHPVa524ZKXzd0hBW
Px09LAzM60V/eTfYiMB139DOfiFZJRXYsciMuLRCmRy6s8QcZiPqkANxXhnr9uVe
ptPhzDAO+qTuEw6bgs5ad/mhwgiwJapm9Bf8+7K0Ue/rJz6B4eZdXMcCjtwX+2hX
VV0mLYEvjaWvyekxCtKg8cH62t/IKV6yVNmsLYf+VZlVeI398Q5LdLqjYIWgMaF+
GitpZ6cK85VfTB4U+vdMD1cIiGDq+ok0nhezbAOXNg7vj+XfvOVdOz6qDVrGCjLT
udftt4BXZDfSPiGPm4pEnjeW0Yb1ZiX4pL8b23Y8Bhkx4r/Zasn0ilLFxwHK7EVE
2bM4ddh4Rzaq22qgKeEYrF8fvTogOE9AcX48ujurblJ8jlVZaZXu8dWhlLl6V/l3
Vi3iLLeyHSE+78QFglPSnUTjThKD6JfuFA0lCSgxUJkC0Uy1Og0cTHCsbvX0YtZo
ODnxyRu7w1Er+FAz+NdXuaVrKc4gy2O5ikb+jVwBuYPZBlAk/w6+6QC9vsboJhA9
bQAdhgzpmhR3z16jQHeLfSuAU8EW/acWBBWsI15ucV93AB0vyuGJySmQ1sidMMDX
9OS3RcN/SPV0N0KsoLMyHqvV3NdaN5rOyTXdAAA1xVpXDN5Mns6AwuJqzCL1O7fW
9uei9BxUHO8yhpuf8NPp8BliHfUyQ0cMjHYQoWYlLBt34wbTqZR7SsFozLKrj9MS
c3lVJMMi7VREqzureaVqUonaMjy3u6egTxo5Oth5hiUkLBVo1MiNyngZOy/XJJT8
UttuwdzhVaedia9iPFDsbPz848uWWBS7QsObDquzYwbN6by33zHo18fTLfQibu9f
IVJTd81oSLR5YNW33FTYvj0pUPkQh7p0hkHxPpAzYutq7BsAsZ/1i1XaFnN2/FKd
oqw7RStiBcrq22tFhEgtQSTaZgv/IcFBvm9gOr7w5qCyZM91hr6jNmFhlO3pijQy
3tmhvprtTdLF7110u5p5upVC/sTYJrMm1mtvL4b77c5vraZCg34mm7gLluVDz9I2
Xwnmrs8MR2fMJNR+1nonAZjhhXVKMj7KymfXZ1+/YssvGMcQFuLAzmw14H52vByA
zKksrK9BxGy/cufFA7XUDYbQr1HswAKVydktA+Z4R0PZRGiP9NXRcUSTFiz3WM0M
xlCELf8D/udN220Ngni0QXiX5yH+kwVx32ld4eVV3aXxC/eZ7lOocPC8hOHkEmm7
UQjzxsKIE77D5xNEmWifJnuWXcEfMqCrMOPDLPY7NXlIyr0ESOLIRuq8UhuWrSxa
BhLAFDnunmfhWHVfinKkeAvAVJq4JOq3NAAURXZu6bqzHIk/poUxMehELxQv1DV9
sFZhWJEZwxecLPaV9sFf+tsWfAfja8fJpSZvWe74ABzVJQEFNtZLro+EI1xl65b2
/i3eaoTa5mQ8Zp4s8C60FmcXHViGP125/YK7qnMCylYkFdCalb8CQwasLa7mdXO7
r0C8NmFzae7tzVDRXE9gb6iX701C1ZDjUP1MFYVOcEcvGY3jZ90xP8McNYOJI14H
xsTyusLS4ccRS0P7vffuiU+2q/HLlUGSO5Jd2/jqHdq2FN3OgcdD7FPdzD+H8qJG
evFTjCfdsYahOeG6/bOcGB0erLwU2W2gNl2ubAjGAF0H8cA6NOBoLMsfVNwImDzE
IvRedfAkLNQJNQSJ3rm+Yw/1vcaBoeZX682ngI/8PbNaPP8AThUFCdtYWv+N310v
NBNPPsp0TOaxEWVIZ+nKBwyIBEbQK8UX/jnddKOjc4rH/Z+Ho4y65F8Jl4g0mhWy
ujfYTszsK5iT5+B3shHIyxklqm49ArLjMN5cp3u8Hmg48nx5YhtyFZ5KKi5gqbTe
lsuFWgBFwBF7jumrCqvdzOxSvR7ORaehALqrrU9Frjgv9KdYC9YoVDwZw9WtXU9b
W4wsoSWxIBeqRw615amhE0PvmfQWUlgc+DXuVpDdCGcKVGuMEB0tAQJqzk18QM1Q
8szHpF/rb3K8h2WOAJYbyPW8lXRw8w8bpXTcurQPA1xsFQkLfqJlJvrXUj0toN3m
3HKI3YMMFDpYD0TjKKjCHYdg/SgUQLQN1WNvDC+2efU6swXjlO22XhmR+LADOtgL
zNe1gc4HvIGFgJB72OBtomDMkwSxTfWv6oJobBp6wcgG5s1CPqb1RJnE5scjmoj7
uK1VgxOOabkZlMSCf5hVVpgKgCZhjniq959sQYbwdoJToj9S7jT7bZV3U74sBMD2
of1m0Em/Z7AXQykq4KoZbN56dm6Xsk+pmMM6ZT5MKRZFtf4mOSjDGocf81eWtsc9
VoBl4JwV5FxTGfWM/S6E1icpL6aiQhQpxLm/MNejlPjHTsy5yIW9SdTCghHNfmWi
qg5KCICzU8FOn/gOSLkLL9UZo+qh4pK2DkSBBsgB9v/xZ/NVAUkpMdPHqkmw7+AX
79+aJOcb3MjGDBMSkb/7i2AEjOsJfBC+YU+/RDIm79BsT7YSPuxLQ7sJQHuG171/
SSoAknYo2LvmIKq3LHP/f6fCR6GHzybzp3Fpcn7atv5Nan2FnG3dJeyQ+13eLExy
uWGBhkFDfm9Ic4n5JGjD/JrZ96KiCltkgfWJ6ZKBnbWOi12jFM7OLrQEGQvm9ZYy
QDplOkZbV6rx3f0AcJEP3NBHkH5pvtC8qxhxtLvt4hhtFfLTtE8D46uhMCYKxuPd
C4hrERL+6L6rhF2+BEWEi5/WDxZn//86PrPIBaXm4aGAOtcTWk3zVfw1CNoftuPA
KhpbkOk6jUX4ubsatWNzFf8xZvs9me3/ig5Ms4yrlfMU2xGuaHj3V3u7vujcFMFA
uSF82S9YLwEnQK953EJN4C57q6l2CHqR0CtEbSAzwL9DORIQ/QnDPTCOl2o6AcQX
1vPReBkqoQn2P8UrQz1xV/TOgRfsKxxlbb6gOg3sgzl8HlA4JXCGFaAdNwDHq9ln
Haa40bao6mg9xMDzkoC0Y1upYoZkIYMJbv9EShrMfAsgoRsy2uDfOQ7M0Tftx3nA
7L8ZHxonzAYqNau6kZzpN6FVZt+lHWcPOxGKNJAEgiLBQf1ejAM4KX3JB7tKuBYN
1WXEdoJzayLxxp05MBKt7iOLtYMqyWx7Eh1KDqg60HBP+HdM4vhqOsrlh2MlOG4x
N0dvCQPfAfjHFDrkJzBZ2FQtQHOqynabf/gxxoz3UMNskzB+JnLNTggb1jek3mrS
i/OFHmHl4ovTlqqGeXSWaV7/1+j9HFhDCOTLp9cibiCwlQ06ZCCYWLmHx1HMDair
PD0yMq7eqMeXSsAe9MaHYaXaWC76rGMQQeF2NHpX52pBCGD2Eax73owdXcRCoZZM
2KgKQHzunLh9Z91uNYThiOCdts757Eaysv4wBJzyCsnbno/wMKYnXj9TS2Z+kAnN
EzpDXGEurONdTxHT4v75CpPwY81dUnic9oq5XBXs88JEPu+aHQUqahloRgmTxwAH
yJJgG0RVxS21T5bJ7mfnMO0f4JVhXCaxypy9TwMHTncreEw3bz8gLvgtVK9XPEMH
iAcWhWaNDbWOIfRHTljfP39hPEZjhHvcMxhA+W0WgrCw7w0YHRkV/VhsRSHT4IGN
TaSu509knbAZ5owXok7IwhHrwUnSVias1lGeIRYC+TSKbC2kNd5m9B67NoHNGflU
nfus8FtAXbVvikgtSay3He/qwgLvDLBsZywSczguNZ9m+MzBoYeJqbwcESlUxjK9
Rb3cjJanyrrVZxpH+I49qfnECOsfAVm+WmVJuKMwqMJbsOB06WvroD1oYoTbO2E/
XvXUDby2iS118AzZvBvA0kWN0kDF28UQDjTF64gEvWgJ/pGdii+PZC51nUM1tBIm
t+OJlSsmlYVmzkW2fnnEvLtgmyv205Qwdte+S1p8KvqobtlGB2uIlI7K+ZqDC4ck
ULGef5i5d/53M8Q6dwjlf7q+1jpi+/WFQVfS1nlXGW446MZcn4RenRM0e7fVTjto
jFKHxpQsaXliM36WfQ44rbkwp+2oCcis+sd7KE9IyZBVx+x+p2kVxTeSiuG+AQZ+
T6r1d6k8rqBBCkz/AqF80uUjzCKjEb6HV3tRgJTNd4ZSNEzqMTuDAU7awuM4ENtk
9TTOGxitwgQjh7Wg5jgTHzrefmgRj39Lm0xic6lbWAyOStTx9SjZAqkWJMlPFJlq
OBOdcLKM7JqqbEcXs8X8QSXyCDWloLNUwnhGi8eAx9OOeoU83PfGbYQAnP7xUqbQ
hC/5ANsgHI1+OPwDXmrv/lEQ1pDdded7/YPf9ppfUT0zyycLsJf9WDbvb3O4MAw5
rDgBPb47O7BWhszh7pPYGBp9y53YuBPL7XI0Ws6EQ77FnsdTN8TUzkfbmqJTJA0b
bVVb7WiZeZV68FF4Jh47gNeceAGKEFqzpPP63T47nH/j1nxWYleWwvejyynRsDcx
JwfZ0lwnbz4Bz1Ozy5LbTJY/8MZEQ2B2OTUbsvdT9fXc/B5SuQJVsLJ74tfo3jPa
Z+iaQiDk6YbxHwyW/Ghc9bFxaGnLp+HprDA7fmd6e9f6aA6lV+CeqHF2MWT/VElp
8lSKobrS2FS1Zs171zVADQJjYBdIli/Q/+fi7bjz6TkgU+93xzenxQ8PSd7wydLH
y4bVjvFgxnaHRTSrzEC9120hBaZ7dVL+wk4q4JsnMHxssGLJufnuxt+nUnCr7e8X
P8YQ6FPFwVwxhi7vvSNX67g7WfX3MUejt8Gcuia5gDDiFjwGMGtZTbCc5VMYQ8Tt
wSQDzje9/yS7jhMyuRQ6istev0yQQv4x3IudguSHrabIFfKhPl3ekSnjKphdj4DP
Gjxk/lvqA2EVO1O22xSITEsi9u2Dcc4G1DEl4obiuiP/kRWiu2Xv3YrlS7qWWXTo
28llwwbPmg0CegQfV57CKER90pCPUVk+bO5AAkQXa+uJJuRKXutQeKfuATIvsZD1
rUjBBsz11AM2Tg9WNrRFG8fUmRPP6dgGn1MPEf2XzcVDsGTYuLQGHwyXxZr03r+K
c8T77xW65maWquAcnd7KotOOPg9nZErhuCUGhH5L/oafbeJ6yrvPTtox0OIYYkFF
H3I+RTRBKFLw/TDXQXOhBMx8dhQuOSd4xfcIHAigYmVULYB5wmUQYK9ag9mx4Bqx
AU71npqDUq/2fQg8aqmfdJnCNVAjcSc/cJy5HmqU9T6J4oUnYtOpE0vtBNhm7Wkx
aDH80CwbsXNpVAQZiZBSFQK8263CuUa4r1wOEyBF3DvwvjJjSZhbPb6OvZpFniwF
BtguK+KHPykapl8FDfe4/HjAL2Ht40xVJT9dpPRjVxMKIGOSjTy0Ln5ukWB1F3OP
KGhcusWiTw0VZCWksjxyaQ+9tmkIjbcgyTpHIwTR0SUi+CT9S6a7YDEnm0WnHp7G
Cmw8oQbN+kCNfqDp4O4VQUxhQZHVpR/tlLePu4H5zzqfNZMBWvARKFrlSWzrp+aL
1Z9xNNEIq6v87YBSUJAoq8eCNyG0/OURdbs/MbB1H6US2zRliunqo14QMRSEc4NN
YzM2PlKUhOlSqQwi2SCMZIQM0CHsylPywUesKPUpbfj/QYJBO9Ur5C2dc8pf8osO
wcm/s/prDtP2Gi3aBdfKv5nQo1utqEroZYPdMXg2Poa/VFDRGFn04/UiB6X7OJtd
iuqtl19ZXwis1AjSb477NB6Y8xlKDskAegz1oPuiQ1WGaCm0k74/cB8bboTiTnwH
L9WEY/PhkD1EyC4kQzorZpdDvys4BxaWsFQFKd+3zz3DXMHVAK2sTiMo+mMa+YSX
5qJF9WSpHVNdwOtyriPA8/tKryjiPudoszTOzuMo3MDyx0bz+PSM44pFS7A2N9YS
kyV7XZyS0TwKgLSJRfOI+PkVTpqWV/82D5MKZkSYwwtcHJO9XED/viwZHYR7b8CW
oZjLdsArQ/gjIZyQz73ePQomAXohbAVCxrTZMTKI9j3/V/zPDhXlseIZJR2NIucu
Uun9i/xIgu4bX9hx5daPBP9IHBVqcvpG923kfbWxfOS6BRcY2O9ThInjgsIvy0de
qPsX9ksbeRPAvC01vcRA9aMn5o/1lj9OIeEjvN3VMROQhuQK6oK6MQowj5hob21P
IMqdb4jOKHM5nGVRosLrM7C15cSkBRQnRs3Oyi8tUYeCiDWS2t6CIPTATocGRLCk
pdzm81BO11cf/JdNn0jEnyUepfRP+WrgMztB4TPL2GOOCJDiQa5Z/r5nv6MJA5Lq
Y+onHp48nPzIWvxy7OK/P1KaDlKkqAxosLSvLsLduz+jfnF1XfvsFpeN9xKY7gZV
768PplDDEM/GDwfhynHLIoFuAn5TH6ohXZXWufPbDTWvVEcWF00l0fub3Scu/zx7
27QAiA7kZx5uU6iJGicd8tusjuesuuDUprZBp7vK97UDUTmr7nHOgV8FWFxZPgCJ
LhOxexAGeLzkUymu+m9EFlApnWJJBzTp6z0Z1SJOJFpoYhNsnngIHHiKa6HJxi9x
Qy+iWYSoFIX6jyjQesFPTBPTQxfAfSCMyfvd5gxfLe9rRM/Zq4OgMW/rvgri9MfN
vh1N/VcIDaOaLsx7L1KOGDEFd6bcucKkY6wpuwBzPaXg3vf+RqjH56FvbFdmdgrx
NsMQdC8rwW9ZChXhz0VP6uEyJiK8bM5U5354BsqoyeIDfrQ+X8X0nbvH+v8ESXzA
GyI8xzt/vs0UV3ecrwZgMQ+vPv8Q7WLHldRU+zYimUNsjEFfg2tCIkOKOlvNwL+W
mZyaZ9XsRVJD1QKo+xYECHADFCuAWGWUdi+srIGFwsHYGAdOXCNW4aKZ8CElBhUn
rT1Cvvq41eNLQ+4r49j8AVa6iWvQw2Z/vEHaUBPzeEjdlaGUeTWAGFfsN3LHjcFo
/IHWMgAw7+HTBxP9xGQHDrkO2wQSMgTUI/NgQjV6F+Zmvzzc3Q/QXbEYar0oSLfQ
Pz8NnNUJmkaEVvVJ93Jc/fR6dRGuicejFBDags3hUsXlwKEaV4QXfXtXKMlqFxPH
C0SB1a4tuQ/dDAS1cmdrctWDI4z51t04uVGV3c+Fo9gJzpkiE11D+fVrTy/kyRzM
BJ73el0d/EPXV0x2PLGyIVXfYKPyhqjQDM3mB/uxicV7haGrswUSOWPlyjbVYslp
cDb7k9kJEdpMc3pz9Si6mznbE88jFuD654bTnDceshAFQJnZfFElxkIqZnKTMjUT
aA0Ibvtlob21YOpWEmJ03UPuBNycwfoXablT3rkRsSrwJpk6ZwGRbhNOk19lGcGg
c29O6RIgswOcKe+sPIrhsBHqK4A4Tyiz9TGmyqQyVAfAYEtv/ziDIUrYDHXIEVGE
SEove6+26lK5wyLS1dk82cKLYNEuhW5xZUB2dGIs2RGpDw0oC6jKHACErpYrcUnO
wxRWQV7rMbfhaBTMxdYs+WSLyAOspCw5G0atpNdZZ41T4UTfb73V2edMnOqdXkJf
kvlA4oTBV1p3LxzlsVkCMALlLHqw0T2djx/b/gEJ39J0llviNOgRQIFDokcKH63+
cXndbX2uL1cCzt0swSZp1U5v3lyEQ7awraOKGSQUzXQ1UdMNlb6N2XxqBs3F6wmA
tIPFoUEaVxpxJYLtTTRaNRtOOrEdHrKNAZmatnmy9EcscAVLlUZhVm8+uCfK3nEA
MtkeyjjaX3WYsbF0OJh0X2GddmsWJlBGJEV8Fmwmj5eqTv55646xhP1CQ7V10nF7
+Yz8N6U7H+7EnKm6IibQNq3qHRIR+rYv+WLJxB4bI20n8Gj+xZHmSSWdfnEkkCMw
H9qoni+rDCim11Y97gkzVzHEC60a1srHDFhkIvLnS26IWSrxZhrd/0UzMrn45eih
vU2LHqhwRBfrwrv0iaSi7xHMtiMFbrKVnbvpcVbi/Y5EsPKgTYab0/TFP+H0kK1z
i4oP+wxnuHksSlC8tYRsTiVvBQP/IeSaz0pB9VE+Szns9Sz9xY0H5SYqNMgv0Y5X
/m44aAXp6pJ3dH35iE5KREZWxFK3kdlwZUXG6r0lj3bTx5C7W/RpmGxyUTIc+x+L
LH+iCdt1NlNZlrJ9otsJAhQVW6Khyv3PRNjjjfkpdLhtv5K811vJxY5U2hn+2k7F
BehiLYbpQ3U6Uyu4TanTkjO4EHgTwhY+UXb1s+TkTFFMZZ/SkPsBtoLSqy9QelJA
qbOx8sbGs2ZO9CFXwCtT+CbZ4AvXE45xSJtprIIyAtNupReEDsFGoVxwhuq3sTNa
UCeZ50z+mLof+rVzrvHq1YtlaFNqDXx/xNdRQgzdfN82iOdWoBHGAMpvQ19Da2la
tETDEe8JSYqbpbzruQEDFFr0dgYI471Fcao4x2KUe/XtViQ3dWvFuhwlKKXZCOV7
cAiDyCOlg+z7NxDYIr3d2rz6aJtdXFMDcvhjrDX56BMbdofNv19SJNRL22wbXfcM
MUUnpkaqeLfSkHVpvj/7KmWFyCyHr6XhD1wOn/aE+LQV4SiGWCehr8JJnEB915EP
eOpAzbxhjOKxCpf7X05wK0M6q7cz4YJHcZHMAEYxdy/bfvnFdMhcGG3WpWn0MHNX
HGMapQ0wTEp/mpIxbZcCNUFMshdKoBWPdBurNtEtSfX6MulpWQjL7C0cSp7g2DNC
Y/nkeKCRJA968HtpBz7YxTGPrilxyRcYIDmbBM7RHIDX0sCrmithOdqaJ8Iu6+bo
E5LKwbXFgEXTGWcGGs4gIQfSDuJPLsX0J/JBrVFc/7W663ZH1RkEwRc0ErpE9xqp
dHlktJHWCNBKYvvLNDw3Zzg3OLXCKL1A2p7hiAoLrYoS/QJLS1D46PVN3TDxywzA
JHfnrbv6w9Tuum1pPgD2/PM/n76BPrjEVJDKTYy2AdEua/77lNfR+3gPotBC12Ku
cssQ/zZ+su588wUsHOxkfsBDiUIh22WbZm2dLdwVrTQ7LxYvJEOshq16Q3wzEtfL
jDVhm17gtwDtDHBfGKDVw8cMp4Vkd7txdyvMLAb+e4TgrXzZj9DuoTSeFpcZ7MQN
bgupOxrD0KxCP+BLTdXLPEfAPdDnwvopZ7RxnAmyE4ihlTU5GGT4cyNsCBo8Lefd
dAxT1CauP1dHPzYVaHJCfVfDEVVeHLMBzZ0yonw54UxEdhWddRXbpRVLmsPWgr2A
n4+hhz3gS8Qu+MHbEd9DAacKwDwMMoXZxe/0pkwxPrk+kch1MUTrmqxWXlaK/Bkj
o31cLOHDPIth5wfO30azsnWAJWCaTITZ1Yz/EuT4O4L29gsciqrb6GFVzmnqRJIH
ih2r/QBqQnNVPRchZn4crJ2/xACr9QVZh1qdd2whV06XbWGF29bAZtZOO5nY9IGK
5Cj/v7n8WPDyFqrSUL7kS9+aeuC/09R0N0y1q7luK4eTevF+sBrkenoMgMB8R1Do
ep6NHP1N3KW+C/a9BsRPUMzT87nU4iRKyVRQt0Sd6v46cpAdAtNLH8NRAucf4hD+
gv95lWUUFpmD7ocF+rGr1bPMCISpxABAGnWABpfycT2qM9/3lgnS3+e2e5QttmrX
tiot9Nq/7m0EQajzqmUeUAP+U8+r1A2ZrnVSL3tMIXF6nl/A5PkNnap9N2dyBsGB
WrXe8Vb4N3TSKLNS1hEH4rSdEGT1tmSzZs13TFqg7/KRbhj1yNj4AGHwAS9l+pAr
/3S0r/FQKY7Zc8LFhmYP0HADSnqhxx3Iv1NdauHE6g455TOsS01ri/NnB4FU568l
pkoLqYbzR8eW3STd4PCFj78qvEDEiQv9cdJ5tV6YVUdj9rf4IA0itXEeBfRlwGh7
vdrmk4rOX/xHfTlzUTxEzRkJ2TB10IEXBdsieLmWx8WUf0pbhISB1TEy8hBv88/9
6Q08mEKDObfXUj0yqZlunoYD5S/sPPq8TVMZNOVIjMDUPBp8SV1KN4dkcIcJiFul
1mpoyBKqaIiW44WKzlVNFKPBi7zpvDjdVd3P+weyq8Fw011rlwJP1z4xV7/9LMSX
aYNMjZl5mg5Gf9JCpMLySB3pnx8Y6zeztkS00+WWtjIXyOg3z1rcWY+CJUksYuQY
iG5h3qyONeVG5I6fvzEjBTs+G7t8Az4fjU8l7AKp/sY7et+hAjFcmWhoLBG8K3Ni
uPUzm5d5Yk1iEEhrKjeOVozidMtdWDS2hrneI2k5aRTck+1WY5+cv256Z+85wV7i
MxOdRw1zGStNBQiPelDvOLZtdn5LR8dr4kjIS0pZz05lpKGgRRnDCgIngVaorZD6
bCeJcoE8CM3Gq+BZwODpvhbR9h6xOEyWQfUBgIyVuWO6KOm3GeLJgtCNEt4bNW8r
274zePilieaAZBvRr6tmq0CCeyyjdzG4JRIObvCyiBoctVuYokZWp3RPYNxKecUB
Oa6BhNuzLCpjnhbVKXR5fKD2m1T9TeQWJMazXT7l8mL99DrBe8T4GNMIaTLrsbWk
yHWIwrJ6LAGoyw7rW/cac2FEFuJAJf2jXrUHaymLOtYFSqatX4C1CIrCmY3L9VNL
V1yH7XCX1O7NzYTN60wgfnL3mjkf9b/lkBlnw5LYrdz4D9UqExCUw9KXiyzt6Lds
y5I05XxGdsz7SI8a5Lno+ARV4Towmqtk/qV+uFg9J56lcQAhy/AQyUcDLZeR9Kg6
FLDJP1gLT5m+t8HEu/HsdPLkV4JsH7HXe6ZapSZEuhh4zoowJO+hzVx+n+beaQN2
Ur7o0toWl4EnZiI1FK3hVf+qTnlGaZbT1J/etgorZc5Heg7rQWYhzD64uNaG1iYz
/npvKPGLgxZUqV2u1mD5YAy+DpPOuyykmewxgxiSkzXGQoC7FkygOHb6t2LnEows
Xo6obIl0L3UXMk69siwlEo1xyKYgAlD649iIFsvMAbgrx0wqrGH0CAR7JfvJLkMW
1XntUoKkqTz7srCYBIwXQT2TkFoXp58kbD/md9Q3Re91/nFTYmQHga1261aH0uLO
fE8d1aLgyyttRBXPCTrUV6oMv9tcDhAV12VJHHVr9drEGtikFPppRy2nKFahJnrn
5FJL6BwzDlqSD8A/kfOit1NqClIOu/gUF5FXm7bYTORyj9pN2efjxhq+robv7zFE
kUx1XbIOmtGvcAQ+OvLIJjjI44bp4MbpPjgO2/AgSyRNsKS49shaWD/u4MtrolHE
08T0Lg/lkA01bVIGU0dVwP5JWXMC1wp5k+crTyVOhI7RTZyZBtJxdJapYVud8Y7i
sHVIwL5kt2ZqODykbn+9wsXl/pg4zkK/OSwcbTeCbinsSeGUlL/7ZEvq2fsvWjS4
avH5Em01zreuNim+fLDVRSEuN5Krqh6kJskghZ8e3aSFCaOp7aDFqlpCtWxrEtVs
OIu7A12CPSgvJWkRrH7+XvYBr6ChumjR+fqpaIv9GADjqnEB0E9QjO7oCLL5I0Sf
oKNo9u7y/vq52bvoeBhJ9P+zI5dR5iJZ39hT2TrLMo1FT6GT/guV68zvuNOsCz0Z
aAaJIfFLKhr0bQnPQoykraLAWJPYAPQ9JT9UjGvmOgUsrOKJvdvFJc2UN3J4ER75
jdAVfeecDkkjp1eMu+SVlUJ8DtLo846e38WDNBDsrMI30fnVAqOgMCCT4/HmAM/w
VO2FlcQ54t2wDztRExsQhNx2Ubg3TtWxVMeck1vEueNhXCPkxJIdK33mx9NigaTM
gKs2Aze3BMG5oCYTD77Re5CiN8Ffnld27VLd0IADwK40Yx0pWm2swPftbeOmYXi1
oB20xArGebAyDnIox/QQkos9zOpMMCkCtJ/BEshTn2QN3UxcqcRwFdhGYUOk8BYI
FDL8eZXvjOxS7AgBu4I6ebtgDDeu2qPt2y+L1+mKwcOCnQcy6UDvxRR/RtmkZopX
aIvU9pz/oo9vSnlCjuC0gfmN8vxiFshuZikSmTw4Khgw3koTnqPmdPDUjZDP0Xaf
NaVKzzHUmov7jEUAD9g6Q+SATLZHJSBn6NRjy0Psdk4bCajbwrOicXGxauTETavi
kko01egGL9b/iZ08pX0na1QW64bjvl055e9BHS2PZdShxQ/X3yeEYUAyr44yFRL0
ftjqvKcHVCkskd+5kZEV/cVkMJub0c6SzOptnzXObbv82WHGw4tzRY6OT3F3AjxE
AOvL+4qhl3cosqKs6a/PzG12uWR/14MOtQ6DKZzfB5FfhHYSd5eXNAQn9I65yHkF
9rAcgdzHstReKFGc00pzHAUt+KbzID4WgGqfUQ9QzjJMC8GFll1Hd1DsYNrussog
KGT/l3o3wOPKQIlHfVSTbkRjkBCc2aGEwfTxExZ9KMStAKgoh8CF+JLv4wIWrK0K
5qHATtuhUJunDOJFulqqvU0t+iUgQR9hqan+UmKLejsr77FuE84W1VkCIkAy6q3S
dGq/7kMbeztXp/PS7hjODqaNoNYmdSgI3+/TnBSPuRaOj+wHU/LG9KQw8yj2N//R
WzO+M1hIDp0HDWd9oVpnxEsf/uQJtHB3nt1f26SmiYz2OduiEFB4y5iCNEqa/305
KBUGJC8jqhw3w8myWWC/agRYytr/Ks6I0NfXrJE9R7hE05klIFrxvH8f7Ij6cAXy
LA2IQRdCQZTZKCVRGvQX8oXZF4aNzB3thhLQjYW9RUvOBnplc4npKAMSOU5HeXuq
mwwfV3YEXHj9Wn6JeM+hwAvmoAcfXCa0hF0Nr4e+Vvi1cpLgecoXZzH3Cki1FRaa
MuH2S0L6tjV+0dXC1CvrzlHCvbborHWivDCu4jPnibbA9w2tuXRvGiaxc5u1O98p
g8M/Z91eA87mCII/bbNAAcLiJIGV7FgHXOnuMd47Om7oTAld5A10NRSQyibU4Vuy
inwdYXSIPlvJAjGiDK3ZGyTa2KHroaEQs5pvNx0zrxW0zdsJB86XH6uVUudDWi5e
h1UllUDqkajKY5pkAPw8wv+5FrbqmN/JSVSvUSF5JyA+GwAl6f0OPxlfTVKOWOyc
khFOUWeWAaxycF7l9jusVZwMRclQXWXT4KHdBMmUVXPS8Xg9FQneARawPdMjl+IU
aDyug0Im8JEbMwMCCVRt2ACzJWkirxDHLGhmYYA4IoNHuUUGvF3hAkh5a1Ydoffw
kiG3dUoDurLYzdgCQhNWAv3M42Kk6e46Ee+xE1RTuOKH3Whq38HUkDeKcxfjh86F
fT0P0Go6De0HLRQJF4hfx/0vR+4aNWijqQ3BF+A7YenlLJECxicrQOEqPDmNmyMl
extgEaZ2zQxCSe1ptUU+iHq1DES9m73FuHjayNCJuT3+jn8tzuuAxwJKykgmooMt
ALpNWqlNpHSypbYnQoyrl/NuIm2tLutk7xzWaiPlMjfvFJowkXX4mZXzVWX77tei
maxNHux4IhfGrm/eGssoXE5qyD7p5NYHsRSqhtf1VPLo9/CdWlOu3Ze31u3kMe1H
Ant8hyBfUh8SZCKZjWJyVZH+3Abne6PfSwMAsUfuElIR02aRf2LZ1oXOWHkJbUAd
5s9zWRmF1S1ToKwxNNKqkJdsBtaOfpPxF8tw1dKmlLZML3ZVm5fawDcj7GK1cwLS
inY4cfitEO4EA6AqUUjgQIaFNrJXuJPNcSJBxnkfukQnlXHh+CXT/+nF1w0OzIAa
8FO3DzUWlZY3ANdLM9LgREd5bfqXNqU8Nn2dEFqGDVYJ/5zf8C/2UXwc/ZyaJvGE
y5CgaD2MM5HbHullUIzW5u68ef9SA9VZAxhg6Xn3LHELuIiFisiwJaQdtHHayEoW
p5IcIPzbHHbvnM2PT9O0fN6A8r1BLtMGMmlhxVLcjmcyJCV/E/eywaB/iRvEvYwy
UeEr+cCnOVLBwNk4hZ4XQ5cG31j3snQFkgOmMPdECjms2e144dyZ5oTfitm7/tWw
uC3iaR3fOoWF6Nv7YnnMGV6uf1pGuHDWSDDps+MF18fDBzBMcKDOSiBzaVzx61oN
yzUgaGUcK2vlD/AjF0c/4ZdNC3veqtEAxIfm5OufQZNNm73TRRewCzu9wrI/yAit
qRQGVCzzitGHKweP+W5Xgxs7OsRTi9aTK50ZKMtLlXU7XoFqT+/HiRuBDFUTkhMo
L5cXdh9IZMoly0By6p0Godaj1TEg8GvG1xFcCxUXoH4UnNUCsKwDvLp9oKOCliOi
R7nwJSx9wzvgK8TymOWNfa9JzJziBrB2GPe2E/3H+51KAlTcIx8XzfvVAZGDJmtm
/qEMFP+Zgt3H6N4B+0iOgDp+lzefHwVOEnuOKnTqm5N7Z/aAMoiwt3xV67/oz6IF
CXMBaHbuhzirN4diD8t/Nf6eZj5zoJgK26Qkd4GQwa8Tu/R5tj+lAI4ybkoFTmqJ
UekD94ALztPDYNq/WNYR6eRDrGFKkj/yaTx0j0nV3+Ywf/GZ9RNpVkLH3lPFMebY
ZQVfT5x+1kmajp5/T1AoBeUQfLwFUQCdbz4LKdlLGDKmEXTjJkD84+j9saJML2iS
YRPLT95E5LYaCRn+RwHsClBJCgafaI/2dM0W+4xOX7oaGHE/Vxz2r57YI5xkGUdo
zs3zAKvssoHoCX5oxhwLraHDb9J8qo4f380sANVUzQBqbd6yeQkmBLiBwWEJfn2x
NuhyWFyZe4LxWE5JVFZ4UGkSg264JPI2iw5sxMLlTvp6lcz5yP+ZHjG1RINIze7w
NX4YxP2R92Mx4oefcMf48E+wpVMRFyQz6pcDxJfBNWtHpkJgtDyh9qROjL9Qbtg7
IZAw+jsWFOflqhFZT/RfyugtP+bHbyohnrTb36aHYSSEn/Am8o93zlUhunmvd3y3
RqJWMtxVvfyySoxcLODMif63AyuCOsritO42sy455ROqPlZjGyG1vdVXq8vENPBe
rR20CiVs5oeB7vSW4mEqlcZr+dK90pyoR4nloJBbt3gJRxNGDQ/mtpC/5IyVT0ej
Hx61icPmt3lHK4FpxzjDxrgCTkKlLMEsL44Q406Rl4wjEzSMLzWW3bzD8nNKvNyB
QKiwdSaxW+WWYiAWhvInKijwYHtK3ZdS1xQkrsD/yjvZDNrs7y/rQQJkvOgzY1bz
IOIfLJjgS9wHTXUGAWAQqrzaFaZhlW+rAJwKWc9LnSxPoH0Zefscmy7r6ztKLiYF
VWtGOSyDCxqNgYiPXQuZZWIO0uhwzgBquXJjUb4ZzEdo/a+uw59ez+aihuVheyY4
LR6CFOvGqkld1b6DV1AvmLnacUscz3+anQzm3QYkurvVoWI/608Q0yd4BSzSDChH
zwqyOfa9MP0lfDIS+o0TkkCrQuMW/aMp4wZnoqU46NMkah0vvrMo/y63uIJ3EEQY
+yJU5MWF1IUgWhkDNkbtq6NtV3janOAxAzA736ECAHVvfZtHSiojry43jL0PaAkI
lb++MYRfsheijd2yXgRv8NFiKWfpreGFnyJaMwo4YsVljNFNSawaAKXx53c6r5J1
VFbuKXjHV94HjEsGrxYsNIAZaqwWqyaBit6xJKgK/KnrU54j8RGqiy/o8WFkLN0H
CUf6PzfNKUVOz4TFQGlpn+9G1HnDnbM+5WwcIGgFwqcx/rcLJoXl0qbIxHqDJzMS
8ciA9RZWY7DI9ZYA3r0svCes/fo7oSe7LSnhldrxl4dXO7nQ5mUe9a3f2Kfl2g2A
INERA2pYmDK3DAqFmtzSlXu1wwtzgfliwzg/630jbNaFHiOXXOY1By2wgXzaIJHk
i1iT6g1y2AAJFT78N2romjAslXO2MsJ0Erx/Rg5SzdjhcI8HEQHFo9sGkkztUi/Y
wAZYsI6pjuMbyZiibBwlpTyA7FCKkYWn41+gQSYwFlS82XGcOT3eOROXYYy6ZC0s
ud+HD1MuC3pmSuwUUsHeT54yobudWgBK9nhUF1FuGcnSYoNEvCc+sbpUbr1BDjo4
A9vUvHvtXTx0tbH9k+Q6PyYY8XryXG6nc5/d/32+ztozUwAo+57DzeRV2TA/n+Nb
wQcS4f5lrWPguDsMc+AOpFijGVTuM2nxEcX9OuifcVM1nY2nXF4VnP60MHC00mlp
KIJjIhoKvwE1Is8m07YVvX7H+qTizoF/tDqYRuVlZA67/r1muUCuoLqPzqlbeliP
Sr44HpqSvlpYAsiOTpaEFOYSExY8YVhtDOdIky3vDcYqC9wAB48vVHZOuecZi7Ru
R03qQM2w0AyBXi8Z/FzR+7VMhCu9zuExbbVwQRgIFWMnZOZ6tA2TCyxdHCy+VvFF
b0rD25Nm1UIXJ3WzxP0YTNi25fVIktkox/lOuS8LOC1R18xNmJ6T8DVinRYNdSvR
W050UAceaeS+xrT80nY30B2vl7DDV37V0F+9sTyaSS1YhSNppoZAvlW1P+4BvW6J
XWhDOQYdUp1ZFCM/HXemgy5EUcCgapg0JiKDMGlRax61sLIjjVwyhz+PbsfpbAW1
tyPsImOL8e1MLSswUn2euCO4oBcZBFoe/sZu8GMmj76kWwA8UCw2Si+uUpywIGM/
bgo9VsUCg2iTkfODacsqmSaklwXf0MWmY/LBRjsSFeqAqC7IdhnJSSbNyNyVQDoJ
8rj5VTy+RNxZQQ5xjl3Eadk2dObSwxW30/VPDKSACXf7C0WJqPepQ7h11z1KksBM
nBvt1vvq5wxQD5osYRhhyPSvEL1jo6KGQhecguFrrhDIL3pWr3g3WmYZxl2ih0Dr
QljfeN7Nwl2GlPetUSHgukCecJzQVVun/0yAenj/nRLmFYSEZ5WerRaEaadgneHc
ziXkhaqezR0Hin0BQCaJkb41UOO47RLPc0q9944Ik6lsiPjWY5zLC2GJsH2K0Wgp
nadgGHt5zu5DCRXWFK6z51qKlSSnF4jvYnRzNl7BODFcbJL5MwUufgN+3ETa+F1O
HYsl02cgyEDF04oiFiAr3JliZH1jaJJK11l1Xy5nIJ/KF5oTMK6Sea9QKT21oen5
wX6OSAynKRG3eD9CVpTt7fU1Shx0hrVEhoN9n7TutygKfYViE6J5hrn04MlkPhMz
YulVxOfJYQDJizZLS8YwnoiCUEFCjZbqsRznPWDIRUG3bM1LLT1WMG5KYtwq1MkE
tYEX5cVtlZ8DMtjdTH7NQ3bgZb0AYLdefEo78sR5kJDiJYB1+hvcZXaVyimH/FYD
/ZT8OwbESMU3TcDx1vEgWh1CEYOHSRGW205z1xT6CWTES8iomaABg6lRTkf0nVAW
RncaLNzz1zkxxpAr+A0VhDuJd+z0PFTDkNwmYcssX65HtbQ1MYgcIIqFdb+qwWOB
umJkdKTN126+496xS18gF9bPCP0OziK7bkDW34M7xIE04+48zpP6F+EehIEcoDmV
VT4yjw1SUJPeTTbJ9RI1bhUCPGBSyr7alB9RfD83NdFQvHjpK3cNvlqekgr/fwYL
36CuKsX0MrITB34XpY9dFu5u98yg6IswT+ijBbE6a5aMWMVloTvZxJ5jlLfNvevp
GpHwKh62sjexTAGfDaUqxVzQR/kFlGkrskf49fTpyTLPay5WT6vFKL/wwJyzrxWx
WMfI0x9CUbQ25/VvLBjDHW04dU7W/LFafHl9qX5JcokOTtaB1eTC/J5mh6/1WWlg
jbcowXt+bI739n8DSxUlkEZ/WcXXcC/jRFwmd4CCMbtaR1VUjEEfnYbtUBRviBGw
kvbSvkj91ubSIISfTOYUL3THp9bS49h/Gu/nToCSuAJzen+hi8y1Ai/uOdDw+zEN
gHPjfzYOSrB/bsfuVgr0kgWDFglaiUfw+jluLE6IwFKqO8KyB90kPWEuGwDl/Xaa
o5tzvSY6hRkkRWtYp3Taxp9+QwPRcYf8LWaol1s9Oh7UviJT9Ya0B+4hMHJknvfD
g62fY4hVjMhlh5rGubuDnVa/3fUaMRgz5D+AkRTQ5YUJwsctqiG2PcAd4rT0YIYL
8OnG0EPHuy/Qer+IDjynTaGpcikolLz4JgV31psC4p6uNWnDKp4c3emtmXm3eHXD
g7tL2xlD90+mOnbeJyiPBOTWygYS3TgyqkmR19dItqR3xIADRaKGQF8bQPWvfwo+
3RrMkvSOYbVCHukQkpBTaKLqGQZJK8rCWhNzf4cHyp3DgHUhL+Ouk4Ou/2vOdWN2
kpKOmWzxv2gfq5N63CSgchbI5cArCEf3BPZAvxBWLjTPyZ5UB6mwCpfoWiiySvcG
izC2xoX2c47HqbbaGAGpUt3fcKawMfwghUzKZwFzJNHqtSkso9L3gsDLKVKcEYQI
sHYvdSg6LkxnzeEzAwaHifJ5iuuOBeQQEawlyJaa53tob/YYj4M+XLF7sRWBv8L7
Qn8eHq7/NXFW5irh6jV0rXwIc97hMbSD3G9qdHiQT+ObTV1mS/DiHD2/WIPyUU7d
rUL0RgiaqFEdoaOwzperpaWXwh0/wZVi0ZqSnASu2l2d1qGuEdHBsnVnXKX4yUmc
zv42LVGLv7i/cb4l4m4VjLtGUO0xQukqZ3MyUum5XMrMZ1+8lVc/9hPKdHD54NxD
0FGY6UWYcd4dnGIHmr1PsDWHrgxUOzWItmje0LGyjWIVxKIB3PMQAlT7B9D6XXgD
uHQCFspmbmCySSBvcZiK6kmb8MUoSN2zPCGK8vyySL+M+gMn01AErGn8Y4+WhWan
pQeauf9JhVUMJsnQgjg6qCU332BfnBi7EGTeUkPsDhbOo3pr74v8TTcvUips3Pnu
zEKCTm0Y9Z3mmTm0WThfIdUTFjQTVxM/omjMIzLAxBAx4pbdlQncvqunuwNsEIbW
9a7M0qa5EDh8y4CHgqc40piRLwDdGckBRAM8Rg1CwOnB+BHGSO8gdeTuw3SS0oAl
heURSBJmUA0BxLqqx5DxIptovDYa5qt26s3XL+WL97aIPWu8AAOt9fD3AA3K9yjo
O45tiZZjRwI/bknwh9y03j6JyHgSsw+86SbpeOtaHvS2KkEpi5ipMd0UoriEfxBU
xsUMn85QOgZ9rvcRRNpyK1Uw5JCgjfuYMwWsAPUnY52K5YN7IVBo5yGWIwA7VWVk
1hN/y4FZEVIysqAYhrdOZICfk9hY8Otf+Pz+OWo6tBfnmu0ml5RzSHh1f0EKlVu7
ssmUJypNxO6k4rNeQMDH9+ZX382Gmr8jgPvxH1yMkDJGkTclRS0HpeklMAbSM2/5
3pxDcbySAEFsq3VuPLrjxM7RAvGjrk8oMrtUnHd0NMjs3bi0XasCelqLbQsCWl37
MyoarZ9DoVEKs9ka61jc5GOVVas5r2twXmZdSic0ISihFES17FCe+WXs6J345EiV
r+cbm7BprV5RV20gjeXpeqPTJ937SNtMIFIZorNoPBTRC5zHTJblLF7/coDsBdMb
KAPOpFrfRyT853xDMTEqoIFb/PcOdrYLsVqGINmdTloOz8PyJhC0r0eLteBqhypV
1rPz45pYVP66/qf9F+shiCYWj+JCzMIWLltKCZ7Xz9+V91BGbo5xjM/7GuUZmj2C
XWZENUOZBQMOycs0bnHt1JfDd04ZBiN53T0G5NdaxU203fspIHFrNdaDGrJb3tq5
eVR64D4X0VE2A8fTzx0sjQvtOezqkWZNQlFP7863BB5B2JNtVy0fLAT3xHKgaTJc
W1IBxU4f2S6U/SBnNald3N0IAX6QqaVtwl/lU/4H+SJnJNHzLo1BwQ7pTtcYguYk
iMI83Ef+QqwefW4j6vZheQsQ0BQGzPBpXeC+wgRcB+7ZJ1XatwS2MzfjwUARY4c0
gDl6JYNjNq0BQAPQlSYi5/o0/0Vi3gV7kvUL5jgnI0Zu5+oQqNL6FqHMGiEFTiXc
YFxguAJMBUee/RZETEUfWEtnJlspPSrjnFisrsLQE4WRaMp8qWDfXR/o2DAFjJBj
7Q73ZHKDQwnTBU4ci6NuLNcUjFsYI3Jw+71oJverEAiZGf06EX9ihWQeMtOhSOoX
0c9dM9coaO40c2iE5zDhRTUy9bE66EQr0XLB4ctliqCvRHUjO2Pul6AJ7TRZLGLH
2eMs40W8yP2V/3nR5uvtHxNPlzxPJ0pgoau7Ks6jZLZ/i9tGL2dWu/2V7G8qfPzP
b8801HW1rRIHuXpD9Gd4J6cixgTu8kSqKl+X0DWuS9N++I3R5CkqotR4nrs+9kjm
FU4AmChs9Qb2KhYrERx3QpSMX3q08reWM8IMhqQUH69V8JGs1cWiasm/eLi7XKf6
WZtMZF324+9wnnLOKfYZdNAAwQRvyYwrh43LMsQUAtb7cCHZ1l+4FgIFOv910kJ4
tKe1s3tajgK07w/uLmGPKmrsUsoIQoFpD446osEq0xVs6YPR8fUjAY+dP2MjPVpK
/LPxE7WIAJADq9zB12E/5QsBEyfu6aqsh3IUD+XCOXcmaDTtKe/ouvk4Z5gwfFPE
c+SifjKO25LhnDJ+xnlD8x5Rmkxv51WAXxhuTUlJ24Gi4ZGYaOi+RM0hKPcnjcf6
OCe7H6BWZ8zGCeSDSFOZZ6f4Q3NTAHSWt7MNsJM+I7toYYw9NU423Ez3M7JxXfS9
mn+3eSL5jH0KPrYzyOa9SMEV9NgM1ad9Po44kwkaMLd4z67PAdxFO+sE5MZdf4WZ
/1xSKRAgfghelLcs4Bmrp9M07wqltzlqC2OFNNhzfKzbs3WpU0qV2MyHtXdemrUU
8tSkp0/5oX3mF+hqurVZLLbuqyjaG9kRYBcDkzwcranernjjJqTmHhY2QDe0RYWr
QSnwQ4Wznai0m/DoPl0uNGcy6+Du04J41DxvurdynOVrlV3Dftsqq5rH6P/GM5z5
BYsOJtAGKxEhOjVu9/TOPx/edPNzc2n4Yf1pnF+82I4jPB+0kBDIa7Hs6sCMnqzv
lTBX9pSrAVP4T0A0lSwO8ooCEdBibzocvk0Kd4R8MIcQq6KX0coaA5Uo0hUaK4T0
C2iUmxYp81jxNnk1H9CwHV+NYip18brHScBLhKyaTZ656CHjp+psAsxt/lsAEc7K
1f+miTvaaEcYEX2t6GWz3D3dWEfUPdqNSDf78mggud1JtSD7iEdkEN+SCSgomN/K
yNjaWO2jD+GgEXstoS7gMlQ/hFVTLd0oZCR4mvRH6BJsdGVXjVJV51eGqBLs8Jjg
VduB7bGyIdITrKuVUPFzl1exRs2Dx3BuBifKQmEIFi9nQvgYhNNg6nWxQx8tTLn6
zYY9aW+uMIEAUjIKaAFu2qAuQ6tbBWw3ri7ddnecHtgaFP+XQXfNQo4Jk6S12GYR
ABGkfENKxY+qHUW5cqW/ee9BOex+TUpwXV9l6lA/kmCxH/EO4h7xoa+ThUeg3EIi
ALBN6UrDLQ3oGJWiWSGXnt4HLfObclBrbrqRt5DKNGjuLxQX0Wp1UQ0qujywWxUs
20hwvxcbyIAZNVWAMysZN3Vr5NFhPPsoT7T9tdLYF7GxRRsYPhC2bBqAjhwxZRXD
eyU7lK/trik/P1hYqCDRt1+WAtJr9ndi9Ud5CbrRmMQRHHoLPIosdFoTLwMfrwgm
8T/bIxxZtqru3ihecY1sV2/XzY8296OCrRs5oUsuy4GObbiu+wYD5vDig/0Zvvei
TF6uE2zrRuYjVvMsRS693c/pU9yeK6M+TvFyrQjuZDwhvmGeRNGFv4p60qpJaeJ3
K9x8ZT7zxLi7ne/Av8fbCbPsJe7Yku89pBviXsI+QzaITi5DoSyFFVSUK7dASMJ7
XhK1brHb+5lzxfMAKhehICRF475e3gaUFNPCxhU6NuKYemiXWoV48c7ITeQIkqLV
ZVS02poV73Q9yRIIGYxs+99IzDYjqktt++AC2UokeYUA8vTYmLRsgmpSlP55sghr
Xr6rrk9TqmnQ1kFg7fusMpCGG6Tyu3mRBGWl/ZuGUd8dPLR+9TRfv9WT4IxNJSXr
aXnasyH+H8BY9K2YW7SYjjt8aIHmhqN9x4AlEzZp087tYXMO/1h0kvGS/GTY/yx9
2ZFiPPQaU3+3Izpzde8dtxMooIW3GJd/cu0mTeYkxEMzdUvZmmDrb99CZaQwXRxR
5gYlLdh52oDAHCbVAKMi2rY+PKZGukSto+bzC0zN3hmkeBLHXuP6dMMx2PfePvnt
ZD0CFhjunZ/3x0CtaNwzryQmYJ0YpiUyk85FzK7dr5XUmO/pbYLdLxPFzpn92+HB
z67cmq0BV6zVpbo8VpftomsrqySc3SgA6Ysh3Lqu3EgPZholkakr3L91c5uyFlw2
rQOf4VMyk3Ugyiu3oSzZly0BaPMp+VBsqyNBcWJoWXu6t8ZdfMrFmLYGO9JZKx3p
vkeklZa98XH9hevxZNDVFqMs3XA2a1B75tWFQdayCAyFs3omVDK2lIbYRylPRK9v
4ZtxjywJXEmc8vuhvf8ChCaeLg705SRI/1zxQ+77ZQXfROs+6U4KQOVI0v3c7+2A
M+QhPn0F8f5tXkXE8ENBxX7OCoNuQiBBIimbO4f7tVsy1nJMgm8H9Qdj5QMp85UK
sp3xFbKBXzZJ+TV2hCbkciNFzwgRQ4nPkoj6IK/i4tejZse4SXiSIopB6Hj2GDpf
yfIjRT8zyXJ+pvuFs99wK2K+ra4mPRLTp9cVPlT9ofxeKtup4b+5vAKJJte8L/iW
2CpFdTHBvVdBRxxNl11NPavBiNRwn/hp8SNZoWIxrOZSh2Sxu9kzhbopL7FpO+bL
111dvJ/YshckG++IMsN5ytuGhu0Gi2usKvptibTl08Z3uXlQYvBFE/Jzhc3yQEAf
NvxCZKnVcS66fWvzzh5NyREFmZtRk/3ZoKPUp0ueB7P4qwSYaU6Pa/hiJ9PhIqsX
mYwa+PRVa1n4Sbo4Nzqe+4wcDSu1/vVG84rlDiEuZdwQztZNO0tObuezxxNFvEMa
ZqPhgPNjWc1pX5ay0ziRFMhy5ZzEhEZP2fftwegsMWGiMYCd/skk9cAIlO5c5Y4c
GORBkGpf/ZwklrrcUIv6ixUsM+MUHjTIKYGmKTNkejxNVDCeRde52t0tzVzpg+ph
BFTOWiOUaPghKhycbfBkHuT0hYqCGdzXDxM5nQM3xg5+7lCSIqr6KPE1JNspZN0g
YoeVeF7iHKS6mJ0C20KJ6SJwm9Im53n0eecn6wIc3r6fcbysr7f9XYxxaYDO8hyJ
nfiN+ZH0SgnRNrAhCUlYzHcviYk9ctX8khSCH/JmgEG44VauZXkuox5vfOU9FcIh
X/CP2NQIQVIK4WT4TvlFmVl+GIikgzhEpWVg7GpchTb6Q8Z7XS3RWVXWXaSYKePm
j8D8F2JKPQZ/FywtA+4xvvXlUkBUIPG5fXEjXs2+eoSvF6Uc7Ai0hoW3QRR8metR
bF8xP39ORnU0wiKU199PgoVt0VjML+VKI5yCneEVdfPIvAQmFcSwX3SIljaBRHlI
GM7kDSTxcEF0t6mvQ/7DW5OIyt3tUo5froQH/XGmKbLdN26X5XSOdl9CujVBTVDe
68MKgQsAIchmPWAa5ik3Fh0o1RjXAUKo/TaNdWcT9Mv4UtY/aFU23DHCTabLkQPx
CiyDDriqyjxk1vf7DNygf9+UrkvA2nPSRxtyz7LMD0h0Dlq8jODTs99pmAm2wZyt
z29qKgDOSIX/rz/F/TUlZEG2+Vj6gl+/FtZdmfe9QlX5NMTvI5ouBCv57blDIL/J
JwKVOixAFv8cNjJMk9EQuJwrUIDe23tRMu4X2v9lQ3mFV3X9R79BwO/8QUcSTx4P
gxX1fuVkq8PXb0oFGms1gRThBVAEeT97sZ4ygfG77g0f2J/cA4ZRNdL4OLpzgZ56
V27ybe64a2D0MB8oDv5ampr0UKoyWIQpzolWWybmYgNU05PpMQ1rNeN6p2LQ5Bjt
fNirPoYYF9WTqFi9odMy58D/vYFxHGr+ZeVq59T6bR9DByhl+bOjEYeyczbqDYW6
YZaD2BCV/2fD99+kmM0PaGIYIaNLqqEvbX9/Y54q5D3ACt6RVe0NKgU0oLPXqdCf
RYVShgLuyWyrKNincWNqnFSuzRbn6UAOBuJrb1nSVCQ+jvMcsn8p8kOgstsTKiHQ
cmuayTtfQGAosNQFASmEGqjC0natfl24/Rwr+83sFFVyJQ0/S8PA6bhvpLyGYmiL
Bf76NuxLRXKuFHWPSBL2dZj8vP015Pnp1fwXSeXiHR0pzYsn0DufOFjjJlD7gXtL
8GqrO95p9L4ZEi2Fsf5kWARDdt4W3pnZXf3Lgf0libBVbIaZOrqQmgdKvBgmy1r+
6roruiYWr7o18GxFJ9pCOltYH3wC9o9CXAzIcGD+7BVid9+GgTGu7zqJ4R1PCXc3
8w6/FD/FQOlxbNtcwm7uZZRFqR0D9SixAHD5UwWQyrzw6wEEPPA6nTJ6o62mHEo4
+LALW9UNz6xgVGBe5thPeSJPkenP+mL5QED3iljFG2ehThnm+dB137xUvbroNZaB
Ai8MwOIZmaNi+pbQyy6omOdki8AmyRJBOBVhe1ZliLvhoLid901JX21UD8RYoM3p
th7kV7O5MMFVqnEcbYPtrviFDtyMcmzNTjCcdl5EauWVSx2JKzvPbKYp30iaERpq
9SOlWewHAF7B4t+34SsMwg0Uv1EvkTu6aqc8RX80aYzxUiDgKzlkjpgwY68bx0zq
rZk1YAbCGjylhrBEXxFKKiPW71j+SRnu8aostpcT/PX5vpxrhNMhT8t4ziWkxO3Q
AkueTNvy0PArNdEzltvkiTPX6zpE9lJAbwLfIfh5ia7F7Ba5QCaJJluDf0pnyUeB
NjTLl8jzNKpgOKop2g6wPRKfuz4AbbuG3HM3z4JGPcIejcJSQwvch9C+GG1/je9x
ugNnkcQXk/GPlfwHeHt4lsSXy7r/uMpzO6hQY2GxKDBso8YUVDbCdQb43JAagc/V
M8Wu0QoJHAu8DE1EJ8QFbCwMjTm647lWAju/1dCIs+vP016NfNnFDr4VNdOh4gQE
vl5DQRi0/aP3Rjgkp5vGOgDz11GFOCg4KWsYUi4ieU0iMBX00zfEEHzJ/g9y30As
2bki2C5g6QMGc2ZTuuaWPKcG17HX5bfDcXWRmemDmPLmNf2fP0i2sbYgaKcI48Gl
UNDpM3ggc6nkKOI6WjpMbBMgS+ZE0ZTqOt6BpkEgIsGx8CmH//jSJBj/Itz3W+/5
1T70ZVpfi9G4urTJoqkJXIDcs2iKaCHipgvv20zLLPk6EL1qx4YeDVQus+7bias8
Ao0wLpfmI1vhzFZ6RVa/stK4enYpEIyyANOrO26fX5Ww/xNLm555SOnrn77RhWcs
kbPlWTGdqzpftatZW6+nB5bPoD9HCxaDOAK2sk9W6bnvpDhCUfmpyUef5Pn/Lt9z
1Osl8RXb1x94Laxp3/g5M4Ohqe7rQYI90HA0wwPPNExvKNmyz3pamLcAgKDYLOEI
878rJmjaScYHBcp61SE4CjjC69BPETZBGFRqnyTm/J9nvMVuZzcdgLy+vnXfC8PP
xR33/gWB5g81ATvV4o/l5GqTwIjdg/Y5qzPiitr5kr37kvW1d2niKRyV+gGxfnyc
fmoI11fgaqYp6LnucFHBhMuMXkOjohJroG/Tuqqy+VZe2opAFfvhclqr67APF9rA
lFQ/8G8AQ7aqD40pGkmYuJerhYD5VuEaRlHD25RUzkLOdNtBT4tLGs6oSrTpwQG/
8M+5xaXqQk6/tYzIPiV5X8yiVWr82A9hzLtFNltfqNZDwSPtcdDS9La8sCSdshkw
lSmEKkIkfZbD2fhdi2wv+1aAeqq2VyDKDDW698POhvWnltrLxt50aoLY7H3OkYIQ
DtBP/rarf2xpVhi4ISBQIoNvrfn7BdQlgsblIKxro2Xea1aRgyPjTBoHMjSrn+pl
bhe9vrlX6wwGux8Zh7zvlag+exeY0WIKG20FczZ648jry03MTr1w/WW3WFY92ETF
TqbGdvbZRtwoGrLqsnoNx99yUBh2x4T1FDpVWABzNbJ206NSDyRk5RUlRCQHxz1l
cFyG6sQeqyn9dNAnXxFaKvL4jT3xN+l9Fi8hLY8vT1oa1SAFBs7d4anD/89hQoi8
ppOuxMVDUMyksfDArzuiLCU7eceekfT3PfSaZrAAVmL5lLKNrxNNrKfGYyx74rRZ
DtmFiVue5m6y2Ex3Iepq3rNB/RNdQTdzp+sM4kjcY5XhvUz1fZw5UBZ1FxV+gY4Y
bsAnJXj46gWZ9v0lDjLctL4KuvaOkQBgaUxpkOAbjiCtEPf4we2D8lp4ALMXCj8/
04dIvzA3iTfvrCa1HS1/5MQV+llcPuDDDGc6uxi8xY3fMUQ5r4mJzv5bV9ntnVVz
95WW1Ooy2dDpJX3dW9bCK0wzlIShPRTIfdjjxcT12+Zt4SYUtdT6m4WNenoFLTof
p6tO0v7vRlq40b9iQpWbjuZ2kwcUYHikZVCEUaKibcFAj42uqvzPUmmFofie3v3d
cB61X8kVP6VEa745rSUEBrMG0JBMaYPQvLO5gTMtVyuqEf6vZSI7YEm/FyovgmKU
cMfO5lxu4YygnAyvKoW37tvVJn+hGure3wqq61cN3XfPueTr3DGTKi4bYoiwNOFx
uP3LbLQqr0FFVufX3FCy7Guq68/QIWHFQk70oyYDdZTjQrKAzesj+gQtHO4nVe1K
18tZ2vSCMKJcu0UqS8B8l1dVLt9QJ6mjZEmeRuG4chmHGligQ48QegS5ou1QWNAU
Q5X/zsXVLDyfBFBPUgup5Hm/LnUQ3OHK3GrMpO2RzXmEI7zzDuiyXOmEIkIjcMrH
hUerlIzPqvg/zgJI87z6zkIspO1IJY+9MMMOLOuLIOv119cgtX1y437HQVAgC8RL
OFouFtBzB2jvq4FkJmJxjyvgLN/OGZDg8ZZ2INNvn3wyETyoRyHFrnpTmxl10joU
WJztn9ow4pNjChEg5pXmPtl4KIPi2TUne6M5n5tYP/uetxfz6BGMPJW/0zlNnL4m
iLFyjzTUdzWML4e4qUdNNAdOcL3u4lsncREM2iJCh56oDIjmULSYX81p6pG1l4q5
DLJecqhlnSRkj58c3ypqnuiRBOR5Oe09DFBrpje0jwu4+LHtpfNci3kffMq2p1Qh
2mvHTS+Did/ft+hl2rYIr6YSyEXs9TizWcjo7n6K9GsvNyklDF+6LIZuqdOaJsqR
YgQ+A38wqLFf7Dc6gwNXlQ/7InncWufYdl/ky8Hbrioykdl/j0muga0oDBpQCi5Z
DlAabMCZLNZXPHxagHW2I7W6hGNt/P7fks8K11eYkh/kHj52hmB6effZoVCORHHy
B5oEPSlyN2dGP67+VULU28ajf4xKqGRcd3uKKSQJVtIsp3O92wLtxJmHTKHKNj/W
BA0dxW9Haq8UFkgL8DYx039PZ6Lr8sBYKUSXXU1wFsrggEnlA1kwRFfEdkkJiomg
3/HvuuFj2VbwV5LFMoa42LWYEkN4mMsUmCn4TEaEYJBMKOcQQeqlm75OvB/Kgvc8
181t89w82O1/K/8m6IyF01MGP+U4lMA1vYKURR75mXbcO1F3IBEtJ2R0hbMuSeqD
PYdmUaSPAfedT+w75Wm7Ntp8Xy1meI/lc75rufYfLNw++C/DU3fszZsxHR9vF0FS
W+JDTEmToOI3ck3OZAuXTidaAh3Zh77M+CGmTdGiAvZBfF8EOwoqDCp53pZEs+gJ
M4mY5//NNZ3ksH2FfYEAg0Rrc9o1TrbGEJ4kz1Vjsf73FDDjM8atZuQGBC/A6l3n
9FQJmvWus0nvXcCk6mnSky+O+jEP2Af9xtVDrisMk7Zf3Ey5Dm+4orrrg7ipDdPw
7zVYtJYM2ULrrlEymYQ+WVYAd9fNGDMwtLEFumhSeiom2E//qpQJ2Yehf9nnxp7Y
2OmU+O/hxlxdGBiEnq8AEvzuBo84lOiAT4V4u/FNpycros1eyey3ELo61VYvWeU5
UYI1algXTm+RcKH0pXQG8ViyFEyRMJHQoVUxbkQ5+WdLXtGjJ0NMHHjNSUBhlQhH
x42dvR0icicybRq+wBvNUFopSRn4fjOBUAQHSvQiwH3jDAp1D+/FJrjuN+Bv5QEP
3n9WFAkywjuEAvEFiwZdDP4JRCtTwTpoiAugo04lFnqNJ/se/4hSXbl9QxoLbCaE
Ml9FGa+KXrzCDpG0ZZ1OoYFd2VQG4P7RffdQuy1bLuC+1JosX5uVOF6YNQMdGJpd
WLnWS0dMe1Hv9l/St5ZIpLYK4iSNXq9gRF6nbi4bICrZd30VFq6PH0e/6Hmt+t28
M93pRhmHHrADHuwj3MDYd2FFt+b3OmXEDJ5KDP9rw1AG0oekQcSh/oIjgD9oJPMB
7gsh9uSDVE76hsbo8k6SrqrglbbHq/2iRjWdE72O8evEIbbof5xU2lhu/i12kyws
E0rcAuyHpr5RkQ7g2VZioNb0ajbpslg/TZykJ4wkbbtWnGaxwnNSih6Ncp2xnFER
8jsdosRRscFIosnKjwKogoyNB0JT6XigoRBWlIQya5y6wh9fzcSxsASFDi7H+w8Y
HKsmtEkoVmvP5QGpo+LJ1KBwFYcPEwdraeyCawRu4FBTzFx30bY0zUjzhSWOHRyo
nB+eEIs140MNvmqxrz1RW0HwYVZXACYV5nQAMQCzrGUim0+yIUoMHwMWCQXziYkV
jPQxuGRPQSUXydKZBk1Y49Q6xkezS1yJlJsx0QkAuLri9N6WMard7ATQX3CvJ2pr
SUNHIrJHy80YCT8UWh/oeQB4hwRxZoopAvLeRhbWoHocvKvwyjtomx4brbhY6nKb
DjwSfgzZ7cYMW7Qb+EtfGQzISAFTvnnOCrRiZHNI8xWoTYysOYMNYrwZ25ehLUTz
fuIuSU+FLA5EHZ7YJl1RpwNxuFzOVIXF/RRebmPcgt8O2iCFHzS0M9tJWbjvXgDg
1u2yCTW9zZ7/xKDoAWhuHSn3eK+1/D301Rn1RSTF7Wcug9IEg/a4bmpjqSunPmho
KMySHo+kZLHeDnjW7y4h/Gy1OLL6jNbHSkAURlOxXZeCNP7/boizNVmwGRRyv7fl
gbcdMCUsokrErUBu2RlqZhNGiWyX/SDvm7n6wrw6MG4zsFadHLQsKu7xBvLN1YJy
1g1HXoYDaz8iUDEm2pEViTsJpQCSb+F+GXlB/rr+OGmMEmGkEBPWZcdJIxS9Ql8f
v7+pJQE3DP7EudrIZ4x6I88/VQfsQMPBv3Af9ib2baZPZ/TBk0CmT2IBY1iLNCaG
5qBFTBVarGkK+blvMQJ+GQbPmURF86qOd2SwuQCryhS8b7L5LUAze6aNEymcyi6r
D+d6hixYI/NJNKhj/klCl28N+XoKYGTGRu+UJeCG3cXSxK5WU1vJaydudU1/HQgV
AbBS/d0h3YM9WvrBMD4YYGH+tQHzcPqX2jRIFZf77+K6fVMvBo7/xZUE4vdFsdNh
UwHT5H6sO8PlQLdwgR5VZy9f/dMuqheMKWoccJN6eqH1nlm0VLR0TVr0F53TUZ9B
xWbm+cgXN65sx9IZIktWYwN97V7tsTxX+BV0qZVCNvD+9Fw6YIkPYDrl3hWiaU6E
T6D5mczzXM3pq00ZXdEi0Z638aHu6+KNBQgx8/rAE99JpnXCIYjkb2cA9Ahb7rVU
YumaYUgeyMPDAmZ71ys+qN+kJQhldUNO20PPinY9X1E8dmWBQ3PM0zzU63wfq+eo
Upi70xJGjw3+KYqA46PrijxTux6qzA4BE5+knmL3nWATJR97S8qjzed9EP1kAHcn
Cgb+ZzQVFwpCvpebWhQrK18BQ0CKbWQvGhurvu0QksH6XFdeht/s75hO/X9mCJ4x
K7jqlyu0c69nrqyGLDNcWO1hOTJ8rht13kTMTo3Z+nm9DLR7C6csG/KRjVSPLZYh
VJrSS6cl55OqgnN05yctl60AkbpnVsOQJ4myKBYrMWlZmOgxbg5x6emxu+DBRLdh
sSACsEai+Guzha2uIdb0IC77rRusSH9B1eeP0HSVZRxddm9C4Dx+YiDmWOtHAM/O
3vGgxNPlvfLV7eQmVNfGamESjwkiMuWPe+374P7PPppP1iiuPkX+tJRRbFe/4U8i
pNbCCYqvforW5w2/XX+iBxqm6eYBpBisxfIwbYofSTqhkoUs82fbtcyQ0qlRoxMd
Wrx74UiHAvJHKQ9vlU/yTflA0zS+37sBVycnfLHuZ9JXX8dZMNHHUiEuoRwjKDpc
0gZHlasdiYNBcSk4LPYtF6A67KoxlpkJEu7naIl65DVMsWX2lQTquIkO5aCPuZya
79tLt+ughrx5NOXzgz93AMhB/U64763QvicRWSIUMDDJPMTdgAKDz6yN5AlUcGG6
7XI8Y2hoHJUZVmlOElczOzBoydJfRlgk4GfClEBD6DUmJbK/L5CKAB0FsQvstq2X
hoZ2oSJcxocZte1SjaRAVKQgNx4jcI8foT/d1D524a8piKXrGx0jbbXR5H8W/GAD
REu2PcY2e3B4iNaabeOj6NrJLROYV+tNWJAb16ihh7AyI5d2TBq2cbr7KYb0Y62k
SXDu3vLyYyON/ikcH/vm60vJD88lZ4HF9tjw6YxKxVzWFseLeNs3BU8cG4WITeax
LQMr7UcuOUnAJYppb6zO6VyCKwOKV5b+q937J30fdRETdXUtxwOa1wxyzAVitOM6
1ctAAI/QpcE67ijyJ2HIvmLu88RXRqN0aF0vrDs/7hW23uh4G0NQb4+KE8rkydkS
NRaKjyO8pOaqWIs4rbkTwv4cPl60o0uAO2eMhEkmluLatdT353N2LMLAFOQTIg37
ipaU1SX+HmNNgz6ukbCij8TSfTUVgvKUryz3hlOQunLmAuD/jG/r460qN8jwNZU9
cAhbedAG1XYQ+XUyPBmJmSjSpArYwRwAysJ0lkBVvH58/nSQH/YwVyIyIsWNbfXp
K6ALoYWKFzI6KsmGxaBgJlu+V1PA9cnHNQiTfDpcmNyljELgQSJa5coYMsa3E//n
UC+Fq4wJ0b5DxYiQQCT3iVhPl6bN1NgdwqC6sHKNiS270Vmp1dBz1J+vGcvgc+Vx
y6ckB1ki6/AbmvY8D9cxufwEtx1Z1eQVqTtTdIJmxK1+lZGVpagBfhsmVrles/S1
7T3RGW+mSKZGyQJLxvO54iuyUCZOKlyVZLwYQj7ka8HV0zMw8LcPJqo3aDVLtUZR
g+aRqaMjv7ownMUTsRSTj49d8C89D23OTGjleam0oDV0ZhFVKolvfUUTOSOqSTB8
5baBVU4KbzJPVLR73eiCPbXvOFAe2SFsMznEj0zhayqMhyQ3zImMLjWhX5yOm124
u/4jwg0Cg1ngk1KSgBXtiMZf4LtXlbKk9bmb1jzLEv/MLEUrEEfDWo/HEJVSJoHj
N/8l2r2x8diDSj3BQZzMMB4McA7yc7dJ6hgATbjMVtqRFl4xKljE+nrlcGJcFSPb
Q6XkoW2u60DEGJ3wuBvEyJ0ZhRVJtab/TZvsyFuJPEq4udecZe0Vn76+1Zf4dpFc
WpLOL3IzRQAv/ieHOf56MSKAJPWzc2nfVoEVFWN3CqB0NcnaNHRIXL8DaluCjOeF
vjw+rSZ3uj8YNdBpFe/FpGxH3qkfn+fPmuFElk2EGABlK423xDWkk6m9+N/2Uf0/
exLFlsASaz94d4bua/CxFpiiLbuLD4f6L8npmw4effeER7QM8IAuJaH/CI5oXnv3
WfOptotdeKd1U0RY77XmDaXgSZ5rgF1ewqm354ZVwIbvMF5wuFhUQug1Liql6anX
iaESoRiCqHZPIXFgqe4Yf56zxEssWJ5jRlBS6rcJxjM183Acp7DMrui+fgfW6Kh+
mvUSq23P9ewwJypVKRBS3FRTgbVtnghmEYznG+hqDino+ZJo1RZZJg3/21pv4HDs
ufIfkjO/NdMPmu8+hxnzpJ+d0wnWflNTMpwH7aaU4qClmQk5OeRZuUy0HaMdDPZA
1l9YsKlSiH+LBNu6YJd/22gR9RxHrVRaN2CjjIc2rYH7i4CKVikwze1qRJym3cpe
pBU9zl0Ww09Yn5doIDrqcG548KsR+mu2SE4UqcHTS5zCwILoOHPE/ViFbGB9MSCZ
w30D0Y7vRw75nmN1vRdPVVpL5aMKllPy6Sjr2wU0WhztlNDAnMFhKc170HBSo/bA
hgyQszPLagv5PbXodOyXJx5cq0wXPbik3i/jKBhfG31Nv35yQCD44rxKPIZSXFEF
G5J8A6B+ciUnzbWuj7A/nEIU77aZYauRk70KlJwYuW44Dh0612VOK9bFoBu/e5Wa
iHXmbMaugk5UAnB5JESAoq7qMXVcH5zOEJWzNJ3gm1OvSHhAzCVzXAkwhC0R4NLy
zWv71uNdla3l9nGgYZSzEY3ttGEwpk4UeVzf8qW8pBWG9lEK2iE/kFca4bmmAM3g
AoCgNMFvkMzW7gRfr2iWDpNGMGrYBKFyib7YnRIhkyEd3Y2D/y6hvFbGmrotBIo9
Hun10Hd4hCOk62R9GrLU7R4a4dXGk/UeniB2BTzd1EK8TqDITHQLh/lTInmaZkDZ
3Jqin7r4vZx0mGozRWI6l5767nnNi8kMf0fx8i13ZEfO7f6yQ4E65UANaZky6UeD
+xX5FX9JxhdSyYtipEwOFFr2so/2AvR7JM5+uhHFJ9DEtS3SR8EootDBHOM+8Riv
6WB6N3VS5h0vvviqzhHsZxXwJ7e0GmtbpTB5wEpxd31Np883u95PujF/Xsgpqc+M
f4SJCQFn/3fVrRAu6wIQrlITlPMNS5IoaOxjM6UYkGkhlJrDfpcQyRNvLLER+wtU
Nw20ukqROSmpbLYrHkhFcIm+DEISDr8tAjnrZ4Nwaj8wX0RaIZ++Pjs2STrTPAdt
Rcv1jjaYOY9ngjlxnllz9s+a8UA1GyfZ+M9xeWM9ovyctOxQHoJ5d3fFqz+v+aai
ri+wCQrJQKqXUuRtmSBDIdMD7wWM5G6tKBhg1J7J630NHgubf0Mpody5bWaK3Zl0
E31T7e9zR+zGFaGRrGzdXVC4roVA8fl4nbEfn/6heJQgm1L+votXCrBGmZAdQwrf
urhJi8z4AVpnlEAW8w0govjdL8yFZN9WYgRGlhr42ral7dSZwUEUIxZPoLhJCmoX
zMWlwQFQFNSsl4857m2b9bJ/ULYhK/MtUgueQDRb/vecxmYk1FPyogl8gWfh0jQa
g0+dxsVYJsMR7I+EmhXVbCs5NrQuEmWUkW6IjTLVsJ0coAKH54ka0IKdlnotoZSc
rXmUemDmEICnmuGWP8atGR2STRLG1F/vgb1k2DAD5DGhNyYHlicdVbQ3W6iIo5s5
Zte3SNfD3N/ewTUwQ9artjmrKauX1CETqN92zS0ByudzsJJ34IhNth7uv57KJ6Uq
NndG4hvKcjWe/cbAo7Oxl9ULZNKQ19koPpP/2mrM4xHcMeqU+tUCA1OvEseFb3sw
BcJPSj34jT5y+O12oBpqX7E/C1pDPTAQxrtyEZUaVq0kV9a0hIb5d1+8tmldkf47
XmnwNf5nDWdMjnVLmcFhUxKbByuArQZV4gSQpwBFB9+yZcaGtXCqBLrKcnX5OHzl
8xWczdXs3GkubXkHfTWKGPBajySwhiMIO1epIvTiCKkwr2TMKV45lkTs1ZmaOTTq
89s8t3EGq6I834E3Ju7WxMNA12fjXS20n8e/QetVsMhCPLMVXOYJBLDp+0WtnQO3
HNZmeibNv2Uf0AEpL1rK59SQspEXmqLK3TeQd+dhTl4lGAUYKc81quxfwBuIgKnZ
8l5jmSDlpq+D5R6HenZA3PSJSgz4xcnCvfro3EkjjMP3vtnog+hwAbMrbmwlI6wo
T7jOWUqnCo8fIOmv8mroxCbkxeB+O6U0YFioIygfHZtMSXOsFZ7Es+Yq5lYibWmG
O8hfPtLeQW2FN2uQbbWDX05tlJg3BK/1obfddqETKPkepdWnUCG3JgXIjjDiEiUQ
rHSXRuhzrEYDDU9SMYGCAyocwKyKGp9Z28Fi6c+UzBlwCjNXzQpHMpWB6Kn/5WHv
wiDTlxDt5FQwheQLHYKuhQgiFLq37taeQQQdatwL73jn9COt+JD38nihRtRQmTYk
RSE8siS8Ntc4H7oh9PFageUjbBA/DyPvoao1PCM5JFZ8zAf9itMPhmnROREu+tSR
RaXf0iG2mPxdAVgiYARSX83i/m/GYVVANhZIdP7DuOTB3AGk2eUbSrB8S3Hnx7Mb
RCdvNRjEU2L/CC9aJzoCxJ9cD49gE2eooBdFPoB9gFuTuj9mtzm6ERSM2ioJiW53
4EYKM9QoXFy5UumSedlR6RPIoArsHdXk4fyaLb/4GPK7q0TLQLdpUz+vLCNcJSMP
ukH9U28xqdSx3AMS92Fv7/CreVOdTbU/JezuxOW2/JUw5TpLelBQOG0dsgc9dwAv
McpL/8Bgq36KURNNrqtv3mD3gUyD1JSgFkEGXiPQ0cWv2LNiTYFTB+kFKXIPwpxe
eO4Vm4vN1tGDS6SI61dTo77N461Fm3nmJpVniP12x8BT2C5WxU9vpt6nBbNHE1p/
iuXUNwwKvRaEkUI0oHf4caFkHMskoBjtckI5Zsix58RqVhjqq2cgJGlewF9Mr2y7
rGQYpuO83913WQE6+3WA30cpr7tLLJ4S4eCfYNEndKs1Qn2DhiR/fyVK7q2QHk1F
AfsI8vydweGPeYGKkuqZETMHzVkSzMhNUMt6akm1HDUYgNW8Rf7asXwk4gUR74+y
zJM1JtwmdCuBIRhhe2w8e/rtSYeZpSaOd5Xq40LxrfPhGZJ94YXxugQcJ2HJlp7b
fjdQtcutXWs+rpvbOPcKvn8uvB2xkfFppekrqesoasp6I28fbebjttc8qEq/Cfqg
yJflhEPG8DJ7rNw2Ls7IjYE8iTDwQlvy4Hwvu03DE/8s6gR/a9d6k//pyba3oNde
CxpNX5pLydebxv5Cvg08F9ugQuwadjinuovYvd4dvEoTHX6Dszj2+5+nXeeQpJfl
C8EdTqdI38lkzUXxsoAZE+pwz4lBLMOWSQ0wDrxf0w7GaBZehP3pguwmtp7L4hWr
EA81z/wQ0e0fA0HSGumrg/b1YDNqb+EdiwzmrOmimQj5LooQL1ud6lYx0uXIx3hX
FXuLJMDBnCFfCINU/DLc7LdP0BjEvNXs7nNSVQ//ALYvXV9nds517OyVLUEjHzN0
zJm24XKedBNvXL2TjRFAjSucWCbIQ0ZcOO5cRQuSL81pSFemqd7HGgeC3y4GlLQB
mu6U1zvVKl+Ok5YiphZUJNHx2lc5QuyLhP4XLq2VmGGqRuD+D8Xwo+hMk8dGHO2i
G9Mwnd9zJVeiaiR6Tu8WFFXNR40RkAA/nNL9gEY56IR5ez7zzcwI7ErhintiL/Kw
I1nDahFN0Rey10FBxPVI12iEPNa4fjP1MAJzrCv307T/+Fh0G3Sd67wKpmkGi0qt
XFXioXIDvDpWvjbcDl43Wh8idZso63z1bH55ZvODXeVrTTXVm7C+9Jd124/CjsIk
Hno8v458NPsPIY4vNCL44fdsGDRaSH/m06yIw4SHv9LjixWNsPLNm0QzvMgTYNZo
1GGyPnpZb9xtvWvJRKvGRH788rY7/tbN+REtbe2LmhM3+ESgPifaqS+AD01O3plf
Ko/lk51NOqoi24xnQQAZdrrqvlUVW4WcloUg09eVGSUwBbo8zemxMzgeejDLK+D6
DubqbHjc48vqJ2pxXp/1loE+ry/vWl3p1FpfBuQNuHv5jnSa6lSy5GNv/5axvZMp
ny2DBuwc3Wftn8COkBwiQ5vDY25mepI5YUZKn3TPlS7xMQGYuNrcCHlW7a54Wgmf
h1C4DA/xp+nheTdv/7VUvngP643Kw8CfmRHPjF/xLcQAUwsdADS4r6DkWuRrUZ2v
IYACojwlr/TVdKixSiZReD+IhphsaalY9maz2cuvNvkUHEhO4XnizkkUmrifYtoG
1wmJlqDKRh9yMIpx1tMiWyHk2GwbnEC4Qe99Q3LmQjbPyt0Mnl/nwGGY1OPki+0C
skHMy6T785cJcEk0R/bl3GopT9kssCJStJefMhfeAGiOzbdlbQltnHAOFwR6mXJn
ig4aqIsQTuf62DKHPJbYhpRntgzKmwHhmjcl8WOvHzE0cOJASQiBT2IyB9KQg4oU
aG9h8Lg9lw2HAhIsLF5z53TO5BC7fDlU7rkfZwgdvLHbiXAJge79aet907kKnCmc
GFafPAovw0d634JQevFffr1PgUVsThpVPgNw2aXvm97aoFnFUuxOa6HFn7kpdoLc
Zk6um3Y09Et2fK3koDiShjXbXu5codLZx4KTARc6eF3vg0uKZ+XyQgCWMF0UFWEw
Yj/TA0P93SWeE5dyMTBBuZ/oYo0Y4hbTpDDt1Nb8M5KIOnV82eaGiEBcc3s+Zdt2
w3dvQHoy/iMLlootp68ZIqmI71/a8/JzwRWpdIq4Iryhp1TwLyZKwvWHhipqbsKE
4iLt+TlffxRU9OdC4a8VLZs+65m1b+L1Ix3TEAYWEXeeNeqnwCbJFfUuiiaorD3q
NqWj2NDPXBpWXU6H9daO+z1XhKhsK2eNqP1haOjx2rcy4JlKXBNGjXCHhC27c+zv
CnFvSX6aXp0+fHtWX2wQmOf+9of9iIi9X5Gu101kAipqZ+42URKVweBHsTdrfVt8
vOhWp8bgVB3yParRfB8K911Eyyd3WLoddJ7ulXZciEJ6yFq8k7P0rFp9kfvBKO8S
LZ/4VG2rz9z17CvServw6tDg35+6/V9bZnOMEfVCE/nE4EepqF5rr5F9U2sSnxMC
t1wusaZFpTCDQZQQzdRNdu7O7w9uWxi4uC1knFDR8k11m4MRvRymYgWePz34VRmE
TAm0z4J03XvyhXYD34TQHgu+YJ8YOKz7fpgre0Ko4kTDAqbL42sgTA5Rg4rwAB81
zeb+lObCeT45dmMdlEIVoiSfsrFfkOggnH7hSMzaH7Dfd3xFtYqPhEaaE/NLIVn+
wuO33FNzJeqvP0jfytv7T5gweSlWMTZdGkQuKcFCN1t7bLbxJCxWApoz8iQcpDXi
frGEMBJRF4inaqaaeUt0AkzlcdlecIUBh8S2zD7w7Wfs6o7XVPHRRqiozjo9HWxZ
SW9pWu5TAJu9Ygxa+ajbWxal+De/P9RfzzuGGJGZAO/S6C6gvJaHMd+jb7bWcGgP
v8DSExtWdjCLXtUhifEFDoQ3bQVZ6keG6HYUVUn8un5+PjKHavOy3vxO1GxwBLB5
lAcpuel1phrN+N9+apxWYnoL3MgjftPM+XLf5cuRKt5RKqHbcX041sYADQLWNhl/
049DsaGleKwqvXOajCBCtj+cDJHKQ2R2n0q995xKp3G7JZxwVD7kMtxbnPvanaFf
QTas/+/JIntT5YnJFfHyNJcyRJ/5XxoWOyid6rdIeWkou+35to0/1jZAjwnptjvq
WNl8iKQns/X0ToG/E5ifTwupCpAhTGF5DFYLbn/4YfXOqwlmC/jyxMkpr7bYPKvr
49jqW0u6SlSVVM1+j+HC9hUEDu3vrD5MxRFs6zgQ2P966bESrx8Z9HFIqjbT9rge
/4N5fy7JKemBUm2GEL/M24JRHJ782Ol35ZZPyjTDmrKTPlwiWPiJfzNXnHHRdxnM
y46fEt3VethDEUu82WreirtLlIDFsrq/ASKhHr9gjkii+4qnSEBQrPpuA16fs0zT
KQgQcwhIs6KMmfLRafnADL1DUkMYZksozzG/z2ZKeWt/xttILY7xo9rkC7MweVjl
To/eROENZWt3xqmNhT5SZu0USkQaGWbBG8Ld47rk7HLGtJ6ujOXOCXxzZjUpKnRU
XCmyWOt310TApoSBdj2W+rjKgjN1q2aCRn1tIPQ5xajwfeujlY59lnvMUiXdSD5u
/0iWHrBWYZNYqvI1nc/Qrj7AkxEzIEaV4vEIxYu6wxV3VomtBVFux48fT4Uhlp44
zGhrWAsWV9AhTn4DTEiovUlZBnpD8gU8Xj+Nw5kWrqpEmsRjBZI29IvW1xVPe6bL
8UDubCRA1Vg9+tdPnajlRGJmUOJyvNtTPtyV0cADU0CJO9jAqxG+8WYuIfhjJVK1
XqGIlGFuS8yy2j6K9Ea8mJjXCnhJd5jmZKzAH6q4+VDF/49F+h8gsDwEY8sQtwCR
lHGjCPUdP7u35a/a0LGRey8QriiDA/4Dq3OweKEQcnGYzyqzlo0u65cBNJHz1c1U
BAZnpHHRCAN06NPSM148e5ctIHExxmKKFP2W9bzu8cl9w0EKUNulY7HSe30L6oUr
lz0+YosDbGGgObmXdg0gazGlqveTHMLddBY1flG2VlhxKC/3g8S4UO7xjFCjyNAH
dD4imGq9J34fRbAMIAu9yYWm1G/+V1q9SUvOVdb9jIQiiA7gF4EpSItPXun/Hifl
Amb6+Kblci5xEpBnWF/cwfeDeZeWf4BraGZwfNSNYtRkM1Xbg73zAn+2IWcDNH2q
942Yrd7GdVG42jqcJntSmoEhXYXLFw3+GRCJA0h5YACUaCLx8krN49ceT2MgOuUa
J08IKBgcXoyPLcscaYFYLriC5yZcT0pZuuRRP0J5XY/4s8c1u56nd0DTw2grwWWc
NOD1PzqsZCU8KpGsPaunDt3cVaP7PmQW9XkgvfRligQhbbWHkilOcCxnXwMHJSp7
VPjT8Q2zFJF9cJrfHfKL+CtiLvHPXT2AGFmwT7JncWsyjayOCqkG0r6KopuF4Yld
5di3u4JoB0m26bvcN6MvJUu82vNUbRmRGqrK7PrfRtmSFhkwQvFKmqoDR/ZgmZfV
InNUxce0MA0fy4wAu/SUlStSx4MWRezHO9KoWzYpovn229kHmZD9w1lzFmQpvYm8
XtsbKl0gewX6Sbk+n37yolEXz5Z/v6Ewb4YDJZvEumMWcjb/sFA7BuFYZzH+yqsD
HqkPGWu4j3tyM/yk+hPmP/SbTqac2XVzsMXY9ERejlrVULmJ3uHmUxsw6IaeUhi8
JjJJMh2usMeA7GCPUAUy0I8NWwmG23KHtTTJbOluCq2F/rKB93hQYZp8X5fOgdrY
9QHAoOMfl/LwnlWfWaRE800BGxZC/URVGh9bqlxdUv4kAkkHeBiIfzYhNSb7hLP6
4InlSzP/kdbMgtnk92akXIhM3bImRf1qo0i67mPkb8Xi0dxrUa2IEjffJcUVtbjy
3SuvaHSTpeyh0UP/KWRx+Q4OAmx/O2gfVERXLrMpe0g72acXUIm8tH7V4QgPVKjG
zp0sfD5J57nygcB8SFZaBNokQRlnE+K0rvhYPF/WxXHGe9MPwZweMReIydV4wtXN
GdLYrUM1rNaAAf5/811el/rUEkkEolfO8XyuhVN4vFG/yhUCp350XDHvvJk0y8hT
j5Iuy3ORsFnci3MQVAOr0NI0+ne03IOi2MIthj5jMgZBjOD4cSWm3Zp/oOlSniCZ
czui/hDp23wy/gLVty/0kzKF3bA3VvIXXmjkxKWBraB67h+a/+TUC7NxpmAVhNxl
F6ioE7xKKvfNcVoxVpYrsb3wR+wkhuAMXrGEAsFO4XpaW4RajJxgyzVFt6cW9km/
/bAiWQ7K8hxAPMU87dB0RIje83mlVu5tPVcfZZtUQZTxvhwP+uBYjWp8noqbpsQ9
e8XBnI602NhOdmNf7hPccnN+Yurc7qIvO7Q1jWgRmVNd3OrAJoTMw6tsAKgqkQoG
AxfiMeSZMJAJjemxlFLn3frCF0AOUnO7XsLS2UQjfW0bwvhqjOMeK1+e2gVQbeFs
SlCE56LIsEs+tT+0wcrFoljNwywR2RQdfzWHm79SaAofQC/E4PHcxFghKBgILGyS
R4be+RoUli0nB3xtig2SfMYxQRv4vWtyaQZWQS0eNoDmA8B2aryO0NZF7ux9bLJ6
mR3Z2K6RrF6TASIol0h3Nv7yFqq5ToCaI/fZMLhNebnEvsl+GD0KpBbpmphLX4B6
TVRHDyn/R6gD0gfay6O2uyh8YdbmgKoDVT/X8kSioml28Qx1VAZ7gkIV6Xn4ZCWC
TG/E0uvvNS0DFR5LJ7gka/wGD0PZQ0CezpCGyctMYKC5uI5e4JjH8WOnC346NWlQ
HWezKoVXmxblIuyo3Z7Xjx6ZX9+ihYRD39ksKz8Z4cnb5fRraYE4f7KZN17sk/bQ
hU9EEO89m26zD1vD2UfP4H6RK/7LldP/zkOn1pC5hT+MyK5dyHQuS0pL/aXPKLtM
Dl68Yt3eQTuAe5JbkoKCLuIk+4wx0fBkR3n4nCGQBMtDRGaBtUPdEK2srlVqaBjb
LX6eGTqp2vkahgGpzcHeZf0cKb/GtAHbLzwkzN2h04Zy1BkF0nlqqOOD6C4mQr9O
CYEE1XzfpxgoYSq3eZgKpT2tfIQWo+jozrsGU/+njrf2jjT7oTKzg59KjwHv10Bq
9IxBfpXbjgiSce7Vpzh7W7aj/NDJuSQDzAIgC8O2SG6UJHuRZIGsdqMnN1ZqTPvu
p85pFqvR98tzHR6DHeDpqXl7wSevrAl44+2GLaeLAvymhsh3AQfWBdwKFjt/81Hb
rAbfqjX7YecXTXj63Oqiun1zX5iRi2epMtgQtWjsvvI/Vsu6+xi6BNbi4Qbi4RzP
tcbOHLUJBTAvLSOV0rU6GjQpMAztSpJZyTCdIqjsysbrcJ4s5zxqkO9NRmlj0FL0
H6nb2b/EAIuZcm40wV3Y/BpAvQkrpUGKnjqXEHEROaK7nnzs5QkgSfIcP3zb5A4D
yskv3itmIkq1aIeKCZuJUxxEjkupWQAS1dC0tyNTO/u9b6cawSbwErC9mliD+UEI
1Jhs96VnhFkn4HUq5vwkgFklaaF1rZvyIiDdTE4du/nmEAINtOWmvIaZVvgpyCb+
hWBHNicmbALzzGqUSf4MwHxtF1rvmwIdfBpCVVgYAgF4PuQIK2y+UEum10c4lKfi
6HAFr3fDvZzbUPJQQ/thg+Y2qEgM/qzWpGvMuH1gs0Gqr0gMgG46ruXoTtZzeV84
HYRTBoQ0vGtHhhmzlZsvL1JZ7kbmZT4ItGpcazgRx3gMDZive1fnQknHoGKJ6vpo
BMnkOYbi0dzDcgPhLZLwOrwG8IzL0W9tmHZDFa91XObkA79Ud1EkR58EaNKAJq34
ww0E9OLGFjviuJUqpw09lEsjfYZbXei4uQ1Qkiys7eIXkx5K5bC/Lk9O4oHuAHsE
a5S8htE3dxnqWmh0UHwitl3HWOgljMNGACsuP/mr+0SFJjs1GFXoK8O6jl+tth4M
PxusnSx9HBTDAT8TI2XpxtEpKm/4GSwp7uy2WetXPaPcLtrKMJ7Zo17ZWItgONoP
pr35d6LlgQ/kcrBf1XPvjeMjVnqJch8I0q2MaqW0MGReD81eWYd5Ex2GCcy1bkQ+
Oqq8XLqK+JuOTEX3Cmflt0sXJv5ABwVCdQHokrNENx/OQfgSLcJNbnSJn21JikRa
elxUoupB7R8s42qQGOMuZXTxQ6afyS5i0gjbYRy2NIHwczIv929oLgrIPyTDqZNg
4c/KZ1EHyTPu4gC2IqqMAhE5rLoc1qIhQkiTwLAiHR6Go5xXvXHoE9EVGPN9LCXj
In6l4ZpZ1LpXDRPpwozFVd3qGPnzp4BK4DzCJdfacxC8m3fUmV8LYP7v2EGDjUAZ
Dsb29L+O/lmzMlul/v4r3vXOYf+CygOTEkF6Cg5WOJLj15tPqkvyBGVsmZrTPj+m
RkHfBKxPt3hrU/G0deH+JOBiV2qcMfSIMrbhRLg/+y3LpnQ0wXxuDbrfHa2q3QeD
o8iImYC4hMBdeWFk6u6azUwPh/3qpWIIPNHeM6JmrMDVqvrIdKUlUrCq71R/szF7
qIjBTam4p1lOv4Gc9QrhCc75s+bFNiMTm+GlB3rHef0ROiSTehYtZROfHtvp58xy
VdscQAPgsUauiIyHhvSZfMhgxWtG6SYMqfLnxYp5JO/Gtww8lv6GCbuUcmB1pqth
+BeuRMNbqzsE+gSrCFHHEs3uzZPPxKyIpATGwmjuHhZ2hvQN3kIa9N4GYc0BNIuw
nzc2J8Y21gKJrNKqfoRL9+fvNtWkoD5yTeEpOOwJ+opX73Qv8mK1y///AGWK108m
HKhip6flz4RGjkdy3nWn/OMxYsh/Ni4P7hWf74w7rZ4gmqxpEG7VmaVu9o43yT71
jNGMauNzYTS9BGQZnOxtG0uWGsBEUtM6ts8QpcgbxsHcoe79YNTMqXbDcqwT2FsO
HTx7VHF0igeacCmPITR3kCB8yNMZlx+AqBZbjGqjifTTJ84X9by5KdAbUdi/5CRy
S3YI9+NVPNiV3VVcKlLYj/iGCtmoriD63o+aHwd7rUMmI46lCBDCyfgO6kvfzZ1w
t2GBEjkoV0FYUzYBezfL93W7YSbALVXWHsOephTW8hUgPZVJtpBDJkn24WNwihdp
bV3/JvX6rXauo6oA8xg7fKH2INeqyQSgY2+tTPlFfz7++KXly8IHrH1SiqU/mPmq
Zflh91L5m68J27Kz8J6WY9acLZjQl2wq66oWqKGH+K5s7Iy1qvlaiiFcAmjXV8Sa
MVBdOpeRefZkh0Kfo/2wGeLUtXstVQx6IiSglGyJhgRVgqo9mh9eTE48W8nhrP8x
bOkv8PVQ6/M6PwjGIqmmHsCPZOBxx+Hvlrs42V6mOw+SHtedOqSvrXwxMWFWPilF
sV9vLbhzhXSAvCYT+ww8I0QLsKJUAAv1qSVvNKHhZHauJQj8zUVkAQKCkqa3kqHd
U7jrZnMB/04YzqAvO+3DvcwEZ7pWjPLPvP2dUbI8NqHwhu1Bex9HU2OVck5Z4fEb
t3Kc7OSjvvzWDgcHJ2z++3p12LjzqpcpBgvQSUby0IVO7SmEoBZfkn9nxVQyXEml
mb9Xoay1riQhDQ3Y8VyrH23EXcE4Mz7V7uvKypE+SalQpEluNAFLEM4nWEg9nVbS
gEwfsAn1MpFDF6ELvEMhmthqGUH5H7WK6zCYOQhg3wqzEL1vmifpwxmjdmIl78rP
VUhj7Nvk0YD9GVg9DmmAPwpwYJa/xB5Xyx1YL0xYb2VZyvz8U0aFwkYOrj17YDq9
ysao+5RkFKnLS7grPKmp1IvloBY5KGAqgKkjqE6nSQG9hAsHV4vYs4xWa4oj8Kql
uPlEOOglPQW5ndJaGJHdd/dGBZkg96wFUvOeWHvq5h/GqccgrR18dlFOi6LkOIn6
Bp0EHWj0Y2AkcHEIQ3bGnpP1BjqekNT4XDR96clTTfvCBMVdTgVO14MoGzM7ZRYW
pssi4uck0u0gxkYeiPYKGthc11hhlF7BTUlm2iQ6qkOFew6+kcuEjma6U8RJq1FI
5blqUxQArTAzRXu9WnY6c3bsORvQV2PYYNKuEqYN3GhnCAbWYmJgZWECz8FEy0In
oA4ldhQf3fRLCMuVnmM5TSqylD4pFActNeyZb8DwgyTmoKcrQJtXzep4D9+M3Id5
bTk780vOHMumJjD+r6/g2LCksH0FqzQg5cH8U9I9IodKN2RInS1QbASC23ZJbXU7
zduYOcPZ5EG4N3SfnY4eV1N4BidlWWpvsmyyDhYpxU/LX/AZMGaZ2G1Q5bCs79JP
yJ7tDvMrAa8nC4dWcml5JcM43qPvcNxUNvGUsd0bMf54bQOvyGm0826a2A+W2M1x
aYsGH9HNpTQnW8M47ysUW2Ey3I82qMtmn5tMw8VG8KEg1hKoA8427AOMEsHvT1bD
xsufucCbbAi+sz76xuqrtwphNG626o+Q9nr0jJoisaTzgOVN7jpzX7hYilJOIfsV
tMEzA6CFBnCSdVE6GGVtfuUuLB8P3ZP+taa5dKVkhsIa6JaAEZiAbZGOg5FbYixe
SycmDTNTA7LrcitdNOEsTBcVK4MtEy+8844MRsVX2Bi6rgmd69S6te8yfjt9w22h
xa5jUjszEq4R8hk01wwekgcnF9osTMPpqGzVDwxcwfwKksBra1kc1Q/+PW7gwpHc
23oAN9r9hzJPoX+v5xcOkRNiyZUst28GHyfutx7PSLwgNThIZOIu0wliB3rmUJnI
dESDe6XlBCXMC0nNJMatzOw5SgiOCEWP52GsA6oW1mkKEABstIBY3otwRAKTFOeR
BoJNXwa0vRbzIpsWNQg88ERkOlIwm9TDOOVEn/4IypoY5AmWSdoYK7OW24R2MJ+g
GPIPZslypNaUYB8fKT1YJzei2wl/J2PEUKQ5w+qKnrZJO0zw5o9Ho0Jvs0YEy4BZ
OfEluXX69XqDDLg1nZOZvc6gksWiT8VY54Pk4zfDgMEigSf1dO8ePyXoxlD5CFZ2
Zx0VfYzBcqntTVPo7s6oXTWmRk+tSml0tnSEgvB00MzxWXccVOUGYnpCK6bYDHOL
4BchTINu2Rqla7h1REtH27k3KFw0GgzPs7E8HwFOdq9+MRl9ZMAHkmOjaDMPmiLa
pQdobNVHLWZVrc4ALiOxc7yIL2vlfhJEaYobhuS0eW0WOblb2S1CIXZAgXkxaoq/
418oVOx3htH/KIDwftP93k9Wmyt/9ma1YD6yIAy4JVN1EBS95ntj73BumVVnmNJr
M9TBOmGlJd7amzZVgWW87IyX82B78Z50LjA7auUhx7+3RoXwj8drIjdyvXAV/Pji
aCgg32zyrydSEkeQ9M2jo7MAjEfrVey/KJv0TP8GOiMQFhj02VzM7aQ6bCa2RTZ3
C6yuLZfi7ygdH7kbVC2p0hVLkQIzgwRaikvBO61ILchOi4cpotm95n0zGkjEg4AG
mCmqsScwPyf5ZMyEYrRIWwtWp4EDQUsRMAoVgOMPyS8ku2MS4YVb8AqmMGjFDNNM
6JZ2NI0siXMYX/gY4looiJ06yRzWs4F1/9/PNZWoHJV6SSASZfk7vxTa80NdvaCN
WRHDrjPegUny6BCjVfPPoYtc1dL23ImJDyOSImNyMiJJLm6W2BOYqF+LJRrigSkw
HZdYRvL7jpeb5l4csTVsv5vGHY7c1quODimjzq6gXkKelToMb/3Jf1LdKnGpyZtX
sm888VQ8a4G7A10BP3O18/akcydXz00l7JvzENmWYDqd1v3ZbsXDnXK28sqZt2uz
VdwCoWBJqnd5TNc+mOv9nAUpqjNWlzM1wju29Mze74S7XA/LchtnG9awWAb94tfa
1ovUqCGz/xZEXLojzWwIyK7iO1k3WWYkAVaniUgw+Pe0yp53sf4Ts1BATsuKZDAo
4txFQguwllKbeABiHESZ0SQ1T+8l16RwF72EX9nKMe7S7S2h/g5MhSZxRAi+N2K5
OhBmpGIqzWOOnWA/0XRv+nIFbx6dh4zZdYX3saL03HhtWzbo5e13h5RJbcG/KdoC
hklmQAbX4yLklK52O0VflsFwHV/uJ/aAEY3A87vAe4ZRkUNXuJZyR5vljPN1TnLF
PL1d+7TMoPvqTFU9fY4mHmLrgEfVTQ+BTPaAmUKxwLYvbap2SylvoHtkz55+5/Vh
fNTp6t9+cB7J3iORphQo8ChbjcVjfFywaZH5sJ8jwHk9z22YpCzGmOkxm0FfWVGM
hu5uJ9wVIS9uye6eOmAH5DWdxogIUO2NPruvrvweIEj9l38KaVdPkz/VnlSWNfU+
v1qEhXBb9xzFoqeoLMf5tXwHcValxjz2+iapr30hb+gEuaUeL4Dh48ArzSe2ePVV
Gr4hekVuKCze0zWEFJiUbuFIUWJ8V5vIc3stSa6BDclS0429EECCeJNL/xyXxwkQ
nJuW+YgyV1quA7ZIOlHZIASO0lcD0n93dmy1G/yxIS1t0laWrA52OiBhyJRa4Q+z
ohw6kf7K4/W/nggaZoyl9GMEVLOQz7Z5+10AspgxSu63WSqU1D6AruqwdRYMnNTD
9dvq9ACg1MCSXTwQbVaQqF1wFfLh91gvCwo4ts803uXez5LMjmRcyF61j5daiGYE
4+8Nm9/FbMyoasHHtDMszH2WO41cKg1HoVth2zZl3pqv/aUTwDlc1lbItxEzCkQI
HNCiwnT1Wh+PS1xIuJCMQkh24546sfIF6JBGuYhsGu6D993krd7lgT7WWe9Rjb5i
z6U45KSSqtS9GOBy9T7fYf3yyAykDOsUQUk+3YvQbNtRo4NGuQdaVjqzlxFL8lRg
/4rvKDix2ztsntsmPcRNZCsGjwc3ZSAzbBmuh1YIwAhS4IEF5Xh/ugGJ+quc72/H
W1Pb3BMSjOClvpwtqCI8aysiY6E55FHzWI4V9o0WYIHJGGyjVdb9d2hFT0qMx3ha
diz4D7C1iUiSgbTpP/gVUmjiXHiWcgqZ6j/DPRwMsr1n6uEF/G07qpJxf/8shWNk
WbkxDNJJNQ56fp0jerS6hcBL+K4n69hK5Qjk34MnAA3ZdB9qWnZ2oSD+wdtL+3EK
p1i5cupAUJ3dJSC/Od18a43XoWi3UavgJCGpQg8uqUGdox9zPnvzeRAK6sKUeHy5
d8fOty0HgZl8VZG5u8dU3FcEvnkvZjTBE+O+e2UUmj9FT1CSXpHnQGSXLsjewX2U
DrmgTX9OqDWHj+H8efEPwHJs1dRErsgN3cCUOofE5azy8L7hO4ILASJmFAYzyMa/
8nVXJFXsk6gRwsivHvQKcZ/fTnin9YpA2UKrS8YJxB74EhRhF6rvMVMydnPZPVk6
6AyjjxEcAQjsHX/Nqv3P/VixYx6XN6cfRF60cGIPJ+RN63e4M+UCQgZ0lRyAz4Hr
NaTDVKKez+apbZK3xWZucJCtA6b/UJfpaVUliaYBoUCC6qnMH7CA7Dv4CM41oCQ2
L3ZunJzhRdDKE7j1bqxB3yo0gQinvX6rVNR+qelXOGngN191Kn+h+kV9hKO8HVBA
rkG6zHTme6MjhTZqbHtdcfQgBQ8DhiF92uFTysYW3H9syk8Knsd9PR0Rkq0+88/9
Aa+HRjmH1DLHOqRFmLXUZwic5Y3YCPLRwEbFXdgY3UlUn+OQh9Q97lyPhB4iAF+0
fcRL8WBJSPC9cjFQCK7q8iXV3oFmEDu7l8OENGQKUDfuaKj/VgDCyHRwDbZoz9QZ
U+79MVl5+Ln/oo1TWb7wV8aiYesughI7NLY/Rk5ROvmjiWCUY2EY/qoKxUwsGyiH
kHW6E1f5j7mlnKcO1uriT0aca/+nNrG1WReyRdLXjR9M1tNaNywW/XJdxpBNM3x7
mAvIssqtIi04PJa+nRrFWGoMLZMZaVPlJleIYH/iLVAbl8KOyugbQe7GcubP2zhI
wgYuWAiD+jr+LfEhITlWMowQ0YE8mXPY4n1UUKsGIv3vhQewdbJ5/Pq5JgkXMn4V
6AHmgYV+cf++4kTQYNhBx695KlyYNJgTUUfdwgqkjVtCScJIsuk4TYYUW6j+73L/
YsApRh1U1IVLe95l1pz0hqKPIMdkiwne4HNkpOGNJygFlOaYTjcjq6y4wj/6TZjh
bGsMmm+Mi79V+S+lkbhwQ/j+myy30zSAV0HzAUFXKXZOmyvQQZz+0qIMiVHt0bSj
iIM4uQa6VmQwjOCq+ETO4qdbL4nzow8VNUQhv7O81vJ28ctjx9wIDxWf2HceP/eI
dcC0RDkT88XjH52yI9Xl2UR4tFfo8lQx3m+COZSfKRrs1AqGOBaxxqwhGzYN/FQL
gn+qVyOwMZHTOlHiJ2oO4BMY2/LrDnV0uJm/M4Sf89X4eHjCZjkBnvTQ8nQ5rQtL
MhrG6LPcipxh2rQWhGfONHYelakxhcJqYd/HhPAEtsKIjButtzKevhQHvgs4mmFd
y2WyvqB5NOQjCOWTWW6hIdh3G+T7oNtiBaecmf6uLuYEJjBQ5bpjhwFogMbPnCrH
SHqAmVlixRZqnhL/EPOepjmyK4Ytrunha+/9wxBaeysZ1+EaV/hq7cl7qrUE3eXX
88ilIrMBKbPf3AtJvgrAhIgQauIoxXqFshEraBhaO480ykW3YPqFmBPfA40YT/o8
jvDBQMQBruC5ieJ4hcJBOfvRQUXkhGJdddqs2vEbJ6km3VusM1e028G5Q2N8YoTO
z3dRpOduZm4Qd5V0u90c6zK2Q8T59QO8KrUorbGp/825aqFElTWAXC35RsxEL57c
LXb3S3xHJa0Y6YM4aGeyMZUcjOCifkIYYvdVJ3DliLuAl6UebTMOzrgLerpKK3Uv
zT9+1ubKatSzrwT/ZOIUsatmjT5KYqPGYS59OlYBfDY/ryLtVqWqqMJuJo1PeBSq
t6HTR8g/s0h8zK2Jxk4EEuNQ7uLYYmQTLtunMNDsZG6LYzKn19kpSUdvLbOLvVgD
kXgK37qKqM6jgnYCUkUIENR0Kw6Hvz+g40/Lui9ZNm3g9CwmeOwXkhyWAyHmySpK
ODjnU313Ln91bDAep5OnW939OL+/gACMq1jz5THX//28KBL3WVQIU44FxHe33UPB
psHrT2Chs+JZzhHXNkAhGKFNOtcsOkH7FOwVbLKn7GCr/xWXYfHm325sLYwF1LSV
lqEyjQMdbyki1Z04ub6MpiU2IsUNzb2Zhz0LvVT508KxMs6FfykRmvgZ3DisX2b0
lsUajDeg1UN70xPshGgvfrbLP1aIb53v4g3DpjbBoe/tJY5wsED+9rbvdV7IBQS7
/ecDDdml7yZPHfHIZj+Z4bhs8c1qvPC9KDJjb2NiNWr5iREl4IMYFOdcpNSf9BVp
vkscDN2ZlwfrvwiFUBnMdSXHMfqaNnd/XBsjagM7qUors8USOlsLAmN1Y3s5TLQy
fYPEZ281AlRkah0TWs1hsO4q/z11GJjndekET2JD4oMNSZoZYoXtwahpRUIfoU7V
xuHY1iF1dqtkfMrDwByOvnmyTtkoHA6cgIYrCdx2FAqsdBxAYatcLw5BNn7keq83
E3mgbZJwdL1Jl6NJg4yGXO8WeyFwLbRVC0pIlTCrcboz0ECzmMGofac6QvqHduV2
/P9Plx1+3FY+3K6giYuTD3WihUULcT/aGygWY45Vyq6hhKENMQihdWedGr3dGZJO
bWs40ZjBVb1qbai+TssLq5gfQjVxkNMwmqaninmEx7GuIflGn8Dy/cS+7PSCoBkt
PR2elR3OFtsmAnMzTjKv8GbVb/lmZtgHUeAGgmtr6jwXk1xD86OxmKWT16pSqc2v
2xkYc8hJ6buDerGznJ4JEod0sZ9h+0I08qI9UW20AeYhSt7Vp5FXFnpfT0KVq8hi
E+HhkauyPv04uqK1bqutJBhjnaNkYk6RKwBYBihbWRRVZZ16D1RWOWc4JB3TZZXt
oIYrUOaxb8FvAuZzOKAeeI5tXUYmoOuqtDP8Rm4BFURk9jBpPNoHJHJ3wNSmbJOS
kGgUpPcNhyKpvSAZml/eDVxP6triAT6rvcD+XPo5HEDinocPMGFN2oY/gvnu2teU
QHTMbrg3Cd+6Yv82l9eP1p+gwkO5aO/X6RJRBfiL+ehAJcq8wzb+fVx/aK+FqRU6
dPRnaUyXTzLscZAzmVUx8oK/4eg9Rqq4epuyZlXrNfMHqnsCqRy7QuK037KpSwBm
r9I5wbRfXKCSun5KdFrrnATc1WRHDAhmjS7L9Yn+enzHMvM93GNkQrqxss8M3Q5j
uSgEQr7PSH45b8b0wO4hkMB8bOy78Bzn4gId2z4iuOHqe+UrxJAeYJJqzxQnhv1G
DILRDa+lKYciUdp9DFpYuNhTrVmvi+iPVj89QxidL8i3TQ6TnPjVxzedaoCy/HmP
H9ayoBBFvJqscPb8Xm/7gvMpP5x6BCBGdarP5PqtgMc91jIwD8wQ0B5H/Ytayox0
rUx0UZcUDQ0Y2um4ehPN8ap4ldpopGFt7+JL6A6cG62MfMCIa5NVtaJY6eZwoUA2
jXrc23BC36Emrh6JduEnBqc+8JrGf7rbz0hEpGOtm3k1Fzce496kBI0w3cpVgB49
+RzpS6q6+UwAEbMUkz81ozw8MnmAeNGMoENpndOipZrhc3wk3SrF0ZpKz9xq4sM/
ZPR4th2+sFJAZmpv2xPvUEsRNeMOsVerAON+0V39tc9ftQgIN5um3pzJ57z+fJm2
o+117kprCnkfVysyvsxc1umPPdxNQBML2cJvmz5QE/SIAdAMV0/4MIanc/VCrF5J
e1ryOjbQnsmc8PpCm+KmcTCZZUcA9DU9GsuRcAF+xpFYlOHhijRjztxEHQXDoj5e
B59VwSyA2GVZI9DXUi1wlIoNuxsJa8DRvYnVatKrZH5vPZL7WjuIK/zdC53f3DlR
5NBodSb7yE9inPU7TJP//AhODOXvzMqSh09K6LQn9VxC80nqJjyK709GMYIpFDvF
GVztt0i5E01kle0KpHqfBKSnDDdY07apm2ycg29C8JSpKCQa7WyUCKWKAdPt6tWt
gZvP5TygF+q2CKasuZA86jU+4fP3IfiPCiBWHr7RR4js4tlGI1Jty772xzt537Uo
b+S6wxY/Q840W9JG5UrEFSJ+10Ys2cG2Dq5MCHFEgOvMoJM9dIErLo6lKE5GuepW
hWImt7jVjT/YvLvtiChT25LBIslQHy/P/yCLN0/+A9fKzteASfcLuv5RSDGim6tV
+O6XhGoKXf52+j1HSt6Pc2KyzyPsFMGFz17RMI9fdOUsejAf61hdPscwTyFnFctp
VldVoHLAsM4CmBxhznFbgvnOmAwLVXVRuBmRWDlv/nYdgPL02J5+zycUBusfbWHy
Wk4qh2UZ2VumEg9sqZZwnzvh8g02qSN7e+StKB99bNn5pHH8REJsu4hsNJVfhOwK
XlH1b6hAHn5RlJKQKz4kFCIkdOKhQs136xXSVmAtV9/C9R2nKp3ZuNNBYMe6PZKw
GWBPFlVG/jtHjwnMwRM9kkaBxwxn6OET/dpAVDYSLdyKADvSgNt+R48njX6quiLU
m3WmP66nNsJT4UXav5KZWMUeXad+GQgr2IHP798kCvW0F2W69KKauyCtYMXXKcA5
EiEFLtVBqUNrdxswTmXDNmjvmrKfSW5k2CDAeJALmlzZcrLfooVaTSYx/u9xaw5V
+pi9q/q0kdujcuobkN4Eeyyi+EvXjZ/LkFbq2DSTgQlVF1MyIKNlupMYdHsQsJwO
ZHUzaTec6uuwKME7qHuASKmnGVPQFKBm1HUNcngh6YNV3wnpVGDG2HElyHbCr3qp
Wx9m6ID/7fLq89F0mEmdctGubfzcqiBfvNehFNRam4dofkhQ1S0H03Hf1eoEcj/p
ctbv4vqUUte3vZxJ/hb0wOId+G3Iburc70vSn7IEn8uvB/8zIk03Ty6ia738SOVN
tqCJdYzPeJV7a66t+4Q2eAiO0lLvSLmheiaJSK29ZVZu8ffHtfsY5Jugvou3Ox3x
UzBSw+pU2gkCINtaj0BXoE7pMl3SVfsQATncXehcxtZLlWHdn+lgi4yb2dvh2rlr
ZY4awxLyXSPgblNVQWwV8B8l16POiP7Ytm8fjy1TF2mov8Va4aIZcZ4MZ6lzzBMI
nBG/W6owyc5+DrTO8+j82jKg3V7Esct6dizRIJIsTLjNTqUqGUsmcCEh8ZiE/gd2
ffLZM+KtzrjeYITQJSrFP6KPtZYMPkBzFO2OwLqOR6GDKnTAl7XA2Fp0xcVOOux9
/TTlUzmAm2ow0K/m14haFTA5td9fmEESl3Np+SckBzs7u2aUd243WXVwrB/dpNd8
nmMTuddv+gXF1AnPUqgQBnu4Q7SChp49mRWh/GlNqCaDyshA4eoHfnapLfoD6fpR
/EPNzu/1qhhCa8BqvVpREzwr9Fu8WsSeE/7EOQHS4NgO347dcTtAVjZVIu38ub8g
/qhm/KUwWgVB1hc9lc8SjFZcb0JfEZF4BAcqWm3dzrRgCVz/ifhyL+xRoMVBBkVI
m8Vt9JzV5tz0NBa1tbjW86GBWN8JAglgR29f11JtlZR+uz+v6eBosPrEWNCPYFsR
HdQBRTvnsZ0XX33ZIkpQrusFfV6owSEQSuLUwPpdQM6YxOXEL77KwerxuvAjgL3r
mdjMvjbvWm7XcrKP3Jl+5dx9s212iaaKTMibgSRXC7N+JMBYIw/bmSzK7UXhR0VM
824pNJnbG2CzkpaPu/WPhVVULxdHzzii/fdp9HrCMxecAbIhSmfMhn8JeorY/rVU
gRCFG2HhcLN0TDasyaf+/3FSNUeE9+KZJkN8fVPTRStG9wK12lYING29crgj1SXC
dNuz1evQtCLu4EMkhrvf0fCvqRwyqYr/BntdpjR+/DeswQsKWrPWNMwWZuHmrcg6
DXPkW0x4I1zUCRCznv51QlMB28ig1OoUuY5bPVYkebSOho084nv6otKwOaHNCZOV
LvYu16Z5p+e+FRoQtAnkdFMOL+omjPojZ4+ds4pq88/9195FxloOftp3ALJTyInh
yyfcQLw3U2DW8JCkugDqxu505OaCSV6XpLgnrD4BdT1GRZZbCyh7bwyHB7WTXkl4
A8k+ljSf57KgNOB6CBzNwYooAPF9fTIEDpgO7+H6zMmVe9bnAwD+LOGRoQ5TIbL3
PQZ+vnALdBbLcsIuDF8v+313kxnF5lEeQmODyOU9Q45dFDNZDt12SSxmzBvXMcla
ZfDJr6E+JqZbB0ZL2PWXsQSWTeBQAjFZ2XP+Txk3tjAyCjzuGP8Ws5fIxm+3/a/l
N5m/WU0NFkePRCXjq95N4ye3keXEIzn/jk7o++tE0ksx7IDxe3aQGn3xmnSb7dsm
xxyvYsiC4sXAOXnJLgYFDRLvYpCUdxo91hNs8Sr7jWALmqlDgsFv73qQqzZt8N0i
6SA9DW6xg7pQFQrbOYjjNFHJYdJ0fbXymsJPJbmdJ5WRAXetzB8PAUX2dWWs0cNq
xfauUqxXPJr/tW6V+F5ipowMsO229BYa/ivGM/U31hjWdPEbsAYheYr4xiEGcy36
1xSpnRcAXdjc0FSpm2oYavsClz1mX+KSp9KY+LdNuVUVrJqOtqLTActICOLDwfgE
6lbg+VZh4ZMDGVbncMa7syVmaEtUqBfbj92fvlMpmUTZ0u06lFw7KR1bkcnpz9vD
2gB67qRyWmtC1SlFR/lQh8pc0T+5HdnSYU/0TItNXSBw23ASmX9u7uA23uJhYf4T
APndgT3Z8OmmXOuUE5zWRVPWSWPuweWsgNvJ9qRB0xY+fC/uncAZJahDd71hMSaZ
DRk448qcYXWgjsLzSROk/FLcld5gmsn70FUjIuNxGR+H0st3l2fnHtjXYsm5JC6y
ypaK2c/UuXl5kJsUzvdQZMxXV+JZi1nYssppZBoYl2a6kbwQj2G8bvS+nf8zqAgn
kxMETJX8KmIhIg4ZU3bCGeb/Z6Z10EzptUkAhathBKPljVJnRwvBERkfvk3BnA6J
rVRQo57fGY8I71l69nwGzK7wzn9dU+v/cpxSCkqusTFU5l8xuhhDJ+4xtgfHJAh4
yz0FfjfCElJyumT9AiYxLuckJri1qQaLr8q4JYmsIU4/gtsu1SlQDMpfHNAIiTZh
5O+qYlq/L2wtX7b2r1aVSd4ysZ0Ncg8MZMAAjleHYA0qypOY5eJdPEs4TAAJUKLM
wrSQeKFDuzv8yRw7htp23v59Ls8Ctlbk76O+oN0rAU5Yz653ZSKY3AiUw5mYBSec
wFJmd2MVHuaiyfBU9oOyV3fQp0G+0akPgrWtQhZtTENPU5UfP6Lg/HyEPyi6/tLa
TcWppBDy9ds7wwqbgSjpM8EwNtbr3o7fET8mx5qrZwKgdiLWsnJR4avb8CCXPa7B
ovmyrlgATeWNJrKzs9Rp8kBL1f5WtbebUxC3LTfdLIJ2RTWsDgT1l3QHRYBjmbk8
8Z4f80zsF0viHQUl0RxQ79PN8XPlO1xo6Yu82ZwZPeNw2MlkvkbnBrJg54cLY9yI
dvwAxe3zijAfEKeRrrJ7NbNG+CPOOWtRO3MNJeR2ICFh5ChNWmRjrqujDbUP4nCX
be3T07sqgVjlU8uhc2e5gOxF4ULStl2BD1dLDhNlh9QYfx5nj6hn7qvUApk18xc7
968iwpwF6HOu4JkN/mDdPmjlV8/sGs0ZMEjb7S35B+GnUpzcW5yR+E/rkYiZoW2M
Wlsxlt9ylmwnLCy0eNFsB9TYImW1GqHOf1zZvrgb0yMG/9UJCI9on7CvmnNkD614
4TC+voJ4PrIJRcYVwwRyNtuEVZWp+BX4ScWSEvvznuMmM76B7ymXtgq/LxX3czLV
EWlvYtQILIHbqbxL91BShEF6ZPXwE2gz+RHtg/nLylLzWlUnyGorX9kv+gQeoq1d
NOAkHZX+cxuY9WEBGCpJe9wjL9C7AkyyjktySCuB1eaWU0JRVa9kK5dvDv8UyyBn
Zhaxy0s6biPygR0bQSRiGbZyXBBf4HOG9GtpDNgjR+h5egRnt1G7zmwcZwM2q784
YJ1vYCWlaAtkejcZRHGPvG3+8CTrWVHak/kfk4O9oBlTmiTrglTO2igllQmNIxu2
q1q7PWaBPrFz0QBj/8BetBIguptQqEbwVbatzNX/XLLbPwHbuloiHuqCY4dLVCt7
IdMqSKgaN207zQ7hJQVLU990jy227DgP3neI5H4g+4Ty/qVBUpaFDnDNpHOgt5ke
2zP+3H0a1LmZCfpClbEYPZL1PXUQzYEAehD81b2q3nRZWoTsP5sSf1IMAAhdKPvN
fFu2AqO4zDq0z4nl4Yecr4qh0tt6jaMfues8j63AVjU9LHGKbyP06aX7ZsiUyUSj
Z1daq+CgxZJx+7UTJwgIaykkGHrQnmBm+UKVSVDoKAhZzNvYki0ihnege0WfA3Hb
fqn8mycVmyjnaXAyEtHE1mlQC1vpgo7vprezxvxO4LCsu9blB53s2ap+ZwGcEtta
uowqMQ/oAyRd8ylAc2UImg1UU3/WMJzj8SQUahZPULFVpsB95jOv5kmDYwMq5Af2
lk1gricfKig8dSbEMgL4Y0avAZ/EN7lPqFPqb0m4hBT8XaudpQ3QSosPvtJNp6ln
XWmvjOVK1fyimrWjYTzTxzS0gfmRi0X5sc1/gsMOs8QyVHcQZ3T1kW1XpHHj88aW
ZTXFRbeiqO01zO04YGL/GLAwehTNkK2G3Lx1sM2iQ+wuHapxdDgJNAuJt+dWrpfW
40J7ybkW159Uqcfo/gk9OUJNy11tOPIzwc1PVJ5r2A+IRSbxts5jJmVr0L8/kPtI
XOGHTapYHUS/AqDEvWQgYAu7X3ZsRuUfO6mKblcprb3Q3PrEbz9KSQoF6vmNdTmw
ctXuuUEfikVp6INHgr95UANq6Y/8LWaUP6bsPpyhDiCkt0eUNlTNMyphddLWLHkz
3vgCOFCg6ms6wYi6lUy/tcS+ygMsGLIfZJrj8UjQC8NTuOAG6uv0stzRedIh3He6
loY5qmhS7dHk2JymXPmwuUiLOVqOcgnY+lJvBjsJARyFPatE2XrM3FZehmnUj++L
y0Fe7WbXlW8inSCoj5yaZgM6RoB6/SmlliCxWhrlGwUrT8LYk8VQdqaWQGO8YVpY
34g6gAP9Mkl11rcUsAGubfi4h/QYvt02COs+kyh+zfWcKa29uFWcORscUR2PnWx0
PrylmGy2Wst4PAcuNVE7zW9ZlmqRtpFWEnYc8AEj96osXzdRDxz3K+6u31mENGWE
/UDVOIvUib+Rp1YMucn+xR0gqQyQW7CP7AWYQP+busMEcl/R4b+BTDmRoTQRgLlv
NcPeckHlXeS2s6GZ9dkjG56p+POYlTWqZDPO5yNTiL7AywEMlEBsCa5RM2QNdaVO
jGecYYZ50Nzy7JyZt0eG9jFBjEmUSZca47haYdPIdykd3lYTAaImIyqQhxrEVfsI
cLqpseZvuND5BczYgvZgKc95TCRWJeKFK2qdKTGP3liqW8//4sjvZGV8qgC1Lv7s
D0ALZLlk4Z8WGngfgTC0dFkKyek6fO+Ry7bIoUYba8yn/Qp8uuHUvKNQe+8HvC0r
X0FDa3SV8TpP4wJ9ebtOkGRcd/DzzOaEpShBeRvAu+koYh6V7aX3ZlwNaeqsIkrP
Pymig8TSzrmVq03nI+Tc7Kf8UdjKx0nMt4O/6GLBKDOvxmcWbBx5oSET5X6o4d73
3AJi8jBuANsgpW+fa81gS9mHx4fvXQUcJysMm0LCRZXkhJuJbRP0KueBHPvbBeTn
lmUZJFi9r5HlOc9TpxBM9vJUXGTwMGiqx4TzYk6n+BvNn7JXJ5shQ830SIZqBQvU
Ek0jTZdYMsip5wJDlLgBhNlWFL3Q9kwyr4QjZ+xzhrjMOi85nHvbKuI11F8n3xaH
ugq2aQpWIOCHMnKisHcyc2TlxuGx8/62AfK/R2e6kJnTeNo/EMkvJA6/yjtDfpzs
fjsw03jJc1weA5hxV/Mw8mb7YlQVaB2JuDsZerch4E7SpAfcmWCVqA3xAOpxG+Lj
+k/T7tUKAHiZfcEMreUyP61QULvdJ/FJW07sOa1EQyZoc+5gcAC1WC5ji+9kjjvM
RHsXWKR6+yb6dMU+t6HTty0GOghPSeoufQxocCN/SF0SXjQQAF6TpSJCeqymcIjk
NVJGFTU32ECYhWz6tAHaTbGfjSVTtdgOHR4nV+jz0HlKTAlLJgaQMivPLjTH+Hl7
LkPXcWobtUm2DQojbafHl0ODTxkFUCHr+xwnjHiCE3O5DwBIg+5QMihUF4v6yu8m
bWcNRfod/KOfpKbybxpl3U16UKw12c/IEiGLKMgt4xG8oIHKGnAiLpuE6OpcAiLj
1HJwHbGRrQ+dLOK5ToBl5R7rDCrCF20vrdKPdgCb8VHVkPIPI8CDG5z0fsI05yOH
Bvx7wAAbbMf3G3X2PJ539kvKo0IU83rZi4IHcLsEYtMd/MUpzP8DP7bvviJk4+nY
RYWxAjR+ILv5g4phwp3/IA3sAzv0ZmamVtVZL8UnDxqONKFXlTPUXXoLc8bPgoW+
vmEVu3TKQ4wxou2dpIKaDiUKV2PUzPfCDrkmg3TQoZfRc5HFENACbAxTpAVXlUdi
Vn9Hxo1bFI4EHsfmOegZI7qudf+zrUa2HKIW203onwUSHcT1oQVbVi3m4Exc8wDB
v6nc1DunPbJeJn2VTVnrSO+ZPVwR7XCi3IifNHTScNqACjjLo5BcXuAoF+R2Igr1
qUZ0ejaxh3QCxgcGRGHQiX4vDZXjx6zZZkdVFnQgxIwVHi6ZbYmZ2jYM5GoRzXhf
MRdlXRgBEziVoa/12r4IC08kdl8YBxbsHvrQvYan5ZfYrxuFyySn/5fbCXUoT+ON
ta7L3DeXNDBhTgutEqswlD1eAG8rFlTV06cGAvqMrhroJYQtsDZzmraPAqoip9xy
O+rtu2mzYv+Sq5RymtUtrcT8IA6pcGRpX8YbSC0REPsWMTb6nNFh2MOENjsP3+qT
vijkH0helZ/PN5HtvgEghaVTaDYmrPm571O0oPcNAnq2U0abVge+FoECvPkPsUR1
+zWZEBc3Hf+bD1VhwS2GhAG9y9ZPBf8E5jeXuexG6EtyJ24cpJyjigVUr3aAY6GD
IpfDKFSXgP24pXsPd28S8zyXhFGiYkRYYnJEAooJdUhUtygZQaBYdp7dA4hbJ6hN
209ouV2idKyt9Ga3FW4nDKo13UVNKUaAEpJUM02yv13/DWPvdliS7TtYS2hhAMxX
QqOSXBjPDH15jU40GfGhsd4q/Rx5ODm/utHRb8fj7CzpnTazD8JGBGIYblPpAbWz
f8dNJ9TvgUluwf0kuADw7MemUbJ24/g0TXUl2RrpGZeTVUK1dGpFYGUBxx4KSLBg
ksuYpb3GlfQpdz0COVHn54EyKarmz1e8XvTr7T3StwOtDbTSUt25WMbX5/uN25Ns
FYs1RO5j3fAgivNVmrDvWJAEXPp8rhUeNznlJ73iGfeyqjjofk7GAaKMcCfJwOVn
0so47SqmLDldlR7fWxTwhu3ZzMB0iW/uxv8f8zliwXGDoW+vqJaaBJ+7zKxsJAsV
HQash2zMmLK93mVFQsNhc7OPk2z4FD2YxopsLuj2UJuyspLtJ5jt0DvLwfVRns3B
BuEx5DhlIkLGSZN0xKkO18zNaFPvEB+nUDr6hhOVHbg/JkcelQFN4JIzuoFd+mgP
mXJCUIXtNGFmTFTXy6ivz+zK7vMiF+U2s14BPg2QQYVV8Njb80dKLBpSWdt/UswC
s8RDAtALgGHMd2IePBTKznqgpcO5PhE+XD7xaOxX6E+L4eHXxdUYzNI+HYqw1+Ox
IpAWG3FtQ5XgI0Q3KoJfw+L3XPUvgWcvKumrQawlU1ctfCcOjgi8hSvJ9VtkdYis
yEoFWSVenYlJqc6BBMwIvd9tFE23BUDPMV2sjyVGBzVDcX2g3awp/B2Z3Mu2SS8z
TPU3aorTVv69fDgDobp+SqcUrEdFOEJMf8EmZE5ZuQJVGie7vdk5b8lSXIAk9ABG
WwGb8NtZAVO+gsB5ftjOmXxihteXPY0znPmPBrlAxs5DOO3vtF+ZunA5qufet7cj
4CRQc6UN+Eon/GV9j0NeDpbgu8aON9T6Yrw2DOFtnkv+7oL50fCGKYzMDIrFIWAL
5kvgCsvJ5LiVDiM12u6Gn1VvQW31DZrqp+sWySUt3HGLrd8C10ysTwl8oJrBUoYT
pnIbHycis8TydYAFM6idXQYJNqoYj25KQHbEXlk+8sIAc3vtqAk0ZlALQE8hwRHs
tdsAofWlm2lU0RHU5WePx1QIjGGdmO98gZ6WI05KDb8+7Op2BnXR/LT4vI5p4ruL
sBAzZXR/cVSpNPsdw/ANnAzY+HXaoNfm5JL+/BD+aynXYISavbF2Ng4pU/RzQe9C
LBIMBYofENvB3W0x2U/e4eprhK25XxlJmPRRWqBgJ4fdpxtmoxiVV3KAHPq0hE2q
3TH0q1lEWKUuQd2QfyKB1A59+S9o0gViJH34AQGujTzpfOxjge/0UTlF4hvBViOh
A3RSzQ6FglKZzVlt4E+43Htxeav951A4gm0RBhBEzUJN8zY7r+5aR6OwRuRmoCSJ
7iWq9eU0g48iPykPGZFrfEedz0418LllafqUd/kVtzYFfANNVDR1TqfYYULHvN4y
wf+k48/jkK+A6aj56hykCfpAvtnCrebWoLOj+BDrpIz+zKEywoio68hPp+8guCP8
XhdYLUjkvGiy+DrMjmGb2AOoPik5A2EhgJGfKx0pF0SMHWfqEeMqwct8ATS7P4qb
dX0sdwo8Z9aEeZzPX+HrzDTeMfHPc6vusqGM8xt7L7o3PQ6jWl5tUCML//CYLr1e
7E2Z0/NgzUMOe8Yd9Co9q+k1MqszdKSHah5bZ7L8Mc+nu2tyl8FFJOQHm9e6wNKw
iBK/g+J6oertkW2WluLz4Gfx0OC3c4NUtxJ9TKxPhrCl/4W+COKcctq0SujvR4DI
sCZNTU9J9IZX2Tz6l+BxhRSFxiEecRYaa9YIk5UY7N+4rG+xAqqkzR1RffbYn2uv
sUll0CdFclBZf0ss8BcgyDOdn865pMBAoxpcxtKn7rOeD0/V7n4HguIMvoEtBwLk
m0YhcQRvSNWGvhcadYtHYExmZqM9SDcda1AqsmGSyuRLxjXVcx0HMSMh9GpW/ZP9
yBENwl56fX7j9Z26sbHNcPaDFbDa/aH5HTkwE7vJ2TdZV3zEkveTSemZFAFN+lih
2hFvCJ8M+PgoDa05fB5fjoJKi++2e2ovbIkPhGdbwsYplcXaQ3tEhmNUI6azFgqE
BMB0Qyr/+DBEIn6Y+NTM6nY2oHYGW+OIqMp3iDX1cy0jfa570YppjTJUKEXNqxgY
VAgu+zEC16JGwIZ8S+OwzU64uJ12qUrHzxfrmVLILnEr1/qYZSDD4McRXnPx2E5+
lL5JBDATK0Sj1f6paJ84BmXGOoy4cHprvCIpTDIVWRYP2bzem/zQyVuUzYvmLq9Z
nUWVzCLCGXIJ8oYYUXWyIHh7ZsFeDU/b83iTQx/Oe3XifzXQTqoTa4rSbV1Efsl1
pLNrASHztK9CaTUqCO/+Z67Vnwm01NaKcf9pF+THeWyy2O3cg6rHhWxEBnhvihqV
ywTbB4Eo4j5ger7r+zIQq1EJALwjZesr3NPa3VcVr+0dAeUy6Td13A1HwD8ftU+L
rNM+WYuURduD7J81bdE2pxycuYbZptU3AILsgA9vqsQmEL9vWBxNBACd9HpTMXtd
SWLQK77XuIkJ1vKycx+BcnyQTFGHpdtg93kgE/prOTE4AtWLH7do6BGMbOihxtfA
1g0rPR68Zw1l5vA9OjomYIMbgnc0BwJhqS8NfK9hyZ4AtPNESFmpUPDwPUWj/A7Y
OoqQsj6O8G5LiLXReD6uzb5Gao1KWEn5LGnuYjJ4Nsrs9Kv95xNQ10Kw/43FsG1i
YUN4X/pa/niADfZUJVWtvyaP64E7bCf2XJM1dOE1PHx4WI0HK345L5oVTbGilVEq
A+/9C7EQhw7xATtVXtXs0UVQ1RYbJ97wCt9yvRmgdN5v+y4lAD1Z++7PpnfRILa/
LeXqDvw4mDQhQONK2K3VRQZ+oXM5C325sclazxVRFarXD2HqpDfSVZtPuTwjTWFF
IeEg0VJ9QpeZmVd7Q4Xh8OyZFmija/0z1NMpOuUqlwgVk2GTNtLOtTew+3RTHgG0
a9xgNWpLobDeQMphXjhhNW+GrlExQDIVrHFOCwI4kPoJEvz7E5+kTea7STGEnwkL
93exMbWhitvwYknngP2hezA/tCiSETN/RlDdpv0Z4i3nEkWd62NDckDsP3EBoJK1
jpa682BD79Db6xv/2Iy5kzBIgxcbWjhArELl6pjVXU5FhPtsqUDfiZOG3Ct8d3E/
+DcUiXp0ILiyK55+MP8uQAqVv8ogk9QzfKTZtoxSWv9PAHFYIrM4GGpnMfbHS6sa
JT45MDIFN5I+bkG7UcgYHf/CtGYoJesX+ehk0lqBvWo98NS6wVGv3ZYqZGX7B+5G
3MJBCF7fIE4C2ezGrQak6SUyoUEc2AftJxxbzfBljxhKeKy4JMGi4xW4Zf9wtQ58
RxSOPiN51mboI15x0dUw57C98z/TALjh0U63JSoT9E+zJv/qqLItUoFSh9zGNT/d
RysSah2IXYWBNVHJ0JPYezFMV59SFXNxrqrM7lxdwHnpmf2pBgV/eIrMABZpw7My
bC3mlR0UyLGwZZGVJ+wtvHmcIbSVTtCGmRIAA7qfRKakQr+WYp0kli1pFAeiWl1n
7bw+IvkFtTCMkkvfHVVzIB3L3Gp6CX9Jg8Kc+I4+NnCAQ3LUV0sp9sSqayg2tBlr
PzoyvIdbSa7Xz43qIxHjXOt+m7CYZcrPlgKZ3Nf42NsPxaOzekodywwjr2R46DQ+
SxImNtPdaHLqa1j54dSWhpvb23kyc5LT9qWH03hNz37NBjS/7vUI1yVGZVEqJ86O
KTOaU8BHWVOc9YOdp5rb0i0r6VZIPqfLrsrBPTcN2i/t2Lz3TD62i/RswGoSBp31
1xc+u2J5zExjBaiy2kglu1W0dE6CBMv2+AkQHe89ZutJzc2CkmDqMPinTxAYEQIR
GN4WY49WzppbLlzIKTH+G/moV6MzOXce5Furvw+VcqRs37l06UdJC6y6h3sgXBZC
IhCiA0c1TnZWzwYoqVqiOpZZ8Lst/Kn2JqwZNWVM6RH99C50Fiuorzh94BA64jqN
WH+vrOJjd1qmOgwGw2PFAOMvlZLbUDQ/77FBlk3F096EZB+DxFeTsobO1XXdGRlB
vqbtybM3W+y+5GUsKCcM+jlCna7MjWBkjllkTCGkgGKerKcWFXY2TO8OaPkIgyN6
KizojZYlVHg70F6WF1iec9uwqGjBo7pYKjquDTF62MyOK/NLSxt7SLX2rbnynwPi
+T4aZgpywWf9uU7nQMUIcN6vFczYLOVYMA8givo8LHXExBhpuu/1kzTHFRoaatXr
VxfRoJ+nK0xzqykwVsKD9k5jZHt0d+XYuDyNpYXNBZLxTzM+j3fvYVeKAsmpAzW5
mrSQBxNA3YXURSOxatX7JuJ44Ak2/ZKGccmk9rTceyJvo1xSr198Vy9BkA/xqfp0
LsM3q7154WluMES7SLJg8nklbMQIyIr/AgEbtsMehMS7zDUNWtZsja+XmHwcpQaI
/EGJwD6SbTcPklMWWSmmLA93GrsBBOjObfpjYnShaXydPgCPYFVf1UccGLDTHRiC
kzh7yppUpJ17UA35jQVyz4U/62TMFmGGRxExEV3kAY4mEdCeKP3U4BoVdi8rk9pg
Ct5M5BXDclma0mFyhhiwlQ/tXUX3O69kopRGBgPASQgyyQ/8g7lBPQqcv+VozeAd
yVEfzHNfUk80xy26fzsEbYdnPVUVIjf9dKJFImj3VKeo49s9xgr8fUYiINtY3UAt
iToo+zt6FYHs5Y+5KmefnkrnhYIFdruKdd4NbOQGlBqKwgk7/v/0cnUy7GEm1nOA
1m1n8iu1zI+Kx6+Kr5/6JvDcJsoh+3CI3s40brKp2xlf80IWbZkadtuAdQetQ8PF
iKUMjy1QMje3krdKlDDMSGsw0GmyxvHZ+sUPgD8DYhSP4TqoTYuX+KhvWxR3ltCm
O+Ybv8RtN0n40Lrmzr4caKZH0zpAPhGTHqJzZDtjWnYELmhuRu86D/zwAghJchBz
kBcL3p/GfxeZhov5WByvER6A2ZUKolvCbCHVD+qbB/rK/1cJMPpDzO/Sd60RlzEM
gfd5HdILxAEdFY7Jti2h1f2wuM0LLcNemr/j0yf7fEvSJY4pq/xRQ2NYJIgaDzql
69ghw/7Fpejhwvww30ato9bm5y0QQMvwdLTPXj+4MtFjmTfbvtJW9uOOmyiGGqsO
GKXJ4GYGW0kfX4Lmlup4inqaDxRqSGnt/PuPAy5UVZQ9PFhWER17dD0APfY2cz40
G76SBSVXPmc9a6alG6dPCTcu9vu3/+VyFEA4/JQrG3JPd3pEY7tpoIFWwmcZIcw8
qpEfZgGccm/2Vl9yo8fOVzti2zuONVvnl+DiEZZVaVfkucYasDtZl39jsvbCcc3q
fo02/vUwrRBiYA6bMHYctT5VUG3L8Y4SHcipEWBeQfKKYLs/M18774K64Lu+A4Cs
WzCuzgi1PD9J2kywZajpqvYHn6SmPA/FTgWfNS7jWRiN6VOsa1tqu0+ZUglwS6fl
cK3FUwQwN650s5/J+x8LARGAwoDZetuomwBUvjI6quJpJX/5ocZZHAYkK8LlxGgP
ZTybGbP4Gp9DHmAeyOoF6iJSFnIApyjeIW4W/Gj/vYFhCkH/w4tNabRPoy8/C60f
PGQB2GeVFebLsLLUBGtRzTH6wRAQ0DtL/iesUUAcROARMskZW0+GHdezBaGXKUpG
qe6K61wSrSUDuZZpb+F+oeZPCNALM1PnFz8eAK3tgqBdYJuSrfOS6eC5mmcFzgma
nA9DVKyOzezJUUV4xXmNJTf9LYxMwmWlQT5FCvJ03AGvjufAbeAEWhBA1azXzXK/
CezNnX8lFcfd6oySvAcVJHOZ0sN/rwzflmE+YP1IZ08oz/8WeilHr7we/kACU0WP
RuRD2dgkQTtgCn9wEuB8ZS8aJhgiPfT7QJHXSSY0z1YkXWNAKSUvy8ophf87KE8x
/+oICb5Vh9MygbmndMhY+1dy7C9ylh2v7LwjIWLkHupKzgD0Ob6/AebZGQql67zz
QdIAxgNU1EFtmSvq5uADc0berwCN82uhNuommnMXnDqrDjqrZi7uMaR5471rYSy/
7P5p9GkbAU3+WlpNVpFWYr+9+R5TPBtjpPi7VTc+AK20o8j84FEuhQeVTdlX/+K0
RibccV6KXIkbc7wLREMM+/Oz/YJWnsWivEK1RO6ua5wyWAvgz5XOZzs1dl6b9TT8
/sog8cPGso9XBmFoj9cCCb94BrGAXzst/OYOF4EHOLdr2LlUhrzH6OrJShZu5z+H
3t1hpeT33WonUh3Z/VuOyoJxOkTVfXfE5N/PVA8BVN5PTc4+6qsqXVw0WpY6neuE
wGCt9HU2sPEbZpdRyucCexj7lxcDErqpK0ZPfODEjQOF5bWgbN0WXT4wKg7iKAJP
XfkSpFh1hMz4/pKHYRjo1VXjia7MTTDHC+SZo9cGGt0YIxDOAqaSZtpfzuP0Dagh
tN9s8m/q2e9s0i5eZboYo2phidVG6AHKwOXDupBDh2bcL0n0hVD5hOgxsBIpwPHD
TeQ9+U43bbIt9y3ygfadKeTyqPi7IG567bCRHvHl+tT0TdAJKeb6i1V99zHDktLn
ml7W7s3pisQ6BF2DH6avwb3Uzha2Q/B9GbrXezlQzUw3dk8umVGBjXVMThj/vsQh
5U/5IQT/HTwRK8dieYyMWzjJXuvq3brMkX4CjTF9fqnZ+rf5XD1/FCWP1/cHs2W/
wmH16PRMfsDVMZAZnjlmWlf+JLyqtiDQH2YgFQ73qhm9+VgrtUeuRj0knPrWWiX2
hA1qvs2sTARabQ1JARCdjSvzXbpUxXXoGudllSUHHKm+apYlfGNXqSvlkpoAubP0
LGCI3vg2w49RU7cG2jsV5pA3nts36ufbIzSYWtQ3ZNViD36SqMogYPaMoZEJgEAx
Hawq4VaSWz6QQ52i+TdeimUZZQKVe2Bbc4/pW7aE5pldxQSDu3OxOzfJVh8nb7u6
XSJErZ3Uy7qVRrltRXz/jD2+qp3CjY6SmYGghICgK6tekRiV2pv1ivDQ2us9o7DV
X3EV/qHRloQdwNueCkVPLyhVGq4Y+sFs2jvRGUvdxVYxsJDUmsapelPAwf1Js+ad
J/AVcg7/3AGnuwQfLKeGy01UepJE6b0b4ioOQoCDAJJRnMX5cOxV5KYmCIAf5xx7
0DjVFZ/dHpSZrPrGFdCSf37bryu08km1BTmGirt/3K+wPDxZ+2h3Ylm2NhvR7ZZX
JB6Jz6zn42S02H85hvieeiGb2DCfLn9fDh9oodRAqW1w71bpJjhy+6Lmp4zzP/ac
KLv92ymJm1Gz9gzVdmMwVriIvDbGlufq5lyMwREc6QA3V4iELWZMwTcG6SaVHkBS
qaT+sjmu+pZ4x+g5NQqagRqKvCjYH27y5nZLyUwFnAi3fPNxzWlffhid6lWeIgHS
wUCHn9Vt5MBEcajoCdrculQxgmujJSwpgGjrlvOWXZIhk5V1zUHkjimKs5IdNGuB
tfhjxCE0IN8PkqBiaxRc40BC9DJ0smWoIfE0q6jxxdrumfDpSu89hq8PbJfkwRVr
1h6uMIb+85lu8X7MnFV9A1+wC5O82yl28lgyv8BnhgkYmQLWP5Ovb13fZVKlCZqy
/pDY5HgJrbyEzBcw0HP9lXJkqVrMOe6gX2OyO6n/5bKcohkoIG3kW6gpkHusJiEC
qDZjcAB+JYRnYUHdVTZ5PQWB/O8CBcY+7kYygtImj/069FIoGmSSr0C44mHZ6j1N
oKPe7X9XECH1l5nLWPNytT6sjEn6lwwO0iKmXSA1TiZ5Dn6stlWf7/tLsd17BD3L
L7A1VvhsQiBrAKkyAZVh/MsUMMdp1JwKwYuuMfqJ6b71IvNPdTb7P0+agkShVeGQ
GRRDU+GWAQa83WtNMKSYaAyHwi57nmj2FFrsG0NRX2qPpUXh+VOjUwUBBFjHvw+5
BAsIQUqadCUkoxGfCcbpPudOLDJ8OH6Tgs86h97XnDWqLw3q/ZxtFq+g+zq8oNmp
2W2c85bwfL15cEBfSCI8z3KXL6w34ZRbVZQicot1ISQZ2dxTE74f0tZxDAyChrp+
u4U+XMHWjC6T9e+L7ZcWHHr/aVHQPX9YmSehEZGpGiYHfg5qypwJ8rmYmKEXIk5o
R53VaONuaU/kshUiPjfB8w2HYwSsIw4Q6mgpvOfmW+1bEjJog378utZcEeWNqwHG
qzNKw2uSQZd8LzsR07IrDW0T3rLlXp+LUAtCi0fcH4qg3ir6UJnaq5HLkC7AedAv
/BlK0ZLipxyXkJy4wl129QvITuJSI8LCZMxf6o5HcRZ3ab6iMCYBfRCJdLYvlVXi
BwQBCk84BphtGoKTGZm6TSOI4bDA5oh70dYAsrNH3kVl5jmDKUyqvKy5KzKc5C3e
etjJe0k6WogQev4K7Ulo/Ja9mQsJjiKKL+nSK//irtMa+irXM8dMP1RL96eOVQVe
VeyyQZeMhfcNzHrUsF7jzZtJeU0cR1r+LxLmSRkhx2ueT0y3jx9oE9e+FL34bZdA
gEwhhvijr0/paW2XWiqifc+dtMNP7XXXsr4GJSkqLCaFi/6aoO2WutL4KnoGFuiw
NwF56yuDVHKovAIwPnW+8BvGZl5ahw7hRAsTBxBySgOKcHqVkcntExOZ40bD8Ia3
7lR2YxDFITbImDRl0Iql3MG9wkUQWpISeikE4AXlKsjOBGmmamI0533E7TqDSIGk
jHGNYadd7b+eUeqxEuPF+D0abyfv5oZyhQQQL1Y8vB5tCYBlD9c5qKYsu12zruwD
bpcd5uyzs+izGJ8gWpxsQrPXyawfaEl+b4EOw0Kf7/NxcAh6VZXcE96zM5TsLwlT
B+Rzq0ZCF1IEC64EpNO/hkz7VisEt8Vf7cdp3vmAim4i8+zBgJNShSPB8wRa5BU6
oVpOqSEx80iRX2gQ2tHvwInBRDJcGh1QmA5o/xN5L9ggClHPCJ/g241MsotuUzmm
tBD4up0V9GY4kNKKnKWqDB2CqvQLGACCyBpGuBQ2nNGr8lRe4/eWOlatlZhY4z24
t2INssgHFFKerZnkjW8AoQSJF29VChdNiaMbpopRn/s1O/ZMjYkbUThDaoVE/LDB
g/GquHqr4yQosVgRBL5gW4SqxtgH3sVPOg5uQS8NC34jfuZM1HC62stxq7NGbF0P
T9oAQX9RBFIVCGirfFXF4ZSq+j3rtkfOsg10Mx6vTL8dE0gaeK4BuF541V7UcFty
lN3sTM7o9LziGw5GYl+wHNidrU7qplKgd/eCUUk4XXukvZ19B65umcy9D5PzOG+U
wmWiiQaj67I2q4t7eNPtVywLnb7nSCNJ7GcZ2HWcMm0MQR+sOUML6D6is0lDKh+y
iyS02BXXHxLfozRq/5IdkjMh7NOUuyrQ3gCO+BjueRxiIFd9dC9yJa6mRIeaGVlo
Y27rncUY8d+Omtqsk/AqR5RFYEorKUJSxG7Q2eThOlSWswBWikvkP4QdBko2Vq/d
su+exHBH4vDTRSreWuiQmW7R7nZcQRpeH1r7KLgmThVJYtHcvhfXKNVc9GHmftxn
VfvhCqoK7DAqU6ZeGrM4iHapYmVPLrxR/ZqOtE+QFGInf+PYuOjnq9rVThnB0HeE
tB3Mf1CwO9vEhGVE5gZU7SE/UnN91zyTXtAbi73K/6pVMymGxCH16V0wUjX5KI3S
L7h9SIT/kDTztnliILde/+6EFPvmGwf/L9ZmS+w9lxen+s15tKtEguyyz4cLbikL
yAB2jqFUprpSyl7BoidDCenviaZr1XDG+BUmhVTZ7qpwU55yuebVfPcE69cufOcY
sTO2vp2o53sxedZ49dCkPmi3XtNHPnFf6HwbkKaw0+G1epZe1DmFOYf9XD3pAQh2
7oLwNjN2MUeNRrrvUL3G0w/Uzs8qJgMj0EXJNz9HoH4maOGRm805hyJHmkKo5uYa
+YJOPcY9XOq6YXXW5gJkSGTPD5Y19QMN5OQqFMQuvnxzve6mZLFGeMwkcURQp3mp
vDx+wGf4NAYB4B7LJHbzBoSK6yFDVdnXnMYpRPpZ2UfMhQ2FCP7UHT+0VB8+sGOT
p9+RKHD18IbDwmI2rNqo7ef/0Uay5h+Gxv6FzRH9GPbolUITynXjgU1QnVhR4eNH
gX7CyYFZGBGF5hyt6Ep5uLXr16G/NIBJi1D0G7ya1OjUG/mzIBMC9XCpG5bTiq77
UEB/JZ8Ln56mpic5D+unsVt09UV7mVfvOzTj8Tdctq3jv85b9xaPPmU+EmYz1I1B
x8u5vtawwnNucBu1IYL7fb25kFf5+huA0822lhjF32QaZtY8tWCO0o8wMK10w/l+
uOIGcqHhnjZp/4xBd5ObeaN5YuHzBf7+etcP+GYODqZulC6MF7KPFDlDq4bqaTL1
gmG1fK2k+z5ja8ANoldR0lmTRQ+LySvCjnvHd5DhdFyBcFICT9HcPML831sCcL1l
6n2+mpO578IMeWQcQCVeLrEYqjIZIE1Na/+pGc9J01mtyn8kbDVI8txORixNJaCq
vLWehmzsXHN5JRLK+UibIAbA8o2hIl9NXtZPD8JjQ9R0Oq+0IGpCChkTwobNCRhU
68mygKc1osx486SWUHZYlVQ6h5q2Q6lTy5Z/8E6Ov3yUCSFfmvF2KtRP3QffmbIJ
EpRjo7ucuY5QT85QrGSJxxJsAc5LEVicm4QaeD6+rCal9uUnVsdSOFDEv6Pxo7nT
UjnGbLaReTS1hixzJ0iYuIqvTqc9q6DkQ6MMaiVTh+4oU+pW2QwDxPZVH1N8pZvz
JNsaaLPjkZU7fLItrVn8nG2mwT8aWDyjjAm4q91RSyjWJu71m2qhsfKFLm9J8P4M
FrTBIvOSWYdvy2pmqflWGBMEqGy8aq6/aJMjH+Q/LuyaTAZdbua2MDUHbfBiU1Nr
V0E/bb7Ag5lsXGFZrAMZuuS+peZKJ/2kEb1TKlnE1MQKgqv0oMXNQoS+fIQhRTDK
8nw5itZFmVCFUI4p3d3n4eOB6Km6Z6AjRJGWScoNenu4ez33nqfWIyO6UA9LQo2x
tUcDkngc26Ei7Vs2EFIXIWeIwpqUoScyixAdKOlpDLpC6qFBwRhkz69OOYn2FlUe
FkQRnWZ21Xcj27pfTR8/Wq68WZgPuWdmeeQJY18ennXBJggn9caTmLfBi/aaA1Ww
qdbEEu88R0M80/iOL/QWuKjpiCWdxLDThfHJP4+eGnkaQrufXMRvMU5QGo83qJHx
I6F+RiNWY4ktRxatZz+8SM4YExCeJy8gR7mGKoaJa5itAfHyczSEdnffBjc/NwQ+
DlBy2qcVFHTN+YJY+BM5txoCezJOvRX1HmL6db3IQnnPybvU/hZ+d9iUQFKjkVtZ
6oCvVgcjEPSimkHCW3oWDFdpuChqbb3cj2jIFvMdCcWExFjJYi9kVTB9RTU+fteT
d5RWGLN2JF8Kze9Sz73/N121x0TmsW9lTfw9POAGPHjVYnLKa1HFW/xhcxSdOP1t
Y6641TmJpoIs3mJzwzUd8hA5D7IMbgm7MDbDogWhOVDRIxT6YFi/02otu4b4WobY
Qx5OXzULfuPr5LUW8FVBBQhy4E3oACq76UGtPXzRwQ2N4YDUmezjDJhQXeWMXBoz
Ua3qs1VK8SLBPCHslQIQ2zc/f58UmqRNTTDEodAWhVSPW4qcqsmRNZpPFNTRc5/c
oCwFI4tbxySwpUhl7it1WfBa8GI7ekjeJpkvzA0+kP1KwMFWrIMcPyqjazBS3Smn
ET0vYRsfXAQY5+Kw4duHvz7Ec1dH6diD4vmYuUcR6Y0A5EuSZnwArtwSdosfS/g2
3xyvUK5xzf2BCPIQA4PJ44MGFu6ukbCmr6inPPRT95O7mOF5ss6/pSAVn9GuKynM
Oak7wdVmDD30FsXnv+Fk/xW5BRsiRI2nA2k2RVR5BlEtpUtOraIps1utIClpCg1h
3uL3Ipjz5HYu+GdPIy/+ERLMTOa6tDqTOOzNY8jivYdDl0pHf8/TEeyNS0JsJUmi
823EgjVeLKSj9sURgo9Z7gQZ/ehCj8ezVXJX8Qv9YMJZln7K0ofQZmUoghQpYHOV
+3M39wsS6GfR4Mx7LYfL7z8GkcI/MRlAO8n9nHoAmfeZjXQdExpRNqsUibCbTaGE
JCdpXDzZimHQRB6gblaQ8tCFRqh3wvHbmW3HZFg+hKph99jvYtL4VwUbzD1Hg9XL
LlQ//BOa+u1bj+V27QJEK7yGy2Wv9Xja99z4lJyt7ucynGjqRZrH0EKhV21gIdh4
mhtyW7fPnUdxMCovnxKCf04NUuQqfaSmh9Mco60A5amsqJ+vOTlkw44sZo9QdXYt
OA1HmfFgpe6Y3xLxtZxKf5NRbWeO3U2y9KyUjTE9VPXCPsrW0RI6vHnHmKxNrDcw
YRv4G4PGe7K500DGCFl2l7KU+odEjqiLuEIncqIBzyiH2/K/Sxk3rTl4s3xyAQxP
G5/N21lnVDlUmnsWqweeGPDA+sdDUoaLeWjEwFZa9WbH2ksD5EkHTu3cTAxXEqfv
dDfy0v1EENhLieNm+ifKT7dR0odRZA08a8KUuxi1Ri5Bcn4uVCgWIQoztdyIlAsk
qNAXdLlKYZuGstPsWTxpM9FiQCkFtvVnNn1wNXRKkXRHPeQrCkUlLdFoMjaVnHOS
whYYoKnqW+BT5XDvz/kzo9E+yz/lngUWDMNCBu/P2XOvBKJ62y8ak+Jz5AZSTVO1
Vz/L23Hpavf3PncYAk4svYqTUjMajuwzgh7i/U85NyzzWQhOEeZ/23OabuLEiuMJ
Z+RuabtBUXimUDeLHmPXwrYECAFTGWm50PE59BKVoG+MWF2d/iCUgmH/GQ4eM49a
Ir+ZLSn7DwhaSSmXvyDHuKMpXoHucvZ49LtwmCy8YwrLdYav2t+TqUTT6vAWbtLT
HncoA9sfNrEv1jzVMieGgCnkv3fE0huqVLQO//Kc5SR8CUrdPI0F3hpi1+KYMjMo
kpl11QtTEKQsLViFcu1aU3q2bfktna9WyG4WBAh3+UrGmP+zMFEWrm9Cgss17jgN
5k+8r785d3icPaWk2rLpxz/91EQOqjdc3MyytuwKW1Cjs/VqqamOYjWQYDxJYt2P
kK9tjwmSVTXNc/T8/ycqR4DCfR7HAwqvglbnJNwqzMMNfsKagY9QY+vOQ2QrwT9N
0sffRQmx+eBj7kX9oqrcx38Unf8VGsshzw6ZjL1ziCAiV2PYeKhJ/ghp0Mlbf57b
xD9/ZXvWACf1ZdDOX9ZJELr+cJoEvXi9b9x+aUWNBGeE8r8bg5GLNmfuBdRb6R5g
zj8ojKpbUhVGwm3u9zLfbx9yYJe7rO/19YanianWeLGiPGt57CiVb8PLLHhVEuU0
PjCb6tFxfPRZYX9jkI/cNJ65Dl2KQSU/Hmy0nOwmAu3u45hGcR7GmADOIW2qeiwR
xQq9I61wWkDRhdwnDTgFoJw90O1N4r2qbKGMUNm5VquTEIB6ZCjeAXOfYVRg0suD
9qtkMX5X82I0XzPuWHy5OzMqSn8Wp9bd3Mg78msbQzr2OQEATXpX1LyuOvx+CWZ9
2UM1sjCGnuwQOePbulz1h+3v3wZe0CQhLY95Ey2MQ3XFdBfzmBiKz0KqMWVHqNAj
KQg23c8+26kjrAOAw3eNsarOBf3OGhlsDFqHYGNVrBl4uhgYg7RQkoVzwjS6e7Ud
2tg5rOB4u4O1RWYmc5xt60joft/z9iZqRvTr41Nn2kumZjFwj/9eOokqrEtUlIJ1
gPCRZcruZ0V2YT899DhGJbL8kzEaGUgO/8apyNYKhv5FlWUhH16zIckf0m8ktuq9
Rb/O3I7p19dvsaBRu4/eCg6n2m2R0fLo2OdhfwHrVww5wZSmM2OTyM5QfC6r77NT
Wp6JdGcwk3hpgfKTtUgl+wINx2/s1I4do4aW8rsl+ypjgGvV2UwH62XJXjUO0Ov/
y9l+uuBK7sHYQjqgeIwNk6N8EEypJ9dmMMhUBuZ26dSlJsvHYd8rldAd5W+rSR1b
UBr4HwUhDPfMzCd3XWdrwqz6IRVURgV4ocMNBDDAbLclQ4Mvl+4M+jFEQCGabRrm
jaAqn9HevWD53esl9/v8Fz6tb3+Yq8h/XcWwUVKap/yoXKrHaPKryIaFWQs6WjAJ
GDvYrVgLtJhnMfupH9iFBsx9iDQ/JMuaIAm8kAFqLbKRfp7XYQEViXyul61XTcCQ
A2AG+adQXioJqp0FgpSSGUEl9VYav19JrzGNTJpF5Z7Kp9j3Tiqj7RBhdS8ULT8N
WGWsTL/gWS0fx4K94i5CM0AN2Qhz8HrMoeOOyexXddL/oHfZTdrAScw+EAyPck+Z
c4Gzp1mCVW7mcG3R35VCYFB7d8kVKhdIFg3ikt07JKNkTmNJWzMJENklJL2QokO+
p3CRhomwGIfr+gkN20Gp4AbxvgnuTW0/8UWB3Qm4tb/M1PtilTOuyqWfYMRspJuh
qqUqN2VzXJdyanxCV7uQbqN9RwvYjkEqi5KntQR/72hpW+dgaA84wpaTSYeI0uo8
hMomhgMDzO0+LPwldR8RHlk7UZQBl98JSSbPjMrNTyCb90SeTxBx7e5u9geZM1V7
G0xvTDyZW/IyZD6bL3Pa2ycQhs36Y+gUrQjXhzvAJVFAuBMzWCsHl5HyppYwCUG4
IEP54xorw3/VDM1cfYpJPt/VgsTbsHic+OByFoIO6bIwTMJAdtOnMblC1Tpvp5O1
MCfIbcpmWGUVp2ijuwzytRGYYgjC/CfVGIcMehZGfaHeoud64MwHTjkFUMMnkCcV
HY8JZRu8nXY43LD3RRCPw9LcfP2YDtRf9RKYsUJK7dPFeXnSXqQuXsCgrxU1zvRl
8KcCBkBhOxcftDeVD55cWKDlQ1NO3LwcRY2lMHcBmVFZgbjYD2t97cFgv4Pb/nZJ
7pmolczcDw8/lABtzJArEEOdCSD84mnkXgl+4qp7H+51zbv6ADG0i/rstDZgPe8Z
35+sOrLyA1179Ay5TK9Sz73+CuRWWQf0zn8w3eB7Q2P/EuabdpI+zcz1JObo2IFa
pcz/u3I6eCtkhqxWUE75caJF4P36OZ7LYYzFgqQCmDduOBFlRZjTJTjLuTqGHGjL
HTsHg2QxEVW7gn82qBSF+4l2tx9aLJOrGfitraMA5Q0dEFFB+utgnj+vSnh5PV59
qXRE5ezfonoxDLXENX3Abjc2HMrxlBIEgNGyOLKWA5lvoLuhdeu45eTKEW7+8G1f
HPlUWLjbo58PYvPuwqiOhX3IYBUcj1CzcQoCjKTFviWhNqRSGQeKyyYERbqFYszh
rMobEKibOfrhQx5dFAyaIxg1KDeV58XVRwg0/DOpHphmAQsPx6ZmI0/ReYNOPO3L
Y4AhjU/rel9kAH8UFIkc4tl8Rq+XE4ZSDeMrz8fy7h32nNhUjTsLm3P9qFtgDNyE
qVxPX4P+cLKyY0i7Qxt5bBCyOJFlouJeph06zKyJCLv25hffHystPPxUQXmAM1Ax
F7g65ArftDKHnuEzeZGPHmeFlMrt5t/oJmOCNshs0pJsO0Kvz1lg3GcWysRN+IZ2
LXpEf87JQVzVLE9ENeG+XEpt0S/WDjbTRqcnJXzO8+RgFR3JfwIR7+xhgxN5QSwF
5dkaq/rPdS43EuWQKf+c0LFNxvzyVChC+MDKYt7LgUZHRVfqf5CMxyyVZaTnZ5ck
O/Ik5GiECcPibdwkTEkh9idR6fy2xA6Wdxu20pG7aPqh4/hBhdQMlaYnq0mJCIea
+0mH3kx8bsnzZyBFOysaqpp3pbUmEzwifDDvcNt2RLHkve3Grva7nFm/uNh2sbx8
oSRRPc5ZWU3cItr7yk5ImM05F1QTxCDkUSDeS+eNNowoYZr1U188KAmcW2IUWbn7
EiaedM497OKubNZHTeks+hkbNy7r7C21OSCpqFFY0Dr1doMF0aO55vc+P03Bjqm6
WR+3aH8HUPhCeDu7YbOR+S9fns7O6Flw7KlvK78+Jy3owUJolSA+JRr2BaAAnpgi
ASMYnNTaX672bnHJZGE0e6Fu5+cB+GenPbXmF/8bQJ1lYCwU+yZSbsk7OFlIVCWB
yv6rU+2Z0cr7HC+xQL+g16mCz17PTZ2iHvPi5hROLLYInYks2eEMbbfI6XcYKGA5
Z3ENS2OhFmB0v/1M+4GgZr5aTSv1F2GboyeD2GwHpTwlVVbKjDRG1a8YtGEg8dNH
Ae5aWhkD65cjY7LkwggXMa57l+InXtvX0wrrmJ1YtcY3pBtQ/Y09dwptHwUL1Sr0
aJXuVjT8UDzMFippweWvyJiuZILM6fZymN+G74LcQFKubepLvjygCEbvzwoqH/P0
xk/HHGIAfKz70cXZeRvWOR/bZWGGVXCcdw+WQAyQ7ZgP2bIpVgMMThM9HWgdPrF+
x4h2niB+GP07jEWHzuJRQtOJvKyiXwgk+oQP+G2/tC2aXnUuhMTMbSWBj6Buw23/
mxBQ2BpzGCgfKi1gO+Ml7FqqXFvEGH6KBcGif1Q/7gwxgLvr/9OYWgK4W2YpSjv2
9fpjBusyctUlSiNijFhtMEX6PJ47abaN0ArXhAKHiNZlhNgcvCZqFArvFmo0J1C+
nKT/QM1bcFHF3T0CCqcUJoJw6dIpa+EZfBRhXXo+YNC8bd66waGRR3SBRGV/PRMj
qsiMTzSfauFLfDMMiQqO126zRZcEdHpocP+zmt+YlqnW06h5ibyZRYKiK/PUjfWV
xymjinzrJchja3x45gkxNAWOYqRF0JI+QpYa7xB9wjB38GP+78nT5cU8sRBs3KCK
BwfJ3kci4tD6pl/PTN6cZq17KHrDuCB8pR5+Pxh++IQaEJZdIzr7Amv5gTysycHY
PsKAC2GA/6pnRy62ZlEaHsbPEK7w/JRQ07ZhiiTmz++wpTdD4Jdc7dV4efbdH5AX
8ZspckXx1VpNFQJDREGN/dU50yREC0NASQef3gZgC/TsiHq8TZnUaT6Tdw1xhw4S
GYnIAr0lQ9h6mL68K/iKW3xeD4uSbY5m6svDFP7DkkG/LNdA76yTn9dObBD7jpFo
D+oS1IjnZlRCnRWQNb0+BPt3a7rSvvAY2ZftoqB+vSZbS5rV+QA4sNldbTJc5BLL
hb2PWkXi0YOCNE2oJSJ6yWWMrl10Ui9lcrh2X1p0c1M/mzs/gOYJLfHcJMDkClZu
+dlVweGceY9kjOvAvr2lC/DAG7UD28/zY8nJtViEmkQhkYxgnDTzf83ORq1rF+dp
OPwMcrdxj2OCEdnAdmzueYMijd54U/p9Bl2/rbDWl9Z8gKVvvCwyWJvFCkoTJkzs
qjTp/hCgzxYTNLNQsKkFQtA0F7QIUugOOTzeVrsVtNBo2cY8r1K4rCeEsvEKg+7d
mKUATY7/gFO7EycdW+JGzq2g7+nhrwrPMhaltQpJ7k7YAJnFeCGll630zwH6gGJz
LAUjqTLfHy7DgBfedJzTVoKpf/t1V4m85aAL6TpXMwcR302waGUoGtEQW67TnnZZ
JpkL17/7WkJoWQ/nLdE8I8WZYuX/OdYGU6zdbvmmnfsZK5iVV2EtqowQRN1anABc
lHoyWXrEmNoqrWRVkRtn4w1kCyQN+70pUKX5v2AmxWCB3Z+/KpJ0Vz6Uoz3fTxHU
srCfMq/yutIJ0HAGnpoFruR/1iCNtzS/UEp07//Jsbazyaj12R1ZMVoHWvgK03VZ
zrFpWTZseRoTM6z8EFgenoY4mk5Fvejr2nbc3w44Ri+SROjCqMomQG58zect4Vjm
0Jtb+XESa0QFvcjAbJhZafYGJ6zuiryybfDRByrziPahKjmscCNi2Wgd1KwtvdlV
wx6lzmZaSKsDojccbB8y6t3DRwufleBXwsTsZQ9EF7zqU7aUZq+jUTSaR8CRsDju
GyFZD7WfJ8wMDp9fFz3+Gei1aU5Bw+gEjsnsB7B/TOqTFL6uPfEHLqgVqT6HTJ4S
PzTv4JLPGEM+pCUq6sLHbwzCFTm/8MflJGXOowaoGxaxKqgtbMlNW9+gyc2jsH7l
6wbrxpQ19Je5DcEKZnKN2n288fWwKPvuTkUweHV/skdUBZ7hNnKuScDsa3H5eCMK
R2aI5ftIXZV76ivPCKbSM518ox+xNZAsieVEydd6/Wbcc/e2cyhqjhSuBC/B8Vpl
uAsq3Qipd1n9myh5h6Chq8pIpzBK/XJNRnDXjA4yRWOKykF9vFGSTf3lEdneHNb3
Sv1euThT0iuhK8Cs8TiBx8W1AESe+PoePnNcgqz09i5ddyJYT0wmpkD9lwfpRflD
HB4blPa1rXLKtsMoHuxRUB4JoxmRf1nYMbn9715CkpuMRb31GzukD/diM/Ev9ldV
IMhCHpkP/oc+deUlEdp93V4BhgjIwn4zXmZw2eSl6wKf7YWwR9maON/NRtHlrVl5
nrlIl3q+Wa+JP3g1w6ltexjrPRW2XNKUwLQcMuE0tBLCekF0sZ8f7dA5yhhTuwc1
nymXrm1wQfzV2oi4K0HPfK9H6pL2srI/aiRgr3VxDo6J0uNTnlqCHOTb01fJloOn
uffpSSV8j2qfr3cUFe+ZwS6oW8hO2zrg9FsnbUyiO879TfTqLhEqtTF73EMi+sQA
M+rmEuTNsuPg9yByMI0cZU92qVbiPw6nNXWCOUi3gI5zEec70cnwa7cu5riQLAog
SBMuTiij1r7b9GhY4HxMIe826GIi5gRVvofAdbruRrONahb1EprKXIDa6dsOyB6F
/HA6BWJZ9Me5N5rOCnMdXgCN84a7yQP7vnKYW6o6p+k5P2q5nSlDyKEUA7JkmJDz
t3zzTue89sx67LKKpt+OwkKITki5f/StpJNYo3tq4zsxGHmrCkQ2WgQRfUxTfmmw
jZ+4iuOYmIhhem0I4WWM5khOtwyaJ8+mS4zhgz/fmZxm0yhf26nfHR3vN0VCKxM7
mTySy2Qtf5sbMeQYdeqcZ398fp3sxh0eriUzUcVMFLW3ZBJ1/O5yAnTOTNeW4kwl
niA/ot6lLTwAKb+MuqLbFScP5lqbHxvT7mCoxYR+A8O3SykVLXAmKiMau0xYuC6l
2k87yg+kcUo2sjiJlt5e5K0UspXmDdoTniC4l+/d4k+EFuOJK9EgJ2hBC/HlnODW
cdA2FWZTEpPm6xfVNNMmt+h8iMuhWTZBXmsjkiXKtmS9oRFEK/PxdWdZDDWRaco2
eGFeIYeqPrUvIPOPcoxHeElomxU3g1aWfw24ynXZqDw5PInxgD9fExx+mwSQQZzS
8OGy5BYjI1Vh2w9R60GZzrrm9L9/4pE+8kCjsO7Ry7KOD5nXP0YVnNkkW6dOOL+F
x2+ExstgyXtcqy63FJ/Q91k6V8YYNOABJ5i1bxy3lnf9Xn/byWjUZtRHjquwi+5H
jzn97X/gluawPs5AK+BaUPzoSiUSN6TeHraa1IpE1KdmzIuMFyYtZnu5pGUZU/xr
HoYa/sQcyC5XXrTcrlWAA/YcLAa8oIbo0Z3eog4ZyM8FkoVCbjvAx6mnCggDYLUr
ZvAKHVzmnOAqf/3+tUVUxEQVJxF+mtCJ69FLOIHXPz9uV6mGSm+Qkw40DpJlTYvU
M/RZbeswzvhiBpQX3df7WbA0mUE95rVa2E5URY9im9G5pmSfuoHiUh3b5vsHkbd9
pFtSxwQmeBJb0p2wgZ8PHQuMgl4DluTLXgtqlBbADCzc0v9aGmejgURby7tqzp9N
pKRXpfBAH4Lb2Jf7kO2IicMNVRngJXVaXyb8KF4h+x1SGnXIS/axWNJvLoc98LGl
y8uxwotj0bwETXX0OJHQCY88eV+3OAtzjwmuVO1+qpNwaN6gK8xXkbFVVUznRY2H
lwlCCUS4Q5OmCnjlUMnePCb15lX7aZv7l7CD0j2xeF8OqGZcTpBbhOVwO8gJMYIW
Zs5WYGhzE94HqMyvI7YDIADXVmRDccwRBF+8i6JD/i4mnlxXnyfE6oaDG8UHVNoA
hzo1g8AyUtfNLLXR4ttdUEE6NksS0YBCUh5K5xFUSOb0twrwuTqdBokcS262HT0t
C2V9NjMb4NB6eesGDnSoQfLSJmVd3sFVXcqg2wmGzrR9WkJKimr0CZzPI9r8MGgb
lSfvEIh7SnzKTSzGY61oz0mabL/eNdvZ8F1Sh2HHmCoSUHgTpIP/DEvTw0Dh6ioI
Bxa6cchiG0437GWLMD9N5jhjTNicJntzQLO4z6aOE1xnAB1XOuS/0qDfyTyCNJgh
HoboztfBXFTWK/0w+40xu1B/Gmke82Ca4Zi3WvZv6XA8gipUOmkrrjZQQvhmrQxZ
RrN0837wS854oVNDmR77lbBeWNCapwHh+UxFzv8DINasAn6huMcE7R4GaweYZAXo
xR6JHd/btErc2eYZ2CrFzjbJPmy1LV49t51fppna61fMUZJEGypdX4c4k2wcTeG7
FNJvxYBa/PQKJcNlxubXFL0Ip9oP8z7oC8KGn79fZ1qel+a/3c8EPlYFNfa6vU36
OZZ1iCh2Kk+zk6ukaxHoyeIm2Th7SBXu5kNRoHGEVyo8X/Z0NZaFWdU1xQ6b7KQc
hhx0eTMJ/oKAq1f5r1YtLsrou1WJvZNPBgrxWMjb1rgExsSOSm9+U7SdE3HSYD9z
1c2PlBg2CDrHPlLPiJMQ8GkKnLCiIGO2fyZZJ4nnV3K6osvoDnaqbF7Y+ZB2UTdK
GZ2fcXz+iS8wJHX9+uW0Kc7S+k3TzFRflKvEFY3ugaGDB2gER1oG1pQPUx0ZG56d
CQnIliYrrEDx/uBIp3Lee5BLiCCSby44tShrIi+XYgXgZEjx7skgpMIXONq+AsZ7
KljT7WuVlGYqAhC49RKjOiVqSclke4lwY21Md35ntFCCEmWKuP+AhN58n5mKHZjL
ozOFeoG6GD86XZWpoU382e/an6G9KdpdIko3UGHu9IIN5rpOLPMUCMiKtGF67aId
qBT0Xk0slEXhpbP7YEPiAbj+uOhCIeuPpd6L87x9QVb0vhWEfvbjDpJiftP4VSIZ
khiQHcl3Qdcm2hwXWIHOFoonDoGF4mlTXb0nUPlz5Y6cneSZlEj2WkOSKPbGwTKP
SkN2Jbs50OLta6Wd1rjcx41yUWWgvs43SIPIiHYTPJddEqWXGhsbLBCe/rykN+0s
VjnEVkEQEJPvfBXiwX/Gh4kgnZ+ke7nbQB/oiH4axOUXkm+ISKuXWVuIECX4QFxl
JyDDt7ovMOB0H8QTf56TZy7oXIO+jmc5S7g55AiiXRdJyKhLurf8/gQW9dSCaXO8
3lCoi4OYca9hEy6s5+Umusygu0sJiLzeWH/DO4UEOgIVpkIJPNNoUkl0Ur455nd5
1ufzzkPmOBuzg0ePO+ilfjHF3W2JO8QKggc4nti+BC/Lm6XIIk/gEW3OCXvSXeiH
ylm6blzTb+6Yd+gdhhMX3ljL4Oh+aKMC606QMC/lsC94wt8VgUeGfeTCwR3ULH5Y
H9TBYCmYVx+i/ges0aRhDS5xq07DMhDacjdebSjvHS3N++FfICQHJVPmn7+7vuL0
xxTRTumop4FpwH//oxcApr/tmAlANrlYcLgRvwi2Ay/JCTfRwUQn1ghJrSG/+r2a
0pUur3zDJ7zJBoICBZBFZhwfWbrgYqfXC1v1MYdgEqGJS5UDXYOMXUWs99n7Rg5u
DZ7Ch0FgOwg4+50mrd3p3mp43ZzNtnbf7jqB1o3NmA1sHdV/UeEDG8EFqUCP/1ov
cRgQnWJ5oxRK+NzWBQgXFc5VDl7EHz8e7raoTKi+EUgbTuqjsochGuozeAxvUpuA
CTsB7Gm6c3aj2NBDEmF5sy1isBsmnmY9Y9FoMoHbDDFes0a2z8k4zKW+QyQmkqeh
t8hwFcD0zcExAE/kjpqbvam7u1vOF7ST0XFMhnVwcfn+DUoLZ23yci4HPx8nP8MS
JlR4WYyN6KhvbIOyBmSALtYCHKldKzAOxBzTzvg+gBbzOueD4M9huNaBlkIB8q6S
9wPGUlra4vnGkXY6x9uwrP/O4Kb1CSEQCrEXe6lbrChEL4iiYf39JkrYX8gikfv8
lDyHWDl+DBqmtknNbdrxr1W9wB9sschhBvlScSyvIQRcigHqOoMeD8k80AEFcoR5
iVKIadtD39EcScp9sDYy4D+QEjB563V2mpV/ZwWor3SrnEQqI3moic8X/DGgmd9u
QiKGM3GAfkzV2SfGq4hLMDq1fGKxh6xBqqxYE/CbQNrOrrDSCXhwNOYQuHwNuOSx
JY9+6MC77ej6+4s4v8y8UsGo1mc+aXb00GKfb99AH/PpFVx1FLPp/RXMETFPRMR5
yImVPWLTi+M5dYImHgWcK6wVcgTYSLlw1LoEDm8eYjM0FtWhuW27wWooQqGHPItm
OCJzEuk3mhqXtvsPTP3KsbDSjZtIi4Fl7mLJlpa4sKAs6AncID2T5CGnxFdEP3wl
93SSejWf1odVrrkLEd7VN0NMYirtCST85h7QyL+2NFKpxf5WURa8GPYr7AkRzWZx
D916zEFFUGOjSOVQtwan50yEX7vYaPH/fuPWlIljqVii6P/YU/O8D8qEDCpcojmU
zfH3rAk2FWRWNluqO7nPolFxV+OCPC4YR+SGMo4cyR5m58E+99U1UzgBxIuhxmNr
OgPjnPGjxnoj4lqPglgt2gj41py977gUlS5CQOPHJ6TtbDkc9fOreD0pCRAOI+47
DaeUNSkXbYaA0ByORdgERIUjrB4tBxET1UOpGmKKzxDEAhdYHsPv9/UA0qcmH73+
7Bgb3xZ/1XrDpVdwxwmimvPPGNA+pQBOZZsERo99AbE5balD871tfS4ltmrvuO2q
uVR6KVsg23Pk1j4QSiqeGktGK9I3igRqAS7QGDaUsO6Z6aTVGn1HLo1IPcLeRbTl
zfzivqlzjkq5sUALWSAZqgOvZVi7dvz3041Q+Zysd58Cnk3l2K33HPGoWZ2tN3Xx
MPFNmXqHcHslrCo8H/933ajRzuSPwuYaYnsa3v1DEs6bINb2j9djrIAzAokrfHkK
/l8SGqLLB4mDHvaRFWWIMsAk74TIius1TCmg2JcaCOEUKx+8HcUBbc+garnt1iu2
O+clJ8aCfFt6B2nxFFN9nn13FapnePOeDo3iU/NHnu5WImurU5+IM5i5cpKGTxLd
nlSEjj4mdQv0nuWDScBTvpGrToYVPNNg4RnnZz3VJs2+ImrKaEyOWtgDAAB/zhT6
Xd7cKx3aDuPyPYI43R4DDlISq9bewwnbavJ04Gzfc265MYDhOPa2K1AAx/jt+gOG
94L1AMTNa83DAhGtVd5Td80IU0PZOVHZH52Dbb0cmmAUU53PLTQ/IqJDgpf1644f
fllIUbItnJq4lJDONgL5Whj1Ku7jHEO9MkHaFJDrqoTp730HPRfC3y5aV/oOdZar
BFZUoZK5SSn4HUzbkl30gVHAMlJ6ycFvZEVQnQ7Df+yUgsgk06jT6EuVAJjEsWe5
DrKmKtpaj+zo3hwXlOWC2EbC2ErLyGSGN4mVd/MRwMPOmDE0ZcOq7Mog5mtdUPW/
kti2tuYZgBXArzx327gjGHb9Oz9H9cKCcCGg+bAmkULvbf0maYqbySmrbAobh+C+
9S3HiLXDOBsRs9jLHJRhhvQP0LlzYUl2PvAlGL9CwlIpqn7M6nbCOSM10JAfts3e
E6FStoJglNfA7TMHz64dURzJPRQKvGFC12apwO/YJPeYzW2LS4VKWTKVE0eQ0AQy
GTtW52fSEdL0zAyFKCevh+gEjurLJmhbFSt59JMhd2279nK8+nf4IuaAasSaVPpi
R6kRzyy4ZtzETYpckX4g0GLkwIKwj6qL8Fblj12ETw6nthUBzUeQNrTSR8zhry3H
HFEUoLvX5UL0tJ7sPvFU9WyVutH5kxQJfZuxiXGFhEknLQtPkoq2SEXg8I7cj0xC
jBKh6hrOvUCw7h0LJ0QvXNB6FA/GvW5qy/jgTzzVHtG9FRnbZyb7fMmj3Qbxp7wZ
fCuZeuvaKyYoTr9Nsnmv2IreAHJyh4oJmDF4933BpYTnIc7Z3jwrQLhz9hBeQUH4
5mlrOcTQNF0TmxAYjB9pC7PmLCSBo5PDIptJZ0njc7ylyDQhvuJJjOhOJnhbUu9P
tuqHYkVjl0WtXXzxTgIW8Ble9SG7ihyhhjE34rRFoxNuut3w/wP4+zVZNVttLx5U
cTEilFrdLKXlmhZOf4f/UzEOhAT0FzT/rBlib2wpX87UgYU/imdTS2KHBHE99kRu
7nx/ogWrdNi+vLuD4C4lkENxhy+FBijhXc1Wg6yVYxyPNKg9n/Ntvpb9DxgfSEEK
Q5VFBRi3A8ODpkusf35vff4qd5EAyyWholYi7OWTXIQJkzcCIH1518K0LRCIWHam
CUe3W72HXSuoCi4ZKIDm87dClqEtPDlCLsx0lZz3YjIAzDpB8fBhMQNUnmkInjPV
I+qVe6Sf9GPMiedadg40W84Osp0AO3C1DeuZ/KKMkA9edxuDk3ejB1npY5VT3JCt
jEGLzF427biymTbzU7wAWgFdShUGVPmd2bz8Lf2Wnr3SphI13sWS2hof1DC7oLL1
OBVEyRO2pbcDnNEFvVIWTnK0QRihN2scr148pNT+3tZlUx22Kvw0ON8blA3MrcnU
HawL9Br5UbPhfCRCuRsetuMhM550/UW9OpddhS/xwZL0P5eM2esW3eSIgtzh9DUj
UHyZnGbN54lMRf5jsFJI9sju3/5xqXU6ZDh5dylWUIBxD7zujH2cP+6RBDc43fo7
kjAduJz1yEt1LLUy7WXfHEOWeevMT+UZzv49oen9HpufvO2hMYK8hXEC6VVLjLJ1
uLaXaY4QHOql6MvI6aLU+Uc0KMX+ZC2Hvvd84wgezHdFhgaZRYBmqVYcd2HvtM0X
2UPWddNAHyIoVmARUXbU1RPysojtcvMAiAW0fHnlX1FFJlcZrUJAuRiXBoDVZTEL
ry8/t6xZJXhuNN44fL88TKSFaiR9X6Vj2oe7V9RYp1G/u+Z38csIGjO8iK9apUx8
saLMDTmwoca9ylim+yCYYj4L9MUo+PZcHQkxZ77++YU4EHYbqim2vwboJz4ZCn1e
xp36//thKXqaDM65+zgjdVwuSF2iB/9jV8ifEQUFaSp5MDUWlg3z/hZmqyAysYfQ
qY1i4xyvKsiHIEmSgtiO80xWnYgN2D7FNYj959qLw9sH6J6eNA2LfAxKQUUyrlgi
s7EiTZEMiQ9hAOjl6MIEQa77+fmJ99S/1ElAvMyhe1dfmw/h/u/bJbTmkek2Cbi/
iJH8/PyKV9WG6d6xKgrMcguBWa3we5WHiyIAWmNJbdKXa5VUWtNxqDyielX88K3G
SZuWnOj2qj/pKhJlCjLkLqqtL0j1YVl0Gfn9ZCTijYiHxFRgdZjVsCOSl0GGixAx
l4UrB2Q/lKZVqZuTmocB/5dqiw62C5Mu00R8dBS9ucgo9aMEZ+GToYUmWkmqQGzJ
nqDeCvwr38OVMnDq5jnhn5whEraCGgyBZoa7gLq6FYtxeSDlKks/tTqeBYVNSEFN
bsLAmatWRuXUsHiaUZiRbdl41KZlc04d3ZT8ltJimTCHSjqFHaLvKjreLQTTn7Xa
pDfSzRseOTFjcCOZAGofF5zVsSlpX/TRP3a9FoOE3imJy1PT60PAJGCN1qwc4p1c
KuxTBcWsSDOjax4O4/SWSFrNlGa8AByVbNhfscnVsdKA+dc2odBD6Ec8fce8HhQ5
VPZdK2QTdHsS0h5FeHJVZIcJrBDIAVF8rBWo++RrFxqLKSsH2YR63mq2ojnv602R
3zC3QfJ8fP/x1vng5QZ7WQNT+gztLDdTmhkhCsHJ02MDi+jumID8a/+OLj6vgq8E
uL+xplET2L6xfvIbwS+xQMXBAuk5VLHI6LT52GffsHcqeTal9ar5EN/+C8KBJ0R6
hnFXlH8oSArT2FbUE9osFt3zA7gxvWgO1FN+AMbFoZwK75+IonO9JbXMnD3beHQG
caIOWrGC1BZzHhDPQmWUVhbyzZ7Z23cXC7rkqNkQsdLKaGz6qpB87KcPWv1BIk3T
8QEwhdsJOugGUtbZzc0itc8wjPsCBtWqz/TuOKtI4qoMqQZxB45VGhgUEMvBAkOH
ApQRde8pOcXYAm3Mv0E2yFikTTA05B5E8oKFJqMk0HnqiyPYHWslQkUxoASm5aF9
y2pbBNEGWi/NY9zfZuAyALgltNp84OwlGoYkDOxQ9QaST5Lb+NgF3EEysp913s6e
AKeXj7oWE1BwJ85NUf50E/+WXSmIfebVe5oyniEeltJiKp8lMOGEQGKVdBjLCd+D
RPjrVm3RS79OnhRESjhFayNNgZdwElZO7k7AXWoBKSmR1vtVeyQRJitLXPK5ZUSW
Ytr2+1enFRuH5Eo1cEzfHjwyBzA+U+4p5xQ9Qvdla8wCG5IlYLIj0GsMnmmpOv0Q
XApxqAlqLPKe3GGp5MFQb3/U3CsWvbooMwJU8Ya3XEjGuu/BYkXE6yH+Y1lUAJ5a
LW1WyWN0ULLtcw2LOqvDwQvTqo4pfS8ZzEbi7DrjNQabXPJs2CoxALo54v3O7Zhl
OsD2lXPhtBKvHwY5NsWbeqPNVHoOimCM9jP5DdI0KHmpuABBnMU+Gb4CS4H688GP
qTglVkdV5HLsnUAu86TuhiDTkXfFbu2m4aTyL02QSTsPIywcYwwDERVEdf4BrKUW
S5BQhFh0PGHhWjTIlDuVuJxMBh6mq568v8RVdVSc2EoiIhGDKjZtFVzzmwR8m2hC
nuzyr1wa39iPguKMbXJPwrGqj/VZzR6f7tbN08xGKYxCvFiownXcoL8lBKbCzlgw
zMGBKzF/71dBa8xWWnCsh84cJVzTIt0TTllDby3rrniDALIlV9moOIJ2YHHWuwbf
EpAB9GH7CD7VmT4W5BaJypedxw6ChxsDG/1vBBg8J01hrTKGn8PUqeHp4AtVpCeM
8sS9i7wRQpo7o6hyU+MqPxlP/BlvKX6er0u49iC5WU7/A+fDnlkRIszysYzdsscs
xX1f7RlY19PNEkBYu1KlgxGcEsE2g+L05+lBpFPIDdAqs4nxQSjo8hfp4KaTq+yC
AcP4fj1JQtraWY8dkC31YnwTWArhxszsn4vwL5oy0+iKX011yXQb5/oeUuUt2GII
KDZrxHYj1ig3CW5ZYYIl6jpcqw7UFe6O6PPayps/HQhSSib5ZQlmhbjOxJzzSf6q
7QWMv2Rwv/tcZBMT6s0ICFOkIWAowT50znkroF0KjgJe7Ek59ujb6RTloRyuyr7n
Cokf4LAl6Eei4WGrCdbWLzLFuDSK6R3LkQE4LUjjnzhXE6DDvk2gXmaIhd6uzFkt
jfBaSPB5cF/zy+BjGPb8TvbHXV47BDwWci6I40RpvzewMsy25gpY+Lm4xT5gtZ9R
eBZB97QnvTR0ueggrsNC1D2smnIzENRlxB75zBnGRFo56UGBA60O9BURki9AxEOt
9lETIttTJkNfEdSU7FKi/Oi6LcVjfXM3ySE9pBhx1OUgT+TSrHidzXbFHlrAWCqE
/0Eh/pDsrkk4FdIDlSl97HDD0da+MGN0+IzO7mqz9fc1azyZnFrbSY9+s3bJhPUF
IitHntPeG+FEak9ukxKEXTUTdMFjY5ZfbPk0Ebw0flewJXHt71ZcrB3ovcoSiUjn
IPzh8hDRVa3tTV6lOscavPSOVdc+4hLV4zfqr9lstYiieliPsS68QbFiX+vmQBJ8
6wQQuU3KlHybji/oCdTx6wAXhf63wVmvs4ngfOfyTNygzvPw2HJ5H804u3zCPOji
NwwyJPTBw5ZX6qoD2brfwEsUvIRLxMzNTVhy2Rh52ws/2Z1W3Ki/ozxm1afikiPD
fZAGlvKiDpsyZwbPf8q+5qTARjau/++VaDBTEgtjJELIq6BIht7EwHdIsXvrzhWd
A7g1bFfPfRmPEP/W9dZFPLoik/Q/OOuR7REJAehE0HMUYN5hJkapr29MPDNdtbVJ
tLRGSibNG6m/1lZLIPDMFQj67nxd/gNHFvj3NDX1hKY2yOxs5ZYyXTpPupota7Iy
caPznjBtu26Dtd3BlnBVl39QDyl8KT6xXBoHVirAz8fqaDcSKnVK9eFwl29Z4+n3
IJDy6ZVteTrJGqJ0rYCjLPjnLWtEDoyiEWVr4HDzNYnxNHnAk6OA1qdrAYQLBZ6V
cS3cBSsY+Vkbki2Kw4pAg7ZYa0ZyVp6kCgvdy2cUxgDjHwSfn2AkYaEE3aKuctOa
s3yl4BvHqf/LVqHxBjFBmEpAQwhGt2ikP8diDmioAja++iACEx6zvlD1DyuzKmPI
KgY8ZcVtS6+Ea5XSNylT5y1Ei51BpG/2J7bRH9+SG5oP7IbtOtfFGpias5VixDrN
6tCl/7fSvsXG2psdmcpLRyXOOh7P2HJbmiWbf7Voi8HPh6OH4p4AqpgY6pw9NlDW
u0BSsrIVgOV4KwQh8zWi5sNqH6OM2CIEhZt1xfptqJwSe30oTrn+4EFTRNdalVva
0PIgPYYV4TiaPd9bHnMPqUqIp5fnZidG7y8yavBe/oTDvFeECI65LWyCyPCZGpcc
D8i8tgayE/2BuKCkXJVblM4dWu+TpiGZkmFr+5MOeNAlCpmrt8W32SuTXffQkv40
a5RQwP9O9HW/rf5dMaoZFw2UzveBp7AQ6VKV88/xUN7cxzB+ja/UWKs18QywVeAJ
v3JRU0vQegqwWKdmeaatYM3ezSssl1JUTkKwfaq5cmJvjtPbisqHoyLuHvn1eOgl
tskbcGPzxJn3XHK8K+24YNbPUkunx2wjO9+MBn6dxQJFnomB3/3Jg05XaVG1bGao
VylqWXsUNJvYJCIYyoex8yJcZgS51T3a9Tp6Ls+r08DakLXzMn+GbIYwFY97TKCj
wWst8bbB+DjxuJur4rUSl+Vse8fAv3CoSzb6BWdRGhw6t1QdGpQyOkkX3uIheBSw
QyUjLqGFh5fNhy/F01EzK4qU6hUUSv5xnjdV4C1ZWWCszywjTqUahQfMVJM5KYsS
K8Df/qZBRZmsBs3ri1UIyR1cdzaDukWsHR+FaP5A5xT0QW5zkyUa9Woi4MpYVqec
qSEEtERsSOjHLQdigtWoGOIvtrllrZn2Ic6Ya6n5AO1UVeCTl5tzlls+Ce8Y5dGt
I4v0BE4SbhTCCq5d+iDsjJhX+tOiW5DUvCwqSbS1TDkVd2ZGHSGcv1XGa3KlcvEX
t7lYiTaO5H+eLVr0Ft1TGWa5rR4Cn29aXDH7rIhI5a57qYkAao8KEPsn85JgouU9
Lt2wkcbUoRcuKoQFoAae27EktLD8icUY9OQ08xUF5kJg0Zx7/uE+Nmodo9jiCrWf
6Gz3JcOvA6TYzeLcDEI+211FMPxQnHNoJC81VLH1OFuqyCRMQQqipIn0v3e3R0rt
SaLW7UCcXMjUdS+VJB4yrF1ml4yqqsxeK13hKqYU3kDRi6sxuodhDSdeGxNI0vsy
cRYHJ1IssbA9esCTf9YDcg3+/k8tUd01R0U6EI0weOk1JHfT8MMT7Y9SQLNIeKY9
w9jrzrfjijTI0iP8OUt3AUCEvRo0yWfmKG7gnTyBpHJibjM45+N7uv454ledZv8C
nDcHWkG+NMIiG4IqRyvzlLGEcEOKK6JuWZnf9AVX9wM/L93j6prdjIw7BPtxydBn
Gsodkmtqn1khJ2OAIPPsarODD4YMxfEXoJbp20f2gNcrrtfBrB+KVQ8Jpci55E9L
LcUnrEiFfofiwoFOLwTA7fpzqBtLv0pAKEka9mlA1dwGYrl/SONLDkSWdHn0Rsey
jeH1Q/QDC481uV5gTG+/tjfQF494Oj5B0huqZZPCdnzxJ8RtFJ6EiSWOpfPGGOT5
qAAeXINfH0FQsAjnMzd7UqUsexF/Q7FUhfY5xXfiLxshhVB/Me73e/yY9JBEfdVZ
JeKV4mWe1XKts54fdn+TuMCBl+ekzbPcJinwwdEdSGVM4hr2dFaNN8T3Ypm5FrSp
OCe98rMRkdbz+k3MBOzpiKgB6W7kpt7y67d+cAFDr74HEx+VWmmu+JhL258yVq49
dtd8Iqwap6/WZiuHPW2Eqp8aL8cP3XEYOwgqX7fPak3arnnzA1vDf9rGKj7Vgnmw
VNZCK4qawKPm0vYhtd8x/lXWXAqL82aYMJ9QsqnORCSLHogqnWRNsHh0yZ2agn7w
ZQw7xwjYTUXATgaZ+s6/3rZZToEQeYFikQ4uFY1yuOjlt3L4tF3EwcgHLKwwIQWJ
5WEWGk2dl8ng3NAWXRkkLW9IWC5/7Zg1pUQ/JUZlV3tO/eBGOikHme1ecu2QOK2V
6WldmLLk1+CVQK+bpJ++HgZIYTijWeUkpPAAFnyfGbm1mMt/DGi9WhkGrGWd1cyQ
yyI/N2E/rbFZCqBymf2LbaA651hE3+Wkt6ynVQJBWPbTfTECaReeGwo7/QbDv9Mc
850YiPbKioEgKHAN6tiDNNZprawBnorJp+WCDWkg7a0eEmHxYRa+TXGSvV297Rze
exSgswNX/ly1Xvh8/k84Gnj46ZtZHqP0b0DzKnFpiF2qK61SZdI852Zd7jpnxDFr
CZqesHwTbUgDXuTaoAo4eTpA7ooRHJMVNHtpgo7BsocNPQYOjHXlD0jXH/qjrX0y
REu9b2Y+i4Np3fzdMIT6230B7hRz+tI1RXUSi1iRyt40I6Qbl8xx2QD/9/U0Fro0
3U+DdwhBTv47rNoQIBnIpLWr//0QqMG5zvW50hiRktL3UHf7awZDOalEMsld+y8V
owAwFDlxvRmhkCim2DLPhxqcBNK3zk+yZgtZyVHcVTtN8x1NzuY82P0R9T7RxRVS
h8b1wyn4u7TNcmZM4JMMY0ubqLrtd2cIwMr7zjPerPwtiu+xL5wQcctHb5taoPtn
JLDTRu1+UTZ2H/fnhsucEQnhdtcfDx0LVJd+FFYbKyIoxU3c9pzc0ZHzpc85h7sT
4MoRJMwjJREt9QdtJIaql8hZH6RdkTzBIun5s8x2EfU7JGbsM2KzGc5HGsUvW5ic
UrAgH/SemZCBxaPRqKjiNnQpWpBhRR4gcNvnmZy4JqzS50727hLG73lAH1SNYyUh
y6eOsggk/eUljsw4vfjqJKhreGB+vbES5ClABl3hTGASc2Jm0wOLndb72fZSgcBV
N3ygdRl1IXRpJpf0vamtS8cftz75j+yq6c+QwQmiELLeE+glpWYbnc+ANk31/m6U
vp1hZAxDfPq8I0oBoOAscZwMJJ0/S37f3f1g6DDnj1tTQLkL6FL0RSyRYgN8Ya/o
SDccy42uJKs7e89POGAO2dkHXHp8nBs81lv7oElZFPj9JlWg5mboOvGpOE4DY2vb
qoRDmE8sUCaE7ICf4uYtiI/aTqeIEwp0lm/CY4CwN0OwoYpRbWFCuI6LtHPkmYun
P7e2D/EbyPrLoFjtyx7Q9U4tzAb7LYbLdG55yjhPGHztP5Iu3FgHOCza43XkeFId
SIP342r9Vs7DQVKO3aYdEJvWE50opCUdryIMJWWV0Eu+JiWO/rkWsEKA0hPhoNN2
K86HKAodmPCkQZwzimdWwqeLpTGox84f7iWLI3AOrLwBkwDsR5apZGvJ5NOBNYRh
TFqUon4ezKcklwVjv4dX8XgCr5PEtB2OkGYTWMGW7kpu3AzCYFXL3mHCwgV+Dbed
9I80804YYXhFoANhn+xpT7rvQCKK4A4FOJn0Hd+i0sxGRgKa/UNJu837JyM9CdnC
LdFd3N9CbPTPoZ7Bxv1cJRLjHBG6JQrJyt/8VuKyN8XNPyivDp9An+Sr/K+m5D+b
LsHLaq+OJqkiaW2pTtoInTkmKaLy8O5HYSOZ2nfRlZzdYicgUm6dTlgYNRLnIvz9
yGz0TEdr1Stmb0n6vYGQpL9FQNh7OYPC2+fVmUEXUwQfHjoUT7gE/aYyVsUzmyW3
cSdIPd3/ilPgUcBFrr5noeuMZPB5an4+pOxtT4YMcyRZ+4rmg0oN6aYMGsL14Gf8
ugtr/3fuG1Zf7zZK1f4yj4BegjtqFNCPhmukqzYQAO5VefxxN7Ojvd6XkQysCJk7
fRGOFbql0a2IazfJ8hOYvkRMUFUHr+8DCVwPndqE5k7xCFr4fmQrke7TnIw+qKnZ
gS/peLkKU71rbHfm5wCh7VUKg+95sgh1xmlVDmFYEwtDNRGRsb7M9nSg6kAJ1xNW
lcaZzzNPVcd+zjbAwiV55IofHJujkZfAuHBveI9UXASQV9nOcexVhLs1DuOc84vM
eu8fqxeZOqQmiiKqWANy6p5mzUc83jzjZHG8fZVZRc1JLcVZJ/fCC/2kiSX+Q+4m
AQdMZ9PpjcdWuNXEvjuFYQPx5iW07BY9XHxHvcAVw53LWLUYzx7DS5h19HWlIiG0
pjQmXJOZPYxWLfuhyWj7xqNu+C5UoCThJFUzqjDO8AA6s6NgHpe4RlsNKIosXzNP
HON2dvRhSERkuZkfarjKNicoqUs9rBdoQuxH4iUF9Vdp4Ta7en9HPJn+2GCpAzfN
/WDn2GH0nBqlPMEo/yqRKryHXqoJjf9U34wvVdMQF0A4jpXLQWx2eCQWMg0LHZTm
OlQz3d74KtJHCps46bggxPHoBi2F/b/PHRmtrxbWx1P4O5SDzuDHisQlyR+yj3vk
9uPoN0MWjkuvKA/JQ2r5mIiH5PtEJUjBV8OWeAKkZb8h+szFtKlOsKGQXR1PXZ7O
EDkUZnaHl20re7LqWQgVVHOLTEd9twoE6U4QAjhxbs5fmqRZYlJVRAo5L2FSy1nm
xEWXVJjXPCgWYDXyw0vtOxJvhPSw5RvAn3IEBaFnhF+qUx4fo4PMWQn7uQMqoDgU
S/l+3xyC6RFKF6Ez8pgBwIgkXd72aSPqTefaqW7vgHLj1YTpKfJe0CAlMfuBllD0
Ob2smL5kitCMZE9yNsavK1Nug+H0xSvO/O8GbuyzKql7SM72JTCD4ueC/ZWO+N5P
1G3vrDKtPbe2/0h3CMEHZnf9mZ3Zj1QwtM2TNWoI5ui4MK36zMxLhgEOo1VaKOWc
80d05XqRnwqRQvbJ64N67R9zDWMyTDCgHksJRCSTj4x7AhR8TYLCWeMaqxZORVvt
Xfp8947U+z+WBUHutMxKyWM/9UrgYAGTsSYa+TdvNJaSjjWKpgTApa8M4klUX9I9
HVRJMBGbgajG1iPB1MR/lS/+SbMHUqnw9R3Lx9K0z02tKwTcYaZQXMctx3KP6Giy
zivvSikcXq2+NF4/MUPzJD+vLwFLpK1HDbay3z54TczIkBv+ntIqHAmoeQ4D9VZL
3cHqU8qz4Y4T0Mysv2nD9M3L9mgtZ4Kiz4TANpu9OF+hSZxyeBLrIls6BzpejViI
GjlQnJKl9HBOq6nH/OmKUweCz1GEQnnKH4jK1Xm4oIgSS7ZnKOC9NU22U4+qmsVR
dNHJT27tbH/0jYUzRIHY22AJBNbBrEs5QDoAqOtTFsHM7qnT8dJzKiyKhdG7Xoe3
VYys4sbwaginevIrt3Uz2C1jlfEphK9ZlaZV8Y9z8O1xnnZ6W9cKjL28LFRq/6Mk
z82e//6XIy1vk/NwNjBobmqA8rcmkds3Nal44KubQLnby5SNxj4uvO9leKhPLVUt
9bBry8pyYupCfkOevH+cpzt2UI6pkTJTo9Hs1pmojZwaPI8h2mKflodrQE5FKi4M
fi0ai8MNe9JdiN/nQcF3uxtCoprHXIjnWr4YH4sDxYlzeJbj5tWVTYsQGlpT4Spc
Sf01S3RszI5Fb3Wd4pW+0REUt87wEGQifviRS0QpeEG561eJAlqORPOljuEMpHs+
V37MfVsIvTG4WpTFcQMRiCYRpgQGqGugDSjQTLS4dqlai4G7MzjKUiGBfCiJ8Wd/
3Npj55iN/WORLT/VNpK7s+rZrBDIoe6fqtAEwusBn65ytdLUtXwth7ZtqzfAktyW
QDJQw29EjqSMKf0JBo6JJ5wTa+GUyHYd0gpSfn8UdUoVKrAQyjZk1azg/2lmRdkW
TBLFxYhMiuPytHUugqNiIz99Dqo8UvFzMCZDzBMvp9aiJbrkvG9Kw1V9ZRgZ3vzx
HHJ77+NkvQQQFBJ8J+lc9z9SpAJNQs/x2DctZQTGYOYDChfNCceI3UHTpKdzByC0
2b1eUkwg1pLez2VBOQGFGilf3UXBM9plgnM7lFYbOYCMFgdsrz4NsqjbtTXTeLSx
K+0NGCtGXjkcxeIHxBEDq/tX8zb9V7OcaP8dPMT4h9OqSktDWv50OTxHIcpmhMwo
LdprkQLljjM1N50yqlI1w0GtxPd6HPwVoHJiaGi/xqBdBe1il3eUELUum/3Qjj1s
GSyYTRTe3Q1oJbgtPg3EWNGuBklZCvG/qYhFMPCCVpEeXOXYPsSYpALlhgdwdsjr
fYrvP+EJ4ZZ/VSUygJmJ++vMQxCE7483xR7r/Zvzr1Sq+zw1UWIlkmgOAeyND2U0
+0uaYTu2uZ45F8QePheA9842VniXnC0SDYxubbGdTT5azqhN1Q3PrwD78RMeMyjO
ifZAPB1NUpAHA2WUSqZNs+LVKbFBwNNp076VUBc8t5AxgWNFwAEPdc0pVzJnRxlY
Jhe4O+/eh8Y27m3n6OVlHw40BP+qOq8SfQ/33LcnGHCTJcFgycizSUSZ146hL+Oa
QoT9ntqFjiQZcEVQlSW2ZyhFAtwpZXvaBTu4hB9Pa7HgiTRh8RGm1pTV3etMHeF9
GALDpzaoMdbxLGeQvS9v0rHMHPGRIvZVjJ8Ha7HgIFHlkRcZuLORSvM2F19jLqFY
FzdRbvjSOdBAcosEoNNj+Ob/DuasLqm0mBlKKa9GjnzVVYN9TDlFzqUG3Xc8jqQu
Q05rrh962elLg3vp2FryBS3o6VRfDN569g08lx5H7b4Uq/abeF6tjyVgy9xVF/FP
u09pHn9mu2rS2gMa2QsBFom44X+WgzATBekNXsZIQsJ6AO3ZKud1XlN3xp36eNoD
qoD/UOB7lTWuXW4FU73fI6oZMaqIwl1OBwGj4rJeQLpbJ9+cvma2w7L+VG1Yu79X
aKbNLwXaeBbo7zK21PyT05yOQHgVZ1/TBLQhQEUJQp7ikT33Q2zTzikc8+J5YeDN
0PAibOXlN8iBr+GwhLJXT6zY4Tqjo1bON8I0T2U4HsyBFx/Y2lX8yMDwyrJI7R24
PbXdMAko1TD4D+nXcxfuYeyXZ6kPICIKEXNEmY7QfwIObz00ADtfDzA0Fmb6RW9r
6/dmw923pTl3uwgrAxkqKuxaCczWhvWcEY0kG9joLC1OvZaqTRpXldQX+R/N/ccR
eccxA5N9cTWbg6/zhC8pplcLsI8VN1LujJNJ6rfnjEQMaRQeK19Tg3T7NoZGwpS8
Xsefys+rUVcm0Tg/T6a07cRN7sbFNQkFutAb+8Eh+IIdeTpHocJQLTWqQ/XpqLp2
lSeWTkjGNnBX7+gE41eQ6qRkjD6KdisZ61JEGcNyFwvvc4EDHXUQ7ZEb8sXlDazW
7R5+vCZ2knfi0D02yLF2tSWcKtQaL1SdKoeXo34sJ6jjPBe7fItA3wafaAwhtPH7
6G2A8XbZUtC6zlpLjFmdTVtg1kVz0rOMLIs8MIq/KrbQ10qJKBmjndpWlktfl3XB
DCOMyRBt/eX5RCV/FJyMR8KODj6s/hvKCapypm+fYHwHh/Hgv/Z1sLU694sSReQp
IrDJT5ODhu8gpmlJ1MWcMsjqIqyxqD8j77dubGew8LWTiBeT8BaaOCk8uu21Kc7F
1G7T+n8pQLogQO2/eg2AGoLC1FGVktGvekP+Swd+CJJBHIEJUEiM1iKnlA2txm7t
L/RISrOJEohWL/gMCOCfb18ZYk+7y6Hu2zGxIYe8o4wWVuEbOCQ2T2WSntG8VmPk
p/TckWxyEgYxdlPCh95SsDUd56L+vMSWqBb5y+oBMJ3dfq3dGvodrSvpU/a5L45m
kfkFQGWysAxdqp0MH2wrGDJFmUhFiL8s2ajxLjCScMgfKiUYsGkfPbDKVAiSxqdB
76LEQxOTc3wDDm6HE3HqEmLgGK+AxjMw9XhzJyOvTS3efm79S4yeHkOqw4rA58tC
EDTrx216VRUwpN7HuPEctO/JpvDcW5307U8YB/Y7pbER3/yS+OmVm03/8vi9bPGz
bJo8M6cJE2aYq2yf0HfteuhjPlkiZ6M1+0svAPE6iXB1WnonO9cRoRPidX92TCO1
XqCczqi+1h91GBOm30aiiSgxSVrdyQAHpARaFPAvVjqCICYPRSg1wFiJc4PbDQ3D
rSARksTHJiyw7O38wC5Z8x6Q3IKFgJnR5h2dtN66S6QTfVXvrT7mSvLmXIDX0LkM
YA/e6WDFW1JBzNNWUnzQNhXUvtM4+rh66NGQDk2aYckdiR3v9hWfTYR3MkULW6ou
ZeSDWFePzgVss47XxqsljpeHd12GuuHf3xzzPVAZ1yXzY1aFw6GpahzDpBoeK0k1
9P2kfrRHmE/7m/ATh1iMFi5k4KD/3RD1XNLcZD2OKzW+tp+A7Qz276VqY4gtllEk
xbelilUH/YPpbnilOuEuY1kZ3x6GZ3KBHWFAqiPPYTUjhlrM4GvYE4HMDr1S5dE5
ILLJPStwUua2QW8TUCmYoEQ5BLpUaIxoVR65xMfHz3QKrrhxRI4lEpEwsN3SQGPM
cc6gVdxcwrTlFntKF+jNwBiUlQ2p2tzUuxuLBtpITRc+Au+9W0S0w/SB/fYrp4KV
ePniLo6E8BH1yr2BHkweQ5/mCdK/cqsiZy2MT4qQf3/rpivCGnWXr4evr9KsN5Qu
DIjwcO+u0nCPBfeb5NgiWP3I996Ww/ESGBZvuZRs2uFq4Zm+FjKAWvfMNMJbLEYs
fbK1VTjr72iStA13sgUnjmo5+sZAqfHmSaH+qmaypgCMeGRjC9juEXs8I5B1n04T
4qxzkxlW0BC1cyAAhW8BulcPxLuqeU38e/m19hPs1JgFpqd8cKFkGytekTUXrYNw
MOD5LnESzxBX15RD7piHYnw/l7uw4Us1HKR1y0D9kI5oFwFELltdbeef+4fO83Rw
sHMd2mUlEp6AdgAYBwtX488vb2NVOWGH9XKITnYl3tE+4fRu5ENj9ihQRj1sGIzr
o1qWyz5MEhm/zis1JvbOASNZGV8IjVlqWW5GJ/Iee8mykas+wbzR49LW6IYKy+Lf
s7XCV0so4qHlW4tjoO3QniF7+UaHAoPWepdFMZa1baR5A1D92rwM/ItOUGiAUPkM
QUuCtTv61akL+E75VZZsW3c4zcMsybBw9pEW1JQFt8yvdlod5uu7DSKc5PBi66Zv
s8Duh5Ru6No4Vo9k09tJ1+veA7ynOE5AtNPa6Z2rWg0RnOUjvy31rwBQvyOCFCto
Gl7NvcBYZqt9MV7bF47c0b7A9T2H0YlZotLJH1XnCZesZfL3uB/mn/64/MBKTyXy
B9Q2ad34X1bu6doBMvCPpft2aCGWqWDRiYpPExi0bX1oeozgRR389t/S4ufUYuMk
7A/i65glmSYN4P6ansP60BdbQ38LYlQ+cVOftdeUIXmp/bkmi6FzAni0H3oEY9Ii
p0rvcEdXpX1pA8n0B4q/kEMBStSS/M9d6rlIj3+EXBCxHHlxwyPT1HK0gqK7KFbn
7oP2UaxRPxEkDNOqR6CgpL6aJGNIQqmN8bB4U7x43bNTLLm7YhWcDbqNGJsJw33z
sase4EStkXy2FMqiFLk6tIOhRuofZfsTF2iITCCXoPF096VMYp0MQVsmwL+soxx4
wo6t+lr0zL3E7Y6YNXVw9YsrdSpnnvZ2n04WdvpllEtoULsHz42GoEk2pwxQyK/u
ce+MUXf+xebOmlQ2j4n/P9DucXXQZHouUHQJ4gpwMW4SmrzTtH5d0RlqLRj6UZTr
JkZbMHdB29t2xmhIspxNyZ+wUh5i12Cx2OXsT1RGoRtojEXvg3qLPewD9PYuXKeN
n2rYLKuWioodwb+H3+6beHS5o3LJYcxfWClUDoQIPV8ZUzlDpJwilvp5XFN7BvLQ
KllU65ZekH5kTm4yLDrLHHBcOgqqsB6xxzQb7zHzWSobc8mg7Io4Dg4JqX8nVyNs
p0q3s0uV6FAFTyTerJ2B23ZdU/wy2w9yP9d1IxgP4bmMT0hIcDtg/la0oDHxDrIB
NZbunUR9kWbqWlsFfYycawCZaWjSwgzAxNDGCemFYgengnq8QRfi8OPw4x6uSBqg
KeumDhu9ny/ho33LICYawS0pbF+aV0/pVCx7SNfdM5SMN6r8jZcLaYhHiWE+HBWr
+B4DWZflg0QGcADlcX3cm2RBkZB0cONQ7/qkPcAx0YTfikJMwprjFfFqRKcXUKrd
zKIht1/80ZCipHQHmSeBy99CrhqySN2NHz8X6EJVICV8SHuLshoRgJVWFXRjMMut
HIdpYw7HQ2RptFagjnZbF/tCOzoVoks2kmcMN1xtaN9vx4K/am+vvyHqfHjoH6EE
4QXD5M9QZz7oNDkr+jt+2/IVCoPpDSU6mtakWVJoVYgrkIIm1P0faeSAOg8CNmWP
dsum5ex/2hf1BZ4e5TuTh/gMrQjmOR2Vk9kE3tKosKsQI7QEtMk+NikEJeGjprwp
z0YZo02tsMi4KFAw+TQA+yLc8IrKOiiGBbdW35rZTrH6jJnaVuY+HSd6ORnSp9Lw
4hF3yUjMVGOHm1yGvg4L3TDsmVnXs4sI/TL7X6XRH9SBZIbP2FWsg5R0b2QRmANg
fmqI9YMB2hGlJzkormWMw8itGqZ/P+VK0P7t53sAzjOUFwh4R1+Gq8I6tvye1L7w
FvRahMXL0a9AagtbTjRSKmsDiWelhSeXFwmKLT2kauECIke9D6qMfr9SxbHgRua/
k/QHWZI8wh72SyZoJtkmZuEHRGG0GZO1cu9KCNUE5Ru6buNXMg1yvpT5SXEfYyZD
utiNdsC9ZN7rp0JpaC0dbbGUJlndN5P3bHZa9EFBTDfzJ7IeX7+KHFULn0Qi2JJK
Q4o91HQ2Tw6ATSCh2c5nSsSD0d6+yrThhfZ+Wodpdx5Zfad2J8j9F8kXgwauZjsF
WtOfk3S2isO88iYNPkdml4VZ6QRXrkAIiODstdlS16gQFGPHJy3G4V5IyHORpzbp
pOlQwBSWA4sYo7Rg/6g3YkoOR3cz8C5R23PjDZZU3sl1ZEes8OkrhNqmiT6xlzau
DOW4S1aQXqxXB3o0lJLWTm1aGpQjOQP3wHVo5ARo2bny/JT6x7PuUHV5rhrry6o2
SRS1EvwUJcTyOgNZAU0ipzsE+RFSIXpSqpGsurn4cHHi7XLNX2hJjS1uZPTlXSK8
S/akZVY4tg80qsA1l+/kcYvRcdMQVJytE5b4RnOlj/R7ZXSefi2ls+Nt1zBmGu+d
Un6Tow0NoWi7iOZL4W+FjObRpxWvfIokt4P/QTbVaC1S3gngRoIK1wI7PoByX9b/
3q3Q2o/UznPTZQgeRkAfZyk66vTNBvXNJWR/RLEwqFDwE+Fo/dV/rFOvX3Wov9v2
+NAocXxsoOyqA7Qp6C462YbzuMiBBxWLo3BOiTL7ktg3mRUdiq1mo0COO9aXul0e
AU+7dzMeFsxNyBENt7ElXugvlrzMXz2kI/7ST1llsnJKn5tScQbNWbWbb4THuktZ
DP+s65tyKeHCloTiPupWOkNg0smYtt1ZXmV39cAlyul2NuVnasn7+0tkbVJJPUtJ
rOasvd+oU7QWcCzroVxOGvVKOQY1xbpCmmrZ4yWVKdmj6JuitO6jgGrT8Q/Q1maY
vIBgZ1Hb63XBQ4YPxlbifGzNcMuXY9R3CuGDsIMpc+XPmVcT88Ths7PeM5h1SyL+
rI56cneiz7HvOw14i7b4yILIJ6dpT7qgFmVsG+g8y9gMR8ZUKBgu84cN3qexEmfO
72xl5afftwiIQThyl3lvm9EQVUZFhySECqkU39Dcb5W7NVRgvOg/T6ygUxP2cfF7
XTeH7Dav9WItBHuqdjxs2q82VgoulfOQNIQiguT/rZi3dFirHDxEhd/qwzS1cgIU
sCpsXG0EQj3qcDVUfdYG6VDltWQiPW2DFqnEGny1slj5+hWRnEp+O9KZuscMY6JA
o/1hEIvJkxKOe9JDYTBomxzoL1SPik2TjYf6LpNKLVZb/DDjMKI7MdliE5pRu8x/
OpzeUjkwul8iQ0DSy3R2vnpIa2g2Y3SiYFB6QNzc16NeGkq3/3JyCyr35PKyg/yV
c1z6pJ9J7vWhFaM8hTyIB5yrErD2go7KbWPFJMb5hAM2uS4kC48n4hSdyLM3r5hB
FmHmiywRs8saaeDu3G9ATC/M/nIpTUqXRUWo1zNW1PVIwGURERCt9A+BimxOHw1V
qWl0X9Cyi8YBYRYJbYUKFQvOZuOoV6nfOFpQqqD7CowtEcBhemQg/sJzL4Gd0/NU
MHpo8BIUBHdqfAGjBTXff/IM3pMThY8sO7RqBlyMNBRYwCTOPkHHeH9jQwm63ED0
J2pinVjvfGIMpvC455+aI+kl+WFSXYkQ+OK8zAaylQP1MbaxL4vQAp7irGt8S+ET
hJo0D3XlZtU5wj7l7xFzzDEhZ9ZrlBqbOtruJ4OTPbrbUF5jrc/a7nvslforTrB6
SASV6FUngSvl1akadIlofjIk93OwGvt3gLZMLmvpSRxmaGjgUFmlDexXdlFsjeBR
TFfwuSXBkE5gY3qhERUG5ivgI+daTe6gV9VyCY9vxQT7PxMW/nca0zOyPZZYFGX+
yHgUleTfccPgaZyXljrGy8OKJkA9tJc5FskkPtDMng2viWg8zpuQQC1yB37pCrR1
7LYIip9D7vDAf15+yFXgmx5bbxOxuY43qHPDw0cPwCSq2au+yVZcbSosVUZ2WNPS
T6qamZYCvKvsO69Sn4VaJcHz62sHIWlSXibnSVIFxRXaHD5oqnZ8msDnCx1YiyP7
QQxKicTLCyS8bOLaDm3qBqN5J1Goyola8HgXA4NUE//uonv4AP8PcCLX1GIOalB+
69CU8R4rM28dG5hSFI0i4LPqujadpcWZWVgIYds1xnFyd9+tytBX5lmZBeqarng+
MJZW3HC1zPyN4sR424nxl21vlyoFkhha02AoUGEXVAO6pSAQeDYMkn2jAwHSSFew
tn5RSbmKff9zk9+0DSNv7HUC6F3E12Q3h5QC0cY322k1+DGWN6EbWmbfpqkPC836
GWfyR1J1Ns1Db2L/ss2XVQmr5P8ltXImuILIby0dRHKR2i2rLeueHG9EbQjZw/wg
2XCqfy7s2pfJCTRcKnhBW0GVDtOtYlkisDfHNvoNCIWcvmJoCzRe4C3Wzm7rnHef
2Iv5lQcQkMMUykUxBwmXi7RaQTzgRtsqRCxfdz/OudQ8gdwegOwb/ssaCSatRKJr
128BnkunT3GsG0ETpOGIJAh99FbtP8IgLVTe6b2WaDC5qpYblIy56i05NzpDw7+W
JCZ3+4WeUObzS7FcD8tlVC4jNMrQYaUYb3n6GgQCbBQC7yCRGCgb6e26BD/5SxrJ
0me/m7A1hEAZchL+ixY9g5qw4mir0hEI682ws7n8fFLlXeS0zATZldRjuYE9+/08
wieUEsVAYIm7EIzF6U7Kn+5SeMr0uJSXm7l5PG7ePVssN3JreRJAkCnuj1Dfwu+J
Bvx3TOFpk8epiT2g5UkvA+oWbnYIczBLZ+ylSjamfAqphE6ASkcIk6GEgWd+idKg
SkEA5pAOu/svJTBExyjXiF9VIJMklnF1uETxcjGCKQHZXRDy9OO9WDjP8Y9/aWjn
bY7KChtAPGXIbySnvXJEeMvIkQhwvicW0kOsvZ2PFPXfNqYqgLqMC+uUGJqWzex0
Z0Q69kQqEWgpHFBLJ4ILQa9z2y8QRUDRVA9cxArdLyhnf0pPTSjGkrJua3NMpHqX
4tYOrfdOl68a/sItpvSMD5pu2IlA7iHRsef9fd8DrZcS1h8JmPQf247SgaWGHS6m
LKffaRjdiXqXpoDWsMuayixZjzl7Lj9TughHqnBcy1u6McWge1MtLgC5zsAsvRq2
I/sdlf+S7A5cJZTh89eMBYBolFFDH79d9bc1lI/O15Rz+4NG4IPW7HmouYvX4Yru
l2EYyxtQHuj8IpAeQNRBeUwRF05/cDeaXV98RmUPyb6bwXixMrEGFqbDioUnW5av
1DFzd5PCMSKBq+g5OnSxZbUPGnHmkU1GepBrnROyUl996Ak6cUdh6h0027trl9tz
ZWUhje9FwQayjRH9ZjNaJBTTLIWLB2qpLjYPw6mjsdKP6717MIPvFBrbPTIDWLWL
W5Y6md0aynqZPkaB1jWBeiLEPdFTDxxLPWVZYbjReki0GRutCjWU20KsSf3RhCHo
yfz8N7vcddXN3rZVgA/e4TyRW7eYMGKne/9Bj9a41Ca3UZPKXbEpAh5L+zoHk2o8
wOQF/VoyNN2VoW6KrZxmOyl8ObSinCBuZ4eCklbtTocp8vsb7T11OaIIeHHrv1Y4
s6mCye2vRqjAkr88Iz6o93E9C72JcZe81vOHu+yRnWxVxsFOIT9PFE1WGZPPIW16
FMgcXcGGiF6vUb0b4mkdu7jx7Aw2tGJc5kte4B+FtvLuLe7YJAWt2RvYY9n09wXZ
SDh0OEJDA+94r/5Xdfr+6PvdkQ/1qR7i8Rf6eih3Yc6b6PbZad6zWjNCvLxEPHkr
c8jR5essOajGqTkCxSMkg2YOAWtTJzptlKyoRhbqlZ+Ynw2J3xEap5obPfPo9euM
kQcOUZygLdv9L+gU9QFfIfPIgw5aU+MW/zel949ifTWrCv9IibS/oviB1deuu50o
KIrAeOKz071zo0yOBRDxqCk6Da78/m0s7P8Je+2DEk0OrEX0eciyOQmjhOqi75u0
FpqbdL1wFX1s7RGFCV6iDJdlKP70NXslfnUv9ODibjQONzkUtLV4H555ToBwqXcZ
fP6kUdgspyNQQKSdDgXi+fWZTjTxN5uBJSMHJP5uScRgUBuS4QNTx5DT7/oVer9D
a/HFmlGuVOhu09ynJ9LQpXyA8H1jh4+NV5VOxZrRTaIqlLkdhrxvzgwB6CZ/aNvr
2q4wyJZT5Kz8pvR3RFS6+MCLfn/g2kPAaoMtP3tVrVxZmzYxqziypyoqTTGuXTrR
IaxZNQAh1Mc/YVuXSPpCxxZ5Fvq7O4VsCnMhERYNU4IobpOtPfdJXW6lx1WHfS9O
v3Uw7d70eax0X3RyyBOcxhbOjf7WspCVqab3z45xYaqgqs2QCZ7MdHpopAM/Ty2w
1VClsfdNSzQy9yExmAd/pChbJ8kGsc8HBGaVyFemN57aII9h+dY0o96V6BZPUAw0
7aCV7R0JjYVs7bfPUmINE22rpkpEBle30fiCm+VzZZsbFCTqrTMCWb8W+t5IFjuZ
Su2Vh+ViFCLd9+rtX8l6nA3lBIH+TDsN6r7qWD6+7k8zkHRhHoqgVCFR1jJsj7yG
B51b1sx4eNZKXWHScVOgKSu8A1g+ivfKSV6VUq8EP4cCe0rkL8ZorAqG6RtHqz2R
nIEotSGmmrJk85uj0fVf8J++X/2ijKvcX9oTqR1J7jygY9dfr16dE3TSkUDzv2DW
eoJHjbUX+SmqATaQIywzdrIad1d9ktnLRwF0CsU6fPAdxFRwM71RbuTmjeqFyEDw
Q3jts7p11WLtpNbfsfbJ8mmGbsTXKlfMp5dyw8j1WfiDjCX4YBkbXEzXb3oJC7h7
lmdKF5l4Pd1oCoMKWxvaK3Vll1f4wHpqJ63v9Tv9R2hvZXvBk/wo9ocf1DQstQi9
ImOMJM2Pn36Aw1fAL/RrGd/wa7jr7jUNNeQEvPjQ77VNNWEu+7lV5EJaaT8m4ZkK
jCtuhC4SXtqjzdE3ulrtAZ+zLIc8Wkfb/xA1mV65QU1ZkfMvo9WionIu9oAP1F5g
ujPI4fd1iBTqoZKRti49IxXgx7nFVcdiWHEYe++MNUkGnswCFDuH9Xi9jBs7tGYR
TtcUKJLMqbpgXeLMnCTdeUr+uRBTjBPbWkT6MtOoafy/YD5Pt580r4eyYYHAKleZ
+SYPOaEH/YJmc9Owe9HVrgWwifMZz9LHFpjyz1aCSJvFovA6M69iUAFc/0YDN8+a
qIcXp1x9+z1DS5n/PkcW5NzqaK0BuFr388WuN7gtbfJoqjTXdauhS8e29tPgytYk
SCi5nSkgRqwODEACiZoC3Njbnwf1RX6ymGRv474WUJ5W29hetWJuPFtJwYZIQbsu
iQHEi/USyRndRnMYrb6t1E1npSKM145Uhv3LKEqsp1y2zgNRB+N7T0FLKNQlSDm9
LO3JusJVQIZC2ORzhssxHrK7odIrqIXt6yzsP27V99uYgQ9Na6amDxpMxV6H6WKc
A87ghn/06xTdlDpvXyKUX2PO09aZUJqjizTR11Bb4HXGnH4HuIKaNkxryWZneFTW
9AJY39/XCS8e2UqWdsbAIKCOnqM2YWigTVozaNAfuDSvjr2+n4lkHxWUvXuFWxuQ
KHJI4mPXs9IqAshN3E1AOrahaSfurnRozgo1pGfSk053XTuWo7OxPndQPMW7KquD
Eg7L9f0+efM57u2qtmS+D0ttYpbZVfxSF5fJDgL17aSPky7mDxFtf0JO/FgN/7qY
GMGbsutYRyYhpZnZJVQtBluDB6x9rKQnRsLcW/Dvmnfd9ZYo1M5aWnpCYoR22F53
fU+/22EVJknvTmFNjeEftkZ+N5Kaa8Zw1I21wNdSiSNi2pf908q8S+yctsFjKiYZ
JEKl2mhDCWYzCZFDANXOz+jD/JZwTOSqqd+q7/VPoZF0QDZVFHoUGP/6VZ7+iERE
8aKHUkrqvwWhT6bruVcKTRU4Hfl/emO8818lJUYg7452wGCkTREoXXLJ2lo179io
DrfnVRmVB0g14jcnTghGgg2Yy0QkFH7K6nRJwrx35OdiJn+QSVFlTBn0Pw843+r8
Is2myRcqIFwDfvsl2ioWEiYNN7SsJCTRaW/O7J1Fwo28O4f7AYF3j2QxX9JGmUBp
0uXnMChsLMo0qZDcPrt1AVU7Hnki2Cwy6ImtwG/MHJHQJB/Q2/u0LTDKExKi4oD+
dH8rhH6OcVdVAgppZK/imwNY4zMYqcqYnpN5FjSWpiosIXjB50z+vr74MrKb4EIV
/hkLgPwxScsob46Vpuk5pypLIGyPw+frrF1DUDJC0t528DJJzeAvvJ1ujABH/2Fu
jWEqyQ6zq7I1euGWeOXLHP9eml53Z0DT0WePwcSm+ivdis42lhY0Vv4Br8Sp6JGW
RxRuUwm/3kew/eXJdAoFs3u8q4HCBs5QvI95nE775UxsrgPDlAO3NGJ9RXhzJn8X
dqOUKaMv9qrYn6sb8QnZw8etX5PuzLgJvnja8hdWxZIT+cn7MZiCBbBTq59csSK/
aQA5AtYjqurw3GfIFHBwzK5Pm8We8/7LqJjVFPShBSKRg6ratOUDV0HRJVmtiyLx
XLFimRzLVzY/Bq3570Fbfl0Hy1WYb9bAQM4CcMR5hw9Npstx/CgxeqaPsylqvcJ8
8UBt0ZsqULTCIH110Rj1eD0Mm/XeMtZL4s9DJh1gYd69rbd3BfQ2HbRXEk3/OfNU
JM15HIKjN3IB8BDlpNjQsq3Up08gYEJIZvS7ul3hDGP/ps2vb/dTCo47igneUMr3
L9ZpYPbRjjms1WzfWwfY8E9v1Uo1ydSCl+LPe5cfy+l0UBk92sZKbzxjMUO+FeqT
456Up2Lp3hto7/jQf1A/ahLJERln+704zA1iAVFHCpJsAi/HqfrhFprgLLBOCdEP
fT4wqKqO8fw0HL2RzkuZY9mKurExX6byP9P1/90/VQCU+kFqIqEKLnG0Fn4B1mtR
poNu7KRiXaPcYRnZJDhGqiNRgYR8yiUPXB8+2qqiUGieeUxjt9u7xwkb1C7ccypg
/PM2c0vxjx++sKOFDauoD+5dCIeIXYhLzOmwt5VFrMAGePXTmxpFUr/lL5qks8qB
GaAODkaI5oswxVTyaNTUAt7r1vRToQe8Mvx5HBmb6tpKhd5317shLWrrBBZk805x
EhU8ooCM/BcfaOuENw99fxXVaX150FYU/sactEP3fnEpoYeiQdHKyEViTXOBKfrd
ieKWUfktM1LSBZsp6LbI6e1fzE5ag8TKUr/AlKoAU1d3e/+GalpYIWrdeKiaJjYf
3Ic29CoaQiJq+ga7lVhq2zQ4uqmlhgZ50elZ+FN9ec5d6Y5C/uM8mbMhPpNXbzcc
sQiRf81/ULFr4sU+A3rYUNj07NgVUHwGlY4bgaj6nbORVxpI9IqwjBc6MVwB1Qjr
dVT5oPBJwTl8Bf5PXkKy7/ijbeYXeIt1C/uGw3WDfxpjBZCRMtb1KddCp7AXy+aY
xSjqpWtBMwlHq8Qtj0JoR6CMqNEwlKrT6ccW8m3DY3e1JaZkAKTqkOskDYxd21N7
WOqz4q9Qn69LJp0MsZ69iLaYIfRXSWc2LGByY3i6nWgC1EDXh7B3xK6Mxu26lWRf
K1BKsvPvcp9U3kUUwsONZq3aK4XwZNmzbjAuK5bCMGxwdzQKvaKOJz3mejypk+3z
tOWm9HHcpdzlATS0994tBE3fT7ykWs2YFvo8ASPQXFOtXDrUUlt7JR7KuWfYNhmv
7Fbv0Kbi3I5POhk5+c+TZ6JcslYTUgmKTtdlo6zGGjD4JZRTz5+Rui3zsp3+Lzhp
BGzWUHwL1JsB5MHSJENR2TOU4Pfk2WuHU5Sg35jaiz6yaD4rBpaWaGK2UtJ/k8b9
vP7hRg2eZgnyGKXG7NIOWhpCl/D769KJ7sGBtaudy3aSQi+2tRA6Tq1rjLNez+D6
RzUboo/JJS2SksWzhtO1Ji+8q2/Hnpyzfcam/Y7y+zVoo7h+JQD5iJ38iZUUepxG
0FE0aO5aMIQWq238nBuLmLERMVbQSXBo+DA99BXHSUuhyjRcUZBfp9J24PJ6fcPS
Me5Oih59Al1aZF8kC9kCeZUk+8sDb+GAR+idKODt462xTm1QRIowmu6cxqAucMI6
TBN1AiSc7l0nQTSaduntwEIqmvgZSY2cMnNqD2xUtughPdvDGVI6IvptTu3lTMEu
vnfVLOl5cywCOTzTCHFkAVZ6jFZnTIK2KfLTb6d8LFm4qmiJsHN/5Vk21vaks5zY
+VvJCdMysXe4bSD4WNiCcOOaiI2OrmhftL12DX9Hl55BYnLCOWeeK2YPTHewSctB
3xJhZ++tAJdfMSkQzbUhSZrXckFd6+5NGidt20nPklDKUkHrinG62PAd2jDnCCTD
SgGrtO3zQ3Bw6lrySyauokcNvRuy6qkJA9IF5FZY95gyOMorErWlANtFmpZ8nf7s
oHaOgCJAubI2AjRPeKJWxOdH6gHpiGogGj6bvuinT393fIn7BXLsQTR6eI8yWSAu
9ZoP45MeOBQbF6q0R+AZywKM5svD29jMYAeW7vwSB8SqNAfZtx3OwD2e7nxw6/V3
Ykb9kkpO3yO47eOIAhVWFeM5UNQJAwghvn+Z/e8Cmn87tiXzQDOcnY8+0TV8OCSZ
HEMWIvnPbQ1QhGPEN/mQEoI3LJyyKYnV6SWUdHjFS4LAdv0UW/wt9OatrPjFZrvB
IZNcyccSpb4BOCkak4VTeYQxfH8Ot3OwWvJB82NUBeoLzcwoXD4TbJ+lQ3f+hB/R
POUby/5vL2XIb4RfE0zC/tHjL0mm4LcUIMBNh2gkeoCSCKfUyl0HunhIdRSZOba+
NCvbM44Evv3D2D09t57/VKBRrDbKM3Pqqyq1cvCyngJD6dhXJ9pKZW8OmvYBdC9w
Kqe2SSgDFiy6enJ+Fax7EOBROql2eOh/alUOrI6x8pOcxE8q7EEsdBiVsQtmI9by
5xbJglLUPPCO2uvSuT8ccTcM2ZgvvO6VwrxJma0s4TWJWb5lamIRY+4bsUjd55iB
EoAsciJ/3bkYMq0JGRXP1PF1MzPF4LkltANaWPgk/8gQChvm0Cmx3RKXcCJByRga
O9SmbiGZVpm0Hp5XSPnaREPDrYmPZZMU0S3ZxOqbRZ1+bBknYQCK2kwncpNqVpS9
dI02rj1F1200aEzgV4trk00IJj3hcPVsKPNYZ/MnOSXAQbC0kjBA2XahEguIRJCk
+MGSIvcxTRmqd7E7rxnpv/RRuWahARjrecC5VC35z18y2qdRwd+K7s2T9TShxsXz
dQmaAjRPS8H7PY7k/0pnuam6bPSzPZoQLAElnlhb6QR7trWqF7BwR/JF15NYuBWQ
NyVPfYUj8ylJLOcbRenARQiqm57Nl5rktWTfGZtIvyK618LMfeCQXa/Eos8P+94d
VidE1ohqX9Eu78Rz4unpKHZzEvGh9Id3qjT5M+IdmX8J/4NicO8VAxwxNjoWlDhE
ZKVORPLlYvp/CxKtnajdVe7STbMhFE/JeVuPwYjV//ggz3c5QJmLJYGLjP6VToxS
Gg7iNy+HFLNxvMAKikWspGWbQm1pNkqKqN+IlrBheoPi426I/rDQA5IlKD/18Xvq
7WWcDG1QXHuoyVjBDj8cjRt6ASc2IRNQMMUMOFBW6y/OTYZUYJZRdfA26J6BoEgV
EKb92/jZQTHn8v7Eo3l+CvtLBeEBZqeoo8swUJ9Vp1vFHPQ+7dQ66d/tzZEDU7Vt
K2+FN/DLuRKeyA96KUI1hVjtxRUZX0PoyzREMPXcD/vbol+n7cEyyPaJpvPa+zLs
BlFo2LYb24B/mBjv+anONKZ4J908Qqy990AuhVViMXdShSih6aJJCPA7kVdAmZOo
oH/Vr8n1hg5tBCEyp4U+am/H2EzhaFqLD1AQR9rN+eeqNE0g7j5xLp23E84cq3XS
IOuP5BznYvu2+I0t6KithQspahTwcFcikHFIfJnoi+Q9hsNrsLAFDtaYUmNXy8yU
iSrQBrXi0rFjN86fzzIoO5gRq1gltc9EmbuDCSP3KlouOvAzqmTKm0WKT9f/mRN6
X7HOVuHjNd8ePmX3CyMncRszSpeHle4jVGJBCevZEQA7OdJd9648nUSoS1BiqHLD
l0lVuhTcVxifBURBrtsgs9dvmujSgtiUmBBjXE6/qdzq0KxcM57jAiOI4iw8TFHP
qv7VKeAvLHyYYpF+4uq15TwOuXBTvbIuPLP4RkSkBrRagra7sTZUknAQ2oE5fIUW
je5+G1LJAhnAeO51xTiteyE9YyuCQoThocFekGqvdIQm9BEKq83klyvPQEY/Afnd
dbHY+Iw4bZPX3gyGPR14nh/vWCASNCBvOHA02SwVPKf5yvsNFk20L225qSJPqio7
X9u3P461I435KuDwOk5mwy8+6sMvPetGvejQWczstj0zEJmNilOQeSKX4cihCAOp
yYqAmOr2TdwDXHuUKdXjExcFcwm0twb8ZCxWIYVl6htuuSn/NowKAjpiAbfIAvu8
dvptN5GCcFjKxu7VtlaeKEAo9rWyZH6NwhO51Ppy//4Jx93IYznaRu190IuCD4hq
oY98+FaMoxg6hZ4u2OpfYVsckv56ZkdqsXGH16kpdLA/OCzASnguP9wG6yiryY+D
9gGBXxskmWNMXlOhaGJ8jIGzHp+pE0mRUgUQ1jR0W3NxaSngBwQDMI6vI/1doLqM
yrzCPhev4F7ImLrE16hBzC1o8nJDHPrHfX6NPqgs/EEWPieGGyaqnUB7SVGREyVa
RGntOyLa2G7y7znPO2PF2qMg3x6bR2CVSJddWY+2oiF32j1Jty9npx+CB6CaEibG
M5hsbCbcrf6ruu4AVZgKnu5Ob79QwMnQRGC2kKz0blVQe7pS75t/OlsSR3Drv4Pw
kSrYSBrceKB5T2kvEH9TBQT+3S3Rm5qVAW25aFl2UAviFgILm7ruZJ7QrYMUm7PZ
Tz6ZoqqjSnItKtVyxRL7SOGKhtwRVcbzesy4ciO3DNkLdn864Yi5L43q8zNY59PD
LI4xs6IhPAYrj3Bi6GJyfty7ayLEbW+h4J9IsHWTQYSgO+04m3DpkltUIYz89xfq
0egRpeEIyI4LRfj4LTIZudBlULdcbWIwMscfc6r5Hur+LTB0UPeLJDvnLcoXHXT7
YAytPW3cb+eVvV718KC8qz0nhofmiXmyHRQbrrtU6bf6Eiw50oWaYlhJQ5SIGbQo
DZhXbl7wSEEDePhJlJ0IYwH3R7PXXM/8t2Ix82fx6bz0ecRgllUggCJkqGIey20j
4+jazG/BjCVg8/ThQlujDYrAR3QEKoh8RfK40Ui/+UY38eKLWrqQQTeMlp+7VAE+
9bImUebmZhCDm/5fjRNC5DKyUVZ8/+NwZjASbRJK9ZmIuHOiOIXMmG8I9iAqpf2I
0OOZkXiKNCfWfzAv2zxbu/I7CCdq2xnuJd7ZL2WYkxPyy97VfjUvkSzmXkBYurq0
sqFVULjolATw0pRkx2Bg2L18F9gVolZX+7oSy58ngg+o8yGCmFx0UvCoIVHDUpHX
hjnAXDDjp1WcmVf1AVc43O2zQIxK02rTi6cm+RD21O6tkykCPxq/bfMNKn5ZvTgo
WPRgYDOHvUO7nEHW28CG4/DkVPKg8z42x5yvBop7UdgBw8YR/8Ymh3pePYsFsMMr
QwJVtoz94yNZ577Tc8tOyhIMLhTkvzcdt9ar4tvDoVU82sYBfbGPm62Z4L7fXrLk
Tr68eLfu5mLzmEjIh0s2cW7QSRobS3ZsfBLUxuG08ObLz42uWviHxMqCMqpW5mpi
vHXaDZluThP6MNScRLNa607L0Rk81afC9RZBYHxO/3KL0rBevwKNknzrkSehUQfw
DlT7nHCpV+4MJmqa7n7nm8eXGy8nvkqz5z+CJ0nJNppoR9GMqXc3JtLSB5/RmePB
N22r/m4FovQYmDGtS45HclfCjidxvORY7eUct9gyynyQEWHyGE/DaArv5Ev2hubu
A2/rPpy+s71/WEm077KQ8uA96N6I8X/JEWbEkzYWaqv2uJh7U15uCPSVTZUPQ7bE
1qe8HknjPGfWomW49f+HxEhpg9oePdsfOuwzIR4ku0f5t2gqpXWX0MXU+mIC9bc3
6whDgLgrsBdXm+5rC0cUh/YWGxjFqeiDsjD7CROxgO2R80cYPZM/i3M/MIE1HKbL
+9BfgO3D0hjLUP91nVNXJxtwlklJEgUeDUqkIKmKMlWEeu3fXFC8Y7mHqzPhDHDb
`pragma protect end_protected
