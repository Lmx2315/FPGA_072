// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:32:38 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
LFdRY0wsj9ZRkM4wsc9kbthJozxM91//tK0TI5c2zVGRWg4+RD0UB2ykfQkLJ5Zf
7YvXS0+/lO3KFEiA6O2XJLLb+qesSKG9RO/G12sVqJJ+afJa9a8xrB73TR262zJm
kjJMO95oB+F55P+pek+mSUW9joQWi4AQxTGf2pA5s+0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 33696)
q5yPyJayjmwwijcMJsAiIyu1r+69jDjJJdEm3oB+RjTEJeAsXigqcKCG4oZUNM8e
vLtUyJbvFkI9jLw+55BkYbGkhfFdPwOHw7WEGizLB//SbE7nYN4N4r85qbqsmG9o
omLaXdU66ZtE5ZPjQohphe8pSB2NB1wqgK4EuokfwtfE1rWoEJ8Y/S1YkMimBp7e
YP7nqNASnakFxfJFka0VJsIJugcFgNnYM0iiRWifsYOZUMn6Fx7UdH4cOF7quxs6
EveG4qlV90VbKKCofriAtHCaIRM0AmzN0lqimLYqt50rQrg2sNvXhshn9NyFiGcc
6jBQSXzaRj+6+5MeeuSWa0PwlNdEknT/XpKB8/n+HnNF61o5lF8UQfDAHSwBum6k
BC6AME2IzvkqgowNCKbxf41Bz2tJmldVm3j1+8/h6ppYGeCHxnnoH8SorioIly1S
JvoGlKyMsIn1R/hpIkThS8CxFat9xRS5I4SAViApgtGi1G6kDOWaH3JmG+E8VC3r
XqSZx4RAOoQcndQjvhuEt56Ce+8zSSKc2xLqdUyxcHEdYe0MARx58FVbxAnJCUfK
gO6DGpN6gvrIlPge6UNEQbrD07Da86cfTrm6B4PaqOSidEjvpwBSOBIEPgLKMNFQ
fBycEkI+kq+ty/Soh2sFiRJqktuOO9U3tfSayFpp6Ph4ZWkKI2Pgp0YdyJTcCXq0
1azkWgSR5wQpJ+vzzicPiqjMFrW2jk1bf0sW4ZtV1G4vh5GiVMSTRnteqyNWjlnI
t7sJ/+5vqHVRTcS96IR5KJ7gMheAv1j3ylVoO3J1A5eTvOXsmwRMr/b7RVYfsBN2
nDAJ2ARZXHgqGQ2iAUrGknE534U80JHXWWbOaaJseOkyh/5C21Em76s3mrzXdb8x
SHpIChLrf2UINdzFHQl1Ck4cvV4WP7uhuyhvD0W7xKvMiNN9XUTZeBcTGX9BqWSl
W+CY5Ba9hGCFhUaMsWgiUuVehQ9Wev//RzjYqVnb+QCUhCKs3NV34bkLGNTvHt81
rdGGMWni08wzO9t6b/xofSXqQ5klwXViOy9S4o8jkEuxhov9QEotbVoLN6KcEuew
1O5k8HaTAEU7xLsIx/ooQB3hetgqSdJWfsVQrZp8fvro/KGt323Ifw56l3ts3K9S
C6t5fEsx5L5ik5q5X2p+XUyOdwhO5K5GoNwbtvw6ewbMsviwaRljSnSs6XsNqlNC
MNUkwPJOG77mM1fK46i8SFQQ2Knd3a4X667Rfk0PfowsQ41uWLODTh7B6EPxp/bR
XdM0w31qMh00bNDfDGbxK/uHHx+FpszbtTZaPQUvqRCDkrRhFc4pwniF4f3BETpb
3k9pOhIwxssx42bo0f938z+D66+/hCLmwOz6mxuuMLsML/Y3IEFn0iFIbUhgPQqQ
RybEo5wI3O0jWBuOfWs/OZEbSPZvTms3DpBbyHrnAO6FoRuU+tIlvJYdxURMVG9S
3FKSxLKUPJ9N3cO/ecCrYE7ZZhNgUoW8jZFyjNwfFzM+r1ryzF3K9baoDvbbUVnd
A83X0WPnJb4VqF+CxLVnkRI8ajZtglfBAbQgtuoKfCv6M735yxYMr7YavsapR7ry
i6G9qE4n7sJe9POO3IfoJtjXyOZ/Sd0rktlyvkvqioGd0oY0BrL/DP8QyJLSWlfC
kUaNfDEvV45FcTiqtLX9gtR4p5rHvH9DmH0adYe3IoAtej6EBC+y/kws+VrSp0e6
40E4bKUMSMqKKfnimEBJQJGSIx2GnVhiZRFfqI09iHtDVSHBgaSLRojs3UHvq+N3
2zHLInCt01FpEw8A6nmPXcurfFMIBd4h6KTkww8EO0V0abAizlqr1lnIb1GJgFFX
ds11SUDk47M7KLVcKkZjty+6WVpilFSWz04unUgXnrrDK+DHB6aMGLZWbmu7N6UY
67TqFodFOQOqPlPOZTtggGv1tnKfYJO7vj4pS5QLO4LLf5431pV9mpXRyY5lii9m
aJoTb6QS9A64nkKvAbExFB+3zM07nep047uw/tQGH4v+/ihA9+bpSSSJiKLCbxnq
ebonAjHx2rwrVlKivjG4hKf0r7n5C4xjdWDLWhP2NWHiuNIgqN8Dl10WmiqOVnTw
FCQqSGMGfF4U1FJhZfpnoKn67RAXPox55a9Ae8b2Yak4bBXWNO3KilUymXaCZCfk
bMu03K1vamkn5am85EsavKWmhhdmm9s2a2KQXXomgDR++0RCANIj7ZHaZmBTiqym
Xb8H3FGFHQNbZ+PWVzkxOOJx1FsH+VOr7Yt+iGsQe6Cf/jJzcfdc11cSp34+HGg1
R8ccOYJy171/EYR5V0pqg1AxnddGQAK6Byp8TDzNEha52HuA/C90DwICRHH1PnCi
R+cfsZedCfoWJur9+vZJp3M1338nxsH8GUzS7iWwYR5D+/Q+sicJaZLZCxysmfWG
re4FMdgxJgxUMPuKH4B2qNGgyM7IZLBXfC0GtnHma+7tGS4/B+cWVi7m5cYdcITf
jqq8ZIMDFEMuQhA3qCsAkRKxuec54V5S1tAFVd8vawqwBEfAHT4VSsegkeynBJwh
4E9ZOcx3+Ptr9csj5qxrdcLgUntcBvnh3is4TkMskBcR9hg5PfXTx7PUlH1P1tZF
Z7mmNXnVi5k33mNKQCnc/hqH12vQRnvLkVA7J95y3ab2d97dRfL8IwqyaOdbZ5js
Bj0AxrZbGd4DGw6+gFfJ3ofViYrkZjDRJBttUx1iLo6jgXTf4FyUY06MzkM6T8JL
PwTLb1DDnWsVhpCxYCuilCrMrDxn4En7pMCa4AGJVoob8EbfKYk1xnZPYfZtr0k3
5ERrvkgTkQtgRqlH1/3CzG4reOHeVzM457jdljGfkKuezRceJ5LXY4+tIKzZX14i
xnPY//oo/4pDeNCKFp68I/h6JaTJ2TLJPQXiHFq6BwjaPHqorbdI/U4Kh2d6kWJ8
1eA39G4aT+5mIaKZZA30TOiyaj2yaaMuQg2QFRmygvIwbYyXLgsYkd7xgY/Ktohs
aRk3G1+iyjQEqips0xDUHAFrw3+mY6z1D8uTiRV3DUgtJPynLp5s3yWrKgNIqRW/
lrZnOwrOHVccQBEYwz1X5+/DmgMePl2PADiOeDLO7fX9dv4jXTvBek3l+mZjbwPY
Fr/H3B/+bOkj1U9xp7ZB98qOBn14uXAyZvfqg2woNeGFIZPr8OMWPU9Bcdi2QYgy
9Ggh+XZmc6uEvUWqLVC/4G/Su9q+sdNfiJmMc9bDFwx51jKWwO0uDrmuRG4/x3Kg
g465aV9eoF6UhO2SmUXM212eTc3rlso2vFjcKzyDi9M5U5wEjzwQzGewnk23anHJ
CMtUHShj17sYF7JVi/Q8Jm4OdeITrNIy7hp76Hnleqp5IsxUvOcuUkCYDDR2qFDu
5LGoYmjAL62I9PvDuQOTK67iHpeNwnaRuO6fMfoQEZm4etaKrLqoJwfr82/HSg9y
NK0cMtJUU/7SoqyDpL2wY1iJ7lEZwgPxeRtWVviEm4G6oAuguxkdDSRMa5CXnQcC
dc1c/88n0Qc7D0tdroQX08O+ZTy20HpCuLH86Sexbb2EobkW2OG3CWp9551dyWm5
ZtfFX6WhlZBGtfHi707Yy8MepU/ujDm26V1OAbHr6Ef5Q+JZv+SIg5RVGIgbByvV
Vs2gvUfJt5/b6l7SAih3ZS9MpWlXEoi/UP6Bu8L+XdI7MxT5tajv0a+J7D9UVAhS
lFIAdyje8NBzo0i8Lmx+7gX33+CySjViO5JN2ckQkGxb83BNryOZsyr7cO369LNT
qdmJNp2tpB7u4UHfA08UIs1iKUYg/liXz3vf3ObeVuWhEEA2xNHr6o+wPhOxhW9A
eKpjvEmVPzGwYKzqB2DzC/wd+xdWBMcLhQ8EC9R07BQTInfCl1lj/mFLYhY946Y8
F0NAQkMh1di77t9axWWl3ylVFefI5+FAvCXX6jPsHpY57rLAMFiyeEioMJe2fRxB
k86yysPoxYtMzGPkuk67m9aWbTbFo7b/hbJA3MpFCGIG0M7M6TCxHWOA4jbR27t4
kH9V0J9LCr+4EUIa3bI3V5sgvVQnhtTAG7rLofOGPuehCk1msgdJohWHmwhuAVz6
oSaQW8rRrkDpKmkMrBI3cw30t21srvlOkHgWlVgfKQpFIlYMJZna1fkCb8RsDcDG
S3p+oto981efd9blWxtBbE6RFVJhFFFrzxE9r091Bb6TRqkHsPuEcrm+y7KrhCSO
dWOYiLMteAqHQdCqXMjLtCzlhRQyMaF1DI1kqWPpgJKGTcmW81jsKN2iOUpqDmQv
usF20pw2Mi5Zoqdxz0lBaa9nisvH6OyT9apdjhsnUDjonn9wXx4etP1Wxy0Nd+a9
Nr9P10O7Jp0CGq1BlY1Q2M4ZRgJScyhxmVrGg0bBKUV7AZ2PcMKZRLjL2DIoDXTt
JFlqDSidcqFtcOiFhOGI71+J+6Ky6LjY7BOToiaOzU6cQeSVcN4M9TjNXIsbHIOt
2K1ih/ZTXN113jGBO608/hvu0FV0XT72mxCQ1oAPuEIQGZ+nFRN3j1xAPZZju1sf
uijKRQ8OD3oZy0JkcqwfU+sLxL9+t6VpuLYMwEeHMrikeYF5KqZJjW7rtwwpOo2P
9CTmHJQqQYwq9ZEkdQ476GnarqXE7MLg6G2SIvVSC5MGZaSYXXLzO1upVgLtwXZq
BQGE9NjfmD7Ba2iR9f5QsxFNH1alwA2wmTLZH48XCWTiKqGaMdhkMLRRfgLFqtWS
3X6dSyy/7v7Pivgcxr1ZoiQjqCsId/758qGRs7I4k/QXlR9jhiHhUWlPpvFY97f7
kfXgkCWazoqDrXABQ7CxhcYKq39QQLMimh53ujfXdwjI/Jhp+IGPoiPQQdlVChiX
ihtrQsI8qNQNKTEAffuRwsjv7Q8GzpgOtzExbfmr27rgPzWSlti6z7u2Bl3WtBwF
K5shvSHDP4+RpC4aDFHQ+N5Pdci4oac9uZhuOi0Zdl68LCaVsTAv7gwsK35Qng6d
JgoyDadPQFvjAXw+ErMz4zuoidCM3+2LOLFOdlvdOJ/veSGPjmigb4QT6v4bXXIm
EQxQYAaiYqKMQyD4ZqfJGIFWr1cIDrLKMNF0+XNUr7+N6W/6eCkcySayPePTALbn
wXC4+lRjr/NPcGnuBi1mrANxWBiXuXQaccr42/BHUiRPnuJtErdhAVL6zGK8mFpa
3yiJwe7xXOI400vJ+hUDl+3V6MMz0bJB0AieyUVzQTAnyTTXMjvH9xZBAlEiydsH
xe9dkRy6DdrmyHftUwvnYWW6pQVfcvEwNQaxiSJxIj5ZI3kKxTjf4DAL/EybJJLO
qvPUIs+4t3pN+WqgTcWycpNt2FmJSYcE1QQ7VUpv3aF+tH9y/7zZ6NDsJDrk7Eep
O9xCH/xBV658wcTa+XSFVztpoRMvYi/0+d1b6UfjvlTodVxurRSKzCZvLng6D1bI
4Q+cGiSTbDJI8GucGXHLVcU+04KtphXmpRGOzSnoZMhPtKg+UrddcIa+40M21wIL
pSIbROshrGrtD+KyOmc3wAHq+cRWLS4kl1z4JcCEojNx4h6i+5xgOL+skQnV7Fhh
yhztPR3fFvUWid4SshVX/6SPdS/RoGBMCSy3dIdGg1wvidpMBf+SVFCyxdXxR98d
gptiOruOlssqC/GryjJHVA6gUGpuFSUFzhH9BT6c4qFmtukc8e5bOrX4Ffh2mBBo
U1NW4P+uvcbbKhFVdDSvMN6KCYlbu4ShysQ2lld3C0eoZMd6NdOCoa1qT+lSK6Ki
Cx2UvSNFB7v/D4K/F1+FKBWpk5LaEAJXhwyzBJ4vHH7AnkMuPEUn9mfoH7klAdoa
sUQCtY1gLaE9F4aE08sEojxiORBFXg+HgU1WOzkRHg0ycsZAhu+4Wd8bN8DoHSIE
BxiKFR3osJr/gWu8kONewtrXF9P7q0u5Jy+55c8C3eDgN2rypejN8nER1llekcz9
G7/+uEtUxWd2upCib6ePNNcMOCK8rE6hGtNkaGvpw+QofDYL/6FI+JtcWLDFM8yG
E5ipsyxm8ltVGSCh3YNcaYWlWiDGCEatFAE3Y+YCG1h2F4vSiuEHmPPeRxuFxRko
sWxbAe26UcmzT0e4yGKYO8EJhfPdDHqWYR2aBUoPVlyL+iNdGMWmy8HvV04oQRah
xxMmbY9+iCP0Xr5FplQ7MLju4ZrCQpz8NVILk7u4JavshAAwjxdXndzalPAQx7sP
dz7M+em3827XXqFzAB7alsLZUG7cUPuU54Z3SufYWI8xS29FSDQQeBTKP/32l1xh
5YI3dQs5oeKTdtC+T5ODmkvehe3fCYEFJHz1OBaUK6yeGthrgyVh0w1l0PXSLtfj
4H2m+meq6SNSCcubE4paKcInJZOJTpmzcqwv9339os2BtHhRjcB0T3jebQXNpeVU
3/Dxue4LPUxOHAmLtk+hsS59BsK5ke48J1JTtZyc4Q8LhISV03hnZm2mEca4QJ77
FwYxNQOPgCSo+2odhOKYaON48fzjeyY9LBVClgqswYDOWVcIZAKMQaG0hpqErMsV
RxYChBfbr2jHO0JJQBkYtmjpG2XucuAQV1qGdtmLaCMPYGSfD7ll/Z43LUiGF7Vh
wpaVBIF49j3QjG0SL4u9zWUOVWNMmscuWnvsZs5hhUX0eawRwMlSzVdPHmBVwd6Q
jOEhCNwD/CR6UKvNegS57iFQhYeA7j7vMeHQskyHDMaJOkfFYmdVVSSYq+QYH4ZC
nOyltfeYUnOnNJrTRK2wFVP094STFQDBpd4FtUAS9RUULA5NpyBaf2QwQoN1ibw4
ifZr3UBE0SkOsk8WnjqD/OZq7Kvdpxv/8dwjrOBV08O9AC8BSXS8tApfizJTdGyv
WmfsLjc4RPxb6+GsinZkwLdJaisUtuIHVCOmRFENsrfZHIenS8L5rGhbkKsr3x51
Cl81LKtEjnuvUDnOxBSNhO+bWq9jOta2yRUIYFhDYEE6j3+miP4G9wgfTubKuUd5
zJh7iMeLV2EC6RBa1+o+9pBuuThpJhHVI19OIomMxrVUd5f0Rgm8zb4T3Gqxr+8/
4GF0ja2OGgCVISnYH194pEglyJ5rBUIhatweRZZmn1Rh5rP+vB2zai7OLBFZ+dBk
SHRuSoVJrD4jmiWXHcOD/Bk32y+7ffBx2KO978HcBhNRx7EHyidG3bxkWPR4wlPV
xSH6o+8VqBTDi8j0aXVaBLDr8oUoq+rgqU6CBCe2ENCJfXpORzLguqJHRWhdEEvH
L3kaZp22Uz7LO4p7lMP6Sz5MW2WGaP28ZgfjzOzipuXcpqOw+VXYlNY4VBu7OiFV
ouiWA9mzp7nA6CrW0Um7ydyEylFR8fIh1NX/XTLxxYqhT3RJU0wkn2clO45z9eue
9poW+qJ5n4jL0HLZD2XbdIuKRwkCcEtze93vgYNqaLcT4UEfIeSGqWj35mcwHkT9
eqAmuwjOlq8JV4jHLezJVB1xXO5AQSOHjCLBElQSLm4oKXcukyT6n+34xY8SN/Qx
/A3fO4LmxnauvF350BGNdzq9PijVkbawako5hQBifdjtHLzSlGpylyExAy6R9PTW
zia77u3/6j5ULyFldvZM34bdEcB9lHXJCt2+m4aEg+Z85pnTgky9umz+2OjMeyuN
owKQWZ98uD2bwrNGLRXFSYt4zjBrKs0XblzJYzr8l8T3vrOsA2SXlnDl9RTBf1+h
tNAgpMYA2rNfp2Pez3a881EFQs5gMy2hqG+mPKxd4SrlfKe0nTZRMB3b2mKPTVJX
cNh+GcRJg8HHplB8Spfe9sBo0QfEcb+ENDeA850uIiehhYM7ADtwAqHYhDIyrBp9
C2Gj6YucByUkBNzkgBe2wPU7vV0GwiiG8jSc74f1AGgNbinz/OFO+kxX9glTQPC+
g07LLIPYhkCAobZbt9scLZxiicKiZn6F8g2NoAlG9UaKcuM9afhr76hfpdFCVfLo
6iCnBMoXNQ/6aw8S2/keUXv+cXEANlQ6lf8fz5muvdYok88NB6YKiUrRC3tYmMl3
ZtM7wxHzpgJN7FuDuQiQQk2WBJeENl3fLhiSNz5emiMy+1KlJDmx8vMqW8SuNqhq
nWFPWM+nqShDRclc0Hjl+/nLWkyM3v0KdnnI9G28HHpxFfloxeSVZQgFqbsqXUz4
g2BhIGKCaGQGZ2o6/z9qvlNKl2saP8yrlcLq2VmffQNVDqRE6fquNI8P9ps4rlD3
0G014GzS1yMCmBGicCaLbcxMKtQXuXc1OqrgU83l+nQur2UwN9mDA91Sw8BKYN+C
fsCrYLIE7fee+Qkg5Cf3Y7hUXk9h24Eat7TghKCRGcnwMVxPvxfpHKZxiSQSrLVa
ALDKkmjgZ6WvhyNH8oOYuTZVzo4HoxpZGhuMAIJeW62YhsZ2awYTS20s8eMGIVEO
ZLtGZ+qWUNEugyZKnhYwpKGWZyaKsCZ5AVD0rHGjbIAH4S8A8zCWzDcs/27zIqOL
LBj+mDZ6YjVlAKD7X3N7e/lWHrxjZyR9YUGU1dZV0zRmrIYRLCvuY29bPTzbxqah
cMhaXCPUdX7Q46pxbLDT+RzCWf+cyxAxphCnxzyJsUHFN4G0xvH4BL2KnOD65uZj
JjBtaavmMEIpY4Q0jw0Xp4VJzQ1VHf+w8zXbhrF8IhetKbRh+SZ2uRvF3jVIZe9W
wB7hkn8lbvnvSvBugjfP9dRvqfoycgHG9fNxfn9oEzat5DF93u+jy4T8x/G5nPqb
0wIYPXCyq1SM6mfy+Bh/myjT3cXXjxS/9GW02wVAEmGsAJMR37GB2YPqZZzaG0U+
YLuIhVWC1+NpQZrTRQ2Q39+/SGtYiHVU0+Jo3fejDlkkspXkzg42xcTrBuqbdT/q
jlxHmBYpSpgiZ6v7oNZdVKyH22XUY4GaU3oNGfDZigzcEbpQv8SGTJfwe1JVP+eh
Ig4bXllYt3oral8uway0JG0IqKjBoQZ8GxIpadSMb/x8t2S++C64O8XbiIFk7kW7
oS489VON+wtoHuDOUTQ6B9fuYK2Abm5Omxwu/KkwlQ7p+wGPZ1iAqqUkVLZk7n5J
NKi7zuKWctV2rGfI6F6+wn15pMGGhEWjKkAhVj8RJ7panlYSki9MS/zldWNPEHv7
xH2OCZsxLykXTsdOjiRRYRmiTzd87aoX7diBiGP3ySZcZQbfOfnVNZHSHrGB+O0s
pxXy5LdKsAGimpTqj47Ti1BSc2GdkuLKb9dYU1sw2abhxu9hhSWg+lrV3W4yUM8F
QRavWy/jBA/FZeYpwTr9zJqJuePcNDVkYZvVCoBY6VF9R5IxFkYUf8cX37tWiTYP
ZdcI5bHSKuVtCfnhp3UT3aqfeMdcOfgxCtsrQ6YBvH1PM4eQmTr8KC6goLK57KqI
RKh2Z/fuYNQpSDLaLyMaf5/WWEdH+UC3KUIdvndbckmOjKqbLg95/HCOrIJV4TBt
v1sirvFHclTiJZswl4bykSVS8PcvjPn8rkRJGOlX2XJIK8ji4y68djOFWDpr/ZXE
4pl+KxJUFzZ44XOpiqeQwNRRcq1Fbu5WyDH4Wicd20Arq36VZrm+WrOwjRd1h8/J
7bgCzXK95EkUkY5MUbcpkjKnkF71yJLKN5ICoTF0JjAJrNFx9dULUA0L/f3btwqR
c19xknx242nBMvAZ1DIQxC+aNn5LXaOiRvhE3D2f9ctGTGVtC8PO8PMm9ixtVlfN
/6ZERwNVfTROcEYJLSl+/XxqGhICRlcLgCJ4UDE1gnfv41eZZMMEN3IcAFVs/fpf
sWh+otjLtk0vgdTfKOlKgKNICcQyOoFhqKpto4X3q/FAbuxiIoMXE4Y/mGoO0v5P
PymL2IhZgbx8H/0zFI0pShyezjUCK/zfYwqs8TEpw+BEk8V0FoItpivlKNHRzHwq
U8+5BjdaOrwxvBuPBPUG9NI/gLSiwmXz/9FWLTIwmCQeIP3O3Qay5sGX1cEBzbXX
sUmnxANL2yHFavD4h7FgeOtEdsLp5VsAZmhJJ2u/7/7L+awEmWuqIke6W7yqo8dB
IuCfV4mhQksQ5iuR9YuIC1p+9A+pRtj46HYWs6Ci09+FtiopMHHGODVPqJdnHyXR
KYqZL8mFX1FFmzrsYki6njScYwcxRXtjdfgPiPIYvZH4c8uDkZg9evzusWqVjWuM
cycx93k7kTvhc4mJsvXwx6jGkJPvjhS+MFMGUe9a0j4VQ+QW41aGL5EoEhvmBQy+
v4E+ZA7SLm3ZudywOF1ta4NRVx3rKmy3taUQAU/yp8uEI/A7AbZBwxJv+DdYw+NV
AZsFEbOkpwJnvXc310dkUPGlsEt+uPI0CQE4lfajqOt+WO2E0SeTOT9fapmZaUm5
mMEUufTToY9wEZ8AVZ2plkfd+UzmUmx0eaIoZJswObPXlgiBY23ekkcmfDKy+pYW
Hptpv6yfZnhAlTRuasatJ3wWghPStrNbWJtE/dgrxGyrWYisKSNwPI+yIDpS5wYU
Jn/soKW0O1D2ALfpJlxBqNxT2p5J1k9SXz148ZpoYzYEnsd0AAshemoKj+IGVO2g
adVxW4xCmdtfBZeIwrPQneYrzw8qJwNVRrpXIGh0YderZ5cK9tmSfB97C8LB0oqZ
o+MjdwGfLknbyGAa/HJ2ceUluGe/YpXK32woXyVBQANq9TPEeHcU59Iueg9KO3u0
w90Wu9MCocA5I+UU1gujXYqxE4uBcb425T9V49ch97HucSzUdrP9VjifYXIwQgsK
uyJ5DKdUb8S+eRjSnTfYUlD25hiLZOZI1RaiZy9uuKBqH4QEjJmE7cryYlni40l6
/8e02a8dsT63k++8j+wQ9829k+O5lNoOvIaL8ppSvZEupPZ+TYSxSFF5JV+hBQxe
bC3zFbpZvAtpYugJ+uY+/BaGJIUR6KK9ynP7P6nF0OqJevYCPHuV4vUaHNvYfXw7
Z0yVMtty6gxYuz9tHpafu84sjC3+I1TQzcNxa5CBLCIt8lToZ19obi5lMHMnPFQ4
93wOZI/RHQu613s2JRFwZ2JiEPryoqCAQLBpVWbMdDnEH0poSbsyAPqJGBC5XwaY
uGtis3mxz9yeJ0/iN+esR9BrOEeL9tC5Jz+PDKIpUDVUM8Q6B9v/Gvv51wSwmrix
KW2Tp+8Ky1pxuSPFMLnf6vcXVHZl1T1bpIlPdLgtKm9TT9fslJ6lOCo7alWiK7CG
Kll8UyXpakiJPHPRWqXrRwiaihDa5cYUEFNTW750XDPYQ/ds93UAHTqPO7dX0pB4
WdNm6jv50Xdq9K5BcWPn240RMHtfF2adOyqbP4ho+zWUwchDrUi58eTSYVRS4W4D
bKyHw+P1KTFHYwlhmdglK6oDG+QtBZKLelc2zj/4XZtEhOfvgTL8/egzeaeVwNUn
j67wYi+Hpp+/Gw4lItI9HwPdUo3SFmodyq3Czh5Pi0fSsypmv9gMOSoxpa8ZLOA5
BSxgFMCVeU9345isU3Jum5o9VKnSQtptdJVmN2ojsr1cXBdu1I0371eU1Z2JH/Lj
XRM9+7NtBlmoHtoW2EXgI0fAkgNlwxqzIAnGfOn9RJlIEa6d7cNEMl/QfnV/WQgm
Pm3WBKhCIbwpMwQdFv86GH7P7KWATqXiGYRQLBCpDRTU2ZsN7Elh/Pw31HgC2AUT
ULU++PDyBG25UH2z4HG4MRhOr3X7C6LUdUgETzznm1TB8xY0AJyE31a6qACCTCFB
YMx2+18KJg3gOLcqSkJbGrDtk2jDCqSrpk2MdIH8I4iP6OIFUO7F6/SjCsPUMLQT
JpStt8jYzGR26DEVJZTXicvRWNAkqPFK/eAAN1zGTXTkIqPs7WL9lUa7x5rXPF4L
AyTvGW71/krWK4d8SVUZ5MIL0a4YOSOzmUHpkRr0eZPYeGeldQJIGfOwv/mBAlqF
MX8/ldKB8xiig1E9rPBfCV8anahMX0dfwCT8ncclIIc+CCvIypbr556wW4dj2JU2
U5LDMr1/IeqlE0vaYtBhtgmq61sVepZ+/I3QVB4Bx9osPrhE0ttXHWJrN2DqwkUf
oQ9dAoBvkzKBup7jMi3t6sWxMFAMN0PoorfJOCiDMpiVyfSNZ+AKsiNcvpQj0UCO
3fzU5s/qPFGUabsPcOHHEUFm/cmbPjfxaITMO61oWu6I4owCFRCGVPW8u22SNcCg
tSeWKiCqI1Qrcuv/1bpY2vYt8+dRFHkKi4+gQ/niFs+Vta6JzxY/w5s2+eiLM+IT
PrtzzX5CcWIJab+wLvt45aMVeZPnKU6i2UtSGl067BYNiwfiyYIz2DJRc4hNRBqK
foya0zMIDCm9W+PTXbff7dpdiaG75sG++DxpJX410wHLhm1qcGNAsUDIY1LriU3Z
Pk81QmY4bOlW21CgRpnNLLOnxmC0RG7x1GTdi8AgZt6FRd4O3g+NNUGpe3sU7RdP
/1+q1U9129eNGJq0p/+Nf2Inwx+XA7JCMjW9tBzjUtWhPEC/84PJHrJkH4yMkQG7
eZYjhMFrfeHhY6sif5X+RRYRQIJ2N6UmG9xwFV3yHAVVBwmk0lb931mSS8YPz0Ak
y69fVbDhg8atGDKB6llOK15e3H6ad/CCnpWV7LNyPYw6bjjTkcvUtFLF2b0yOKa0
qHkqmpQ5FwrmVV0yyhruLVSLgbTk9hNhUMXhF18wYKk7YPJAbH2wmNA3qTAx2EJX
jd+PQhljFZKi/f6+Jse2oIGXnZqeSXQ31HMQfo+FTwBo2Mgocm/zlDD/SW3g7btK
tBjyvRQvWRkLUeCgAm590xvyc8rao170SasoXXu95XS8be2Pg6q7+9eJwFjSKjyO
L7bEw+B7idpQukA8iiTwu33eNrGL+Veq89esxoOiz2lvNPsnwPEx5dwLQtGRBzRR
cLmrHQFXUcr2GQ2+SNDMj7kicPsFpOeEVduAhSdE4pZkZt1bMq22qSwBE8auf76g
Ar9eto6VpyVdTAZRE+cM7O6rl0rAU4nJtrvpcrMKSARJXfzyWGd1WJobcTUnP4lN
56bK4g6hoj/0oxRily+P/llq39h2k8c18W+mJg+xcMPDVOTyw4iN9fejzSKu/M7/
pDBSwSl4+klfkSMkTqfWgjVUcD5iYsi1SZ+2HUHWYv6XMD2TqlEddJyMKBXwRx+O
lVlqUfF6G5MSSqzisx3xXCT4OiuyK5qO1GMhSOkY9KOv5l0idymTZTvTWn7QYxzI
589uOzLH0me89Dvn0k/CxibHPR2oI1gdJcZPhalGYKuWFEJRBNdwz5aMmMl0tfru
EF2SjXn6bUxeqaYIcobSTKhvUWc8WQitIYGVmOb5SGsxJVS67duDthPZbTati3pj
PddMxj0Twu+rxSLL90ZMEnsVk+6l/YPumnO9flSZHAgdHhOquGngxpFvBKXMjOoj
V3V5j8vq6cOE6Bey+lUfX3Vf5Px7CUgWZPE7w45Dthj7EdM8fBR7fAAZobTzQGE9
CmKlBdZQwWTqMAS1UzWEBnKIdXSLI0OqrHbeeqhkbT661wU2BuVxFDurZmw1NQEA
XcA7TD+vlpPqDI9ZD2E2kFwlO0419BUzk0eyzElx3WHuriSKWKamsxMQGocZx0wl
ntPGGCR5NYSLS2xfJKpfC48Kwdvi2XihGB4LnM7U2oiDd7KC8zzKrWimCcjDmAUD
0+URQwHcyAtsvyNbVz3sh2XqR5KwM2t9+gpNLYphKLK5UpvKcrbWRv712rV9AX5I
MQL0pvibcicRUGE/m22Q053uLZ9NR/+ioXOK67D/Zzpi7sGxOn3Nsf3uuhVwJv1B
F8Xyz8xXd1J1gR62EvkjyD3PN6gvag90LkPIcnkZmWYrkv1os7u8+Dqf/6roZ8LP
AixXC+VDFL0cdNAc3DlqjLq1tVJx/RMUG3IFXXTUnzHWMBUPhhGnZuY6764MoxJJ
n/B2OVYLmCplid3KIpYlxNf1xNkQiiUJlqNKp0gmcYO4tvqRGzcegvfa1Z6aNHCB
MYOzW6sMJS0q7tNuH9czVEBewLb63lMAlpSC8J+KCqHVTS0uo+ZP1guO5gjVAzkI
S36YpsWlZnUCRMXt2WSB20Hu3Sv5pgmkIKG/i/VKudMTZO/UJ5aSjOt6Av4o2/MQ
s78Owc+uTC2fya4w9Wfri4kwKEL09LX1VDLxYGd+/1YRnRAdkdewv0/8dl1vIJjv
y0yGzg1BqlWfL78U7jnc8IcVe4EP3053xpnt7AlptXA+KRGiYvHUuB0mE9ieIsA8
lcJhBWCKvlWi3YygkNPeDbq1aIxTbpgIcxbs/GA19d+35/cnD+ObdU2p/AoIC6IH
J5IZzZo3VCZUgP5sY7zdb2oQWzs58+VbnuD+Wu0U4Cy32ONhh4kNZbsizP3jjLAz
0iTaxqdX1Rd0LawiTOF7obMPTBU21Jz4D6YrkzYgqWPdehtfiYrsWmbd/GJ4nVD4
Th5k+J89Nd+Cvov4joObI9thmkFYKcyeHr2u5m+gH0YI5TJavmXjHiRoffME7/bm
iFCgSU2GXtPX7m4OPafl4fJKL2MnNq6ZAiJa/0f61z7e8FP1YrqOoO9C3B6LoLMv
oXn/mfIQlIeRTkXsUhRujefEBNZ3AzL3yb/9OPHjxcwdrnNZerEVYJBm/CdMfXOV
bz/BOIwYBZ+kXnn1ntNwr3NoIWhXIcm3LCZjF5J82TLsT0mlmK6fFW2AFKTuaORT
wjx9k8CqITgNxAfqVzFsz4CPV+r0HD1y8IaHrp/q7ymGtymhUxooGjgJKX4CXleI
GFuDODkl3nZYDi25SfHiTXelCB68cvUIArCVPBcl+2V5cnQryuaANq6ppAFj/llc
GRJr0OyUqChKF1G62QyjXd/YHwtPFnMeRt0fKnw/32n3hmHRo9PVFBQlWxMIZU3t
3vlHxIzFOK3EHBKBwyOfoR8NCkQolMI9ciX4QNFSVRPKP0qT8Z1yB47SXQ4M3oBP
eQn9SOX+bMfiD+LVWFmKrOMK8zUWmrWAYOmwnoV/ACBqlin44ppTFuDKpPln8ODL
0A7BVpZhuauHeHoZuhpgD0mRKj7VmQBhGYHoLP9F6Hg4kVjg2MCkcljmpl5t2anh
qIAiUZCaOJT5ku0kN4TVYw39s1KLX/6f+Tv73kPGAA/jFDGkcmyWNeQb+89+5qiI
ZAvrVyP78/F4V/XeO/rF8HP27XrWrgY5wQjhpvirklojBSnGiv87tB4d6HoG6Jck
qOfinVRf3xZdA1QKEUcf6Vu4z5O46ljMIXHijgdmWaf7FggYMJzX9IeUYwLhRlcT
z1h0lt6GFVa3ypVqrdPKvwDJj9J7rOG2vWADaMmYeks+RtrhXxUd+rmkanDQhk54
rmDGi7zMeRywYcggj14qRfI175xJVC/F553Fgb9tDow8P5WrOZhQJo4MOhpR6UV6
51rjJWrS/SZ/Fms2IMIzslBsouWD+yxgXuB7ogFVe2xYVCjX4aJUyosUzTMt/Kx/
FbxP2DSOD/XdK9Av9ju7KjxPvXmKlpfgDAfcvDo8o5DvJWuYy9vwbzq40aHtlems
JTOWXerWHqx+tKanCDsImwrEaZvA7W/XIrTRZHubbiFe5zTKk6MNNcTPzVYfPz22
Q597xd+Zu6qAdaZPhkCQsZVbOcNIVhLXaO4YWf+DYRr9+U/ZlaYRdUPb7q1zMdT1
SUx03Zl+Y25Pdo1QjDq1YPtYdabhROLWgix3BSF9LO5cY9amtRKDA6DcjWfjPxba
yDCOI7UVhilV+4cfiW05hm7hw2kIZZIVFz+Br2u7BvzdLEtOeSWoHEVdBUFDy1cc
NRQYIFkGgd7ayP/oFWCc1jsyfDh2k/VmMDLSc2kqtJKpOOkP+z6Pt/B9ayWxl1US
hDhuA7cP2bGyqjPyGOnbHPLFyic66EGe2gflURGTI+tQIwF79XecsW95Favto8/E
qXLRBKmlbixphEdGA0BjFRtUAcmgF+6+JNFEclZH+iZTlzhwjjHk/00jiXZ/kdss
NQXq1O/frI3DSExPXsKga+A4qGzWT5q0z+Rqsfko5IkGz4nizy1ruY3jqbuwA3jX
JmFwLK1zGRghQoTSQ5TAkBNNW5LC1jKUQtfvD4iJKf7gj4EJJqeoOTlBUmvlnigA
viMmIyxcVUTJ9ypGwkolwx4LLm6XlHvbJdzgHLY2wgAttnZnSGApZUuhH7fU0GoO
Lih8H9YBkdWCSK5A/pj+tvpjtU66tTQwnFpDyYiLCA8tcbAZ/ptjl0YacQJfPYhz
2CIEVG3pExMNQMF5AYPz5RFiJdVQvkvQCDM1EMB4Zf9P/RaH25/1+jGOERhrHSSk
+FYvEQQ83+XUnvZD1/y8Tt7pUFYV5c0zJf5ifWRpMoWqfWxKZYVgVuLeDvAjTDUI
RzrxnooZZRtLpOqJJwSXBtbEOmInGW2OaONDPC2fWDc416VZZmVTH3Z8ZhuDS1N2
VdRHI9yvgOTpCgm2dAyv56+C5FctG/Dg999j2/Ggi75IHTdt7UjJbzTdm87v/EVe
sntrYTT1z2YQhaY9zosawa55/3fTfBOkTL1ZVmJtXVGDTC/owjbdt3dl6eTJNfr3
oP/sBMqVO8eA67dvyQHjWsjnhuGpxanlEFdJN7vljy+owqkQTDA0svXNY1g4lfd3
xdbdAOQZeEIjrJ8zrKCJSNBJhjM1EU7wRKuJOqv0svc2awkKx8ppcWR8nj2X6m2f
II9GGutCQjEs0F4E+r8+I7OyKUlpf9lExKVzwPwRl/QDP4fqsioUJgterbV4EVht
F0lrEjeEcCrGxRcBuuZL6xSY3qCI1PgB6W1IShGMq8TrlRlv3XhSyG7sbITGQdlK
iKkb2p+HTKm7Zqve1GQR8tgx/wwW4+SEwAPv1a117E2tp/7FWNSV2FI5AuMN7kju
Q+2kDgrYPQmFBYIq2liDlV36XOp09wH6S5+Mtf+GJMyxPrXjkvAMoVy9Aw0VQlUU
Gs+nr7TKvdPCi8H0yRYe4Yy60guzPlKXhvXMAJsK2wtg1Z0u9GsSX8WJglfqr4IM
iDQZUXD1FXAmcWjbPGjEcyK+Z/LpF+unxkGzPzpz0DnNGIAeHQyEg17IZaD5Zjg+
lRC/Ux0eyh02mKthbwGHSnfhkQQKOszaSfv42unP9of0ASi5aCaI221ry0B9+49Z
xrRddUoz86ML8LnIyOmZJNL6KFQP2kQHNnhIj3iiyUXAcQioxBr0GJUL23+veERb
ytxTxBvy0LB2WijQnj18vv9+8+j4YWwKeCbkzIRVQ2Nyj3InSNTGfrapTInZaoYr
rV8MLTWPr70rP10KGN9SqZ6iwWF1nrYtUBXnD14aB3/4Ae8Jp088JCJ1ocfShgc+
4E5fvLnixeUyhvHiViUu03pzWrAIujh6mVEGp77fSX7L10ycxlfVMNZcQdVZfLAU
RFORqj949Dh+GzyhKOaMYYGqN4VEBXCItAbyM/u/KBc9i0lxwN3j/RHkAkHTyLa+
gvImMUVEwX5YbGJ3TNNYcdxZl31Z+TjuoBN73UMCGS5QqfK4oIB+HMKwK2LLlbFp
Rt5fn8y1EIJvw3fKTcLzPWzWEdEguFLiqHCuA6C1mV+fH9udNTmLRCJlsCBv0Bbb
rzgjihrT5B0QAqfZRAUcctMBjmVMloMiSTPVNQPKIMEiTVXc0L+6v+QDJwU9m8UR
VXBwwIoPNUM/2tCkLKYU1vF/7DZvk4tSq4LR+D+j0Jl20lSoQ5W+DrKh/Ty8MB9w
joTWef0G2KWACwUHW3gqnwyzATkXv2FZviKyYKqMpi3d0V8miLfZpN4cpH6BK8RX
RuOkNK9nHQO7GtsQV0ZsBwbi43bbV4MfxRAZzstEgBfJ1u+lJz7JtVst6RBWvDeW
aD2Dqm8ptUWlZ5WOnmK0bgSgXM5pNWFBb+RE47PtjK8PwU12vXI3efTdvTcF8ZmU
spg4AulRrwHwwIy4rrvmfuIRAtxKBejqeg/qiyuCdFrbM/yx1jhgzNq2ut2ml4ig
qY6Wkne/1JyN0B8+ER8AC5s+5c1s7KwDRhQvlo4dp0EILkQTShuAAFin+z3Y/nv2
iJQsQ8zQEhG+rHvh7IaaNueMSl8LsBZKdYgJNhx6QDhZU10Q8RgjG9r7EpGXaYhu
pADSyYe4JdgX2YG8l6T3SO96dqCdUBl290im67IsDLmC39QT6yXr8CRmoxLPMixZ
6a7941xTPxQYUjJf8UNlbeSXekZvfbsDPNb2Lbwd/V7FFESaxWja2pQZ2wDlKO6e
8yc5RPi3D4s3Zrl3hUWIS41mntd7gwOkZRempaxh0kmXc/cSEbx5fvcp91CUFLM9
jwwTUesRoR//+nf1cs1gOImSgUvoDeoFA+FknOxw/Ejz7h/FMF6bCFdxl1vlIt1a
t5ndA9K9s3cd2k4/mggHM9SQuU6wEVItm54jTUrubK277YBhxDil3UmLPHQKGfcD
xEvA0OHEHBRcyznWT5n6WBa5EVrtnXR0pVMZN5e+I+NY8gsP+reXXoWclD2VTWA1
pj8RE/nkT2RplgdqNyU8wyA9RvfVp1HdtET15JJPr/t13KrWSF0YEjoSsOLRAuZ1
WzVAdFxg9jZ221QOWEE4eosom4MB5/PnYPoF/jL5EgMFf15vjDRk6A8usbXOmwVL
GHZNInsy2YafaUAinhOLh9dkPqKEYyltKvmPzB55er2BmYe0NyI0HpX1NycS/fxN
BkXqdCbQUJMUiLVgP30P0P0h0W+wdFmwl+gjRdWXVtYlk93VC7MDkx/N5nYZ5KMB
+0cYp5wb0xhISrqotydfoB2/1BsGmMBRwRmx6yJdtKMpF17e7owZAxupz1xPAjKh
KdN8gf9wv4abW4qul2gm71LJrpqJYfcB2tW8IbxEcoZuWy88ABf4CNFT91p8plvD
di7bNET/nHeH8jWFZlkEcJNNrHUSy9i9+LPtiE109BUSn6JMFZhANXXptZxSUbym
otiYgUv45QZYs05aaYLOjqZyY4OYRY8G85KdzlSmRaCTtjcbO1QLBoQgfUtZmIuh
ParyNip88f2hzZOVaaEn1ev047C35yzinzA/TQgGhyCZXbd1w5WCoQFvbYHZKzyK
aTDeE5wEvP5OZ9YBUhdnkppbNkqIFINUgo2G+rIpedeuqEf6z9I3nw0DKtcPHI/k
SIPUeq035/BsAIgKMgN64lue1dyWfS54HKTP4f4hmJyjfgLrQz6id4XsxZCRFyyD
w4dBlWYxwWc/v4W/vW2nAkslohvVfw+sUcpWYCurbRtq/ADAbKnTAb+LUtzjHumG
Xib9VlKSO8lWNA1OZ/BsZdtKJB/dHPhCfh/i3ymDV6UC/aKU5/cg944DbQ44bwnu
hs9KS2O6VHOlBdoCafwqkEmayNWgVaku/s5MePnTVftD4TDtArMmDFD1jK07mtBb
wqnpo0G37vN0KUCnc1FVrmEM6wQwJPBM4PzIOp9fauufTtUIt4oTUSkwZVZksAAS
E9dANMqok3MaV/Y0GBDSPJTYk7mQpHJlTljJ/zdaHHPctSn7U3yXOENCPBLmomF6
Ndz/xDL+zvnhMZQuncoGsT/EWLlGKf9Xs7vGWhndv8niDtsqIl8O69LpKHcfHFyv
cj05fk6Qph38P8wh42Uh66AiZOFOeN0YmLvNYfUjzGSwfcHdm88MF/1W86uRe7oL
JEyW5j7JZHT49OJKuxn80AcMjOpDk1gH1lMV+/bTbn77ws6ndG5RKN3ETy5bkQJb
mHd6ZCi/oQj7/h/s3qdgYlAv13g9Xa/g42Cq4Xv4MiPkmL5fGpsCT+ICyp/PrnXt
SygarqalMDKqv0DjEnNF4U/i2NzGKNpkaehWsvFRWrLW4GGW8lWi7iTmQHvSKJ3Q
Zom3FKW7LgliH508KcjNKi88anB4F/HSRfgFjpewmoiVB8e+HD6kR4E6Xw+pea8A
cvnuL/C5kT8miiLr2WesoPn5m48r7z5fOWJfnaSrsHOpg1ydW8MQxtmvZuDrW9Et
JWVieCPvtOqXWjx5hI3yzh0C8aZQd7jMUif9wv4yDF1lD74lC4js4r9kfdfxxObD
Y9g+VSgvoYt2jq/N2loc0keEX8yUCYPr0KGrr1Q0pmV15myhcqN3A7g3PUbEedFp
arVGxPvxzbY9Oua0YBsyF44a5xEJsCfRczzJhiKuuiXFhDbwYPd/NJLkuUF7hEts
Zz2KVxwjNOWbdnIReGt1Qxn5BLTRRIs0RRO+9Jybs6ud9zEtMMjKcMz/I+sNXYIk
QUgbscBrtDqVig6Z9AbVk17IwX20iaSnrDC74U/ri/NAT9T9lsA++fDxI1DHIPiz
dvJBvK0G8YgHNLxOGG7DKWtcgEk53j1ZHWQab5DEEzDyk+t/FAuAtp96nDLerjjw
MJ7In4zqeYjamMAdEqUY7zIpg1ZRJprBC80DZleP+KXZ+eLfziez0JzTLWXHSzUm
3fv4qrS4U+DLMLCtQvKSH8OZNlfeIP6riH7NVJ5MRLlFPylmoIbWWUz9DA8rquG5
v8aIkfqu3PEZyR62JkjgzJNMSmPwuHiwiOOYNzK4aHZgzHT+0aDbfNZeOWOkfrOT
Pd8XWUxswS/msB1UCvfEfIc9qFNREuM+q1p/a6tXMTO75i5oZVrxLV/HC9/JwmO+
1Px5N06pw0xmPmMkaVCZx2KNWEgm/M0YjkZhPcKYNjtYOE5JbaLX2UittOrykfyL
EiOLrQw34WEGJ+UOKtPB04VmpN1TnHkpw2JGvpSdRuj6XpuPwmD0yL3UjtsDaoPG
fXdXkh2nvxL4BdXYfLloXpeU5KqciN7bopjoXndSog2+iwqX9SPMm5qFZIJAmT70
8Wv7Gj70AQd23cLaBge4e3zjVeSxyZVT7Ku1aarptCMyRLzeKXf3aMbbtT7AXmIX
YRIgaX2j8Px6ehGRiBViMd6DDj5hKM/AFMxPCdDl9alkRfbA/7hNqA8LfrwrCGiO
+dlXgcDolukrvE2ZLr8DxlG98J34vULEhRIBsGLcLTQ070yfzVpM36ZOXahYWs4m
/PsRqgpScr71YBjXNB/NZzLPZxCb9JsVPth6rFOnFhG6Rip7obC4RCQGbSd5PVda
fmfEAO+S07nFnDloTMunUTQtapW82POgI1R3cj7wSXFdTnimXOZSZ0/HQQ0FD0Jc
q6mLW2tZl8bWDnp3EqITeNoYpvn2mSUUh5YBFrBWoCrZmGvBTNl5phzvsUhC1xXX
G6dLZNL1EJTONJ2+QEWDKa9+zCpoJIKgf2bHJNpw40sZHrbu/hR2DQBey0d6BOvB
4W1ortyYlpKCEIPsyAzzh2e2t9cG/9q3/41iRfPHBym1GEqVUcqBIkAb5qoQ6nFa
ZSCkLWnfPCp/x9IzWlONapPb6XoLdnvMoJCHWudk3uogCSSjyWB+F/wiHdaVNfTY
QxB6GmlYN9CxzSVYKWlGUTGUnZPobM3Lg6rB9Vhda5odiyRBc9UZ6c2oyGCroc3S
EFwaexaIJbcrOkWxt2wKEzp3r/vsYkulu4HjdmmhYsX5vygOph2Yn52TifxHSOcz
MGHq3D8IZYJsvfgNdCmIEKhVLkb3CEq+hGMrCsg4SMbxUKVDP83+VeN45Mo1xmOJ
HZHItjBSx6KU+6RCKmE3yhBew+0W9nrlDpYWnGdwoRaB5QQAclyoF7qxz1DJZt22
xpC5rm922FBh/qsJk1PLRUJQrITMCQPVrYGpTuI2BMBoVheWoOLntxVsqp9tc5FD
/hMF2Vd/jQMBF+BjgtSyzTDS4Ie/vs2sbnxvbFBkWd1fY01O074kUBWBHQ2+dkgw
3XVAWTbY4lz9blVPZuAQkLd80y1BF4SG2oDfEgBxmBKs2AJzsllfMveJt9bOoIz2
/eRiybD+pvfKPak0m0UIobwNc80sDyOm/DaB+G+cR51YP3asUse6jjXcHAPx6e7p
3vbzz/Hy8uInsfspdTMy0fzOFQ9MzMtj2RNu6L96B63Jh3rQ+4jr9Xxk8SA4KtLj
8f1G4+lJJkkUFrQsHEa8d0PNQQ1dVg8dmkpV8fofTGuNZ4ZIhNoV79diMwtUfx2u
BkMqiZ1r4vroHTb7Kfr9QzJo3ekctR/jr2YufENbghRxAn3tdOHe3gzrS6dwrFVi
S/18pJqiDsSs2u8jD63TDw1/BVJHmULuGOzLeBfqJkeWIyAsWAJxy6yet/bAksVd
swinKdkzR13re7PjD5waEHSZLqr4f1tebpHBx9U6tj5ebV3rYAhcJ135OjCIvrwW
OqTnNne/jUWwshzzeiek7lDS5LOYO0RCRG5CZOtdrBTwUWSRPXUSAb3Y48WIW5qu
dNAMYiK9jvAXwI14tS8/EyuzDtI8ZHK3QNrvI+f/75wtcy16+Kubbnw7KwKQyi5L
Zq4cqVp1AvhO4V5ulSGpqcXG5yvfWaSeqAS8EG0M+i2ZJzeujBPifxxdhHtEd05n
pVWtea2utEmQEQ63rdMMg5rQoMoa6akoDlhk1OA0MrZXhGoO1zFbTiMgdNrfCuNm
gPqnRXZNFsIcyPV8mYhw6e+yi2vrinBzzWMlIQIO4iz/zi6+4gMC2BkbSgFr+C8C
6TWTN64WI9+YDRwDUgss9hqSdZGdtzYsHVQNqDv82QsbOB6Ls68rAgxU1u1nd+YJ
6xpBakJHwCLnqYPN2Z11j54K1WDyYy1CNbJ0L/TcHxQICHWTG0+xIWOZcf26DY8m
11QpvX5i8NnXWk0vV7G1JR5MvKRIvoQBuBeZWxSjZcKMIqr8sqhiEDP+Vs3fiEuO
ScKl34b5BGF4XbsruVYIVQDpXX4OSVQmHdlpDhjHWQTE3uRm7kfhGW22C2LdixeS
GEOAMaTsn9jlsuBiN08EniB6PoaFyfa6CPFSTPFfZ/C7RMOwhIyqsIIA4Otk6REh
u3BJvkLT2c8M+AecSbBKK7qfAwX+PG3wsIgJN94NQbPjPNJsYVOr8Kay5eoHtzjJ
sHvek72WSM62u4idxE+jxp4x4dz1mJqbLlyrg4hbFrKQAmpFslyXU03iWYiw7cHF
3zAYRdSW9CPxh4IXexcx98HSeuZvm11+hG/kLivIerHhYwEnTlRyIpaOx7t93sLt
bohbC39KrFPszMiHUVuLiwvV3yBNll/AB7QHp0SW4MEbzkFYEu/UV/Mt5S7E9VP9
9WhyyKL5DKZ5e2w95sGXfYcUqNvqeOZzSRpp/ugF0bNd4tqjLsoAATrpdr/fTyn5
C6dC+19G4oPqg0/2gwHseiXduzhOBqhBT6kdXGTNP42M0Rtug59atWeama+zRYfX
UHfNaQC+YbC2JE4oc+gQcPZdMfbLFcm7RylEcJrwCQnz22N4let7kdIyz/3+8Qt7
JB2LHa+9xf2EPFQSOdd7AdIaQX/pZIl0VTf0Gy87o/bd5cTQKnD2CitvTPGa2U8U
7DKV39FWC/RvF7N+e/7JoiNWEjXqrMapkEfJ4LSD9ailDnB8elp8Owa4gtX2RIY6
s6m5dtqB4XfA5SgwCYKHUCBstsPlxChoYSHWP7qFXCcbGdh3gbEOcQ52iyKaArs1
zDw9b8phfl5su8xS3e1bXXtd4lowShD1fmvT+oUWg+FSKBZ7HZxN9VNjjt3bOAW+
n5DAMvGfFad6nsSfyAHGlIrFAuqDiTFSY4+oVkro5wZEjnuaKo7+9Q6F7VORtRtF
3jXmp8C49IH3cIit6kvqeMnKVh4dFA+evnVFltvUbedUV0lDwUX2MWbWVjw0wrbH
3Z4CyWIET1MPOIoRrPz3qElPhu/TSWdc06gUBRXRYcIZwvgqXwQbfqbd6ZCoF2sq
Ed144Lc7cTpxYJaYxtq8ehxI3E/43Aq/1+9oetAf3B7zGvVNX/ExCxpfTDU2qosn
HhQ5HPKa0Q4e4dCt5jS4jQnuzypoKS5DDk0RgHCjE06ccOzeZe0StOx569+yv/sv
9hNSyIi0h6DU6VHlcRylCR/T1fGIE7/vlDGkmN9A9F+yWTva4Z+wMhkrn7DgVCKN
Lhcc91iIxPz+Z/VF1ZjTitLSRVaMoKM0ty6Lh7EtI9lYlsKhmeZNa6tn30F/FgiV
M9/epOVycinoQhZfHdQvoKTJq/WO/bh784sJj7WeztP69TBAbmgmIewtPxrWNpe2
SqFE5DH1PQMi8bqduBa2KI9Ph5cw2H/71GKkYIOsXJeXsYDinVSq3+HGi4Et7KkY
o/NeRmcxY/zz5FOCqGLVpIikbOge20vRaLYP465/JcuG8OYmz2UrG4sTl1cUz3pv
SATLvXuTkuLO4s6qx12KWLUXUeLUPcJOw3RzIl3IsCrBoYSCC5Xew7NiQst3gim1
vOLHl5F+jmfmKNhXq2e3o+wGqlcEx0fTU7u5FwY4+MeRbrfmp0H2s46220jJCACe
EzdAejL9j70yOSrwVN86a88hGrgpEhxEerSyscU4rkHzipbCApHs9+rE9/iDskHJ
dc5e3ZrndYqQtlZmBHxxNqPOyLUQPNZP/n38zA/LQWoMVzFUBBCJenmbNNpQ1Uit
Zpk5ZrxfOSdW9SsZgSDmkmua09Ps80H6zm3KJJLjghhDYN2r+Br67RTbtkbqz1YV
y/PbB7P3tZg0lvK38MFMYFveEOn4MCis3/3lIQny+3Ywc+3PXP1W26UJ8YZTEQxo
VLIyve8pV6ORMybonriLngqm8cvC+ij7RZLCP8h+vjOqGb6c/qS5+C5JQ0JuOTT/
MGHUWhjmy8boEKRj/4D1ReT3sXPiUqtlmsmwWKJGEeryA+/zmYCYg5pw/r7NpAVv
tGdxTQGfyvWFBlxGur/5xCpPJ5FXLKu487m7XGo+PdXk6EoqNQpWlusLmzG77gec
hU5KVEuGGnr7qppsCBI/3hS3cPfRYjpYiXkTVCtHQTYGtMI475eUljrA7x+F99op
6uwL8DYyiI3odccHC1FBRjcUspbMNB2ebLwMZl/Qx0mP1kT/ZySj35a0gE2vA0RN
nn6/d5DvVSxOWhrBwmGgtywEtnXkeh5rcXTHMOEefVBd8IYOrc3IdNBx13xMYpPH
uhAZuJMVovCheI8sCFjhUhMl9zEiK9qGJB1ex4CPPj0p/gtAcBgzldpH1O1Xa8kB
H0PvmT1aawVRnEht2bbjOvQwer3AyHZxSTZIPYiQKjbyVZq9Zcf7dTEa6/4QreOp
jGd9hHrfPy+QcH4++6MAjYh7s77HYYVpsI0oZpriVf9SMg1Ck+2/iDPqGEaR35Dv
E/B56LKqVuJVf6s2s1vRCScP6Xx0aMjJEtuqCWtceSePQtNbbH1al7qU2dsNq2z+
j3swz6ySlafWFtLzC/lq23Wu3bZIJH9FcaK2KDe/Ndt87BpqSWzcrI2UIuFqeTfK
KfalnHwPRM0yuR+DQxm4KrtzzFoWGvU7hGnKWNzBib73y0NeWqK6KmArdfPD9ksQ
ozWZYDZRMGZNvHkAgF//Q4yVRt8PAdLJU+FtupkCqAj0m+OdBui2B1yg90IHCynd
2+Hl2/3M6TM5CnwPoAwj4y7BGn69AeBiJOaq/MNjDj6geaLxd39+2pYIbcQcnbaI
9wtWxfEn+l/qjUypCB3APaY1pllyhmSqFYVJB6bJBYsEpXEfRntPKSsoyp75jACh
DQTnH/ayAC5s9u4HWU2u4iG1qYrMfXPm9X58cza8y5+la1jdNn8hF+e8WYKoGhTs
jeAeYM73kFkuxF4Y0Kq7WdrR2s6a4WJae1MYqE2vf9+FNAfJJbt0dPMLgAhwn9Az
vpzj6lN8rdcHDnPMV8T04BdR/d56GeE2sWroiwHj4U+FKC2urGX86om4XpCYkrbx
O3D7/t+25B87UfuYXKaIqfpfHsuSSOSHl5jZpFqDPylASkJD1L3Pgl/cyU2eJBP4
EKp2ap2nryVq/C4i2oOFaE0ZmgMhvSCBGMmbaV6NUEP4HHvNjFwg1bcstCiHPkID
0duv3ixN0DT052WVCfs9iQJu7osBmb6dQ2n7qInMulngxMzGrFzumxSMMIuFlnO6
0DAcl+2B4geavqbVcik4XCPKNeuo8rWvISytYfELklJWXqQOZc6lHRHzYHVctSpD
AF8xKu3iG7Ai7DuxGNTm69DgLqcDhlcCIsr/8kFGmYpoa8kV02PsVvnfxgliiZ45
NGViBX2BgkDnXiP+1gdV9v+3Yz4S9iFirDrk4z9bFaYBfEdBDs5MIhKTIn88KS81
oXqIgqnhy/Qc0Ld9Vt5yTHcNlqRgDsCgfLeN7Ku4yxBX8Nk0UUZ0Z4AphuvGLDkk
d1ikiOvZCCJY4vCDyvLr88mgFr7dMGPOAUtG2AJzka5R6xs6BK5sX8UwiPOZMfdA
tzQ05wwveVP8NK1mt2U6o+5q8rh9QnKrldtSmt+VGBDpbrNgONWtPWmjPWkfR6NI
HUROcwoqzyT6p4Ezq/WtJNaNHz4vFFFYP1wJVh6WGkZMP+gnZphqk2KcEyWMrQ81
eb9qLx1d+ccdyEPjf6T4oKFJ8C5XPWLyy6IF9wxT9H5sqghr3uGLTxyETsBaQO0m
O6J3rjLpOx87hQOiSleb/XgfZHRrVOujSOjmE2w8WaXmZ1zsDUq2yPLl1yDXAo0B
nJG0OUCww9SvI5A5MnR1oMV4GFWdz3pmkIsmZGITvsiiUpdadYyQDkMSx65V1fOF
l4EGCfZEqgOPWu8niMbG/I/FIM7UKx6NhSfwYrmwqFi53I6qwl7/bDMJVmS+VBCH
eJnPl8HqIb/zJOuX46YkUim/IRT9OqgMQk7xlVBT2TMe5bnAI2uRZmX8UdDKc3ny
CcydW/vQ8S8Uelttz0DqbNigtZDu7DAeYZg6+artz3PXkFCnz70yb7FBF98vlSKA
+J0e/PiuzrzcXrouIZ6lcFYXV2s5peFsumMVUx0zcd58wIJdplEm+c3Xe6Ytj0KA
Yd0guL6rn807vuFKbyYHHxY84dM8V7vF+lfeMVvELITmOs0C9zxUC90Hgqj7j+kt
ZzSSyVPmQl0oz2+MROuwUnkjtT/S9uWcQFmfVSpf1IBbQ46uaQYOXYbBMSRr5nv0
8hhjJQsEdUYkX2Ds8gIyty+Sl1sjuDXhvrXFqzobXOr9b94KuGD/QSlf5eeXJpM9
eIwKPsgCeE6AEIprme1fGogu+nML88TeBAe7n2kA+uJZ+k2umT90FkdvCDi2rMkh
pn0nYZlWrEidpkO2u+1JtSfFhP23RUVTnVOGRegm4eDFTv4MI+YjvzVnkqgOKS16
vQtf0CUml8BteL3XfnYczgGnxQDAP0Vwk0DJbFi4jbxt7zQFQd10PrnVeioVo+7W
QqzD6ire7jyKaEFt6oD7wtIl98+Hn4ZNpZgo3IdOCcL5/sgCudmxhIZvyNxtbHI3
jwRGEU7QMrC53/VijQlFHDbxrOJmc1Q0eBhqLWCIPS/ZunK1WtoDaddqyOfWN/zr
hBkIgzgJE8ORBdvE2s7IZuKtWRIIsU6GJElMHHJYCLnjwIasUfE08Rcr9lbaXLIY
qRIz/RuI7MpX6lLSb9nfIraKQbrdVmfDMfw55R9udMWZQapMyA1ztyXOwOgQslwS
sILrXRfLy0bI5ICIEkQrdljZQNunkbi/ssSm5jxoKR0ky/P5xmaurhd9Be/FXkly
233BIBJL/HU9yaBkTNnBXeGgUEHnN0XPGC1zGtypLpmzGilHrUw+3jjJGmtBNFOm
388Om5YvEry3m9W5y3syeCozEjf/PGBA+W3kBfOqNC2/D7iuOxDnp2Rf1Nwvd4nH
h1vzw8rmAfDnPEmdKr94nSm7Ql1MsIytRC5wWZ2F/FXRDEDeOIPUShTRr84moydW
T5mxzThhL0pXFdMydvrFoNEZaECQPgAw7OiH/4aSAH4yhn1kijcMI8miXK2R7Ih5
SIcxGeTyWIjnkwRar4JsBd0ij1GpjJlJu3H8l3T0CdUFdF7/3HTtPQm/dvmMi1GT
+vwBd3/RM9lAwWTvBA5sf9P6YX32j1IPVm3OU7AdqDTya0GvfFac64046Z3/qZAz
dboKXGwZ5bGA+7wV1h4pvcotg9bEK6Etc6R1Dsxj8t9qWzlHoBh9UeQGIk0cE31T
rr3wkN2HBitb+3BjD0srU8qNvCH/YlS19CgGEXbrbV0mdEZKkOlVC/6wrOD1d72V
MypFstRlRtCWUxQZEhaZgt58CYsFNVIZgbsXaOSqRkPdXd9RsobYoCKiN13h2RyK
wmuJS2CK4irVjdkw/vdpuVOchE407D5eOCpNYdLEIevGWGviPSy0fHkmeyX+/of1
Y6mfqFUgXg1fsniy/94Cj54d+Ez6iV+mxmZsa5HwT3WYMZLnH6EI6g4IDU/n7hup
H/kC7IC9LeAY1OULP2tEn9LS+pkyQr+dftdi/pXtmvgAyCWOA0l6eA/ootxZ7SNu
wH40eqHbPkGkOIlaqJFOt2gsUy5zC2Lc6pGYPfrBinZlsXFZQl0dyzf7MYyp1gVn
QvKVk+5p/47JKmMY9MY0tsJKYo46kvCoHkhegH0AOGJHltdCoRygwaUfGay7fxaP
RWVUve3x4QYY8QhpBJ6OrRUzhz4imK590oKdxXvRngpHfCjz8hG5j9c/8IWsN/MW
EEW5/4voZZsU1IQ2SOV8E9QQmXsnyZ2NqxGz8I/T9Uxvriwgtmf8Rk+ZfZEcOCmP
KmQhXZvkeEfn4bvwPAztg0mio+jv52u+AaJFX/wsgbhy0rSCBQo9GJVp2qDT2I3M
i2RKq/VJI8XZfA/Ld84h5/7V/6gNhMRV309pJ6EnSW35VCGT21LiaWjrXb/G/2AG
bTqRK9IwOaL0FY8Vme6dclMvAePa9b3sUGaNhNcbB5NSeuMIH1Lgot+LgznN145F
L+DnQHY9iyNHtFfDIu4GXFInU4gDuugylIouY1A6pdsqEevruEfcSwwEd03RIqFY
TFNKKVpIg11Lh7oLUlAJQEPSdi10499eKVoWyfGp0gg7fDUDwMwBXk/OHzlVjiZ5
SdAgx5/GufnyeNl/8K2DEmFZKsCO3A/4cJ5+v5+d1TWux0/bhZFEleLc35SF3MpS
pnFjyFIs+I3SvbBoNcmZSTiakdhOyWA3NmdyVoGoMSXpVk3SJBN8irZ5egeF/jrC
Ww6XsQDCv2JM4iCAm1M5kOSou7gG8Yc5DaPFsTLXEH92hWxXIVYHIfoKM294lTsY
656Guqm+KZLOLJGyZNKwaXXIvXCDpDh6hrwoYa5L7nJX5p19estnUlFfCtxc5HWZ
9RJE+Kzw/8owjcFthmr2ySUKkeIzRq5TjTEd+EGONDW5KwCfpxPxCWQXrcoo0+8b
MQ3H3XChVt2gOtLTSPQn2/2HVJwgkHXGqeTFpoKVVYJvRsVF23lijvjDRkO3NKhM
i6kPfRdCpWtLCi4NEO2I0hnsqdRy2AgnEaNTZA4zaDnBL6XD7CjcqhM0mMqTRNvI
GkJDx8H1gZreMXoS8i4Q1GlDlF4P0tHAvG1k+EAOVUcBfgrUMDXMojmDHEFpNxlK
r8O01lik1DXlEyonvvvH4Qshjw2yJe7Y8anlXq3fezB46Qx1RP+fB9KHeVqkvzjJ
OdJMrU/gWO2bNurCree0yZRe1SJhNeU8oag8JBu5n30o+djZe2ptwgbm+9fXMHyy
qxEH3Esqk/CthxRs4PcMkx8T77UQU06y++L4wxE7dR42fVT9pbDBSSyYfqo08oiw
yegdmxOYK/oUUe3rLGXcfz8S3ZC6lSPIcVLs6+MM2M0VuVKGpUpy9o0QKQx1aJLz
JNlCL9I3M8Rwas3yUYsojpvz4l6CXDT2+n2zb6BQfoH219iChljXy+SgVQd9Ay5/
firkxNdVImgtLGL7aZjjRFusZrJer1SErMB5A115qAzeSLEhlgX7+PhdZFrnozQu
lyhXB3UtnCyhvdKr3Cl7HlVS6SzFWO4xjmWFZEpB2vZHVAVig5EDcZxajTnB4XAY
7z7p8H7DDs5c3TRpSTwI8d8lZJF8Bira/2JRJeHrJO4TU9e9iBTkfSxvIT7bDKlC
BjbwQwdpcI7eH3R2P96N1M/vY474XDq1PNII37zaKgysS3d4H/PfVjxZR3mFrfRD
eISNMs8odwDlAQnojPtBqFuIEZPYXWEFCVilKyAAsoWyIYHezct93y1Dvdraplz9
kpXshy+CvhPl5gVrKebQZ46OfQ3BGfnhkjWAVOnkiXNVtygYzJtBxfxYjaL3Jdc/
r5LbAGgY+5rZnHOyCfxp0gpf/GmAUZx6Tq1nF4S02o7j9e70hs5/RBhOJRz5x44f
yjvDFtzJWOgO8xjbUtjOFFhNhDoGy8tkoxOLMAvo6SDzxS1LYmeCpe3YKVGCxxEf
LmZuyWJrNtRRu39BEm6uONKVHlOPaAsrTtFgtXkXOfHzQzh71a2L8tnm5vGgoL1W
v5tAIctPHsiqf4tPzMpWTI4T1A5hhWduxR6QaxmdJ/0kpfCr20qV/OUafR1rKubh
vxPq0VS8oGmgKmJF092jHH6QkvvP2DhzVzNKgc3e8TkU1tIeiT/XIbbqLpmsyGX1
3eRvIg822kw1MxlbmS8FscsV24vczZFSqCAh8uNs7BS6bGZJTUHh87CEeqDSuAv8
VIHMVRUJMbh3xP5hSOIjYxlOo50ABwLUWWA2PxmBvvOSL/7fd8pSj8GdfDioS8f5
HVGA+EzO9F0J6ALwTDCOiutbG63zuFZtaW5LUjv20nquw7E6r3LIbNguag2B0llH
0GybYFCI9SAXahK8PY0cFwsk5EaD/ZapWay5109qeqtgZqEmMvZ11zAIROvPWATB
2rlqxBA9pWPQ/fLtpwwlJEAOH+zFV89+v7DBs/PkyUQHgM4eyesHmQaYpWPJigPA
TQwtkHZsvIYlgSVSeMyTaVAVtuiBO1AScUWljlT6YCEWdhluGMjBhMj+ZEjL/rlh
pAMPMKkm74C4AFMmivU0voYDbNSS5Ifp0nzYFiCr0glbItkqyL7Pcqi/tPc9PIbB
+VWIe215Xx06iQ77xhreFeAKhnY/rmkJVRLLatSVcPI2Z/L/2BRZYBCol42J+DbC
unKz7+2me2QqPo3ulAcNgxeYL83mHE/QjNt/g3FFxUWSOefgBPoEBBVCnq1Efjdg
bBcWQhMhK2M/n1Rz6nHLE7ztDqm33E8LOtjfAkDmoCCQ42wvcfogRThyuwrsbf+t
ehY/0a6c0PLige87faoyS+lajzsA8XNfDzs0yZrcdyeI/8VbK/PpCQc0Po3/j4AD
Fk2o5PdjOmjezNiklNVQXhhiSZTDbr7qEkxbkm/337P9KhIUTtqPugn+QUqhqPay
18xpXTvpyE9iPr/e9roj4GcCv4t3IghEqB18utmnFq8XSGsMhkFhYWH4eUAH4/Vq
pRjlZf9RbZMFSDtg205bEvY01ibcqGRe0khRN1pquOhNprJbGrEbDU4LovVMnEwm
t+9o9pjizQ4U2ecUqZ5BHE00hwz57mrVHOyrZuJfHZVk405ZthH3G2EFlzqOKy6N
57kLdBolF3woZJivovRaEUMM4JpeAV3yxmVmP8QG26ulDwSCo7AXz6FBrVC90tUF
MUEQzOKe/y3KQghy5s6mr7JHBRPTbs6BPf/KO2ZgaWx88U6unIRFK0mp1M4ZV+4U
YpBG9iwUG+LhM72IdGNs8RGfIO1hMiESSnMJ+D0aRKW+gimu2GtSsSO98VVmh/Zy
LQTg39DOhSIMJr6doKdVbYVSdTyi9WCWg/otIHpbS3QQPEchEc62oR0gKz8HMeBN
ysNZyLh28RRKB0SCNC/ilw5fJZ2B4exdyDk4VKcG7AqVJ8SNYyAuw1MrftfIBFjz
rgv+SHETJi98oKLayxLOsG2vyKZ+eu8QgBnP+0wbBmTxseq+xdELQ1t39aes1Vby
r9SrgEXc8ZNVHjGDyukjy+1cEqFTqVsiiY9PGj3uVi4YeZJPPJDu5+yISss7cLOB
mFtTvk6u8jyTHTKkWYO0oZKI5Lr1sTO1IXXb+HHZG2xA/VYHPqdbyRBVTnGwKgWD
nM/WEZTF9t6KfTybjcX+hycXOsK/Y+wc2QEl4/zere4W4FgD0lWLw7WS9rq/px1u
W24+gBQHGnwaCV2rnY4qmY9G976w1CU70+Fyrchb7YWQp/OPR44lwO2Kdhi82Ku7
39jpYbIbhd9q3PBIN4j9+GdDexZkGKGWPFN0pZJuPV3NvqXFPLuB15SbgbO22ZXb
/JQpoifyqMOI4+4ha6mTlur6yRsxhn2VtSixnmKiLtFVE4h583WAVyDVVDPiYhOU
d+1/U/zCFx4n59pH0SbPEw0RxXy0zekrc0ihVd/oaM/PvZx8re8vrvR9D6fkjtzZ
A9b+/Brs1WeCMT+kzlx0XhOSRxg3m1LEvvFao7Bx0Duw5CR/dQaLLpLmx42pTTf8
iRNUo8H0Uc4eq7wL0w+9gPbV6Jh1v64dd0JicOlsbDEeMHCOwtyxDUhmi9Ok93iF
Cd2QTYK9amg5V03lJQg9LBV0hCTwzQrU+ENUo/nCFRJ3jIfnlUZIKJxR3DK+lVKZ
Rbmw1h4RBeNzPPVTTwquTj5GhvFJsYUGihj4cEyH+ZCM3SrxuTLT2R1+HxFpu9+Z
8qUUjO8cdG3fq5p/0MY2NhKRmSSKEluo+pHDoBds2bEY0dYc94Sk+Hs/F/M0e5Xf
Cd44VzwaJVviRf/NcxRQGrwYlFIqVfPE9tb2KAFfJvRpXFYLjaXbKgfiml0SvTXo
cungMa9QLLVm8q2YlIG4jWN+jOjnyQ0RQclL0rfRbV94V0TM41ggBjbAnRtH8IFN
9Yxl+g8E37zCdNWP1MUViI3DoVuCN0eajrJpJROgpk54+nZ8TPqBLNExTXg2WEvl
1coyMslMp3tFWH8NaK9dPjTjyY4CF1AxJsjY/9TPxSCeay5Va9zZCZryvxDK5C9N
C9cxxfOOsKr3IIrcymt5kvomix/Z3/scudbgUNjfGExRKf96TXxGjXACrrOMuObM
pUDy9YbPzEE5GTTYcoy1//bO16s0rRa9Hme4TV6IyesMzg1Ms5HWhwroJmQp2DgD
/JVEZcAqji5InbMnqKDGA1la+aUe83dB+qWcmED5jXt5g4T6g7s64cCqFuAh7e9N
cPq/57dhlH/OVr35tleblccA1Qa82TmU0tM23nk48IUjAKPadxPL6c/Hvc/OjKmP
8xJ/DtNYSdWPlpqBAVt8jg/sx5JwnNMwLhTIuEw5uuYKSof4u0A4ltwavl99mnTV
G5Qx4r/avjsNxFzJqO8obbWKvsswhPnAvq6H2UzxwuxggLpMF3QHEHw1tWHckwEq
3DFaLpOT5tNccNPgS7WpD8LWf5AcexQs4WPuxpzL3oz3PGCO7f/vJT4gBhvhRGWD
J5NGo+34hUrQ8otBMFQWXZXT9ndw2nOjpF3S/D2kYqg7He/DGbLJIDNZXcBDxoVS
BX2ERFyiv1asXSMvfglnRYmHHhlcNFekNH/Nbwcgth9ZfqmV+LFDY2e5X2qtYJT1
G3zPG4G5xwsYtK5ScVREpyhaeCYZV2xaR4quyQD1RLZtbem0m+sFvDI5dcAaC7CZ
RXv7MRhAJHxRCYmbf4A7U8Zc7NGRwsyQVUbdZuK9xxrvEvhdmzY13TZbwMwBNcih
3CAHWFBnbCEs1JJMopaFlybUlZWb5Mf4bfh3S4wpeGAMHKwstaORqojvm5V1S3xx
zXXWt/ANDoJoyuFyJaNujBdj9Joa0iv7iGEpVgU5fdtVo2LcljcTZEyBQszPZIdk
BfGsppqKnqnWizxVpdbEPoHFzcpENLErquAgZAIhIzbjcqDhINsZv3iqqRFkVyaF
MaMi+7M1xyl5+JqXEGkRwgCXjBGh0DYBegQZpPTmCCBzIrx/N8nAUpD4XJU1kIdH
E7qVUkLkA1fjQoVIc6Kw/7J+TCvAr4ekKWGebegdZhpriLurmZbF2MJCxS3XOkmX
d76OZp/3LQB/WHtJvV3PmrglIiK5b04bcS43FJpXdg1UFuLtiGpmszXCRQkFZljf
i3UM+D2Swc2128ayrOQ4OZ/CSxBJsRQ/9fNDJ/IwmNGujbP3iczBcxYTb1Eg75LK
Rer36qWtjYPLaULAEWtxt7t99lUTUsFIuT8eDNTZCMVDzyZOP/wEop2I6SFDF634
/BNCAU0vTb5K+87K0bLOGaPleKQ++/yiF6Ao/Ucvsq+qpfCp+TOKaXmbI/uuue2d
RsnkJorXWvzQsNicdY+qcuabmwpBn5n22dXKEgsf7U1CjLEWqafs9Qc/Ks25Lj+y
lhlnsPS8Bz0SILiULFS9Tm6Kvg5H9uR87bLeefgqD43rPBiZrtZH84BTcM6Uf1tV
4rqQBkHbkMwwOE4uryHEDlN50RBYCq8fT4RHpgnX9XrwM+C5suGqzpfhgnDljtDZ
III+hOGpgFW0F5Y4H2sYIUF0ZH4vuMv4Himk2R8t38IkAOtpndEReh/m00ekmMP1
MRkCC/E9qFeMJ3RHOLXUMKSTT4a3OffFdy4429A1KOsCJaVpKof2PXYZeYTSyy6J
8Ros4ODCCAQ2efvGwL2aQ6R2pHLnRV4rW8XHA5lrJARCjX0L9EuomRaVOn/DmJDm
JKgdPXfupwMhFCgy060dOq0o78p6BxZr2KVn0xUc8ZxThUNtnyXbxqQP/DrJTzkw
uJojdDtjErvr21YrRQld4LJkDHzIkLuE8oBuWX09PxOOYtqNejvnmAsG8HgQZLk0
CYeovp389Gt8UxC/PixFMYVelhDhJY3+d7caUpruP8G3EQI26i3OfVqeP6SAzFCb
20+fYcweyU0xwIV+Lwj7W7v5Vq1Va/hOF9z4y+0B2MiWfAwXxCwJB/BxFtOZHGHI
KTzT+V6YwbCBkCfQn0VpBkSBOEs+VCGC48DZkW0LxTRaRsZ/S/amK4v5izs2LO7e
GtLLu5y4H3dJDhd79s1WmgpVoI5z0usBQRjvWjzQko2zpiIj3Q1kcIMrJdWwZE26
aZ6tdAuEbvc9OhGaMV7pjqHx+le8FQ8mO9UkfIW+zvqxqhAE35uLhD3thhssFnXT
zxtiUmzdSWPnOslyvdy21ew4JkCeUMKCQxlMjEWKQkMbcZ8N4f2+Tbm+uwXWQMpk
2GhQBAmx4E1GNoJmXGTK81yG+QjRBC+QxbVzIryfjGVa/2aXpBRMNnrrsbUUG9JD
Ugd1neuN0QQax+tkv+yCGeXgzyctfRuIXL63y/A7iUxY1y9XusjR7rlF8YphCQn3
Y5mEoR63WwUdSO3GOOTX9CXd2iz5eW7hnr40zKC27zUWJuKMtT4vBH+qVpBPf/ob
kft1kugDrA1dUGqcoT9CIBB1XhNlWwrTURDaF9DbZr6BGnUSSVKCpLbOyPn6nuxm
RVs5zmsoMyGhIA7+uZ1b4stebG7oR+6Hbyw9Wb+rYhbQdbCJV6kPX0mL/7if2MeJ
5lqknTOc24N73WBknXJe5psn79RugYyZEunim2L6KoOzK7BmYJaS3orqDndelB9r
axfV5IP2wBQBUKekUriCNs2rhDj0T88DAH9o0MCUvKfruZu0rZZhw33XmfYhu9O0
jMqWEE7Lu585tquGYGMyrYZcyFX7qx649Vyix/LxJg2kqJAbL1K+SoOgZcvWpxoq
V00Z9oqp18LYHzbhFEo/mscUkiOHPavrruEKxzaaReJHv8MPO42LFJGVJoqU4Rck
dIFE0ORDuQuUoc+qgY7mNjcHF5FizE+Ea34tUFITXsI196987gWdpx+ciR3tI2k3
cTT7hsoD5VYN5jXIW3FghF1JzJvXthsGNj7ypLwT3ibrq6VswAuBnvKcikY/ySre
ShcgVV9BwFITmVWi5s1rPmM20zUaWxLqxImOUlnWpjmJRbFnQRm9/M+rBrLnUXFT
hhnupF25ozHUEdDcegiYc3AapDHvqMhTqIVy5ljg6y8xg/9u7KOX5/N4DchnxKtu
ss56uBjxDNW5nzCW7UwRUVV2AHnU+Ca9UuwUaoX9TTKrjqq7ek13NjHrcIAShro6
dAxim6mr0Wk4boVv4Xt4wd218lEeCgyxzZNniobpEfxHuBgY+jxsolKkypRxYgx7
ZjNVL5pmhkTxOLXAyycKNMQ/fJVld7jsyArCX5fnKzfrNePJyOCkwJJm9XX8DJyA
jA8b2WxaXp12ZlDq4B1XQEQbzr95ap2Pf2N/4aRhCSuf7GS9f35fYv2E17krlnWU
XDu7TnpFFXgeV730zs49zb39WrcMLfSZsmbrJZwtL1Y+D2N0qg6aYjzGw7TtImc5
+keJCDuMV+wYgjup5LH8z0rIP4tgf1sVxRoeYVOKTNz1eNUAUT5hkEhAKCK5TRUo
ouVyX+dTrentqCgRq/q3dEFVQEcp82rRWyZMgBbbq+fStZpyw5qxFV4zOe9EDOso
wvSzlAy0t+Ak35NUslqIkQpl6bnXSYc37SRtPybSB619l+ENbY4prclNjM588hKk
bkq5pt4OPuSX1RYb9GIrajE1Ov/PElKUlJd1oigFImRol/ZrHHHyL96VUbLWQA0x
thURhxeaEx1/q2WUX3NUnYPDl+MAn3BVdD9J2R5O1BYOTJZSNyNNbZkXqnliPLNt
X0yLhyHksYt5bYKXqgWA+HFMYM0RnBKC+1OsfXq1Gm9ySN+IMTXpczwHcsTUcyIE
hd/E+Sc+J6ZX8jdObldvnkyXZp6+Xqmr2qOMg9prbnQogvapWGV4ppOX5NdMokcY
m7p388BqBV1zOrkA3xVWri+6sZGpie+1na8tZZb4wT5stiRiCUX8qg4vcSBVw23Q
ynnT/dwU8vpmW2UpLagwmzWs6Ewf7J1/Ps1cQmcmc2thCJP57J30s8licy5qSZia
io+FCTsFMZsor8pINO7qhZw72DQAb9UuXS0x4OTKw6tsuFu8WCmZCVGtToV4VtdI
u91eDLS+1EX2dgQiXfK01Q36OPkRkWlhIrOgGEPzEk7JM9rESho84RpXxJn9K6Vi
MXPqO/WnvQ8B9Dmbjdp+MBF7i3THRlPsZkzooRzwzYw370IdQ3MewG33mtcBDlxz
U87iSi5xhN7zAai3YOMHUbXqDZrLl8vJRGI5XJ0GvzL1JbgBAPVYbSd5QReILCBN
21kA1uy3xY1Wt8uZ9VVjdzheC0+ywYKcMsr+9uwdYLd+ojZizw4zBhRJ2ZBET18i
3NaHn1spvbN6602uV7zze6cElwfrzYQO6QqOw0y14tMWIS0kR3FALZcQPNnc0RDF
usmE4ws3atYTFDfyG98Uqr0DLAUSVLFw3vVDGTleb9cIvaO6TIC4/6piNRhAfV1R
EQ/4EcCkn1jfLgaqBIZHGtZ7ZRJ6/9m6eKBmt6btak3xffwJ7v+xMxCDR96UXvZs
z5D2uVdAF/urAEttg3ePXwAf23ASDbNY/7fbyb3t9FxCO1H/EG7PtNjR3tfyxsi4
thE3CH0UAYRxcZE+Q6hR0foY495Q7F/qehRbk5lms1g1Lpx6uhVpLKbfw/Q4MUfK
X+IEvo3EPDEM226gPf1Zu8JOoMP5wsfaoKsy8hFa6Ih7ISDYBeHr29/rAUUA6p/d
UhfDsqGLSfn+YcezgDnMZsI7mYYDHCG6yLGOEYSjV1tsDSovxabwfTE/DL3IPbfI
Bjo9cz6bnsNdfC4BQ1SAuNdUmTBrKcMt87/rqfErhLGtIPdBD+8CgJrN0fmMfhp4
LtF8TARPoyWmR+cP7j4XBekaON/fS+UK27QG6PETyeIDc/bd4EwbOgCCmA2Rq8Uc
xiwdxDKUcrplNqWG+sQp/NBIfonhfv9JZzQdqcSc0gkgzYRgPZGfvWZjpR5qIpaX
z9nAtLwh2w7KgJw27PgasxYcv/nbmz7xeHATP43D/QJ6neclbV41VXJlvABO4brP
LPhr41O7a1qviP66+9Tpr59oMRw7uaFa+dbyjtEHeCExiysvls3Xc+KCWRabebJt
xSAZk3RfLvxx58ZYNauS67BV4ZOVM+LP2YnJMeRZJwfUd1/Y6ON3RAig0XsVAEu4
TaSiZ/J7GIUmh3uf9tzKOzp/qNdq9AL/dwckaqIMlZjTcBxSi58r95n2OnSYo+bu
O+EKe1fpBtuhDxq4x8ty0kH6U6sIX/gm5V9OcC8aVjBeHjobtO2FKzHLQyPAhdUe
VDsIzeCYGIkXyqe9o9Mj5dANKMVBn10LUmBxJNxtKnfX9KqPHnK5A0t0Q5kgkEg3
1T7O5aMI2fzHcU+RYn0puO5/8rrZ8mmKmjuWXRTagVB4eS7fmQ/VByfqsepXlqCr
wwEC3kQdk8Q7refI7gnc11C+uCUYlmFp8+9285fsTHNf5ceS8wX8aZolBN9hjImM
GrfPcRtwEwqRmKmlprD/jT+dgYmQfUhP8RpGl2V8sNQqdIzaXd1KHUA03/MwGbHd
qLqefcNehanGxb2ZOuhdzspGzABSqQ66ge57KLbz0ZVCMrvNRrvwVtfesRdEq/A9
ugXdTgsWgTsoViuBwQPqMK5VotixIDhV3wqmojBjMNyU3NeqtCiXOLfRqTkOxeyL
KIKr4IUcIVRE5XMrLDUEH5RgyfLObGe47YxwsVXURbAuTzua0fO4qLTX0DOlSPE5
BZOE/PR+/75FNMVsdzzxjpldfpf41Q7rUmgyxs904IyDUjMBXtggdLdkpGivjoh6
/ibWY33IKPYzHjZFM+4EoRILuoq148zQuf/F5NRPdQr3sRGZ/CMflt56MM+DaRpk
A3OoPinNKxvWtCwNbzmZKd43HmI3zurOR3vE3F7pYYF7KRCCWmeDPpRU+Q9uHvv6
jXMXFtCFG+93NVAqP+bzN6pnwV4eMHO3wtuQO6/iQWHW2oQCAQSh8KgyXYv3lW3q
rcguyYyQi2cRM330vUP+/I2T0BNwDqeW0zsoHwR12jiVTSFqz/jRdkiprRDPdSVI
pCAwriKig/ol8QwhindCxh2v1813phxoKqBOXj6ggMD/olfMJqILdbhMvqdCKG59
B6chaDn9CJR2dhOOiD0AuRKg9b6Wz0XPbJNKPkfh3ovzwnRfuvYXR5jN/KCPvRud
ogl5ubUJC85RTD0QXEko2g891JoZl0HMEelGXvs/Z5W2gDKn/+SREUTodf8oQDzm
wXg4cgDjbmGAS5e3skhlo4v/IxopjoQEkC12r+aBM+xkGquuIzxF3kgFmRPTuUZt
9MbBecJtTdwfuzBQveyXPCaJ9CY6Hc+tZw/NMj3CJ4/gCrGJspbGx98Bf1HKWKAd
FPRiXkkDbTA8MJMif/1KhB4dTkEYHjgoM9ZyFh3u6LFO51It62P7wilba0HFk9CY
8B9aWH04HXCIp8v0UlEOYy7RoppqTGdMwLsf5cnccsl181ib7NwBWB2LLSq6HoH1
xBYQIdt1iwwIAGgT0XjGYVvwBj37QoGDyT+BgtdbVlzyqFYsOoGmOhnuCtgVuDx9
SEl2nIjKQRb07IP3LB2MN0M6PBZLF9Y0BFSuQZWJYi1b2akVZxEFWmUONKgsluyD
1xCSqXQ3cJXf0JlDZNODkO6Mz83Bmy9iMTbqPM1q1j7C64RLbPdZIf2EK6yNYR2y
aPsnT6N5I5orxBJnDTEY6Zsau2BEN9g7u6H3Cr/IwrIH/xix53SdSfXjC8x5i/FU
kiC8cN4R7+mWmkrS1jQfhDdNTl6AWjgmrIkUKJRiD9eTc8uhA60GAmjv+dN+0pSQ
wZOso67H3FILrQWg6iz/dwDPOtUyBG47QklgPOnn9ul7E5HYpZ+heW6VAgx3g8Nz
FKxpLWhLKBPa1CxsrPcRze5BGBa7mtsMaAEIblq4sh3PvXm94J9vARq7QrGAOx1A
5njHQmezRx6dVADQhMJpq6pZ6x7t5aqpCSYT9e1Q6R6kgI+w8COWCqHD/euakJXq
eAx4k0TG/4mLUgEjplqONTsfVOscw5q5O3PqA7//P2mSoHG3Xq+9HdJZ1MvvOmO/
XHUPSfA0z65VQv7Zs7p65KyE8rtjxVQqzI0sim0E7MBlbYbha7M8AVKnldwRFoX7
G01qINRXWNdyV1NhkxljCNbrGTFV01mwEHF/R1QQTiRbNnfL3tO79Ncvr0WeGm8t
cDQwRrTFOvVUlaFg0AknP5awuf+maapy37Va5mT1ToduNBxcBfKDNsOlPmsb4Dfk
aI52dK9X+uxtWaYEnpHHw0RTGPIpTSuW/PPnBp4Mx3aYEhT5ThkWNzuYx0BErfcT
H72XPHNJ3X1F4uyCbk2KcWLndMq3uvVyZAOXV87T3GuhFJry0a4O9VtDzmDSZI1R
kLX+WN3Qu63JDNdE4LPXJNM9DPnEpdqYULeKuIU50Uu/4O6auN9FfcojUW1hlgoA
a18Ok0RHA2k0TJnBYLq86x2D/FX30BQN/PN7ckL9hi/bcxYkWU5nLkDqMYQXcd9a
2riBtcbImjbEM7R2C+aM7R2YBzKpYlmYVLYj6JkJMEbj8u04LpqeDWzo/v5FVCj8
813rfd3T4zIx3uSsqSG7uUe3qCcBRvNlJe29gG5sNsOTKK7WJhX/jWPnT9d/eX7n
hYWU4IBeEWArdC/AqJCpIEGwYwUgRNFMfNSgK8F6c6b9gEwYlGemfS4Udt6Lwrib
zzz5/UzBOJbs+TvOPnJSSWutpnnoUo6r8yNRxC5FFW0WITfZKO0xPWhtRG2Znjqd
4OoObJaMyQ/yvBdzsrC/bTjfcSmH44tsPsxPMZ7u5J5l1qoHaJ68e7nwRsLZyQ3T
3ex7Ts14Zu1LX+XLcm51Ny9NNKvP4SbozEHkkVr2M4BoQZFr0kQstLHwsJvLXPIA
8NPDURhpltWRPkvIMMV1IsYR3qLoFapesmG7mn5rpg/QjCtceHBdY/FNWHHRLHFH
XUp8n1EPeKIlStOnnG12RbXlBn6yFQuvH8jcHvhxi571fXE68+B0yDZxWC9MRe+h
Fq8FuUHR85284qnE9rtpnl5kKYjMxBzsuKTuTSveq5vtqiudqAvWAQb/gYkHWJvM
LoVFAs4jqmVytImpVUbbA0sP2TIIobCBOttSeh4FoTy7sEHupaQDEUEf38mqTlk8
SoNAboHgSkMZJMUZG9ZCaMUUFCwPIQW9JQnwyqJhpFzbihvtHUpZ6hZkM97nlzst
4QX+ipjhBL+Vsk6jsmbdB6iYCvuOrIv7wS3uVuHTtyACc9cujGyespNuifpk3JfK
MPAFKFkmHjSbY5Rzf47m+4p/29LJYTJlqIcN3zNJriwzU/xMCHzhWrYml62N9DFd
0g71mJWWwYe0oIVstt5k44kKE2P/1Hbzc9bVrew3NgVfxtYwMhsO23PxwIL0C0YK
vb4FnyTdNZWx0OdtSIX8yX0t2d+BB+cG+/EKbrtcx8cwZTaubekJwSRjP78AMFgf
2bHmhAy7+9djgosl5goyBfrwPjnX8YUcLCoXcSsF8cJYEJ0JkE6BanHWhHczus3+
BIH4kZD2dRP+epoSIK5aKS77t2h5KKQtjphYMMFHIXMwTuMzXsFUKCHLAVL3o4g7
8JGDhveA1YOzZhAtiMA/qlOTT9Fx/kchZ2SHrzRTQjb+IGiMg7Oa4Q7IC+5ycHXT
GkhNFemsGR4hgONWElF8HT1CV343UrvQKLfkowCOmIfowhC1wv8edF/RvHo92XZw
SzxQmxccNfOnKKQjbeekE4rA2+EdTqPhjFrW5VTbkE4PxgUIBQTtWvjj/WMAb+Aw
Y18CRi5a8+in71RDcEcLB0It10sAdnrqC5niJpmmtYMPYeGZiIJPtG49hp8i6/PY
wGYawNrmgoYR0czieDP2yZz5u86N/Gu1HkgkRRGBhwAZR6ldumIA4/LYeA7pM4m7
gYX0rhzfU8mnlgBkbobyUb56AJKLWCIAqkKUfZNgcwsF3WAEMai66WzBBlSCi5b9
ajMKMgoOlyAWWHhjC4gOwes2agThiXY1aVhuvzRVMsfQ6xDybVVLMov0eFlbRMI2
yegmMM04UuQlliMqVioAu37iz/eXqLC2yy8JUzuZnf9CIKR42pxQgjpe3W4KLUwJ
E8HT+HGlyKg1gaU6SSMklSHsZkHAxWQQmI7jBPjptzsPtm3Q9rFUp9ur7g96zK+J
zvYLjeY/bKzCaEOblvIrH0pbIt0sLeF/q4oZrcOEXFl9z/nNFalBGsVuRV5g0dWa
V2iTMminN7PJoABQ1umUEQUwcdchmuS+AwPiXkYS7JLua9H9skaUE8Jl6rqOgzRs
Otb4P7JNSeaORKsGCwqBsR7208N+hGf4KpWmW2BT4y3kdHwoxyqxGUGo5LmjnLPd
XevDT4PT9LmJGS3js2JSGp0BK7ySZpC/cDQdS0gB/e8n6GZHP3cLCDIJT7hlaYlG
yalOCuwR3kJ82kGLFwZuy1QTPBCCTWEVxSnj0043bKlRIFmH0j4OAKvHhrJn02Y1
JGcC33lwgzYgX4Vl6q+NwlhKAuHwDeti3W1xbRYCWrRfJ7vroh5cBN4vWlb+p+r/
8JSXk++cgPrU0DKio0D40Jt4+rch1XuIjjXTcFOcxjGRbx/s/tI1Jk+btocKOr9j
TizwWcYEL2ra4T7oVAi4ZzuoTetms4QKqJv25C5F9NQBX7hfcG5Z+KwF6MU+l2f1
xYu1S14w0h/GbKOCaKBIxk2zUA/dbN6X/w7dedYocq9VuIIoDQMWhkgsuuutP6M1
LADcS0P4pdxHcA67E+uQxnYnGX57d3sNGLiZUSGhY6DYPJp5sJBNvBsZTt5aZu/V
6JEh21NnKBVLVP2Sk3++8Zkd4SakRLTyT14lfKjPNmWxq0eCFQDktAyksBkaQjkC
CXwiKL2pkOTIe7oqntunDtpqfEXBztmGDyph97zvTyKdDt4epjnacWO4DF3ikTYc
n/Wf538PazqNhaYH4gga1yc/h8lrTJftvK+BY0DKkotSuf7WambFeco4dF+YPTxF
brEbBnwxWFMoT3yzve7Y+8sdk3NVjNYMjattwFFY3kpLl+gqFqulncgQ4E4LDaSx
tdU9DeIWn6sAKYWn9EwoSH/daPgy2YdB8iCf1gFCtFHNJIEwWBGRTP+D1t4jPE0C
H+p+i40hPzfwcuBv6+lCZL9E1dyYtRn77B/69hnhmdnTP3kReXaGGKcjS1lR5V7J
P/f9unOmMGRCIBNNpJ8qegr3mmNibfHDJrMl4R8DWi4LC1WFPxgPSzhXqBfDKS4t
giDl80fL2r6mYuPJWHRc4zh8EA8WRdxswyIG/MpAcxHApYCgJi6Q0gCbrnckq5xf
HnRF8YEDp/j6ckpfCN3RsrUTQCL6E5KxYiC4RI0hChubGDU37Zi2fr/OV/YlkWt9
Q0s32B/333Wb+gxSQzXn+xhjXvzbI3V5ravY32GnI6Zpt6gBmnlrSitljNuYsOJs
5RqQMjzJgvLzYQ4yqJUxiAgvRsy+Qa9ix80pFJIyuipHoMJduZqJ3mxqhyTF674q
3uoREX+///Yh0wTl4RX2SlJSzvjivmernGhEsPWFchCR7j10TE+7V70XoBB6a1D5
qM9BAVSMHNQUlrxYodD9axcT2wZdOuzaUiyy9v5beeTFqVuNsO+KhCEU4CfHo3EN
dEqjkKculoGdkRRI+8MiOULbPo+KgMK/+9SZ1k1FZDeFL1ehrTZxf2BH71ElQr/6
/2OZK/G87d5WCyFiQTLi0Yjawk7pBfELxiZRVcVmLyH+G/eAgRLiSWeaXRQvPS70
1QnYACOK5vF0/Ahmote2QxxhRG268AZMXLVStPB7UsQC2mwEvR8Iyi6LKoeP3rX4
xNW5BYuVzj1Vs4O8Zms5b3OPy/6NaAozKzgplTgTUaCYOFdHVsOmiJOZriaBvEQh
E16dPDq68o6lGnHl+/39I7uchqNWzo7vnjR6rpN2I1xPFUuZoGKp/O5VrT7M843j
EFmXgBpGLiE8V6QKP17KAeYb492LyoFTVqV9cb8HjWerMBxs0HTiF86wOc7J7RvT
tf623CXvkJ+aebgpEBSi4uYJGeY61WYwVk/JdneLbvynIfh0ZT4e51NhACIk7+XK
E2XAEI6K9eFn9ALVPPy8nXbcmoGYS+pDxdG+o+GZFGE00iHhr/At3jYOGnQszfuC
1tdQuSwM/gkv4ro318RlMXEzdEMnCpOPbyshM7c8/KoPikIJ1Ggh9YCWt6m9wql6
ZTTpfXjDlGFz+2vF2jiMYzO3OU/nZU1VaHjUCZ5J7v0YDiv9DSxjoAQNCYL95+CU
z2dc7QynhWtoqAKi77iNQYPpOR3pWcQU4tNIjNTZVRrkjY53yz+L14hcCHfjPaA9
nlCYyuksVkebzsesF08+DtYN93lu2rwl3Do494X3SGOgOc4qanEaBO4Bo7MU3s+u
uwmZZXZ/NNsEmlCf9Cro6p3EUjWdEIT0vCHJOlADeqbBD1XA1lfnG5S79wtvHP9h
R+aEzNmmG8fjp3vfE999iV9ntsxDaZSqhT0/6SoNe1eBA3sggLcnLR8PgtgH35xU
Vm1rCJlnf2oJvBay2C9+oCBQWHJgARGm/ePbwNYt6PonHZ9x1PCYrWaMfpnhpN2t
eWb71/bxBo2EfJEEBAERlDBFfVEQgUO464H/ZD2Txyp48h7s4Niqt9au0bvZGZ9P
l1i2eOG7xhugJAAx+x/77WkY5DBSZ4FhjvNbad4ut615nTER+SZIr5KqypLumzU8
1yBmXtsNYth+9GNXZGb4rsASKGT3ME8AcZfscMKDGPo5oLNNPwW+/iYkNdmIByM7
+CZOJzKcnGK+M5CzT9SpMLy5r+joXHIzMJoyMbD21RsBWSneYhwF8W5Y3wmzwPUN
ZHFuPdLG/q9Zx1pbf4ONVxD4oDefNU/YaO2FIY9F8zPOz6Tz/R0BdIIEH03BKPyN
bZpTby6IbfuaHDsz8i6MpbBh/62uCnAC+o6qEJIvwS6M2o2Aks/2bi+fEef0b1RN
8lpun940VTd2qkM7JxyKZR0P6aGHjR2rWjEWsg/yrXNGB4iY7nNf1HYuj7HHi90s
w8uHA3MhSXwJMZMuQBUw4Wxf1a8lqiuLtNDYLfxtYtw+jYGGhj3R2IsYALR5xI7p
DA7rYNPV3NeYVsODP+aBf5EHbmBSy5HQmy11qyaXzQSTkCaaizaHc+gHBYWmsgKJ
lUyE1aKuuGinLiswa/K9gXe7bJN4NGPcVgurgQrc0NUjlG/D8EiUdNVXeP6rGRAG
1q5ipZ//rqxIxMc1SrNuiG9Z+bd3exghT/ysapSAGKgw9VXcrSNppNSGa6WDm90o
yu/VWwDKe4ikfGwhnfbugBEAiLQ1XbUuAu20bGf9+rp2uqRAQOYFy8XU9VeR3X8L
`pragma protect end_protected
