// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.0std
// ALTERA_TIMESTAMP:Wed Apr 26 13:33:39 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
tXEyttYJTyXtjKiEzjyNHh+QJISXFjrHFE83bd3CZKDl0RfNVMc4STasIxuBJRml
zlttvSYVQHAzhjeZ1ez2qplSC/ACS9aFe/V3AR4CiUJEXv1F39vxgWm0cTDGnxP3
VJ0AuGR7zgn8dMb0YOohk9Y2JNKpluqCz9O3DXzjHAs=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 57744)
K31FKBua7pYr6WujiQgRX37e6ZfWF8HjS025RyUpBnXosTmLDQIVajJI59ZDnNId
aFtVSxu86iNiLCkWBpkuFZpetQSnIRVo+XpnIfk+iMjrASnKri5N7nhl+aFGyIZY
iozBMx7ChK2gCe8cl8Eep12uPs348E953Lwha6sJD7TC1eDQ+v9rsuzrldPU6opH
/rB/Cu3gsxjGbo6zHG54tf66zfptQvRhBNgxTGqiFP5q68RUg/tYhn0miYbp92kX
hbnSsnYs2rCAOMFX1uoa0f36tU9w+64LKx9l6vogKKsypyP69hVFT5AFvbddilce
eFtPZ0ZzuD+Evg/C4QuiAOwB9CZq1uEZWBOFSE5KwDu4Q2yKaf5m/OUnVUZiAJI/
iRi/ZKNCv/osRL+6xFV9DvNAOL9n+/XPDx8phWygkbdBuTlHeEkPMXmB3C2VWNlu
oHsSgfvLzpKpDSoZMklHIjFKQL56F1k5ushiImx1/U+60uW2pabwhWjnYS8TRbVD
XdkrzmmjCb78q/eU5zdTxnHCpdEAuuw5YmR2ccbtoytO9Kk7r4PM1hjcsnVfp/d8
Dy2gymenP3Ih7Kzvysgi5jMVARkZJZzyVJXOUe8r1LUB2PvKrj3bEILMCyvr6/mt
0FE0Q87G7LkwZveWIwV/uAyLs3fNCZm21frpg66uubRZbwV4XvGTKiVCV2v80jPo
kDLMjs9euGbxfbBYtlZznu8CKLwxwcMe/qEqI6txLs9svMQrDSLHg16OwQZbJEVG
fO67KRd4/cOaGJsrGA69uTSCuG1x1L+P62Xn+QwytXLmZ9QpFWlGfrzu/y74Qb85
CKPHKlCJ+79Ppl6/LKGOShOY9tbwcqyfnP5iNW1jWjt6oKMZ5LB6rzDg+tOrfnDq
OkGjp8GZpjdU9enBrVpoED5dPHf+saFMk6AYBZmYObar5iunTwlwvu1H4P5Wko1e
SyVOKE9S1y+wPnlxH5x0UM8onskc1DzkK9dTLq5GHxhsKiFaNCCBHbf8XapAAzZO
+hKgOQpjVb2ldQDUrBpI8rSNoZuO8ZFkKYMlYI/JJIEHbrI4mwrGB9BpqhrYJLzd
5fMBde51PX1hQPb/y3TLrTdEcPTzwrTGRZKA3Y+hqsJOTFgZP5yU+IZ2LGr9F9EA
Mw7BZURwhzD/R119IT1GZthVmVOCREV0B7BG4/tTe2e2X9JPQNlXL9AURwtFYDDD
hsd2y0NEvYGb07SnfdIkS0a174zlUrQlG3thov+cygXOFOFr1Z4HtNAPPRYRuuke
yQsEYv2ZwFhM2dOu2LKV7Rf7Q8BFPWEr/7eAFquNds+V8ec2V0OsHyOYSSST+ov7
xMqYeAhYAzgwlT2dn2txgDZolynLO5E+GE7wb+8OpwyQc+2EM8pDqie4VQ2QSS+n
I0QWVGWidW+jjAGzcke+5ne8SCnWW3pMKqAwJ6T7aWwJJiSMPSKwFgMcWq/P/MYS
Sp47V7LKg8nOP/4xJpsklOBdr1uBCcpjGEg4naKPevuWkR+shnlEN5fDkgMgjBfM
DeGcyuLhYjEVX0iAc10PKhCRJZI2+9aQxbwD7IpBQ+M4GJXCUUVK6zlGgaJNSpBg
QBDJ3GceHVhgpMMvt0+tFvwmG8wIQ5a44zrom33wmPO9qTpPW2ZBhLvLNR3k7Ih1
tTcpKxIJfML/ZFyDIXUWoR2cY5Sat4Ci6gMPLBbXjOcwPB4B1NtGkNMaqkbc5Bgy
WCeCR8Mi9hmx5XHX7eyPYtZZ4PLTK1ya7pv4Fw1/5dFvR4NZZbJy7cCKIRjwLVAO
UcPov3Tt/lAB4vMz0IWWvxl9tv0uaOVBckwSqkvAzFqAbfd8WJ1xzvPHrfFsPwZ4
JWalHNeYXcWQsj/bChPUJe0HxjNY3GZkikdv0GmBar43+iYl2u3xpOqoqXA3+9vE
/UOwmQce+7Zigf2fJLOgUHw2cUaxVkzQC8Qu0QtWz3Gtbsye+Bvl1+Mxzsjs91qx
+m6Lv6zLb1mdWsHtFyG16CQ2CbwpCX+hjGQ0dZ6wTxUjDN0GANKHDgEkEOoqiVri
Az16apUC/wc0Vu37vaVo7Q0W0FY2H59LAQGMW4gojFlGdpZ0d2PC/PM08/H6InqY
Wj/Sdwy75dRlJ9C95GTE7303A8s6c3wyH9uGfNlL9+J2XCm9rTErkMQ193LLa3Q7
KpqvM9N8og8ZNI8t5j+/KfZvJ1AmBPmdOVgLtXuSqDFdr+qtZjlpa8ZK6oU3vioh
JAzK19OYHGws2mt0oIh5GjN2LdLcrMpVzhuIOWDrTCnYHjODDtR1VqbaOJ/xXzdm
vOX9xwbN+0H0fGF1GiYyKKrRspB3Fb7JJsrcFZYXaznanAf9sK++ohWjho0NoZCh
1xdhI6wnvlhzN990qMYap6cVebosMOnGwQy8T8h7PfkDZXz5D0chwHaWGD+XQKDD
c8E+ktswbJ09HUNGsVpo7oynuSO7hbmSWrfeB6AUykjw1S0ty7H7ZeCzvePPKUwF
mDZYoX2RsxneikGIpAdk4zhzHL/f+39KIcy7NloJdYGIULw1nqEewyqNrmQ2VUFQ
xbsGsUnaygyPcJe8Jklp/bLEeyhIGCdZQLIY6UOSjto0tyLuKia7nGsrRJT66Yok
QNk+7XJ4ei6U2QjUI2N/eZRV9HnuZZI5a/NnPoHIFyg32joDS1uIVvhRbrg4RDNZ
rxCaPycuu2tlwvUibs1zcLHqSCX2Y6Y1RaEx5bI8Jfsui4UCyGBphFSU4RgmkMxX
72tLfDAMy1MLNzgTyl+dIbsy0iy5wKqW8oc8E9OryGEqwnZn132g1Nn0wzkrntIH
MFLQDJ7lH3/FsEeq4LxLLs9qqWYR/45jOp3Z3cnTBIi+zHxw1HIabK5fbBYQ/ZUh
LxSFwHtH/XUMZrk0SHj6uLdwxoCZTBtFdm1HwyoCeOi6K/cGjtQTrf6tw8DpSItl
NhpMvViDZbf8WObLlHS/3JxkQirrVczU1PkoX87grngj2caHUM4a5h8r7XPm+t7j
djrQJz1iMWEl8atBk3wkxeqEX4NA3aKz8hT75I3URqnJwwJZtgomgkbrtZeyK1j8
oOKZqVLSYvmabF8J8yCAI1eP4VfyTq85ygQE4hNctfGoAfhMf5vt+ipj2hss3W10
EUarkl4BQ7PxFhoTPQdidG9NiDEy6UWjP3T4HgZ6RvTHnqf1ArYW6ctrE5qIRfit
7smPwBw01AD4x4wjP0vau843ms1yBXJ5IpNBmxUpKzUDMlmZ8km/2zo3mz6n9o5r
ObqZos3VgWMvcIciPrsE0/TlasJh6B7kvmG7QBnxcHFpNrNH0MDtt/cz5vPkL8BJ
53iyElBZE3IM1hrlTkOZcnKTC0d2lF4ZQq6Co4LevifP9krLsLpWdeIAy6vk1B5H
7KYFiQ7GMgrE/QffuxYW+Gjpi5fX0etGqhH5z69CZ2SxfJBvY7coVsupvo3CudAL
aB9v813Dl8omGyUKBfowwbAolot+a1JMmCkt9On5SSqzj1J39fZ3zoPj9QMCpTb9
UOlHv3WgUex9iIgFA1RXzNCY59iwCjEypC52eBzHiUW/kZIF8pSxw98CN+ST/ZuS
0Pvp1EGC4BZ0NfTOWEJlcEvzpvsHzO6pSSuV+jUjb6Z3jZj4DRgPC4GXKnzzIPdH
RDhcSmrocr6ce2vpNBjsHUdOdFPltHr9Id8muaBBF3K4gRBTUywnucdR7VlGqUF6
SvxY8DHvcJLwbTYJbOPu8YA8hcqqDu/2To5flV2AHrdXN7zXlk0ZqPCk1KgrfACi
0DfubNYLz/D7i5RVScFAgrUOzCC+QvtTENJvYEyyLDwDDGG9UnRT4syHe+3HHtPM
3PkKn3ACrSyABUnDPoyTmFmjAUMYSPG/od4UQEk4Cq30fI3oIOxNxWOGu8l9pM1G
K8bALInv2O2hDMQjBdQV1/7kuMzoRB0hmlEcfdoLJjo2jWHyxEXCcbB0DhYTZMvR
VGCponKvNNWdXUvJi/pm3nvmc9mHYKoWzEoIS3pb7iCNKInQ/P8H9MpYsLJE9R/2
XonQOVvldd6zZXowR67U7PN76+/C5TCypRLyn7owucLhsIoOCr5MoQkmz8BLHCnF
CsfPb+C1ZUZwCSfbWw/HGGUjwx1Lzb+9s6NB2l2Tj/8bEyC8ZDoLuO9FsVnJjhYN
pYyB4V4bbxJLwvvSAV+OoP6+szKCl1zVozjR827Tl0p7JlzjpAezOgGLFEjyBCXi
icocqq2gYDAN0a2td60NMsmukAjIyZygoHUCUwfZ5VdE06lIOZQlCQbGfvnaqLgs
4+LYUGorZFlV4Xg6FUk0vGNExW2+1ZjB+/5ZoffD6ym5iE70N1AbeEoV0rbpYSvS
7l+cIismzG1J1OdSuGwL9nf/mPKgfo4Ena3Z10/klhvTJawfkzFBC1KgkbXgVE5c
nkGNcKv/XC1qQBrsnZLBoJUrooFZl0SvHpntTzumkuYTMZmoMW59XkvzVKGZpoRC
lrhdkGha8D27XJwumkSENKpwE9zjRAoGaDy22Y653SvdW0BX2Nrkaepq4HHdVOTQ
it/+DKcRzCQN6RcZznmz19Y5NicQlLewNfkTuIt+5UOGS0yauGpI8kpX8Ps6q8aT
PkEunYlGENqP16qtdkLvCRo0YcVefjbtQCkUnVN+S1lHehCbU3q5iYHQkuKp/yvU
HYWltRY35YDLRwVIqGbwgzQ3oCb9q/ZQE6nOW3IqV1SKkLIGZPVmUG8PQg2god8y
tRpamTqrDKlpR+b92PtjleDroTvlNG4zHHTh/u3rqM233sNDTis/em5dM6PSLVEF
EH8PiS/p4qPVGOA5yQP1qcx+Fpo3m1VaMZY3On7Njbq2cxsJ5S9rDSRQ28ajyPFV
aRQo64TUADCR1Eng7QGuSB4dp41uGmmFOU4nWOC7FjYuYw/EzezgzOQ2bHUIsHDj
uKOgVfwy9yol+6eAJoup1hQqT7PyQ/os8s+FjcGJrRty4dtdqY6QUicwR6vftw+C
r+2/XHY9tBmXQIr9fZd9Odo41wrwsCtn2FqW5N77BFRC4QYFmNh6yjBZaLmoDgXc
rkd1oRcrAEvLiOoaHWeTphaCxhjm9n2kvyDeA5+N8k3piUzXoRJpADSxVsYts+Mg
gDusElXre9pRGhk7OAdlm46r4pS6BK/UZwCXMRJKfdLt5KSEMF1P9XtFJ3f27aPu
xuW7CtMppB1VVEzQ6aP1c5HPvkoKd+92X8baIP6nhGYDZh6cza3VhTnLXV/hjNsZ
AshnP9g5bthUUPEZZ7W+/WKdNoY1cZpoHIZycUY2UXl59ryLeEDFJawd2yF0hxHf
vFRWqUYoMbljqifyuMoivXbGq1rNN9QWW3xeIJMkOSeCdyZ2g1j+jX34NyQzYwjs
W0yaYbrCaTzkTZPeX/KDXdqpRVz6iP/NEAMVAGAmRMcWEX77ufbpT25mZAO7TrSe
Yp6PqP97S+6BRom4PGiCDzSPxL+4fcjIjPRN80QVqMFGP14pU9UkEh1q7sCfCFGf
47oxcMSjQXGNJkAJD9tAJTosco7oJYV2sDRCWOiohfeyeCqOKa5AFe0+H51E5Yc8
MJP+r/BDCj78ImpJCvQGyvmSjxVHwg+n/xnl1xbMq/a4rU4v9nWHRMGB2Dw1kuiX
TMKzAw2CJ6WPptu775BtlXQpZe1x5uaAEQHC4OBAoyphx3VbVbd8+fEg3nqE0laL
81OIxB5LQdtOf515FucBwOIu7FZOpbjHPXps9whIyf9431pv4A32Wt36+jPGDl/Y
817APFXw5vrNphM3ysEukqi9rEIZNXja92P/6gIwi9SBhIlCzKSs5l1Pr1Sja+lj
yhHtrlGCmdpvnQtzRJRbl2e/art9ZJwlaXA+Yl65zOY7G4tDzlkc0I/G86xQJr7r
9pnXxQr4WapDod6qHBJVkRKdKEVo6VIpv43sJi/17SxqPRJTHmd83D5nw+mFDe42
UdNoYqm+Q0dXkbVVHfpWD9lQG/5BQm6cXJLpZ6LVj87b9bmxJJwRF+/D206PUEAp
9Ec/2JfANvW8RgLymmE5s6yVfvqO2g6mQJODUOFSkGPuXoxSmceojFocyB6iC4M2
oh2IhszeMNRXqcv3/Vd5YKDXN4mjQneQQ1KwTxIX/V3dC4oZLyZEof6+DToHgOhS
fbT87IT6ffQrPyZHLGVLDl6x4FPtxeD5DZQao0+PFPU5k+FWE00ihLwG7XEOGqVJ
tiZK8ZBh2nFAiwoJBakRcDLzcu7Rs3r2BpxElp9cH3bKUVe5EyOB5ewku8rYLehS
sKo+pc/R+bZu7ZknIV6bDqphXTGGudwnqk6iLdaLzbrgbDWSDidEK6V4TtblZ4Pd
0IuQqrZG9rtzkQXpew5VswDBEk1HpEXY8qUqMRuACz1rrHVjOqYo2yl2J3kS/0L7
K9rgzYOH62jUgdT77HtQjTOvUmNLiHtmU8hwf81HW4efJYGGxvv804wASDvRIF0+
BEfmRop9mKkXBIs2U/LCyUwe7qDfh6/tneNqN16FQx8giMwlnUhY30sA0b6bmh56
tFo41wm79pStC6A2l1KfvvhQSotBJ0RzV6iUejD3SvDJ47ggpaoIncTbEsijrITw
7Hja2l/FIBsCFNprdJmoMOtDa5tQyF+dMmD9mTayC3Ie8p0jKa6peB5PkD2f/O2Q
kodRaAFiYQV064o36KlSKyCI3lbS+DvV8eicM6AWZkuIj0IKjjmMn8T7/H0/W6Mr
rfmd2PNU7RD2va3ztxvMwdWtKVTTAEQZPaZywpK5bmm1lJpAE8oDX/PZQYaPnHWp
zECdzBelVQcuilbAw7JWWW5chJASLRxyvoGAXLH3sLLIa9HzrSmGOBkMAp8lgM+s
aYx+oe7IbPesx/v8vbG27r+ZClJIWWabz6As3ZAYJPEE5ioFFk7Y5n5x5cxBcRDF
BBo2PPOfUJc2mC17bqYCRWwh4jhJ7X7ZwY1fWjjLtFLeoBemGQ4KaEhR8xaKAd2Q
HuTIJxzu7qQ/vcwixKOER58FKzKVyyU0ib/ZEamjrUbdbvmDU9DkZTf8BQfkX8dP
1mtbc+qpWwbCTpC3Pa51YuAGlOGr1RIM/emZklN7jWenEtecqM9M7V0RQFvljP23
xutIxNFyxV6xQZhedl6NvJcB7bNf7wCzy42A2yZshFqjatW39tNArzKSe1e6d3Rt
nf4tpfsCh1wZpXwNlRviGVaWy0F//ZVSL+QnV89yWskpp/vN0mCt2BPBzazC3hcK
DmaDgFj2Teq+ckFD+l2WYW+m9kBxrO6X9Vh92ASq3UNPOh8TraEhKi6HeJNwfYeG
2zldW+BdYn5iJ5gggPaYkhEpzfhoarJYg+veaEq2z89q++7S2u08LooW5i+P+rvF
85df1ddvYLf6wqaO7Xzy1WxagBNU0kg8rUSCPhguNeVy5+3ayOcRcO3NVQ6OkVn0
yefa1Hu8Q3Ao/uWZ0dxeZjHRxFngf0S/h1TcjaJtknJQ9/ptqejMYkqNJdOeeJ3w
nVAwgjRn8NPPQP0czJ47bbNiVkyhonqOyH0PvJmM9xIaNcqvQJuBoLsZwNqv12kL
4mvF+xlEowXxPI2Up2Wetw0+ZJ0q5Oo0MA+rHgw2VLagFemwhoJBOftw246CFo/j
AnFU57JwnnjzO4BFaes28z8cuJdy1+9ZUbJKgN57UoGATnoAiq1j5ET85DdBPwus
2+0b5F6RSFc06wmmZjtPxOudIv3ios/1HMKAzN72whCl/A0bBnIJlFdaVQeePFL6
1SnoAJnf4DlnmCUVM1kinlAXUkoMxc/cvbD1um40wKp91YGByWaXxdQJjc3NDBJF
PUonf4WGlPAjIhcdm4qA6C+6VSW2uvYbQ3G1yE4QgvVO0sPNfuV8orpYYbLNpS1N
H3okZXZMos39ZFdvuEwDyYeWkWKW0DuW5yXAf/JNaGFguNp8bffRv+vLZcG/8whV
if4BQl3KLJlFzftC5PbvbiCJPOrREA1UBOYYE6USSJXOuYEKqfmXX/QpmC3F5tvF
7v8MQlRgSk/NJ4SZRGeQcrbi1Jzm8ztJmsMynVwi8tG5vXg6xNklJ4g2QhS9joK4
ITTbL//OjEd39fuKl3dd7Ju6dlMXbfsQ7DMY+bpajD/oZAYH0jxnBrhgkiMdUQLb
a73A6vfyLA/IsQQHH83hcISi8Yz/sfNDB6M7dkrjZnAcW+fNd+TCi/YGX6rLJLUK
m23NpvYgdjGUcd3CgHRD2t1msXhqq/SPLUfkd5MYEAE5E3QrpuwTNcJUmIKT1dAT
6MoRrDk2Og3i0vbqiehnQo7MirXM0EQFuLQbGreqBAftVHiLAQ8V2Ajaxk5IRLku
kHdOsYgZvOnsZ0E5R1ybOLZ7+qD6l8pxy0z8yyQAoZdm91qxnPcYbfYa+udFWGLu
i+HUom3agpnGxqyucA6Y5GQb7RRbHSC4NNSrrx9jzDVD+SGFAKTz1f2yfEdEN41b
Iy6hSHqw+O3MqKMao4eYVykarafvcm8b9bgnbI7dDBs4TA6rV6VJBPtzc3P9oSXy
nyq4ofZwCLoRxJmWNlrgdQD7V1zC1OtuLVCxO4j1vAwiX8o85/8tvcPSpUcZKI2J
SBPZ+T2FBfGLk+va0JrF+wl9/FEm7pj+BpIfdYfcz6bLhJ2w9tGUEvN1VwS5Vqjm
3SR4bPFB5Yuk9bEzwapzPjmxGb0QDjWJVSs+01yAywaVXGzmuC17UpDRosuuDRgA
gD/+ngY+s7p+o9uHEECofItF8258+zoJP1C/szlXOD4mD5jG2jnJK10VaoKLslRl
8uq9DBko2YJu0CXEt30tR8bGsqSK3oZq6jYTAmVC1mF4JzzeyNXWCCZMlq1r5HHQ
NtMs4uVikEKwQWxTyPv96p9Er1bAYJWAYuvenEF+cZEub2FHgTwz/yuanlkGBwnB
ekPEPUgUD165Wp1fIQCmJJr5+NxyIabwkS170+WGfQ7WFgOWqYcwf06YkTWjCdYU
RVaibFUHVqb6wH9Z8q0v+jM5+X+FnWDwR2vwC65XsS3rIdSRNcRnLngDIEeRZ5I8
VqecBraSQOALqrKtaUxK7VkCkOLgbyBpNQRTBIA7P4b0HYhXYnd1BlgOB6Il/o1i
vjpGWOxzPsPpFNe7+WGYJ69uS1Z/XpQXQ7bbJk77Wa01008GzUKt3CEjdFTDwz9H
19cnGEcx32kYRV19vQhd3+X4yZ+4SDM9eInqBdM9EVark/cx+PUh8aPfAF+duLg/
jot9E1L+L7YBKqZy4vm+EeP4EsewvbRFPqzwHXpuIYCnMLS0Ey49rOtArpPdzaQp
kg9JwhwUhXgeFayKEC+I4WMAcXpGXR9N3iw4uKvk8J41SdJ0EdoFomAO/mF8t2K6
2HZzFrFaer+R7dM/Uuw8OcuCzI7jQRPqi1oyWzJ06YIpHuhwzwIvqp8znw3HWv9r
pwAk484MLneec5D632aXlJS1xMa40UT2O1B/UUXfu1MnVgYxo3DwztJv5PKSGch2
ZP+xQVidYulocXcyfqikyhA4zlV5KMLHmWbUOCMvk9aUJhvUp7+A/YauPdjuv3IM
IuVZdra9wQJU0a3BQrLE+GaSA++ki1jE0VTLdbNoCQl5Ba2esZ4Pd96ObhRLfeCw
Zk6X+bB6EokohDPSsXmgT8NgbJrp/WuhfyXiVs+ORmGZ2RHzq6HyKH99aqzkReq8
6IIFrmueCXlcg6XnXrJaaz09uxIHBUaNX+ZSJoEFukesm/0IkN4syPW6SDxSZb7m
ZnRGtKjmm+yC2kM06f+wla4G3sZNzhhUYCKvIRjrhBjsqoNO4RP96KOPqZ8Rak7Z
NrGHL6UG/b7ZoqmvgctA7HS+kOOhHerbBQ+gvWZUoShDMzBjqE+3/z+/Y5GgrDt0
QmQR0fsin/Gekgm9jotK4lGxzBKo4EbF/uIwoUi5W4tfhsxKBxQcJ1XAxgtu/vCo
5GOcoy0lugCkuJofnAlgqUT1iOIZ5Hzh5iTyo5N47A0Dc9X91zXrJY4V0dvoCIfI
jJrD1BLCrwBQYlmr2Bokl9B2ZFbT5o32TOpyp9sYuJFn3kjF5tm+WfKU9rAeD6s/
Icgr5ID+aqvXJXgv8T5YquRzLp2lzWT1Dh6TUXkrYXEyy8McvaT6CT2fyB7tT8r4
4r8/TpXvmSlkQd3s6EvQ3YVqASR57d4TTjJcr97di0viWCi3WBKbpO66p1VHmpkx
zc5JgC0aX05M07tM43DoUi9um0SOOSToAS1OM+ZfODiWHTY96Dfg8Eg9pS7PflBj
8R4w9XARBN3zOcy/7oGos1+nNWQFjJsGeflecXU97t6ggSVYpFpOhuAn3Q16k2FI
qqG3FZ+H4nqu9eAtir+KQXbWFtk/QehrKUETiat9+BSPpXVyLEdFTpFy46P5Eb2m
/aMFpQvpKCnqgJwaNqF9QMDpEGxZaLg+t7C38uQLAvE65NqeFeXpM+ipLP6usyV+
LkHiDHTXNwDhdHw2hzz8+bWY8GpmiJdS0S2vEfveja6tg0Br30c5XDVuuRza578q
3w9JFnJMxx6GcSiAaictVuMAnqxDBhX12Pdf2CkPsAFWhrACchBumh3mwTI4Rdhi
vxIAljV00eC/ZzbNU+Ihz/MLt5J1du9e4Dc6lCGYw65m9l/JyaaumFcm0FDOx+Wv
9xb+jzalIDN0SRn42Xnwpvx0GRDEy8Qv6tCvunL1SPoCUKzrt/BAWnrcsiXIgCF2
T6+gexQJi28ld/qfbjBgqpL/zx/TvY1j0r1QVV3Gzeg9KpER7MSYwKQ0udbTfjxc
QnWVS3IByH5RoBTqrg5R1YpjoNf+E5fLxTj5XrC3CrjLVitwr7k/EKszjo96pq4O
ZQtMO5D//iNtlmuhvRI7E/5GlwUCAuiwtWecrzSIdG2aMn3FObT5tR1Enb4CwAOS
gKxlnrfF4lXzPrqQH0JblQRuIuBSLxOVRpRB4kYIGADYtwzSljZMO81YMVAFrtn+
vFHylNVVPc96yh5BQA/Vw95rADnJiOoTiHBW0Rhq6WUoNYEh/r32vghnpUinsJxy
YYpZNfMjL6VYG1xnY9QJZ7LQeZ40iwW3rOurs6yd8NE8dKC0UCaEJy3Qyi6458W2
26Bp/4sELa00gLBDc897JRZQCNexSRyfkNiGOzArqNCX71ho7bH3kPPQ+DtVvkcb
69LZspFa4E2/Dl9EOvNxXz0rZjo3AxNVY9bpPi2S5nxN3jMm3/t3mXOHixUKNB6c
R8QtCczygSXGKt2ygoWMK3FoBTXo+Zd+EDM2szlgTYQf2kJ5DNsElL3BT86eAWF/
8t+AawCsvhhIh70eXWYXC+lzlhNmjjBsHZ9cJ92HLeoq9KTlbh2RvK9hSQj6R7wR
AgKzma927daAxIlty+8vOn3Y6/SAesEs8mO8/7h9iouB4raoOCl0yNK/ylc9Tqyi
Oc40TJk3FrktQ9hyWbCnRN1CvVA8B92abQERqMvXIhEPvvYBiSqKDrWfRychVuTV
xos3jUiOElibBlpQQYU489glOm80PbMl3/euiKwxujEhtbUeciXSGqTg+KOn6S57
1JOoZ9mjE6WY/JpFLwjprkBOGhVuVU7xx84ZAmcNbnwxeqT8QgAowwGJomBMVu3j
x1C/ITRA7Qfq+qwprF4o+vUGkzvaxt6/t/AKxeyU8aKxNw6NB9YnhZWX40JWDw2Y
7l71+uxBbR4ttHzgSSKCi0Lwz8z3ytvw/wDS1d66KWBjTKVPdMZx9c0RmKrdDCj1
e4fZRQH5YEa6LHWseu3UViWBT0QQN+vmHTA4pakNpSMAcApiOzWpXlQIUU4GIQlA
jp0RT33OMBnDL1WdJmZ2E/Z6uXIs+q3ktnolCW7uF9pzg/rTWgd7o5qLkBYEJBK/
hVmJNZR6obMVtijeTF7N1AYXdUvtaDn8UXyduPNlqAFcPBCFwkk1jXzKz0ou3ebJ
yVBrvI4L5GyjvavaptISS30wL2giCU4eG4R1TV+NuQzW5cLmoSIVwADqVn5HVFr+
r8hKbBcZZKRfi1ESb9dEcZ5op37/x2C+KsHC3X12HQozR0IfExzf68/BCt7mOeNq
k1pxVqLe68qLvdftQKOevaK7vT0Hg9ciArI30OVHJ61Ind10V6ReEC7Eiqy1VU7/
m/a8bZmbvRMdUXD8yydQlau4anH+a0SrOKMWlFAtoKc4Pjzm2lpNp+gNAv4ktg4t
y45Dg/5nMpLiXDUI+gnOsfsGb4oTcM9lifG3iZl7HqteznPIM1sAus1TFFqAyToG
zk9NTOB2WOmyIw4YzoIrNX1bCUhwY29Cr9HgfvM5yuUjvu5PbQmVVlk4pQIFFHs9
tdhGxCNEcoreevdhOEKgXU2iJemIc0mJOpt9NSnYihxhUUqoSP5QKf3ohODOUxE8
eDjov3B0T6XLf0AWpQ6oCQa3/h/ccC2jybI4xVkP3qtdJbdBhuwotJUxrI9rzdl8
49t85/qluBJER2P2M0Opviul9u6FkE6eTZNBZeUVBeiNny0G6uJ3hZvnEzzBuJVx
DFv6BMBNI0NEDWqEACScDqldx7ptrubX0dSxhk6E/S5feMITOYCShm2W92Gce6dz
VWYmAZ/NUfPRxY5UnGSdhETG+hoSHE+b8iaxRly2Ew6KX/JpBpbjXTGaoc7KvL9s
pIcR96QJF7qtfPcEQpKAXxSbpDRUc56uAk/D4YEYaKnSeW0WlqtGzdwe8uK5j+PI
x9beUzVFa6lydzncG0D9RNWigekfAxZgSqipBUBk8/Tn1BbCUVSmLIafJWzSVtPz
LBD/IwmYQ/JDnSCqlIOYoIKKMdbmfMlPU80GNIePOTElcrC8Zk/QwhEDJuhO8yw/
rLlTVI1o4flHk8wQvT1e6wgGpdstuxLFw+gQo8IZ9MS1kqIvescLPTC+IB4Q68n9
g4npUD2QedwS3wmcoG5ap+0aTxu7lsSo0CKP3DpPz0vwBDcL/r/2bBxmj7Gg0KlF
78QvbJUeWcZ9nGRRuQUi2k8FhuP746IKD6xBZPm4LUVuxegN/UUph9NjhJQlhy+/
CzWsTUKCbx9xeJgTbiccLSDWt4v7eVF8xs1A3sHbnMDaCLDRTGO75Vy5qzmGicpT
jY6Jm7owjvd1F04CN7ImWslG3PY8RHnku1rxJ/uQTr3p6wnQO7X/xvD+7mHV7AkW
IFePRMocyhuUeE0ixxKkocTKNmfkSWCimaN2OG8OIKYq0m5LVytvjKy7kWVGY8SS
cWj2F1op/j6xjsrWo335yPqK2ek/Azdg0AzVrODR8+TWT9UAt4bilNS30xggmbYk
QpTrPdgP8EOMtata5sZ/h7J5Z60e67+Eil3l/txdnNj7cFXOpXnyBbVEvHAFbHGW
Z3XtutbE1/smQMwYx1rwgRcbAPqfyejPoBnrD5h8y/xID/Skdjwz/9BHAYPRnBke
RZwQL1uo8iOZbO9ou1lNTbiANTTPe9upVz4X1CsTNxToj7uqHLHEXbMxJ86H1Va4
BR1JJ1Ci6wsVLz3KJZN8PnKe7GDPT6IcTB1ncX9BYKEYIEsk4QeienBObdGWT/bZ
qQ8uL8CMoMG9+PbKlYf5wUErz8GsUrE9lczyLo9L60cYiERp4EpiUUxQv6o+ccWc
uCp9L/3HgS3VB63JUcOU0pKogMCU9BnNksd2YgxTD6OmqzUWgyyItsD7ouJ2bWwN
YBZ7LaD8S0HLq4b2ZK4YAthjQ37jB30viNYyJlbBJuC1qtEWcIFkKg/+hf4gobFA
0BeXDZa96JVgC9ZsqxYBbex0TXxQ/KhI6sJwPUlow5U/EyhekzDZ/R/5Vrd8qkgf
LiUF5cLblfOx/KpiF7aJkE/4ESHOnxBHAZa+I8F+LD8mxYjH3ezyAKKcZeJVLHY+
ds78323HllYBiO/LFP+L3E37Slus4oq4VXcQXPf9qzJ7pk8ltpyef4kfU939+CQb
yJApBrSTZAAdAKDPXja9dA7jmn8mqpbgo3F994ieL2q4PTAGBsKsnEDApQx+Wehn
lhSNBXwavho3OlAjz6m1RtXDhJkq2e+tqW92e3q2EAOh7XxhAdhNMHit4/koLFY6
w2Gq8kUV/AS+6gJMd807J7y25tFgSlxMYVNl5cKxcDnuL1ESufHN5VJiSnVqMUYp
ttQ8kdD2Jx9ugL/Fk3h3UXpLYxmM0QXiorF/1HxjrgBiWQOWLI93GpzJXgc2fjqF
lF9kHnSVJ+DK3RRXrdfV2CUWtMkgbf760KQUT+c0beDB0mdImKF9fmEhN9X/bnjz
Tl6UTURBpp408KXBVltvmwQck3d/mFokvghVzONYSFfEFIWx8R2zB3pp5F95Prd5
fXt+GkkqcrHYTybKhqSy1dZuCHCtm5G0jqsowhOwuBi5tUytD704EEpVVvJvIaUz
+q1him1YXGqvuZ45myHkUIGJ7T7/nUUefoTstGilAdNJpNx6tu2r8hyrq0dPeq13
hR7+DPS5OAJH3I8xwH0+m+69LmUIP7sUxRUgF764qut/NNV0LZxSv4u9QfWtsWxW
9bR/dX1a3vqlNB4soNGPfKKoH+9CxX3/51y6Dp5F+M/2V8Ba11NyD6f2MloJJYDK
Kf71NGCMtxGw+8+dyt6GsPjRVpvJv5XJ81IvHCftVb4dP7TLzJnwOC5bs6grrtq8
L2W5ESPCOUE29Rtbs4lBiyCAbzQQWqlVZ4R6yp6gy/sKS1nTr2fZHyn0Dy5a5y2I
zejpjQJJPx3hR43ubbzZUmzrdDwpLOo7Slq0WsUoHEbp/o3mGTcRsecLME6mvCn7
WO88cBh+8nSBabYSoVCei96usdYN2e0zEqRNwnYZ3q2pc6WenR6GtoPGBNPRJcTw
waEn2/4XieKwOZSBawWCyx/Q/i+Fwn7x/XMCJaEcyACR+BuQM223RrUxMMt0yWch
d8ptVAelrrT8Mu8MiEl81L/WDeZT74+4g5nXyzzC3CYkJ03jmaK4muEwL41WG5VY
hC5J3M0+VJPpcPpvomhEVTdVMjq31aSkZ18KEutn3RX03kG4FmGvDk5G8G//+D/e
FZPv3DSpSHfJ0A5tOvyu9+pmNGlC6oVUWoYAo8ggSdldPx/UBl0lKLnbbLTVc/Yh
GwysBnRN4+0ujgHcY6fQUKSzjC6fcuP7aF2kUpKXIdMD6rILqTo9PVRhmO2+emY1
VXj+HWgKtvc+/SDM9OHIVP3cIBloX83pU00Z+lobuNf58MgdbByC+EgqpJqnybre
Jw9O+7gxbyq1EPiNiWuLHSIXezQTc2wUhGVjWdrWrXRu4sWsC/A1DGa52K0JUr5C
5b0AyQCr0zOI5EMFidhGQa/YsWiiqUZ5KBUYlgDWZC53JYlLfSdm5XDWK44VRIRK
YAqClE3BKdEgOmlv9ll0SMCLh2sYjyYUjjj4s6o6DCRzEPgtpWK9zhl/TaTjxwPB
jC/pUE+2FfT+Yia3KxpxsrKCKdxuFEG5UtGQ4VwcN1iNG+rtQQXbsY86MslEKktB
eCSLyBRpfDljd/AGcOxScq+rxbHHO4fznM8QA4MJnWcTJEDQGZkDGyDwhxqHOXHx
eXlrsHvGvlrifjjrNIEwCz+/pcfHnYa5FXnJ8FpdPiBlxTD3nOLsMr+feEm6YRpO
3n5ePDYIv+rasqKDYbuHPNEQbW3z8xPjXuDz4diYX6JQHx+yQ5ANG2URg/m+8R84
/XdCNojnya+SjH84lEUYyBH5bDmhl4w+iZ97dL3hDnnt5/Ie/fHKWbJQUDX3nZtN
iB2vRAdtBHKlMkPvQxm2HrM17Huk4OhyA1w/HMkESh80kBVX+9S8gTaqyXQ7SGsZ
vhAAxbfWIlaHJeMSPU0rMzU4fL0bOfGOMNXAaBtzPX8fEdgk6Wx4lOfoxMoxkSEh
nwizjCdtzKg5DYNUerPTGGYMPjZrMnEzH8S+irqlJbb3T2uIk9/wAyHljo1rfKeB
BJnBAeks2y56wD2NwsM1dWniikmOja+TZeTBGwxdjuwrMslEFkTGTTCba2nQPC57
eoZntbLLgLKRaG9QozBr6cLL7+mY7EFiZUSvM0Y7bk2eSeWPX1ldFuNz3tSpi2xY
pzHG7f46wXDdfcBOxWehk0xSiHBWTVQQtVufcPgTrcVwPRI7puSdrGpz85lSnYfn
5oQVsHpjefRKTQm55gjgaPqCWf+b1Ceu8bJ5bGYVvRDfip5mMg4IjiwOGhbzCK2E
W+VixbC3yyfmNJtwRODq/MVcplPT4RtpHL5UI7ro0poBkFCrKPRs+FxnoQfQkBbs
fVnVwyJ1ygK9YQB6ALcIGD3n/jRO1sk0PQ21WFBP8K5wXLRcxShWtE8lzW8yIOop
3l0bjlp9L1MJNjvLAVlC72KxGDzrpWQfUWi9FrcUV2HLfo+hWqinyhmiuoEN+yfk
x/Rbd1ZwsF8VHX8TxGB8uL4Pun0Ss8fVZJMhvdFWtgcP44C/yBWgzhp8A00ZUKHA
uzXfV+JD3UTpMh56drVAFNn+cFBDEPu12997vfVRj+3oRBgDUUMYyBj5e2hxu8XH
wclqMy/pOTmiMtAi7zc+miEEamu8uwZQ77BvdBKQJXfCyh/YhU8MFDyZi4YSdRbF
bYHDdRRlMBWjHVX9nRjrKBr71eqzHVBaFlr+I5BTKe4AXrJMyLef8t6Zttyhcrgq
Yj60sY0oJPXL0I6zuEDItreGnDbxgcQgfO50bMOtvnlTdwQMim0ckr7d4EoqYu9g
fOu3VoFVtYKEEY1GYf6A9lM1FO4CU9qNcTFGHdie8wVrv8KNVDfvF9/zoFGvOcU/
ehX9IqttMjWEAiXM5gghOJMCrkIiueZ43VIFpBkI1FM1d9C5L2t5kFNEJPqrm65h
LdXOfiNA1ZHOCZi3V1C1Hz6aq9v7HLNBkhgY3oq5RBw7vnyt2N0lBk4f0ELXt8Qx
ZbhW4oWKJrN/e2nenwkVBnu0wlRve6mPrgsVRnoAcZt0FavA3Q3jl2eZ003834jR
aTyDPP6JbsuCSEpW6JMZ6YKw4GGI5YDvTxdXppIH56vExocsO49M81YoIGbn5MT4
fKWd+LjD4HCkSGXZKVFQzIoI19BOTR/PEN8BlzPGm34hnPCdavs3Z88qA6v0/NBY
Ik1KZA+uZZfz1HTMpRy9m1bivvJWp6/EqUAUxVB0/3NBUdQGQypwSplnF3bFPsGB
Fd6wRx7Nio1UBcrixPMUTDmEmb6zdRwO40u+wHlCkE3VwjCsutDeS6E1VadG7uay
jS+VA/paWvxX3kjRia8cCGONQ5paNtJ1ZoeDnpSGmM6DtYrR8Z7oYuyZ9fZw6eNV
ef6eczQfk0toSCyvYbSg/i71X1NOK+nPnnwUcLn7Dzpe3FLL1/zPwkosgUCOEj7Y
lbMm8VGT2dP1g5ORcW7RDFpJFhxAL7IvBbbfaJtIpaMxqtT48Sj1sPoWyVxrB6GV
FzJT0j/t+uwBaXcP3MZ7wPfR7zsO/Z4L1qG1/CyNlRN1L+Q7sETYWAHATbfPWw6s
lXuAuD041i3e2B9kEQ8JK9ICp7i85WgMEMcSksFsU35N1rQJwtcEmQZHe/xm+yV6
8B6uOyK4//EtWSqBXJk9TKmh9vtHG3lo+Z8tnITjG398GcEbrlvq+F9sYcvv0Ohs
26psRw4vJAMLPB0M1pelujIifxLbq5TGJsR27Ya0KywF1/1RzYa1WeP3q+HCSIkK
TDDOtzEXde/Fw18K7lWRRo3hHSvR/mDRuP2iDBIguesvxdGa5wxQoDdp0KYojyS+
DmT1ZAIALK+WqZG58AcA4Y6wUlUkWb/w0i59kT0v4TJ0IkpHfdEESTbuHAbWaoaB
o0jrruIhJRIxPbm54B0fj6WpgrGPIF4plSJbkyqOiGLFnlwKBpEAK+duLzMWxSXr
drnygK2+znF8PPixqog7lh1f/qhYpFCJTKlKY2VS3cMDxaPW7KcLiEX3B7N3CPvk
qthZdP3WUt8orhk3cI2TyeC4TtgwopHJ/jaHd+1PoCtRQhj+s9DBCCocfqSf2AOH
z10poDSbUE1LhDu530KcczR+OYGwtZHOF4ILEzD4oZni4yxDwsVITuVGuI551KJT
crJ05Cth9nqT7rrT/xdhN5gk4EkFNrJqciTbZkqjbUEzRy0fwAy3wzG73Exi1jOf
tv/cvUgmSEdsNaCz3s30hnHaIRiNX7+SyWbENA6shal/3ZOAOU9+9dhCZO8bfPdu
oEXdX9eEkVQzsRl/ClRC+LcG3qILvmW28B2eJTZzBOIMCD+61XSf7660v0Q821Qv
5xPGpVgwPjOvotP5LkULK5WWlrVOaCtlM4YqjCp7hv1CvLXXNu81zwj/m4VaOXMf
/ziAkVae56wPxX2KYiKAg9nDqepCnGiV5f1NguIyHYlEdlq7NEtNQcRvGwphHCSg
19JZY2KA3YxGgaawTEXhn+C83UvLbnik0CBFN3+mR605V0zy3m7fYutz/ZjfbdBm
BKOVxFkBDNX8uO6RHf1v8HV/iJtWLyxH+J4fBuuBMKqCV3Zr58RbUUWyPoT9QTak
LIp2S85jvdhxsOszBKo0aZUpOvuFnDpT+VsC+/NHSawTaPbmlEs5HYb3kEP99VYq
T1QK/kTLQT+SDh1TI6mVDxgDcOefShiB+U2L+2NyrO1t1ltz5RFmXbP3NymUjZ4J
0Y44dQYX8E/x1WIhXLT/ZmX3z1W3TQwN+5M6FkPcvs4wCUeaSEM+c/Qh1yehoKHg
PuikB/0ec3HQmbN425ZVkCrH2S5YzMv+31yMBvxkRr83R6H+Z0DfvbfocFjdSMTu
RaPoGH7aijXMa41zYA91HJmPWAx9UClkP2Zuv1jp8uwaCzV/axqV96F3gYoKXvMh
hE54Uw/RsocAy0U1IN9OWfj9MmjzXyaGqzRNiz+T3i/JskByo8CpZRtyngErJhO2
MHBgUGggHoDxvtVkPbb2qsebO8QgaOVEYc8MjR/hoa9/jVk7Pm8ejcHNWkul/CS3
Y0CCRp5jciADTSQRuLpLVVNu2Ds+PKWgOH6bR7aeX8HInSLa8y3wCP++smgRDil6
PEG1l7V5bF/ZN1gkWXRGyrr/YUS6VKDKVdFdldMlgYrW8AVzi28wPSTVI2vnWZlI
YtJZD62bXUzwkEStuBdSVwRUPyllCin+l1O2m9Y3VVr9cWV6BRiZz0j7Je06XZJn
neq6i7qv198H60BUnpynrMzYkQS8m/9+LbhssN+qXrirAEj+fBGzP1ORB8UmT8GX
Uuq2cMSJeRmG9odqz+ATneXT+hs4y6mAho4CGIkVkkVczNSM6hAuzZjUM24s7l6z
YI6PPgmeNv7G1B+3r8XokRE1mozSredlq9HOv2EQ0zHcai6NbGBzMb8lWW0WjCRY
JSksihjPnBdKmUuDabSi8MSWkb6wqfAJjgywYraTuL+u398UKPrML6mX1bidq5so
edp3MQs/RO2+eAkrLUWKp46jWw+jGARleZfbPYmSj8KfqcyTujq130n8oGW4bLoM
rtaw/6f5Uc0Yv1JO/zUJSDsEMBJ/hPoNc2PGSzyXWO0CdJkJMr7Nz4vOOW3dQrGh
B1Ke7kM5B6wrm4Lh/WDfMbihKZLaeLZ0b17gHuDHsOGnmH4YaTpJK/hafG04nCz1
uTxok26GTDpK0LMug9S1muoAMrQOq3EgfcS86dZn4oZxejjBSvgaeM2jAIXgZyXt
cwuOADurUH8iFd4gZUlOJA2gRpRcMepBHVs32I82FneioIpRdVQ8V5cdSovWWkbq
djnGUAfSfysFIhQFzE1lXhOO7MagnvXFs3/GKr8Nmp0nJNbBsa3qfG4QPZSx1j2g
teUTsCicc4T9PWdhWTGjl3W01D4vnpqW3zSjdw8vMAGxsP7lXZnToGubwZs7h59d
PzltJqHx3dtMSNbM80NWd+T2M//cWq1X5FX7C2s53DyssckQRCJn4e2ocWt69CoQ
l3xObQbGZGgSHeEqcw+eAAf5ytYlLN5hm7fzQ271pBDrVpcJ+fK1Rduf69IKrJ/x
Plgi8CTTXrawPXTaMy8FdQTRBHHwCCaSQH9/ZTL7BLt0Bn4pwhvTQeKH56AwIHxw
J5z4eqjJexsWl8yy8/vdqOHYdqQ1bLMlTi+6WWWEtSv1rff0Rw3IfcoVDL2lF/0r
T9gXaRN7JkAJbn4163dilO9cWOQxLsBotwpZThOW+XdfO8/HfGIlGFkyu0WF8dBQ
A7z5osvpeS1Vyi/mlxKs4k6ebXnx5PyK00gDbwmqFCceWb2yOmnBE5rzt3YnWjE3
BFzO615zKbRU9+uaET1vY4WY18X07pd4T7TMLFxLcNmP8djmWySY8SCwqmlxUHwC
7pxGRvrz5fH19EeUHfT4viKvWnjmJBjt/0SIMoy/wJKQNIzZ/aScL+g05Z/p7KSL
1QYX4CFMVHqPOZCdLlnUmnxsdD43QFfUcZuEDTgVjMchvbm67VqnxbvxZufUgQG1
2Wqmp3nm1U9crMoHy0fDU3YV/GCj3n7vkul8fjTA5FWSqRy4jMkmodU4XdxAUgOW
7rK3J/C/5PdSLkKboOqBLU7jq4cukZXcTvkuxYFgqDxF49xXaDyNwE4ZNewcwPvt
I5hwkmvzh3mrIk+TrHJMh3kBcQLLYwxkrewDhWhAWnph+CO41gyw6Z7AjVGMQqbs
EdSbL/2ufvI1kEdg1iLmCnqVhOj4bpsJ4VSPhhlze32iE9oWuITMIZcemHwO2z0M
QkyjXa69vRmGO+FD1GKr+XuZJvANoi+KRXFV6lURmw25/UWVFh5QuW4TcVtuX9zI
EckYDbL3c92IdKzhkV7Fa7iOpiAiG9R7jJH+CqBrnbDxAat/4h10V90DNv6A4E4z
pv50jj0X/OSNYI39NmZTW8l5qZPaqiiz68eyqvw61u03cRduUfxovSGfDE0oKvp/
Wr1jsFwF5ThKqOeW+nLRfThf6gEZRBRQHfwK906TvXG6JEXgG59PA9HvAp+Oasz0
tlyuaPLHvk6TZ/ZvunoM+0nPldXjIfNLSC9xLfUisJNsBYYISBpCAp9h/oiIr0R6
pYNNcKYQEVBOK65Wqvq363CvhBdJnBGirXuYptZHx2r6ZgKcrPlEbCC32qevP/pr
QXaWZVPN2qHuf8byz0dX6Un09cHyH1KDGFAztcoKjlH6ib7cxoNCkJHCRQpRPI9c
fJ/tlQ69f02ybrOgzIVAU/kq7XWJqZXhJLI8Jl9Y0ZphkTds08ydvyamEenMgx0x
HhtAiBCy0YMn8OaTBhlOMA/UbpijNfk2L/U7/mTUzdOmjNcNZiy3XPO2Fq5IG2g6
BefCTDBbZNJP+GZXW0oSsQwqYbb2KjqQEdaXIEZgDfSYpMS7dlUIvqHwz6GdA9/R
11wSBnVV+4Pg6n12loeYR81GhQpGvmeDCH5vg5+BoJzeGdHHkAKYj6aN6eQKlqpT
i8INqN7LGXGx8ZMmvMapfEp5odtrgARon1S5AI+JUVRpzw1YzlgfebVeyO/8uTz9
+nCBhp2dAghf+C0UMDZoag7kXPsTw5wRUsNlIKmBUNkRXM8j8EIpt8u/DEbaCNMp
dSGVY+Tz/IakGTrH5sYVGY6sAk01vRYtLRTzCRoyGnMc3Y1nP9vAG8M2iojQYxvR
dSsFT6GvqSooZQphdjTTgWIoC0uSozhMvvuBSdy3KvtTDHa4kRCqrnI052fv79Js
bqSr6xMXE+y55qWYIXEZu5s0mroCFnMhF6d957KfYY0gAip49m4NQYBQETmnkxZf
4k34IPBfFt7GDG/syqncdNE5bLOwtwssNVW9Rma3GeQfRIdiGY/zvUvb2UO9qioP
Vcf6mzRYRWnBLfO0Zg7z7tPNaKbLRqCMVHc3RZtIcpJrixLbHF+2vvqWzglBFdhF
QjqVemAsADVz25PIIctqwDEUZXmNcd5IgNhYB9WX0xlQY9D0KKaHsTbT41n3uYAb
OshSAT2aDKmp1CLF1PUSNwStcEtiVypTlQf2uFXfeNTD6AbQktg7wTx1lmJtxrA1
IrKPhNkhUGQBeyZluevNUDOctSmKkAl8jRER91TNvSBxXrNp0gmYlYVN9oFyg3OY
tsx2wKnCOKHSTiRscheLtZ1RVcz5SynnxZrf7CALEy+G3J4wIp/iJNWciGnQYBMv
AZys52FON+eZvCW12XijCNGxG2TbNm0y1XcWOKAd0gasdpuvkr3Ge70N4+YjoeSy
64c4xpm3Ag4M3uRyvqXEghMK/sy9AA8AXIzDBQfkx5GNgH6x1EcjPtieuJGkAHo/
JrjCmtziyDPzTQfaE/OYWT/7vZteLOyZAwgH3OQmxEjh1iHkaTl04qaH2GZFHF69
kBaU1YgX8JYPtQM8HdFkXU3/C0TtxP1jyH+q2jqCMhCC6JcBBtVYu2zR6+uUeg5F
NxPdZw3nFbxLtOYWqfplhaJZIJI/ZTNFcxm2PuaWAXZg2asHfSKoMLrW4pe9HhEl
DfdRTo2AZHd5D0vYxWE3dQatSDdCWAOoD3CEaE7Icl392fD48/jMhS/s4ODBe6hn
aUQf5Ame+SDZRYaBcUZxo+IpY+PHrw6XiRtSxIZjpOkFejJAOlykeXN5oSWcxRQh
Ajl3ZGkCtpEFdwnXTY8BvOJU86XAUI39hg61X5XRDb6fxGJ93pxgSMUm6roHiley
2Gt0NqW+APT/9DAGXSOELQyK8Kfz/jV8vh8Lvf9G0ykzuGlF/7D6wALbA0YPVkQt
4jGaGbVnJgWazQJAiQnaisRyouHojrP4K6hJ4JULYdm8jZ1XDdCCDFjpL1qlQDjH
GFY1d1tbfgXOOB/Ru4iuZBfW9F3KOH5ix4sY6itFoIYGODahhF60kfeLzyhBt1nl
EfKDXSlXm63UmqT2bF/e1iKYc34ywnMCZhNHmhW1gZU+7TwPhDbnxbyzGAvBrN6z
leDe/tGRdHrIryIImxT+DOe1nK349l/F7a+CmAxyEn8Fb5wGPT9JWGOOoytvVIRQ
frsvoRL5By1un7JRWIDynyS9QL1OnOkSjSljPBIhfRTI9ZHOeHExgbI8CFQvWVvh
EYqqJHnSYCmS/l6b/xnlqu6mO/UrbskTxoyhnd5RgPqnrwCF0DKvgnfmeYyA7YEm
Agn8DmVXzUtmdiQKE/0qzq/h7ITjIm42lz2SFr86SrwVHVsNdTe5sCdl7adQFBEZ
4vKxLToIH52bb5wO2+ACz38EnR36NQRbfS8X8WX0jWDulQMf3LT+nwpt0LDk8v8p
lQg2xe0H4vy+/m2tSTE1KBvHmr/3+UZLaFSrEzfC0tLfgfCuEhGDRgfaPBbGjsZl
cJu4HwhfCGdqhaVIP5/A6imE2wOfq5VXN1CdmbMsqV79L+k5OmfO0ouHNFaC/zk9
MDYxLtysLgvtkiMOgHew5rgLs4oIXwwwMuANPhUOUW+XhtUCvie738Sfw+/MxpH1
OrZ5vjEH3FbAZvrgEExO2ENe91pfFjjrbgkBDqzfZf8GVFyOUF4xuDuScsvQMUTL
t0hIYQ6eLcULy10uIwQGr52+uuM4pZxYi7SQTo+IIUFtwCjg4Z/mdw58sTMD7aN3
SeBxwwnpMvhfImuQpT43fPGIHU37dXoehsPVdhBXL5yssMI2PohgY+qIj97PIi+w
ret+xjoxZsqQb5Oj1HJbQEnZBSKmcUqa5qmAcTpYAr5+9H6FliUD74apThR4cLOG
19kxDfU94YDjDLqA4WAbtLa47H0EQXPPavGMMzsXz/lOcyqiqW0oChIYL1KjqP+l
XCyIAd/gVPMQgy06o4z7SvyPCSqjj16PWnXTsYjkQA5dv5h/OwyeA5audcmobdW6
x4RlEAzixGhHOj98ykMgxe6cDF2Yk3SZG7SHttvor2BI1Q37YKzaykSj1ObHVbrF
u9UlsyWeh+VQ65MO0Eb7CYQsDvhYa5wCTVcyvxgP4q3vOtXLZKDZkSTBnra9kILE
uLPEXqp2aMZlk25rqzTux39LX+FZ5Guu/F26JFVJFdQ/RrLu1y0QOVukQKEiYzxx
ZauHhDRfrlVhDy7TGblMZXINeoi0YvtdgOAHF/N+3iWdDTZ4nIMZ58WlLQYPbFRW
eEukZX/y4krWpmbjYKBUiycgzqJqO7WhtoHju1rxrhgAE0WOdU+43Zk0owZnw03O
owX/Xmv/9IMd06jddGzBM5/H6y56PtN9xxNuGBik5vy36FRGyVTAZvrh1OZAsxVG
bLaSpBEv1w6zxjeCqWc0Vd31iCAw5HvG17Y2Nfe0lxIZGq+jIT7Iz8wtMuXXmPln
ONeRWS5E2kD94JNGfjRtaHmpkLpZyBRgE9zOs0bkthvfajS9SeBs6CiczwJjCk3y
PbXmGNA5VQkuZgU8Vss0j+3BYcP4uun0y/8IHpthKt6MrRN7NlWrU9OvKy2tQL7d
N+BNtlpeWYncwmGXicLvQeWYkaf/JoMU6aARMF99Ex2DbHLW2JANVAt3kDn3vbsB
emwejiok2GBGFYcG3h/W4jmtEa23PwGNqhhNhp3JPY8EbWg2kwd5YhNQNVjFM11Z
groWOVXyKV80+tvbq2AlqWCNlnsRqZYqTl3iBhro58Hgp8LI05giaZNV0+FQeap1
4dBjwoBcupWSSBnQZ1g/OdKBbkmvriwSOH1ln8i2Le7EtHv+pAiGTPZsnXVlsjCF
fjBnZb//oiCIxIHWHaZa4H7ZHAM3R202pOk/gx05QXEV4PJONyko6m6Zpxp3AXo0
2zr/ANoTpP+H0CofOCeQVr6tHkLL4LOhy3nF2C1WxJ9zvgicVFFk16NkOIDexCyi
dcjtI6Q3qbDN9UBUc7KIE2UeFfLfb8DDHZyGbSI7xBM3YVZcij3kBXyxjn2ztP7S
g5riRIRhjldFyHGo5dbxp9dEz9Q3anCG06KX+0C7jz0CSZKnqDeKDjnGR4IXr71f
zSEWfYGebtcaEZyDohyj3iqsqeI1Xeefir1JHQ7Jmq7uaDw/qnnnBcW0yPvYIyyo
OH+orp0iXafcry7E7Fo/GGvp/6AkpN0PjRI7y21p0sGSInFBCZLHMpfI0O8gbKPu
mKvvcigZBE0fTU+xshp7521vNbMiOMzKiK9gOkxW2OzlBSeRz8uTyoOUiLgGlTRu
mjq0Y0qlfIX0QVNwGLAIwKLIkPEaq2oglTMJKzP8sFiKPlw2hchLb80cnv6Wmx/u
nYe3wd+DbNugHylAN5/sQwp36U81YPdcg+6MDOpXvEcfCVU9SdEAjohtD86+6l+0
mVcVs1vUPb1Up/nobCAHbUHaT23sNk3IaqebE9NHFd6QYxKsKsPISptgdZwZtsaF
PZ0jd3xewBDyjcbcTATm78bmL7nrcrZxfN2X3+ffqT1ar4zVBXzajfc/AxLRH2Q1
USI8PYg14hlZoUKkwQ13D5GPNEmzjWBl8O2V3FvramDJT39/hq5Kf7EYpJ629cs7
avUP3k9TpI0DfkPJbf3pnNZwig/Lby+umX7ajaA/OVSBn4lRcv9twz0DMfxgSDN3
xN2Mu/tN4nZ91IvWunu/77HQR+yKZOk+CZoE0O42rzofiBKufXBJnZ0CHxns0zDw
3N/BFQhxxR4uxeDoVLHZH1+mAApKbQg++tDbb1vt4gky722GxlOBgUENfQNG2sVE
i8iqMWJFFPyEg3FAKK5/a/i9fzzPQgl07DINeFM1sSUWtqoLnwOTjtsEiYb82CFj
CD2Ep0KEJP5XCO6MYykq2mZralbxLBBdghZZDo9nAbz1VAKqvxVTIjH9I1LDM9JP
dt7LcqeYDrqpbpaRK2fARIrXo8lqqeTXc+Y0TbHcr8OWtKLL8/DXfpVQydXIXyYY
E/TlyCyCoLsezRe610ztMBl9d2b2hkK5QQ7gGb/xfD7DFwRYp+rhzPr29j5moNz0
nUdvbtx54oqfLCpThPL3QMgTsA2wcBIqaGlJpkE5Cznch3CCug/hJZ06yyt15a8n
LCKJ5hxmfK4yS8iTwtb1uhRhp8UgWNA/n9AIDqyu/cEQfw5pwjlp+VwBHJu67VpD
fHFoY+unjr7HuS+VGb6E8dxFmAvf+QcvtwK67w5uDN+7753cujOYCIjjSba5lv4L
NjyfbyTWXNc0fNfObu7yYd+RTTorKO/AlCrd2+H6gJoA6EiV4mPcAgJpfPUA9jBh
HiR13R+iJbsSv9AqKAVXvqUH46pFmyIMMgzJVgA7sqyZ9Y/uPca+EhomzHVwBhCy
MLOUa49Ptwm/oM0N8MUA471jtwR1XhXpU1iUWEqz5WFCBy7yetlY4ejXVdKOt8bw
LGXjOqTb6EJvCVl9AjM92eRPk2SPxTmKKXy01m6IN3rZf95LjKWFAZCulJ42Stfu
VXh6hY8LxihoXutQTGIlDpNeH9qdoPlQsUTbI4Yyr2aMpSivgscs1J0UQo64oRrk
805PpchYulW3P2r7WgJzVXiEQgLDmyjvWKu+CEp9J9HD9DqWi6aHCqBpUq/nitor
CDSuukiBas+RnWJKGVqRFyS93gLXkxp7tpwuMtfB1NUSTqWc8v8T0YyKSNzm7zQk
tkY2/uFZYnRjNxTElnam0IiNf4LcpKjnNlbVMVMWnRmhe/Uue6ii6NHmkUUPXtb7
pcM0mT3Z5HHiP5OZMWSZDwlEz86nhPOpucIC7PdvkPIq0X0IzIDHwVlx1VOplUEl
bkWG1KRqHwxmrisjyX8ZB3KwtI5G6cJ3f8v4/iaWtvFcT72h4QajYS59tpEAkMNO
aM6jPh8r/P54nrI2NWMu/AJ3RStt3Pb9C5WsQupBeIebgBs4ByP80B5w9ukT1YyE
iD4eIWJdnIiwepiO6eM/Tc6Au4FqxeXKNclaex2Qp+YKAttvS678wPg0KLJH+rU4
nALsx7HuO/ZohU2/bOg4fvBGORBDGSVC+ZrclabkCw35v7MmJLcgeNF5BFdb+163
zn24L/Ey/+gwXP8pzcX0mlx88T8AG3fuqYYpKLAH4qhtSBRLeGQ+qRc5kbsUoflN
mA7zktHoDynGpbV1hw56TMtQraiD3p1UysJk4/WXpIZcsrih3a7JBJD/fjGoz7FM
rxTmfknihMywYJXPUUURFGy+qcZ4EBLD035mFVx7g527OeSeIuoUWwmbUHb8fmvV
a/cLp2Dz8L5ETVPp2Kq5eBQc3Mkb60VsuaPZbyuICzj+s0PqUJJphdYdR+8EQn/R
x8scniT82NiERKk/lbGHsOoxMYMZEdpF95RyFlV5rJAeHwFnUlgmSwGNApy67TUl
yCpBk5PBBQtJiGeg0vWuKBXKLcfXnjrnicGfSRv1Gbm+DSmlZe/pl9rAexfmm542
dkBtnoFRLI7NhhCaPOAPlkj85TJ2tpO2nLjpD4Vkka0IEdXOkt8S/N29nGZmPj3b
zM9GImFVEy6SbYalzhWyNo9neR8pCs6AEXmUr8tn2tiVYz6pWzk3M3KXFqZv6CLz
oMQE0aceysQev7DjMJA+eXVylShq01+Mvrrnwc1IBudryxvdr7BmXk7OGFfV6xl7
tX1zvDNwC6cl6W3VJhfuBm7jh+P/L4vI3ABte1FMHmHoNtkMOggX+N93I0RMiRqK
hvY7eyNw6h2TSJmlxWb2tFIiBdbQ/dDKAT4n/zi7iRr9DzW+16Gv1N1Qcu61vemX
op21VoQ9WMvgaO5aj/SUvZiot/Ues9eVql3bQB32wSOGYuGmjg6MIQ4H/5xnVNyL
bo9B0rD4Z8NDSBTBJk4BovtJrBqh1eH/LEOHdTTXO28vAp/OaEjgGQkc3k4zUdKM
TL/dWzVMaryU/kFR4TJPefw2emfwUEnGGyWqMXfLUxXxoRb97yA3/QnMrYD+tZOx
8bH8uyZ/0/bDgrPAkdeC0hJK0TmAQ0OBmT1qOkXfhBHP77EX+KO2vNK7o3+qQoKc
qlifVHKHUTVf7vUdz+f0dS9WSFX4STiN/ZSQwz7dUvdXRWBCwq22I3uPSssspaT1
DMZlrnQ2Yp2X2cYNdQfSIGrOMJGz+Oh6jINeERc2guzYDsodRgmTb2nLVB0y5gML
nwFOgbgDOkOzd38Ar/Cd7z+TXj10Qe6RxoBhlfGc4BKbkUXJGi8PW3S08z2z+pfs
DDw/U2Zwl+r3cot9aEfc5hwiVGF8+5kSn8qK5eR6U2kJDfeRxg4eRXuCVR5pEOcP
DBPZBZ1uQReILNoxg2i/UPxWsT3Kkb/S2Vqn0E8p3CAxUhsGbkSy1cl4hmkg05px
Y8D2MKjyah63oIlL2P4rqPqH2z2zqyreoZJNfN3S0vFrRCo9kMJcECUi1lPxHL3k
E3697YKDj6AS8Zav+A1Y0VDlealXnn1kEDiyBtYJAgZsz+RY0E/iE8XfzAH1TSot
MTMRKRY7/b5KLTAHjGXpVM8ToNas+byY3FBRDpZyRZf/CKCKt6juJnL4A36mWCFn
FWlNShMcQ/sXdRKOwk8Nq35ZKf86YWOe4Bm0JZNqunnJzI4HdsW7zID3LWRO9jl4
wBJHE8V//NZyqETklACU4J8zZLglMtZyCo6FNFFqXMQ3n0Sv78yn68D8rReAh3vX
k1hWlEH6sNjp+1Q4pRUq4en5lESrLPaHsuKvwx9S4Ik7TjvEW2p2JnkJlLTYBUj+
DIvdpJDAUhxx4uyqDxie0GKiAGljA/puLpJI2LQ/iOHgFz+TN4ko9m6HRdOaTJWJ
rV3Y3zO4DHSow/5JFbCe3YMFyQCgKoVlCh4+AUw3qvvIeohcQmtl/4awX9FCNSuW
e0NlJkSgYuxEtISxvyZOLC3rzLuaTErsNFdEKGvikp/LXYTjVIxef2/M50nlGAyN
FFV1VXQgw2/wtYST3hF8vtTnnOVVMWyjjk6RffPnwHnt+Jisv/ppV1dqmD4rEFEo
S+JRTnnoRSpCiCMtAsVxaXRYFbp7zqlnjj7Wv5BialUqU+HiEBxxJ4GeKM44jELj
4vMl000YfAG+LT7ivjA+Y/RIu8I0TJUlncc/xAuxP5OsAaRY/LNhxRay2d38B7tb
m7wWynarXNDHjgNwEwdqka4g8B6eVQme3aWbZv0MwDnZcBNbaByFOPMnRbskOMFL
+juWqMr+qY/7AOV4XeHNoTXW+Pc4NRlvZjA8QIkmxSnZYDlISOf7Xsz4VBWX/wGY
UShqvvAiIrlZdb3KAR31tiTONCvRupI3D5thyelAzpHFCa9nhJFeKmGAjpHa/xeu
VyuaM2Qy/tdaf/Gmxl3OjOrUrAxKYLCz4PiW5NsjzMaXquKQ3qtpzgT+7itZLgML
wOe3XGkLOUrYDw4Gjo3T1X2r8k+bNZ8GjeDOV4OxFU7slIPxM9pFV/YdTbx1bgFf
8JoiF4LNAjSbDoWwWpEyNfntUQavyXinTie62le2za+CTB3O81MkUJ+ifrMihCY/
gzfd9eIEwDru4Vy6mpSla0zBr1p43Nq6ybyvfy5hNhHZPuojpA3fXcd/dPQcDdx1
rjz54GNsttkCz8fm/I794R9MOy0cOak+QHfQFmbkF9bB5eaqHLM9H05C8mux46Y1
mGd9QfAe4JPpQ5cGVXduCWB7lyufawuhDizWjcVq9/Sog7fYeI3otlfF6qjKjP2o
nreW+z4PPkIJ6AdCu+9Am64Khtuc+MActV53D5j/LshCYNIWeejWKLeMKTwwTOdR
BogwW8Gq8rYTphKNXwrb6Acuze7EhWo1DiwTul1D1m5fvR1DRj5IjY/D2xXDe5La
8jT/2jcq7qg4r/h/vvbw8nJ23XVC5u6K29UrTeVUqqzsY9NL8zHM5Fmr1I0pNEu4
/mC7gisBAsZLwRUDGv6UZS0y/ix3Wk9vJcTpBY7FJ0idkJlrZUIw7nz/UymVThAc
ZfRUBYAM/r+GVt7REQFiNrdCj0/n+MzSM18XF3Ftzi2v2ScAAR2OQ+EBbLXmj9eO
rVTxH0FTVoavgq+Ky/pQhSV7twURqcMMyKX1lagIb1XE6ONHnqxd4t3ePgQxcFxT
pGjPa6o0gzOYWPrTnYQm/yuGF9jCb/TfiHm3HQ+N+5XvTUbaHfLO8ba3Ni5uJg3A
ACjRpJFHaR3wzZDV46RBWU4JG9mMbAPasF2U2Migsib5daDyNYaa/0imsyYVl4aT
wIXcfQ56D9nfluRlBJM/BxqC9cnLFLGeT6zZqfpYaQB2H9DNZvLYhivMgAIPq4L8
Pn3HZhpfSsaK+2ZZaRfyauDr0ODQZdRZRksQ5pigqIdtBUee3Qr77t8X1Nw5eqE3
gQIBiiMnMd0hWoihkW6/R8UClnt/i+OGyYTzae3BZK3cRFbBO+tiWAds9XdnHmUq
iRtkYZLjV8VaJomoeHPZxqpY2d1o6U9N2joA+gDyWQ9mq69lzfi6xvSuPDec8Con
VdIbMKnvqCSITdTlMPhXM2h8WsSRmGYvmjrhwv0EInPONDNoJVngxhLZI8nkOSjs
k8V/cCPKeOi5B/4sZ2TmhNvcpAthmOv+6DbFudr2Zt44NUZIx15bAKmhOsw2PMpe
Yo3NWwn3lLm8tqLv6XCFdm9PJFEQxnVxzHdyZ8tqFoFE8ewnurLDAFOpvdkFTcFc
MVJMiF8bOZ9xdAC8wY5SdZu6y/kEJLGNuCza82yU0Y5qiZMReHttK24k8sEyINpd
FlJVntiwYoRNeLWMctS5wTrAyFSI2bud1TKRlDiiLWx0OJp43N5ieCj00KspAG7S
a6/sadg+6uwxPOvvUQdiSJhtZpfhNwqpMCyCQlrc8yidoY+Qv6RJ/0vR0yCs6ycG
IuT/P5C0/GjNqn+kJ1mJ0yXMFSuk0tGrqXvGBo2WVfRrAjEmigX0YtHHV/KDvM1K
XqoCDAvfUyxPL8exRBXqtHCnuuLWwF2VupZaY+aQEnSuozFIkK7Rs8CKT1slLCIu
pW162MmsVddVdO1YhpWXsxt3l1l5KQHeQCtbWhMXR7hWNRsXMDbgMoYnvANkgvmC
7todx4XVjwWZSTmHq8dwlIxFYUBjnQ+OJ/NX1i+8sH64pn563/MeSEtgP36i+2ap
eSkCJgHPKEjEzHZTU3/t1XledG4qrZn8a7KfmFfbv1SgkN+uMihD6KwY2gX9Ywpz
kOC1x8zXBNiu942aKdTjMf0s8PE4F+lO4IJSC75r+BResDBGLF2JoRDACI0096To
f6ogwxiUgGvj/9T35KGxJkhSAYMRWzC8Fw77IqXlL3Cgr2ZJaepepywQ3vZaVN6X
9ZisXpUIdMev/PVG2YpzHS+pXUOYfE2Wfx/nQbCQuMqDKyUhu4B7gXYmB/jICVqP
247UXtD14U7fD3WoSoNO2d1O8DPQvr3osxYS4lFMpuYll88mGlvx2nAxqbBystis
eZJqrEKmdeLsFOxL6sA7DTN0l1J3AZ1thqYfxIXU0zaVM0fzaafQ+5Rnd4oCNIFf
/8zkYmc4DtNQe01/KgQZC/94AhWYaQZXL7qz6natxzeGqdXdF9E12le6+o6mKdG8
RVtnSu2AJoCsjLaScOPZWKfHHzJegIfLCqXO1TnC41s0B12bgdwPGko3cTFcSjeM
BC0fleMadmvNuoTIKAs11UTFXcBC3uV3j6d3OvgFE6aBWODmO1gbCuQ6SuahKU/3
MITF5sWU9vIrRYlhHmBeji78TWHk5gdcdOBmCxwbdLNOLFgUEloWIoD1OnMfpfnN
Klrg2DSPTzKm+H2SLbqyCvdzkLOYClqIcu8ZeBxztiO6XGo+6N5VDw6/5JTpFC9o
Q9zQo7+nNsDje3epl77GcIwc8n83Rspi144D9pXS9mkcNHKdU+6AjXj81Uj+iCTW
s2W2D+5moAsVowMphLcavfDWhVQsBz8Z9vaVcpnrI42xeHjVwo/xc9/Nj14CxavQ
6khc1Ts6NO6FmNSiw7CqkAQV/BfN20QIBs0QHh3FonXJvCRNWlwPKq1B8Rx2pOav
XH5y3BzD7HDMFXPhwxMvUDdyKhZXJKFwlkG4uJAZTAaYv9ZeXBI90hos/8J4o2NC
6xUA+bqcmnwriAvy2kd565dfND9/voP3W2bHaMXXRvFGU82E2rfZa6iCuxFmFo2O
Xw4GOivGt3qz4PHHBnfWUhnwnfQy8xEAazRt8kSdMn1ejCPl0zxIDQ5YHjB1Vfh3
VqN/aTDc2whHajBHQ4iCzDPYuU1MP7HX8Qd8Ytye8IoOzIUR8WV4EcRoFqS3WsCn
XxgNNXm5vkE2YwSo308An9QV7RBlVbmevvhCCwGICQ7iA65cRjr+D467KRwjhxXF
30k/tvmCWL5AxGGdvF3yWsEMuAO+cIsPNNKQ4mwbePZq6oWzUKzj3SCdbLK28D0s
dHNVVYXNE1PB0GQtzu7NiM0Gbu/CySkhqW/JfeB9N0rgCIJa+JGyG+2YyvZPWs3h
O3IukrdizlA6T4/TDr1REhcMBFrlgMorUfmQxVZPakyCkPZRz/ltaagaTWpYlODt
GXHp/ucxEXkTBTAjXFrMAZichaCJPNUQt9hE/e426r64emtNX8AFdTmSZUiWTwAA
AZmtxlrqrby4U9HlbasEFpuqbUuq430tCEg+dbHStEAX0pvrkefLZ5TjEyaBwV3a
nzyZlONpakj4N8iEOqFCp2rP/OcnNThG8sleZwxGGx91uv7QSvcfySXBsA4VKivM
UyzAdc5KgzBcyh1mAf5SAKSPGR28gSQpS6rvUCZU9bgYQuo8tbG2BIG4uOCuqAqY
x19fmIImofWDh0LEcyqawR0SM64uBvhvYC5d5WAHRIo2/mIwFhxPFfRxGMR0xkbZ
p/WLtcERTFRaLpgJSi7birkMnTnwb3h3d0khpse/cJujCYqrhnUY+xdcnlN4Fun3
lXfKOp4xbylJAgCrTD3uPXScsBDhgv7hztvdUyS6xIeyf/CthO0WVvEN+p1/dx/n
DMIV43vumM8AL5curUt+71arSeIZHWFw+GdIkN7Pt9YUgU/IGGNj8aQAgvet1bho
ZmE7zegUQ/jlS0kuNn4K78Yrs2qTrxRFYADehgVKuSK1ZeiBaI3WXwIEJg1Eo6VT
aRVKMfXM/HzvayXkMkRngFA3WXk+beh4bhErHhVeqLlhHjl2B+XPW4OPDCcCxkcT
2sdEle5xfU716DqAzRqkOFX1pX8fwivvZd7exN0mI2Ec2ImMCv4ceQyvTB7V6A9i
RU1VS4Qfk7xChAG+tfohHAZl1Z+lxna97jHsfPvFOgf1r5L0kAC0uMBU2Jgp4KNC
UxgN323DedL913wPiBSk5aDE2NO/firExXT7o+10VLYhJizc8g4bgf1qPINtrWXE
l9eGxrIYnMce7IYeXJvp86FyFh3cwMTJAhRtqKJt7gXi/Ac/nPQCUuJwOL3pjpms
cWmFxGIW4A9FP2fXcpHfjKETTn8L5Al/wlmPSbhnRmmD/+JuIJaDTRzofjFfusX8
0TrCJ7ASxmkkmx1RDtr8qHcfYyTGqBelDskg/UpljHYJk7ecEj7fluonBhy3hKqk
+bYfjGzekbi9W9xFe7GfCELRJvrPnOMSBc+1N/5Ycv/otIY3TLeskYJ93Lpnq36O
B14oCNL/6S6gMkdFEpFBuuCg05qkCWad37dx4Bmyo8SrPpe8g/ikVrSSyu1yjvSH
Q3eCtNoJdbPUjIUNEIaHzAoigepjqmPzRpQvpc1JCj476h/By10Oy9e/96mNcQuN
H41zyVuLXXnDRZYS/whXw3KCgd2jp0XaXWL07/XEoepONo1vdAqXSNskjzCPUzOa
Oua+VqknVdCE/P8PD2VpciLPabtZ/TNHBBUhDrdqNB2CTf80VR4K5zum1zlbdZTS
uZnjOomhFAPIhftkXmjsMLjWamk6Pk8wJTEgx2Fie9JLbxVaSlWfPvCjEWBx2blu
EoNa/6oE36FHLFvDChmWn++CqIkaKzV1KNCOp69C5du3/tXoPQfLeHSVNrrIczpy
ettXvf4I78/6DKTuGwb/eWX0CvLz1t8aSMOTEW7uVOoMMC8E6Bbdy793aEGgLpIR
2pPwZTtBnlRYaKZHHndsHMtOiihgoYABwysG2Y7Ba0xlv42ECFXArzz97YDQ1nJe
mmBR2JlXLGo6zhHkRbDJndLp4dW8W1CvL5Dz7FK6YH/OWk+qah1lKxHWYexksIXG
5kQV19EtVuRjQZQrPqwE2Uxo1X1F6gCiU0oDjicPoGnYy5rc/sZ5mPbs9c5lJAN8
sBA8s3AEDzlIQ4umaOFqOJKzf1MImeX3lfgdTgt4iBONeKWh6I3ixUfowWm4lUsa
We1Ivl3KRQ11SDcHNlM9pmn7V1sGtrp1xFlyusyOFXXZ3emPyansWOPz1qGJt0AV
f+bdcITpolZ9DeTFbxfIS+hZbkH+6QdJDrPiVjjyoUjyKHIqgQm36DhA3AYJpc31
F/dmaB3ZinXYZY2HuWwVj2c1/myuB3ujACl/nibeqqNh7PSCp+o/ZxrrMu0Nmv2N
V4rK2ba5vKThZdmd1ffHsxC3Fc/4KO1JiP5zXwrdWoLGgwkwwB62UBl2azOL69Q8
zpJAO2TBkWPGzHDrYcX6Ol5kun49oUiU7LODjEhkv1a7dM6fuU5mMACvptLFUkDL
S30Fb8U1j3OoLmNhs1HPmZWOlOJ87rgfrxx8vdOyBBtuqEfCIIW/EpXJ7D5Z9ana
FkpoESpvRcQLpSYvrvwuUD+PV+v1Qy/OfTe7JuXBOTnwlU7W4JpHEmRdqo4PjfNI
+3QABiVPt/YZMJPX4vBaqyz2TfrIL06gDnTANBlmCjO2vuYzs/xbW4rhlzI8KN99
QK0nwFefieGuKZSCBjQGNGFGhVYacdS7w5R8jZmNqoSaJwT1jZGBGr4vuEvbZUYg
DMX+qrrgSnf1BGs5kSMcUcKaIR9G0b47n+zeBzsKFvAvGfgJzgiVpgIvaejvJF57
BMg8p+LKuUamm1J0oM1cv68HlIsJspfC/Rhgi8ob/J+KvPSh4PaaNpYO5y9YTUai
UbjqfE4SxzFELY9D/691XyzbuO5hnBI+6reaWAjhtkmgG10/qjYSw6bTcuzeF2rq
t3fSyZeKSnKGRSrmLgNW3NQbqTqgtgNoFrz726r3v9njnXPXn14XYEbxSCMABvM/
/K37jK3pkRHHNobdonow8kNIEdLzqTmpaAz/Z+jnGZR8j86NNXlAygTkGmlIHKg8
QixXP++iF4bdjxcmJgEvc2uNzxbSpLud/MPMi+g1vQe7Alh7+XaApnSWw5lsBFxn
XqCa9NQ3/9me4Tw4tdLM1+ovrd6hS4JwNL5GlnVarm2y6YO9znYv7pvzKryP+RIG
Nhp0gTo7jMsxenfSPvWztlqvneOIjFUcNTNA7ZgGKZvsAK3pQ1RFd51KsYkme+uk
yvk95CVldYTT61reda4diw8c4p68m7MmPOT8EldmhAspzzq7+YgGDMzs6rbUBKVW
plLSf+twoVlJ42tZe2WiT+le8crRKpoiOoGR+gLsA7wEAqJyMo511VrE8ygaCq/H
0AxLegWxfgHVRdzURTiuODpGbGDV1ERt1VL6mRF1mIsqisdfoqP4Ii8kSij/f3w1
hyj1Gks/kINwbXZh9kRYbMtYKL2SFrXMBC7vl/JMiC3aGIczc9JPV5kgf5NzDn/U
hkn+8stKZGsRGjewVrLmccizFII4BlD93E4L10aVlazrIqwtuy0y/XZZzGTjBcFN
Eu8+UCxQQWEdkoAFZDe/3VSqwBHXa0jb3qCAiFvtMC3fX12KYYCRJ436VhMTc/Wp
6f5ZYvQdots7uKAJtN4L7e9NMHilX3fZUiVoE5swJmBTt6JMN1KYkP8zROGVsCso
GBCbLfTh+LojALpfo0TblqDxM7higm1hmgXRHFVyNXldkcWRGU/qQE54rW0U+vJg
+SVJXzVlw/U34SDlBvLXhJ+ByZbCWcKfZjxfx/liObrt/35qy4z0e2ql1jBlsjbo
ADFLHUic9srk9V7aY3WE9zQDxTJgOjTSnOT0Orclhs4S22khBXl8skzrDfz3/fIu
UF3feA7mMhglZcHChCYUfYT6YBoRphaBl+rkkn487r2U6XXboscy0P1Pmo1RfFi3
bvDJfD+w9zEk+MX+H8KL9ffLAj7gz/wrUlIe91+0CH0gZUJYA4m71Bj0CRHEXU8A
5OJpVZsBXCFWdJ8I6GQO4CHIJrDFqwPKcnpCoC2aAGsxQmDsgdaQJv9jXn4sR773
EbD2gt/Fnr/M/jUYAv8K9D+7IFx5vjI57bvMj0rlTdn34KpLtATKDibR8gfXyhwt
Dejx9gGY3ly7yvw9KZFKzkMEWOxuDoQJk9AafoMbEcikqQM6EmItgpSTdJrdNsx5
sVEQKtDQZmEtQOLS/WeoEzzojJmuu+6x6z5aWZgJO730lBstDA+7FByvnE/AO0Su
1W6Hn789eZqun4gBC23as5uD5aL5vUuh+412AqRyjFafyQcPudNkrzrBvOdcT/nz
dBBCS0ZIv4xiy8/gx8eMkZts23OXTyFIT6WVConAxN6QMa4Icl9aA1R0uVb0cCLA
lPMAICb+vqPGnQr1XimCjTg2dOUWrFb7KMGoq27gZp6BNHWh54Je9VlH1bcGhlMZ
gbeNm+nAxm/5LqWfrqI7aCUhHClk+mHWvE9+u1+mp2Yifgs5HvJfhu2CSZuV64N/
54mLaYZvhhzjGpuCy4uhEecLodTlZKZho8hj970Zf6gT4jheT/FJVzuSzY3HYj2B
+NaXK0h2+14QFBZvS+quUvraiuGYzQS11XgPya6qZ+niCulgGaipB2miPkY88p1F
3rzJgtrQVpVrYfmicXW2NcEMMQC0Epdkf2KxAg7kDiSdesXlaxOTbON4ddPcHxho
1IRe+0LRQqEHcORSiSZG19ol1TKttKMU3u928xWw5hd3I0o5I5c4XwhN6YzJx9cK
m4+m3VDztkGmbsaNMorKlXQvjm7a8JJ/mpX9L+LBQbyXCmGNZIiOxfSERFE7Zp+Q
FZSYzmkS4APn4AkiNlF96A6gyPztqfBpNLfXNeicvcSHeV7Pg+Nddx6nEgvCF7Cf
QU4j+ypcteEHaWNyIWRGzBLukeSXHYcZksqazlLXwztXJ2aJJZahrACyk6zasubT
E1hv0CRrKmgBhiU9Vo7GRIYph9CA/JwA7pnY30INvRKy+pxpRlLvsIO/PPB7AzrY
ryyw4Y7IJfRWKX+8kgEWGstSYT6ma2riOzzWZpf+rB5DfX7aL1skfA/6N4YFl4aw
M1HYHjKvPdIkQvnsbKXcnPNc2CrXmQI7EppAhGIBTO+QugkTZax6hb5C6jXkcs/0
2OXeS8tfJXGdBlhRqXU/Rj+255lDoatk+1M5iUoh28T3JMSF8F+ydq4zswrR9qFW
QFWuric4OZCU38wVa+fTFyqufAZvhOr8OQc44TZ+nVSQ6cS713ru5ZgOsLvOgHWF
jwOIEYWA4ISq+eHXv9FyWBc5B2d8LKhEDn1FplHzQjCSpcWjdV9tLuhcSF++mXkR
DRKiPyew+1xutnvJTdWV0iaCq19xqDkWVSYED9T4MuY/j/vYWF41nroJhxJB9MY4
WSHu4KQWDD5f04Byen8iKkYUCP/5QTt1UZmWPXyQoTe+maC/lGpuu5rK9hKeZ5yw
LamGzoh4h1NsJbjXjN6pVahpUMq/g9P7+XnqFGzRsQ8Lem6QUfwgUfnZsgJGPeaW
GN5pmEM81yDKLa9Oio4RMjWyfqqsOKJ+3rIbnD5Zr//pNveMuIM8Jy9KzFr2oHb9
aiTm8BHxLbiR//upeKpkPKyztBrzLKtnefJH4bitE3bS9ewHsHRNrL6EinjKbW6k
7/QtZcA4SvGdiFSD+b0WahVJvMj2ctYtkDkty4Y9QHZWhME6wkYqWjyUH4H7yPB3
mWx90iu61k52/Sj8bb4HTy4x5dK4WO9rJthBjBl0Jv67S3xFY01gwQABJMnMSPbl
4GZOQ1lcsPDlZPGGyN7iD94P9pcgGbr1SuQ+sBXc4EJDZrn06924UUO79VgYWrPa
xke10jBlkVgJB+jg0VeVLFJmuMPfe4FN9tfR8eZEaKoM7PJZtu1zQpFOp7EcM/Ao
DQlTloVaYPN6VQeHRwUqgaWbCZp6sD+ySVtxcS+9M2w5RRvCbGRjgb7NkClSCmVl
+uMa4udfTZ0MeQzTxFZr8frl//iR1txEEJ/NXs7vrfhuf+HTqsLDjy5KBob1ZvkM
1dKxbHwSO7ra3XQsXKhVue2jqWu2UZp6/jSkp/381U40N0dl/KRNlvmOwkmi4J2F
xgR0WoJe0gMymzr68gXN/j/9VXZCv5IuMjKZOvKKrE1mseIe7j78UjlaGaJ6ktO7
tFb1RoqrZUzI8JTvmbKC14549LmH6UZundYLzEL/GKOiO6HzK1xnaWCzI+jo6tBN
nL1jluKjyHWY8GvP4v0pGj5SLiBBOZ9rE8u5ZIHfr9WXo36OirPu6wn037OdXzw1
YokdVT2m8kmEsFRbDaCyVpBn2zzhXYoMntgjwVpZo+ns3g/vUTI0agjqwSMnUkN2
xV+ZYZ5tVjS45UNvY2ghKTTd0KPWiYnSZwutJ5wktmWXYEMua8e0+8rvgPWPANrZ
McdR0JbYtV7L26bXqges/gWgTCooWh7LDidvgH1orFSAo2q6oW5SSNrJowKeZlWa
BSiivG6i7zAWrKu5bpzq40yGaDOOFK8ZYXx8uGZKgW5QHszmlTZyz4HpmnDL4Gt5
E9Q3OdIdVf8ViliWnZdDXuN111nljU3uzf1ZUNAwyN+XltdAn5OWf35ibDv+ik6+
AbcmtC8jQe7MVTCv1hv5HRFXL2IaxQ6NG4L33ouRDOquHKGhGR/Ux7dJtWguNImA
nFNxHldrwc/yXrU+ofKyVb2Yu93cZg/PjC3oS/J5T6nM2F06ijBu9XKqmhCvR9oe
fVq6QQRwDYAl7Yzmj1utqf2P5T+WDaopLLOrab64z7InlVGNiD4tDi5OBE8dFIIG
5m90Ap+O/abR/wJGmLUDuUOWxZ/lTdFa+mXWdS29GcECvUMOr3Xn/aKLE0Jg8MXa
3AOLM7aSLogXqSxh/JOFy87xBlYd7C8UqQE7O0z/XPUmZJim3vK7jPUvdqNggLcE
8qECNe/djOn9MQ1wOP8cnqmXtwv7ymYQfX9+C7Y4tH0rxkjlnEtwKKo3uNH12w4p
JQdqLU/kJ75S2N7UWeig73bgRMax5cVtFhxYnazsJuzCV8mV2oIPrZL6end6eAqY
PBkdRuVUMpb3PFj1tB2mdLNjZxWfZYsnemx9uT1BHYHAQ3zRq4lssVXp6L+x3w6H
TLNDIJvpFIRXGA/4iI8s7LfQSUr03ft07kDHQQvqI8plXArje7yK5eP/9PCpAx6X
I2X05drFpqA7iSRipejH6l68vBtTDrv09bsUua1ZZ1nIpLavR8Z9BvicdvPCmpuA
e8aegzp0dgthYVumdnFnUaP1imwAh6bpNCbQhRLHGR83AWruBNUPbeLv6NrQQaHi
xB59+ZhGZgSEx9ut28nmug4GoaeZ9YHxucXPQV4Y+h8kCwZNldEdPNv0qyHxI/xs
ZVE24y17F5k9+RZAfpRm5EsoVD/h+WI5VpHa1ugb4bYwY6az26iMDmcU3TJGT4yl
nv6fCGJ/mHM4l7M4RmlvS+IcvyPaVY9IV/hzDSu1Y5vI1vwN75gF1jvD6kKGHUKn
heNomszk7faFKfoYj8zSEbvhijIVoDhzeVt7bdc1hQxUM5LK7tYNTkjhU+NossgZ
Wz1V/Rxj4gI5bAWqFI92yNDbGE1ucj9SclPBy7lJoKuUQNj+JNReswV2yq7C5j4b
tcapoN+/YpEP1+7LPvkSUYO990zhoiBkJgcfaWbgtim0ymeDgdlmj1AoyIyP66kY
QME8MhoXcc2hwvkPeb3wnYERvCR1SOZp91fG6Uupu4zSHQrvc1cNTj6j3dMfkTsP
pwa5QDg4UChqAhYPlWuiW2/FbtiL31sUU93+pmnnoiYQ0P0dPnvNqYtZgGTCG87o
1G6iICsvsbXPxXyvu9RhMKeBUTMEBi5RPzgWi1w25ojc6U9u/ixZwfd1lztoS3js
/oQ4tnq2zu6/JWbQXaG1b5d0b6d+rL/JXdQxT0R87z34DDtzq4rq2Q5trzfQkziB
oeErJJvQJL2MxqfKheosfFPSkHT4CX8m9Au86yrx9B2nIPEIN8Zzp6FzUqCgrsOg
cQ2Nauy4qCLVog3az3rnOGBCjmvZ3RlygI2XyHBOohSMeg2BBQ2P2hheJasdv//Y
aF/FZ0YBsWTMb6Cido8g+LRI2QiHylKl6FhNgQ5uIzS7QV8zc/m3LOZlzZ0Um15Q
hNbfntfgxs/l9ly1hkhKJ4vl3Qmpr55PYvKhDO+XoUd68ZsJOS84tHOz3sRQzOSM
vsZpMV9HAUjVfJYucJAwzY/80YJ//BRgbLdFEkTqgbIV3aco42g9t+3YZgec4OAM
ThNelaQti0Sf0gC+F/O5g9vfq1ftIMYzdTj+6/nJ99FEO4PkVDAA6zoRP95m99Qu
0XfbYWO6kL4ASOxLuRSIXiZQuNOnosjZVp2EAd0TfuWPy6VtQn3kc4eeAkWW9tng
onm/jrgDevoot7CHQftKs9a4XkrmCtxZD7n3fdgfYafZP5dVclqmYKLu0WfhTcMH
3fU2zg9gqWJubpr4IalAHBA6zAlQktAig43n3Crjgj77LmvuSgPsEG9B8kMQwigf
YHlreBGXpulsuYOR7EEK43cC/GvwPxNS/CjnXD5ZUZzOQr56/NrfEW+QVePZyJDT
OEEgZd6vjQoxjqL7ujfc3tqn2UPyl471UX1DTXurSayKooDL0QwsG56f0FKTVYRO
O+Ikj7dqnpTZhZ4DOzOu0yksjQ5fjud4TbEVveFlvk9YIvr+E84eRt1stt78VVYA
uefbigTD2zjL7Rw7XFyoM65whLTKvYUS2votdj0Mu9pwve6JcZOAhZ/MXRm8mj7y
nn+/Gyyt99TwZ76Vw0uMcjjRehM5geeS9uAwqbSGPF7fO4wk7fn7Qsj/DrInz61F
umAHA1Qtzi6fYhjtHGJI8eKuMoEij21yfceRms6KGBX5+5MvBkaULDEHa6NOd/hZ
4ZjfWhW9JUMRqm4fIbuVwztzZ1eg7E5lTd9qecMWrzeLB338+mb46ilV483MQ5IE
4RpGg45vghsQ8fNFzKV366qlDbkuY8xxKrXWCi9yN7kfC2ijhRZFPfXH/Rq89YN0
9nji8kgRBChouzMHuScPwpxtVaxX+4Qbi5ZvY0GgwINhLqwow4A90NsANRiPFciQ
0h3euG8hm7VUWfjhh0zrrt43iwJWUcAIcqhLk6rDCl3TpmfYU6uu9bG67+6dCZjF
XKW3Lks1ix8jSV2eV5Ih4szwiWfovbdR46AnlcQ6s7cJKYRywmS7mJrh+/NAOe22
6a4acj7ECZdaoR+7pD2qM76fRTf6VyN9OaIsqsft3qP+kg6E+6aZeUAR8d21nIwh
GI+AeLNmhID/HP3tXiWK3vho40v+lUIcCYHfS32ZubZC6Fvg2oRuPRb7bQtrau0P
ZmKXtRDBHoQ5hRej/Ogh8CyeCIE2CwOS3wmdbOilEzIM1grgpf1n4D4D1T23kaEN
taksXnwc0BiCCeVFx/8ui0FANLeNQsdj1dmPUm9j8YGbdgKBNkXcxZBJALdVNn/z
1xrPAwRGEWjfaPBlFBErLQ+lBzfMvDFAqE8wn0OMDhQ5FreVqsuDA8Tzcy9Mu5V0
mQfbBD5rpJokkgefgFFd6DcFXFs9fLz1lwdLmMU+fkuQiJPrxxYS8VNZuNzrNuL9
6mja8FBi2nEn3Pc0fqNN8laBJA+l8je8mjcV5qbZDoWwHWfjkDRnirIo3qDg2QAy
VlHtT1OMurj8tNmH/KqbzYz41Rp5pd4DYtHGuE0XZ0lC9Al7lLCW3OBNnH0nLifm
lVnLsuQJjV+J8pSeDLyv/5EvAHKR5njBWhcMA5qCJ/mc1l5tnE8qV4cYSXaayVYN
2NcIR3ArHsyXlVRwLPQxe13/5NoYLQAns5dc3ghhMJi0POu6p+d7TuVZRVO39CBc
qrrtoWtBcIS6787a1grDmSuiAXbx+jac1BWFM/nKYjivRyOYp/z6MN5joaf1u1ut
ZWZ68VEIe3T4XRZ7wZhmeutJ2zVSK94JWJ0Oxc3J1V34WWzxuNBpomDDcWlREsqZ
yoW/EQtJbYYskgQZcJUUdLL0qoSr3IDSmDGV/AOmvjIc0rdWEb0jLAxq9ynzp4/A
89D3/Z6CLkN2Ul/IDF34OmKmGYAl5/GgzsR6kZniv+3XX9F8gbaZ/yZxwgrQ9c2x
SPJ02JfoaXUWosK3BRF/Bt+bykMLRy5Ks9XQ0bSsnnV987lOMUOT1S21URdZ8/4+
tFX8lI56YlU7tr4/RJd4geV1vkyepO1ixNS7w9AKovoyiDdwAHrl8RaYgLcHqU0K
BPolZGiZJ0Mb4mWSrIgYuNfFu1JNOHY6kc5b041MXCKUZjKJU9T7qY6NklPljYSM
P3cwL230zBIgTNF95RiPWu3qgwiYLlZ5R17RzfaUGfy3LB/xZigms0hcPBFtYSHH
WBD/HNi2q4p3Zo9zM6qj5wNY6rSG1sWfOONhkSW0SuKL5nuW02xg7cLdobKJq+i9
pDbEkTu6r7yzlddpIYRl89X8ZBPjumsu84mfHMXckjnApT4p5lAF6cZJfv+W+D9y
OlTz1kOk7ZtsPn2R7LweICnIJOAhhPmidZmoqxcMjBS/4q0pyIic2u+rNkHhJ3m5
vW4HGA/EJ90a69FiPm0oA9PQXz2DkuYHCGHAbd9nFTxPD0OU0JJ4TELuyn3JtvKv
JiMfz5wtcimlGQZBYZOAdB0TJo8uLI3xBLnZsWwA3++g4d9hlfNyjTeBnmlUzsv8
zH08LiYSIpzgO2QWRnpAiWlA3JRRpbvRDxZsveTIdd2FZwo4nUGbaIpeb8BQIPbT
9X23I8dYiIn3nD1y3kfyskjQiz0G6yex/zoA2mgqhe02XVlZF9h8stYEJqicwDeF
WPWw07dMQz6WZm7RcI+SvOI0IUHTa0ZLhABPThGLiDcj8D7VKeARIMi3SadbThfI
yf9Pl7l5Y631mu7cWGbcMB+mL95YtGFuuaI5NNFOcUBE6Mb/0djfv8cbvW+ImlPs
2H83tEETNjjq8fbhKFF36Lo+N5AIWwl7eCnvEpt7RuiJBQfiNIt0/9gVIwYsUGeW
FMn106+1b4DSGXaqnArKS+ierDKERv/5dh7dSm+OMYG528/ElIAq9zB9TLpwtUnh
vumIE3buMfFd5NmArxFVPA04vrWFz5e4III22UNKXpkhLd7NMLIuIzzjzPo9Bsqp
K5S02kd/4IgfxbjygsDXrv1A+2OxDFUn10BI4GNuD3yqYmQuOfePsi+xQzHw0jm4
D5HFuqxhGTXLB/lrqaViKlcn3ZNEcIZ9PSwBp7ACqg0O7MNq8drb7NqZNRwizpr3
sR2+oKtzaLCvZea1L5xMF1ZKka6uTpDhQx8TgZ+W187Jp5vULClaaq5cKJqoXPa+
kRVvdjHiJx73dfWe3PxIb+mY1y70i9BgSvOxOeIWuXQ4Qzx3edXlYDEDtkpgX934
Po8v227qI6veFCwJFoP3uHoa3uPnJY2AJ5RqQqDmd0DWM7W39mrhFetFVX0Vn1NL
BVR3yQVesm7uUwdYkT8fZk4/Q1UtAsxSafCao7jd20dicc/BvSm6LO0RjYJ+5O7u
RaBEs5A4hEYWMEzG+d89eDjGPB+yw2FqcDYFFjwdGJsPGCj3gIq5thwa/LvsE6gW
MDNGl3Gm2sl1Ad/S2datp1w11pKzZlp4UKsivrHBwt4It/kAmOqvU0sjL/tstI8J
Zs+U7eLGL1AsGUVuIquZZgqwW3GSQ93e5gg9oM2u9i1eleO0Z9lm3PWs/ao7cSyl
WPQ58xU7nIC+9rw+YfcZS4h6qehrnVENbQuGGcmgX36Yc/DBM69fbh5MMp4NgoUA
muCLyz7Fn+aH5SwYeyHgwFImFN29cKOrDb/JYmSghNDDkNDfXy9YuO1xoHNaEgHo
CxitT0xexvXtDtCclfAxkGCql8qBstkid427P8wrQy02c12gEBbpc32woOef0qLB
37/GgjdFIa72k/D6RogpFUzbwE6MJVOcBJUAdOFphS6R/bzHWW0vIEt2NbEnEMdr
JYqB2lbhou3gZb6FX1XnGZ+fi/CbTUaTCgZ4HiFSHI7NHuh0w2DqAYdvSF+zVBkV
p1yGzCp5g8j5u8rrzhkYQRA6eIFK1PfdSDh/h3XuZyq3xzDpiDaB8U6eW4hVzu+N
nBLZwE7Br6U+4YvW/g0zmqTR/8FUljjcdFghjgJTieWC5KOmCf7g66IDVQ7+r9o3
AUCIvdstDYJBUqnOejDt7BZ5LZmSaJNDwo9p98g7JGZGlmLJeILzM0n2xRtI8IZK
okpT0LUpDLlSXkcsxazsaajVFiyNdU7Lia/5rgTae6tUPJiSqTYeGlbOPSsJNq+N
Rkje/TMN6jivLbL76WIqjOCBKmzHKPM5Tw/5K3ko0l1aYMiZOY6wcYm6odLjmICp
1iu77H/KLlIW00hQ4be2bNj4avarA2Ixe28i+AM3h07HSbU9qs9hssWgG80M9dBD
ZV/XBAbbDEPd6UhTXn7ugWP4sX649Fin8m6JCfqOywYh1aRwEJke+nSOsCQZS8nY
4NStfCtwNvQL4muvs/G+yXILfb4es3n7sLaR6AW6Mo+epGsWM8fLSsJ/uVDWQeFy
BOBM9FUbNh4srvK4ZndBEM+I2i2WXpCoCjVWKtq+KHEZ2OGx3jnUrZokt4S1s5mM
7KnVk+9CuZmg37By/fVQXo+aBf1HF9RkFmmBt+LVTdse2m/Kty6brJg/lvgBjxiI
wt2MYTdRX+3bBRCaBM7dmCltbrOSUxo9KQAQzjTrS+VS1bOCfFwDl//1tTFk4ESN
WpvHuS0lMbCa6sS8lF/RYbK5CS4I1gsCxNFtmDo0BdhNSTYTj97m5Mh5Nl+Hyay3
WBFYfn4dfezfEAzKmiuHlsqmmH/3Fi8V2DeEcLWE1WX6STKr/CrpY01+8H2a9i+g
ZiZvC75wJXpillBrb5a0PxATbMaQ+Rq6u20hX8M7ir6TmRP5vI3ObiQAnSilBbbc
sJyR2OyVUyI0WU+5wE98zUs4plB4nAAspBKGMf2wA//WfanF3Yid4p4JCBNh21R+
a1tu+Nztm6OLVntTPrnuUt7XLDKZRWK246gMNg/xTw+Mb3vkR5HlD0nFQr+MeDFV
4ihM9uc5gK764Gli+vwhBs/c9Y0/oPhH1Z0RV51d4izrU8Lhpib5Y8aU5A+eVe2e
/OHctwq35b+K33RVUD4HlqR8sl5Tk1wOobommo4pzsJ+2QYiiDmR7fHfLvH2e1ir
pQ8elA94IA6LVsZz0lxd2VfU15t2unFC6/MkrWyvEnxCfC31hqZbSYw9MRMl0DdM
5L701eX5JpMQfAQeMPS2LM98daJHEyWwBPWWWJ+C8J2S75XGPAzGIt5u0Yjn2QXz
ShyOERBe3YJJDYp3iyLC1hZyKZSp0+pEHVmHwrPWv5RXwJG4hJRgPWpA4RHvmQfW
kuMATiKKjzz3XzDGh/MB+gBt0F/NrKR7OWHQY7/CQib0PHr3z/fxYv4eRAtVrh54
Qyc3szKLq+BlpEQjSuLkCaD8PdszVbi7t5cBe1NIv2OPu4O0rQNN/0zTebRCX1Zy
34mv+SIjRCxIfLKawdaFicEdB0lB2L7a8tR6yIpiW9Qog1L+mzbbW1MXHXR89sWT
X8+YVQiUZuudvf/fyl3zBuweRA74EpZ9lWyGSy+XBsudj1bfT0bD9W6WVgo46CmO
3Ew54Hh1H1b1AiF2NGvU34hbgJgtl1OWNBaWf7BaH21NeSr8/UNFjOb+vsIN+fOM
lIhLO7q+P0hVygkp5UNowQmHheTVdFr1ZYcGwYSnKkycZ4RaZer1z3ejznZI9xAy
i+IL39VSgY462FIDkz9Ibae4FsLEKMxTFAA3l8ue6Q5bUQNPMasYJdPuoxby9n//
y4X0w0eyYP4P4d41NY0ShJRZ0IDmmtUCV1l+43fM/TtEx/6BHHyLJsmsHyPFdqtG
MVlAegozu/g6HwBsBjCQayYkkEM+U/H3HTwWdoxrF9kQUGYqSVnigTB0vj1g97AW
hXseuSISIuLaAeAL0y/sf0zTzRrq2HbPj+E0f7dd8p4mahgGsXrEGMDt7LezurZe
yNi8zdgCp6vK4WBD8wxl0I9xc2oc7p/ETQf/DDggZRt2jy439IiBIWYCJdhmI6Ly
ajmIuik3CZpX/I5+1+JYaiHaZRt3jogySWukAbm0/kywwk1VyZMu6gK9QDJZ1EjN
x2V0QyW3+ufcRI5DQWtKpUVGDeGZgEYmtXiuoSWmD6xoZ4Ue6d81Dpyxwonq4y70
4FTr+zQpDPlNUNMX22Nnp5/WepgubkT6PsKobLy+D0BwM2BSKk7/y8g1/REID2WM
7b6fkn5EJgqtsYNp1UG/EsDmlmL1+kJwxoa4pBXtDtDcpxQfgWhkIJuhkQpwigKi
KhVPneABf8du644MF0++UgIG5sUUzUrHfWxt6sZ4QHF0uEGFzK8nr+RQVLVLxqnD
dOCFRHHq40LurmEPYL9l4PNslwWu/92kHu2/Crl7IYuGf3A07laZXL3wJufU+DqD
3fAqz4O6BLOOWJPeioal0sZ5xce89sxZjySyY+8JqSqapuzweB8XrWyMotWyOmyu
6MOMkj4bgIJxv35p7nkZ97myXqrXQW+gNFuQLQ2vU/RnaxPM3ZIunGIlrdBIscN0
PsMezGsO2D+GNgVq8bRhHKCCbkKRWLH8XrMle6pccQRliazihLLXhWtQpvsejDpr
QXjKqKmLI4ctRBAR0dWP3TTIXaq7Q57bSxWat9nDY9Gp5tYW3jIBfT7HuT6BDgPv
2L8KCEKNJ9rIaMZ4eqS1+KGkCIlfgXjI7oaQzffOuy4yaFMGpu2QS7gBPVOYSFZx
iWBh34fwERAD8OzDHIoUtuKsVXOG9KC16awrnyuTnPz/30aPmMBqrTOuDd4/bgyv
07fCvYusaAG9utcNN101FWZS/wJqT7SGF8V++SUn/PxtzfFf0V95hh4ZDEfkKHum
Altk6toouFKJiNF/Hm5WGbP2Tme73BLerx4C3yV6sHe32sQ0mV8SW5IK6hqC+KaP
Q7Z1+AXdUd9lnkDJ8ZV0luHRBWswhGh2GYc7jdBMG44+mPhBLshCWFKwY6Rg8PTQ
lJSTXjkIsiK3dkzPDwVuVpNfw6CfloBAG0+Nd6Kq2G1gwv5sDTJYxWoRLy5tADXM
9srDDToWaQFllNHFi8H13L8us/U/LUGJAjIAyfsI+UR1uoteLEWz3FL9UJymNBPY
OQa/V4Jawx25eWWCOGt0nJTFYUFL7+VO+dgFK3ihXurcTRd3/iixCryu9d5a9R++
RSnpSxJjw6Fy7RJZTgUbKIrbeQbgq9gnWX2aMgmLtsmNgn0ynn7YcdHfn59Oe/RS
pLrg0s9xzoHab3A/1nOlJAWcQ/e48QdNJpHAs6K9nbsF5fSKaH3r46kTbe7hDbfc
nQa8yIHKNz+kKm3oipLDwfFd8Yd27UR2PD8fhrUMHnU+MMHtpLsfmf+vQIYV/7Rl
f7wUo9nrprpk3FhU0wAxqYeKl4YTCW61KoC3wGh08+bIy29y31YtC5xQFpDMEHfl
h+nTfwHB5ffJOPQESHIjDEu2rKUnu5LeoAk54r/05Wd0YfPTxIgk/NrmgmLeOSjz
MXhJSAmIMlVzZDsgkLZzXg3+PAWuLjDqYeVTHLEk/yOIccnIR306R+XSYTSoOMYS
W1K5I24RqHnFzNH2l/sgNLsHaGdU38Qu336waXzMOScYuaCI5Hn+O6A1p4D4mIrK
86voN4w/g4qLPi07OeI2EuvOZT89HtSyd0BPCZCBJ/EcUu7vhPke1RHetF5vdxRg
tdwDHaFYcf+/F7CkEGueUW0OEKZnIT2FjibTwXggt0oo3/CZ6j7k5cfj732wvxvl
rA80ZG0HTF9RmdLCF9eiQ9TZWUWtIbFG/L3+bYQT3GU97N51zQ3aFD7wHcoo1zKe
zToK5+uXgDziB20Z8SEPSwB9JJPVECKBqzbNAQJb5bpGpM8vPXOEfohynhsyzvXP
UqiPwmYujef1BEaIVcEaPIf4Jmk8HTh4rKHyjdSyZLPp37zIG7I/Vu29MKCiPSOG
7yU6sf5ddMJSxvdcZ4zME7MJiFkUTSrtmjMPc+HKaM5fB9y/V4Au/z1fvZkeAe0j
bRhgt5mlYsSAZ/K1ZTimQi5xN0DrydbXOhm+ET0l7MAhKnSuhf/eedSVQc83wE7d
q+CFLwjTZtzDu6RWK25bd+PSXfnOCLcrjpS2bUv5JDTwCKjLA1ERqNxdTQFO49GW
OKihW6/2sPLhk8T6AguBNMEUVHi0UVqtxd/lde+6G+2Pz9it1Dbp8Gj+WoW/BrB9
DljxKhO8EFsvnI46VB7ZKZ3IWGF+vkIqgreCiCXY83PrJnVvZU7EFd+Q2dH+F9+d
TFmuH4MzEBFauBJcQkEL1TtX2acTSqsJZYbdKgas5tB1kWo/gPpJkrtdEOAQ7J9f
lE62F348jslNZvTCRYWnlmNUU2yIfusNoJaA8VO2tujFPGfJ6n55/7v1I/ecvu01
u7tBNYgOntvkhNeHCgKNd9xHjvim8I/FPjRodM2yHyeEiIK8WCBXS1fveC3zkK4u
kIQlzLcsc7x6dBiLWSMkGxPyDceGntM/CRZM8FLgd+VgSRPQqX1JuRrwqid0Dewq
ESgx/wUzZ9tGgJLbMieB99WFpWXUeWZzxjVMbe9taKieVt8dRLgFRvVTKGa+SThF
c+gVWE0Aa2QVefcW8hvC+eyO0n+T1w8hQ3LvVUOhkwC9qnW3EFA3RMiotDSTW7wl
1AlfQCdN3PfJINoZPG1t6se1O5HZxqnSVJHmW40ed1A/LYPSc1tXYZHwDBqjsPUJ
Yu2jPNiuSf0BAz5NvLUXpa4us3sWtadoNqw547IDBWKhXU5CSgGtrRUsoViv0Bdg
/XVbW61sj9M6OPwz9ITf0kMq3rlM0CcH7MbFYcle822s0eB2LecYftFgShfRdDaT
mvzKbOY1CwAR2LZ97Ff/pEFib9H3+lCdTLhKG55fM6pRtsu1nJJHqBqm6eJjyimY
jNhXTjtdrT0/01VvzYkdUMsQAPe8VAvofL2syJ+3B03QkyVhtNhP8B0kSXgDTmSc
i6/eBdEeA9/ZYMPhdEhRkxOH+AZZ71f+sh9ZtAvGkI2VhIpphmtvmA61wt1iQ4pp
POLtVl4S76p1JnQUsPkzVkW3tphkGzzMIWiBR18xoFM/UjSQUSnPmKgRSU/XamVa
Zcx5+P0UXQ3XKLt44Ylmt6JCJz4/geh67t+oO7SLXpoP1FF6cBzTTE0oaPL8knJv
b585AoSWcqTxTutVCOnBCmwlu8rCWJ5zAT5RKfnAqVFVUCMOFAOKszsHSAXtprdy
jMbeppHA7/zMb4h8u1tioRzuD5yOqFS9/N8LbSvgyVP7QoLwwkhpp1vuscD1Ldx/
UgyQFejtavV7+WCkha1SjWqA4Nqt93Ar8KVDiNraejWzH1BevbYjZ2GIhtWuWHMJ
g35FPujcksMWX5CW2N4sPswTda9/uJcKTcoHxwGuDjvbYYG/xHQcJZ+ui3ftO+dP
Pl566z5kn1ef8t6h2wkjetFdbbNaFRsaa0y28DxhsnvK4v5YFRLZCnn/atagkjEH
YSxG2xK5N4IZBnRhpJGAHMpFcKN8AC2SYItLV7vDDkiVv7WM87W1tUzbhB+YJv1k
xuiVWBakpbxaMt6oErF9Xk8M7VXT7sefB5N4HuyHlvGsELc4YoQfvJfWfFp13Czf
yez32h+CCLwW6cmoyJn1qSW3I3SxdfmDmRAGxjx9brJNB1BGmNPSG4Nyig4EL/3d
AxeAYkoM/+J9Pn22d8KGVBlf2Mj4CMwrhVpgZe162HrRrkORG7uGHKUn2eYbeZjj
anRCvDTZlz+2fSocKChvC+B+pLKAVGCv8QkJP86jMH0dE+C+wyPmJmUdDXFQGvyo
K4CfI7glsoA/obbtNIuHHBg4eJDNFpp9wgXR5E5SNCaYElraK7jK6sagFfkjwxR2
Bi02Q027dk9s8FhBkDP7AftkkzMmZ46bdId6yHB/+NvzD9hBNF5MVxddLAeS+u8/
W0ZVgSQ0r/eaUfsVdmAt1VAzEweBC1IGSnQdOapHlrBIDSu3i8nu87VXbbcZfSLH
Aw2FptnbDAZ2BH2vZ7nw8jBB1RVkb617zy8CzOtZa+247prHZE4Lch10ssOmWBAz
n54qpAZDoapiZa71/Lcq8AIz7oqr3JGufI11cGHFl+ycZ8PQWa6RwZETqaMo5CuH
rf6fY7hq8XB7zYe5N3sNuJY/Ht6YOQKoHAwgDCWrgYYwqklUvmrYsoajTEUjT7nV
aNgGJsiPc9nS6EKImIicwxYFf5eDvZMShCPu5kw+eVjkQdya2rdiRD70vJkv5uN/
u3uPzdJ0sLPxq7RrsB9ThnBiZzBfbyoFm7JONBdnmFxxXza+z/SIdAo3txmKFP1K
9di37yGwab9fjP/9L2UWs4fnf3bxpFwqsBm+4Uym7Elprp3MBmfw2fGydL0uAt0B
g0WkWgUceWg0AeZ+HvAy1i47mphT8jMXCqcu2Gq1BzWHSJa/DwzPcNDv601Akib5
HNxxlHnVov+Vm8vB85cFieRBXns3RZnH1BGT+NZr77slv3zB0syV+lJZOt6nkolC
7euolGd0oRVuY4j7CytLUrXKm+8vHrELlFhgT09HcWS4vHl1ggQc/kpoD3vJImuJ
/S0qzFggCLfetekNUj8lbxOLWu2jJVPVQ5IwEvyMOD19vYSvqevxov9TBmYWJrlo
1PF9PNRHzxNu7lIXBxPszEcCPHrWu2B21X2EqH2i0QnouSkQMT4/itTXzqZgDGHN
hexusf4gfka/1Mj+jo2+5YBbWEgx+nqys0Q4yPOQYgMUNe6HgVIrKtHw9H4Zxv7I
BUpr9YuwNXlx1oFga35ZjFDa1+IuRlxN8B4LkBPZxw0Mfm76Z00eS6P1dZR9PEUO
TjRvzByTl1vHal1p/apXPYgfB6gKEtQ7syEiNXuQi4py5joHSLmYeMBZjOr6/CoV
IGQr+AqbsSRTETKB+jcUuIZD+LNCY2lARKLdud5/jIHVFP3kHHZ1hc9LivRw5DBL
ggWiRMoC443pGbl5cRqp7fwCkKeYEQNEQjCd8vDL7A+BMoVwjoXE/HOmoT4UpBtV
sEh5cCyhTUUiqBEkoUAeBTjvgpbkAfckVxkYhF8VVq/Qad3NU7cQ0O4x4lhT7ryO
1Xe2eiheOMKZSLZXNo9ibZvOWvcFGsumJIUU0tzhYC63KlZBgYym+xPGij4P8bUP
QmFw4r495RSxFXM4WYj2+/Dz/+vRTTeyKwyJMpzZoeZE6KuSbK4QQMcePt4WuiPl
g6REOIZRCVScXI+qkWSqyefGM6vKKiURT+rikM8x+114tHdVEMMOpcqRMQL00GnV
O8qk0oiulcPfId4SgJCSAI4BMOc3ccnv2Y4aMsPn7Ef7nE+4Y72ZCrNge+eYv2eW
fKfOtiW+arZYiYrChEGo4C5R5bC6zXBV6rQO0jyzGOK8V1BlIeYpTwoe2Y9mFq3X
cEqR4CWjVVALcWdQPg9iEBWJVEQnj6quSXuVVQFd1iHJ47jNx1j5wDzxNImdUtLz
nsY5ES27DWPYNdy2/kxM6Mt+gHET/lYdQNIqkXNTrD2aq1Jyu1vFIxmKv78M2BQs
NfOiPozAN8a/daxDu+nTgYea0dqbrqhGhWuAS1FMdipxXhyH9t86MHykgf9d4rIH
0vRAzEUooIUMzQj77mnhncjxRumy5BzRtWr5oyZqONmi8rwlNkNYsFZoihN6Dnd+
+oLiluca1iCzYfUCmrAHAjGeOy4OtbEAKui5INNU8YfMbJ7GZ5rTejIUpdXHiopx
uM8nGGlDs62W9XiMctb2fWmrWQAXhwxY2AGXvLQ/JJgdL0NzYgneaFCzW+r+k5w7
qSrsLg8nzOE3r2xWdOSbIfp9KVki4UkKkg+NuyLARcwnH/fN0+ED2yenJ+cTeyyf
3vhbfPfkdXgwj4aNZqfKAkLoaa8G2VtJATmrSGPeWNhDX3KOywiCdqMPYSFRNWOj
9I0SUaZJXOfvvaiR87iyl4l6ib6IG6cu9K25o5MdVQ3xA+LySQCI0XbfruJMr5+M
nC/6P4yP8W+2vg71mzV//TDQHrAQxc0vSy/kx5bb5xqW34LFQqHzqp422he8838i
zp4iKoNGuwdBQVfRNj2eKPE4/rqgaG2ec4/L0n3I/j2z7NtLWYA8Tn36M81Q8f6v
qepdsf+5RGgdpuIov2dq3KvuZ2gLNmuIbW693V4gSA/0sOyrAh3YnYYODSr12c8H
33a+o1IHYj2i/YPsRhmegvTIi/Sq6n3sv93GqOtq0by5R48kuqW/6RAD2m2FwHdB
OBgyIcrUMs2mHQzsu79hRIiVq0Amm23U8WNhfHIm8G/dr8w2Pdv8OUASI2LwbC6V
xP461M3MTU1vY8w7s7MNHYg4/BuA/P6G4M3swFsY0nThSnvjQt+ujVy3rsjMCkk3
mimreMQXZlhVXSQWcmnbc4jfl5cD+5MEwpoGtZoX2SEkScNY21EW1Zvvu9qXx/SW
EvrUWsaOtaVdLH00hiegtZofMX1dItWmSjkjPfg3NMp7Z4sbkz29T78RyfWoeXNM
DaiZXUFQ0uSQruxhvDqaj+XK5cqXBmcyrqD+fclJZc6Sc0NvO8WRlnz7M2/oM0MU
jtTlS1MURtdswkktHKTIyCZwxAWP4NKJBlp97DtgB+5TP1aBE58FfZyzRh5sE3hB
tq8zHfv5FeWEOVshQbkqKrog1dCfPsvK1tCq/pwogTgrwllaMVHTkoSAPv5JQb8y
nMbE13deRQ4wD/JNS1Sa1fWQ2Ydi2xHdjMymtqbRk9a1IPlhMbIgk3Cs7tHbmdie
cDyp5eq8f/uGGxRgSK50vu3L9nHAl/cjFwhYV4KLNtYKGN1eEAhVYsGYol7NK8nM
K0xFYQRXtUYiP3s73AiIgLjo54FqmfGpyPP400D9cqpaq5YHVD+AhEg139QaM/vQ
pD48IdrEnCvbvnsBIknax+AgFh+laMc1+/Sh5VTPEhwZmDxeLDwXXOwHQ+TATTG3
w9y3Yv3vMOX165zzB2r8AGEzB9JbyyyeeqILK6aF+vXGit6SIaPQdXyXgnSV4W12
0dmWERKCnooIMHlhy++D/9z5FwN0o+cFO7/5rMhTzwZpE4bOxf2/9GYmXvrPuXv1
kMTeb6nxLspieOHnH3aP7BNtqLDltlu6Ud9RyEqYqXsOvHY3Tin/BOtCZG8QpniP
a8k1SIxrcAVvyBmjiBPy1FqULeJ7slTC6rx+plWrTiw4UeJ2WoKPTAzFeR1P8c33
xeqsbLN3MxFijjOSpZtD2XMR/3ARauE4hy3G6UEg41yhdoodJB3Jw7mykfnjanKB
6aZphrAOt9oy0UicJZh/s0bnV55P3R4iuPr18fmLCnZUS86TSgfe/E0uEIIRU/wU
OroOy7JaqSXfd40mmDPizdbsfuSjlIsrd5FMBvRyqWaEQnmmCIitUapt3lH6EuqA
5AbvI+XyxB9ILgKUEQx/yfC6Fymi/cf09yG/kENV+MGJE0782n38ko+1q528ybJ+
J84IT1AOsAAYg75JBL1X2BdwhwZujxgmPdvZmVsyrJWa6H4li+1cyCafE2+8aMS/
SdnB3/OQziOtdMqCcQEAAc+9O4i1UAyAI7v4Ytu5CnHT//IQ9TnkyIIQ0K0MASh6
gM0GUfT5qznKVRRI7cBPho/HW+Z2CAFjU1ZWhCB2XRWZUsFtR3bfGAZ5GFO9pLu/
CzISnViQAZA7yZIlDGBx38uqlZrS1QAtoc54d4dFhRDg+qiQ6WrMLaItUBPXC4bA
k2z8J60nhGDU+8Y9QpRz1gZv1D9YwBLISW76yILpWQvH4XSffT1+H1ws50qXK0Ge
KamU4jCsvxPxTRnK/uCkQGRvWQd6vMOMY4zSYGkvs/iJ1yHLGzNCqULj2vPW3BzG
cFUHjGN/xZ+p77qWCaW1AuOkVsFDXjeYrXRrqmFah/s4H5ocAhQwKs+im25zPO9F
tojaVPAwDmYVo9jRRBqQQpEY4TVRSgRwmR6DSriAitiD8yBvEXt8Qxdz49AGd8YM
a9ikQ7qS45XnB3q6UzICbIcLA8CAAPVVx81H1OmMUK/gaDAtptQ5BevNvlfVXixY
bO1SC8OQT03AGVFW3TW6SpzVhYTDeHGZ/yUu1D/b90R/1Z+0EqFLHv8wgw/yiTmQ
l2UufiM9qZ86E14Tq9lOriwUEANqSYUGaut2vqpMD9ny4lTGsLeaJb+CXQimcRsU
QLC5q+xVfAvPteosMWxGLiMXNbntCHxYo7aG6ruZ/sqe6NyyOSsBnabjdZEu5/ko
auOyxSKoCrpXXoN+cWVr/KdQrWVmSy+AuvdkhuWE6gub+IT/RE0p8wnWWlJc9I8D
l73S6gEUpaPFo2bF+m8qF7zxGJJf+FpdPBQ1/d+zyzQZfA33E7epOspzqyF3X9G5
60urqlxtwZptMRl/1vQarRefGQ2XHs7+iIrnINOCqS8q3GovbcPeFCjFEz7RMoEs
CjitAyZL88qu1VxW4d4+7PiTsICeffuiiv5/RatzJDnAfMq4IfVbNAuUmSmWTv+M
U8V9G04c+8vc9QCCodNKMGlHapha+I0vGtqYLoeP0FEgvUK5U/xJH5s0AcKHUycC
lGcjqY7dNVSPefJnrJRX8Y4SZ1bA+x3aWFPSVK/+NJjN5OfAKCvVWL2ywHQDe+H5
iShVZtP9EWuvlQ7/tWl4+p1W+cMOn/w5K3fJXrcpu6Eg5xatHDcl6pG4CwyANqq+
GaVV4kFtQ1Tb7vf9ph//HXDsjYd7n9/fu06vQrkgL5UWI2fOqO6Cqk4Fp3J+C84q
KalXm/dcgFDfqfE8zONv8HnnZf5xgErwR/xqfdmP1Rka/QM9Uc8QHiAZoHy98Hbr
JRl1xka1m5MRhRctZBOdqmUY3anJpd/m9pC6SH5gJMYiK6O5x7eMRxWvbPEvSR5t
38Pd/meKEaSmNJaww2tbmot1mtRBwDFw3zpomqJfus6h+S8YkT+M/hc98x/baYNC
9kBoovJnCOmKAiwXsDVmUCjFeQ32rmLba5N9g2XVps50ZmVoHhuasirSXLl0obHr
dCOL5grq8kitO0PdRRInJsCJrmk3DmKCWPzkwfEUzDoIkXzpN04g0v5TCve91BkE
aYw1TyvIb2xEXEJpuOhj35nLJcdePq3g+iEWDCxvD4lSEmWKkYJPV2z7S+il/Zjc
Q7S43+3Q+3y5At3zUmgQQgglwCi0xX5pWPkJ0iWrTjXvJfbsl4MIePIHwlAWJRlh
tB2GrkiqjlaDMQoNsZDr6HaQiixmRgczhkxo3P7Pdc18xZJSYfRDK4E13pCdptC7
Q9o9YnDv9bAx6FKLp0TEvC67IWBS6eYJVyVn8vz2CDjj4qpicG3Q7HbLo7iiDAyy
ZVzwAbDxyuQ+Xzs4Yza9VfLyJz6KOCvBI1sUXUCpNPYmgwIeGXBZ2TQ8Xkqqwllx
SC0bgU4QQrOkCR3j8wwFISWlZIIg7I6a4ZOwGLRcNFqU1hJmNuy+aFN8k7sOuntt
8ZF6XB8VSv9tCEzWUM7gQVAXM+5nRNPP1BcV0s9WT+6/He0fKSBI5XYU6vV6RiEZ
2sdqOVuWBD0Djz8IbBwACPIBSV5c3/sGDTkmEfuaVWIEnbP7r5bHBuZlkf4qMqAz
TkTqNrJvskKh0aMOIuotR69SyD4cJlIGVcfnjUIxNh0O4kIejePjgqlKbkrOPa+5
OUPSeIJXl2ogjMJiFFFCEm0KqA3Bpqw1JBVWTO6xmbJESld+zMD2xQAMKczMD9Ua
0mt5XvcuS0xcN7X2FGjzDlP1ilo6PwyglAnBBWabtdcUKIkSp/PbexLuCn3zc7YV
Gro+5cWBauezs7XNxxFB/relQbNDFFSElEdP31q2fICAqjcMlEM2fL0XCVxS+o91
SC350iGPDJ0NhO790ROn4RfAbOLpD6Bk1357JWFSswDOwZle2WyKyqvaVxVWRD9O
UIj/Oer/G7DAw/A3mrXP8Xu3aQshGuTH5YMS4tjkMkJ7N/TNBQgvY6yl2FeErDS7
kicmf9MM4V5egu4vAoZFNxTrXDZd3x17lbt0ANqORWqGMUvRRUNymq0zBDqn4+ma
iDAbQk76hQrMIP82lRMJs/+4M2udceDoL+BPyndiP5tACED4tS7k7xrG3XklRzpa
yLBSpTFbBzeHJpp5u3+Hfrg3nM5p28u16w7tysn0WPpPXDguwoMJlhQNJF+RMI3j
6RNNFD0RcmUirJwxjo7vunPIxZdVGFt8Ki/AUkySB9VSVzGo0ATnlNU72LCmDbhR
fC31oHMeqUSOOsX+crCNeXZvZAHYzl7BLSxKG5eFSztua4Szc88FBFWnphUAvpeO
9LtslQZuMf61yXpkoJ3c5kB3winyIRIbJBiF3QprzQSI9l6g6J+meptxZgs7gop8
mRplFX4eRTxmLJckaYiACwOFdjhWWu+qGvaZIYXsxHJqgNcke0xqZqEQ2uWq4qJi
AKvHEFhvNS0g/5SAWQuy++NkbDofTDUORejW3DiSJQmpeWb7F4eTMH97V0tyrofI
oGPDGejPWB+dU2s5DazB8HGTuhtvRt+M7mIz1AXcnJnKZ+6rf5Vdrp0ihdoLFEpU
wNAOeIGZTvWtdg4xV9jUPT8oiBGxQmy+utllRdbpzU3lmiZKiAt6c6j29SW/o0nE
OpF7Eo3UL/IUgDwVi8bZquRnsTEDQ667NZBi0ruZiTP9iDYXsYBN4ChoL1WPpx4W
u+L+rw2D2dc3ENSujWvFP/msXGiUHSEyz8/8Ez4xLfRtIIptSLDrItzfSpCkH4f2
Pkbbt4U4kQBE7omDEHfMB0c+fmOZ1TxExF78xl2zlPwTp1leDIEBi6VYzfEHMI6f
Nusz/m2G6sDoR16pvnF3wsMiNzS7aU37LBfAUKgUaNuuCFV7t77e/3WPL031tujc
T/We9ixAYU31y/tPDLGPjRuJlpPo5gti5sSYhOykueVptdtQF+l/p5jX+tMjwtlc
lOPhkM9FtQc2uzNzwx6wy43f/8BRiNkAQKv66W/jRBz42zEvc9ZwUmWAoxgFsntG
5j1sRvX8mzVL2gY7WBp9XwcKmmaDV4lJjMu1mZsP2xDp3KhNC/UmiNqCbqat+h6T
qyNRnodZUWYB3dbDrZQ5SRqxc3qV+1WYM0uMvD3f5hmNNsNzPht4yLZ4BY1Pmrta
6lXXaiqgidqC6tFwQpGcqqm+ScV6IU2+pj4Us80w3HINzStNMU02NbBsn87A5cS0
HB+z88PnKONgSPI5QnqAOLP095V6CmJLB5E7kZKsvov1OY4Ak/fYt7rvi7HAxlYW
ecKcSFvajUwrjgyBSd0HwFggdQoXUfxJl6lzwCSkkfntbj5slxtu3DpG5rBgotpw
ujKnBsc0kiZuNSmwC4xXxmagf7S4LUmgTt49Xahz0i2t/4wBo0sPPdKPMfDLkxnL
giJKWrbgSC2idCgl22ESe1TEtQPQ0Safai4/TOylfwxA69sprl8Q+zQT7MEP/bRG
wHaD/NoPCavsoMICjVg8Fsii9xK6ffWSo8ZUdT3UbZ2Zn4fAb++EmYi0lqvr2BmE
Tn1qvAJM0VUpcj3+ds65Ag987oPfMxIsXH6XzTHaTDTu+aB1wjVmnbC7ALflUwSO
dkSK1mE/T8AhWxQPMphoFcJOEiD9FgW8Mr6NleNhbEJ/Dj86hNeEcfX+Yyv564zD
Lx5ksxamu7xA1DWtCXRg8uE9YQ+ttRGbW5UYzTIFTOrcVQEs+OK3V0TuNnNZslrd
KWjigrx3e4Wc5frIJ2mO04QVZT1li6MBbIKxEeSLzFiAQchsWzimoI7L2JJA+wjR
YBZ+jrKf+L2V36Wch25yffX8P7A8WLDZ3e5WgetqLYe2HyQFOt4pr7pGpjU8XNkf
T8aX1s5Om/hBjaOBbVAhLN5WsD4VF5RYf/0u5FQim319muEn2VzLA+fwOYBS2feV
DGp4QLMXi6NmtixurqWmZQAUQHrp6zUa8TZxVB70jgYDkFOPCM/qHjQ9xd87N+O+
VB0a60lQNOTFpFS7VpL+K97wKXRigSHade8NpVJP6KZSe1IkX7lhpv80yDn9EIpv
irHVahoEVWtV0nDxi4pofOusCdlRv14YbRrVs7sBPB3VJ/oNY2eEqEjjiAuyDhol
FNyRXHSDfTcDmvr1gLMGvW3/eRERXvDepeApLZ/3sFSV2rYzInYezm7B8WM8Jx2F
gLoFS97PgFXj4efhyvBgKI17QT6okNJx5L+RkrfnGMfn5Zyjm9ZX5wOQWQ3DQ6jl
BrBXFgQUSstoyiNeEV3KX1gwRhjkLzMxIkLDsHN/skVqU8Bw1IDSGreNuT2H/7Fm
qZ8XcoXcfBMksacEEfSRE6wRtDRXpDIINTSc6Fy5N46nQEGrFFHWNT/km0SbTD/a
oEAjMkv6x/LfzWWcSOrBMMNPASPu7Iok7hi3u+OM3HiSnV0wez68rgUW36YK3o7Y
2BSZmA2YlzzxCVoYKD1DK2sMvOLjeQD/MyvgLUzyGZkmDHqF6Ku6hZ4g8SuOcSon
K0gpIkzH5liZbEmOZLEcCeyliN7BinlLx8Go97u/2SLHVldLGkZrsC4x8Bf18gjr
W562DfATb28tG9xKcOWQs++D6CywFwAi6WtXlzso4dw1/pb9y7ngpOtLHRBMfI+Q
WgNLKOIgtfbdgDwMdnPfvrsmJEkNB+25K87qHW2dixEORnCtkZI3jm1D3He3ZgqJ
3Lsrc+tQEpaRP1ZnCO9TgUQuGbeLGX6ILVRaE7LbSMqszykV/7l/20H+ZKfeU1mi
TO9ghvna/HoWSTiYSytFKoevhcG5srytOrbLskPBKJTeTjjkErn40wIvdRz4XG5F
VAVAtXlGrxl2KQ44jKt9Uwhk43bXpU4VZFEWTCGyxyV5TbRVG/GBj2psJRQGU4Fx
88lJFM9ZA4F5CF2m3mt0/YU7GTTTQUtny8TI7zCEfaj8GKxiUf8ijCZcN9kNRMBD
gMP4ju6/06i4/aXyKrstfu5tPhOVNJukDPwHZECEd4qw5pmUpUeXyDGnq0axbNi4
fTwjq0WeqP4PO9RE0/RdhmOr319jBR9fE4L/RD30wH/MD6lvIcqnrn3Zqx0RJmbw
CBd6L3lquMn9C+C80VhgTZ6JNZSdzoobxUBPufO6vpKi1hyfGixtE8+NpNOKgSqg
BkNJImtg3R59KZj3fEymi7H0OsZMhneT/jDt8hWeruVaA+6nZcqTb9GkDYHVB2Lk
d9TuOInB+8pffHuISKV/8TWBHs7L7S06fjR93vp6wl0V/ZihXva7Y1iIWL6gMK4p
3sIQMpyMi6I453xxzfnfY7zwaFYtTvB+g5nltMk2Hd6YvES83QL7vJFB14+p6e43
V0N7xlQDOxhpu7kQrej1De3nwDfLWRdIClMUqNWHYmyrJME765yFrvXJlJIIpsMQ
Ze9cNnnPCiaC+h/fcShspKjiUTqAxt6S2jXAnY/U18bz1717mWaJpJUYLAKB3/HC
ngx5VHqYGAfJJawF7Kw0LdHsTfaRb2c4qfSUBB2/YBgaAL9pMx6uZpiZCY75fsBO
EXSUrOJplBu4gwLPLhTrH1zrENXhkEsgVSumiJVFjDZhb3CX79SkMLjwNNKrqW+w
88LNTQcefM7ZUzIKzZv8WTrBo99hA4Qc56L9U2BYEBM8ewC1VW/VGKhSZr/acJ8C
if8zz6mFXzLhuuO4mRMWaxmBdCYodwCtdZf4e86it0qsOjlfIvG2h8w/0jfbptFU
ISVOVSuIbRct56RPjq6i0zeYlS217kLyUvXk9apVNdTg8/T3f45WNjg8pN3GJmfX
XxuIrH3y6AWDMFGgfuNynFhHinpk2lkTsbo2gg8LfOJrE+inOCAkEqD1lM0BOMsR
XOkg8uNW9KrbhyBFY9R+gDDReqd8tY7UYnYO3B5AV8hzbvnNTKQAwIQa5jcazaRj
dT2i2As8pWTO5T2hPVLbhZLGgB2FsN1qekB2XwllbuUNN3fCe87ahlnqjRdJXFhj
hPRiqoSL3rkNrdR/vqJhe6bpBAP5V3RXsJf8dTXUYcLJUjlWagGSmeLjYJhljOcL
Ma71wtylGa/78i+iNagXlbmYrk5scosk07G20kCMJarNNGGrbiaiTim5LqgVktBE
z1M5QEdT1sUYzyjdgaSygmy2kF5ox/5ea7rtuTlMPJ/uwwQwXjZ4Kh5t7j8PjznZ
y0XcoXdFLvlpdkyTMCxzeZViOkzs+sJnK3N43DxOsYZSUCpyLPXxF3cFYnSy7y/4
/RqPBTwRCJwnOdQwqzrbWNhBgHqnjGHpn9sqvRaO8r9AT3hKELDaVdVMek8uTvsg
zQcoH6zAsre5I13oLUfSddH85T696InQSwYZYbZz9wdwZton3hebRikxw1jxpGgs
Mqs0YHinQxILZ8tn/rngBjT64ZxKsn+jbSPTW8dB83q3ABwA9kwgiDoi8/RqvF+m
akGEC1w6Mf++l/NTjPNviCCymcXBwcfTC2YHxexVdanNrwMHj+VvTuXqYkZN+x7Z
77svxjRMDMluWsW9zwxF/FR3Wqdc2EnKQlgwtGILcOR+BNxUuIIMe+ozkX8Byx+D
w7nhMi2gf45Yj5iycTtAEy9B29HdpxR7ppLJ6Br8V1JT7wHYT2mdB7JhDLYN4WDR
/HNPQMQqyWBpnLzmqI8RPh41iOYkGysb6UDoMRzl2d1HXEQ02NSsY10frEvOuPq7
RUL8wia+jRcBuCFrZkOK1qUwCGJ2YjsgTtjMLSQIbJaq0mOtSobaEwe7G/Jm+pZK
E7lzTLQobPqXlUSrSEThIWL5bDXJHUVuMuFum1D+vo1UdagVMcG2WDoBlz6UOdXq
r85u7HK8q+Fz+tF0LwrZSqvCN8vnVR3S0vs+HPH0NRzId832OWL+C2MG4pDeSNjp
lqIZpX/VfPUHzxVkl3LXy8o1miIBNDWPfM7DtQXfZ/WrfGAsUCCtt4+0T6RHTtNZ
Jqz2FtahgDw4GRL+SYXIiTl75vfZaDByDbdsYazQg4KAPdpPOnP9DOHhZlTOG7pq
GPdY9gSPKltdqRP/ivGbFtlZQUjIIScb7hK27cw5LNw0y61lmrjjIlkJPYuk1Ezd
sPbgFxaEhGiesbNqlNe1LyL8icB2Q0sQRBjNNwtZQxRuuFxBXPYr9edVF6SsV0X5
8btjLS7Kzwo8ccpvOA7iHYbErYRl0yhASxbpfRjTgOuAmGOTpsnh+WRVwASTQc4V
Nn0S+ljM7rdzygiIJbRUxO0CwRQVaFwluIax0+GU4QvKGTm5cBawlmRPUScTGBYQ
6YK/1lkfg0AJ6vd3xJqIWADID5IXlsljoyBGZEksYqNsZAPsQ5Z541+esDx24k3n
gL6mh5NIQ0P0VaVaFiH/vIcOzXBrEx9QyZ4tYGBroLGZVgYg3dhMKHRl7gSOxs1y
N6i+tFHBROD79XR93P3ElgqrMsXmveXVSwUniPdkndPk+zVUsYOOyRFUo+GYIkZD
hVdh7TSe0faHPTdFz1+oTcRVz7rqOOoiNMXEA/kQgQJrNuPOT+Qf+VRRl6zUZOWx
IMDxloIqZuxZSGTEgee24jfEy4PNoulicof+1BtIv6X+ZqYOCV5OQUPoEpJHJpeJ
5/IjLi+8gcmGnvJCgxB2HKfRUunWmkWJUmsyH7NX1RKNdDl8rce6OiDiyhdlTu5R
imy/Lm+nJLJtGLo6u1rKaSE7WbPfzGZwpWCUfediyxKQM0RvOkGO1fgMtbC5aflA
xAR1JGsY77xbhymWNQCDJ++xVas3B0BSe7wC/7d1ixXR2B/eURw7Z8wjzpi3W9vJ
vsGunPXQt8ObajkImjBXjRup3JWdKsHPhyX7y+Letc2F8HjLvslZ+S/8qJoQ1t/H
psXjyJRSy40Svi+9wNkQ+FDwjdomTHA6QOVCb0Mz1X0tFIb9fd9KjwBDqygoYVGq
CeUnsXMbY2Abz0vdvf6r8qgxX3g1U7rnuqGkijndhPou2okew9GdpBrBqW4pIf9d
b/nvjvW34dIxsQ2n5aLUi9nfm7owytPRdmYq0M9wSLXsHsOA3qLWvv37M8ON5RXh
yLHUacsWS0obB+hwSHiqhSyPR/WOBX3mL43WaIRw6IVTP7oniJoF99SINg5MJXHI
caG5UWg8xR3X4mnG3JrhdDaeAkLls2DSItnI2k5Ex070qIyl+4fBNW3Z6cA/AYJN
rrzGO4721jN0pT51incmwAFSgi5MlTCV1JADgl0VruKFInmJ3dPGLoC9MB5/PLsk
OSIR3m5fMRCO1AJ8FDdxpU1aIj5cEFDpmTxCMHT6+JQqJe50wAoRJ4po+T+8gW/V
cn5uMMpFpy1tsbvmx4D5tZ77eJcYN0bWZTL5WkJ6SV2ga2lI567LsyrC0nADMwNa
CVPWSwk8c2iRT9MIC2Vw+qb6XyrzDJUrlJUBCxsogJaXgCa8TsR1mhPLZNwzTGLt
jPyF7VGUfSZRuviFa2QQGmdc8TntnkcCE7egJSKbauErokG7U5XrC39mJYekjWRf
AIKm9TrxIWFiKKyleO5GHCX/qIu0N+0lEaz3vORX0C7uBrVyehNlD5JHkpATyX5s
FIZ+1+WDb/iZ6IGKTEc8lM9aFltm/OhUajuFjYLonK/XF+xhgUU8RMUbQ0/bza4h
EBpvvjy8ZEHhf8pKraLWrUzaekef1X/rfaOBMrmnTVvBfU4AassXRTuFu4FhuGHX
EMTVszh6esfBUSXmJz6/8gX7ZJ/8aiWvo11xBgUm4AvOL7kADKodrHg2sFPq2fX6
8X14t+o1RWH4yUefwiVyhjz/ol5ZL10FDZdtzXaaVBs8xUSlia4tlBQZOGq7Ulq2
oaMhG+rnhz5/x2+KYfkccSntHRMujiOQDZZEGxVk19/eofjvsw4HVGlr4QclE4JZ
DqRQ8v5ieEYcUBJVYl6TMDu1+/M0l3kv/ghL/TwVxIXLyleHSBdPO2dEhXYfNS0w
Uc6ErToZMH9ZqMKvI+uYcKoVYcd693e109P0LSOwhBPdweb/4sdH/Sks2W/nSJTK
0uuJEFZlJ68Q9vjFlYjKJeY7cAZ6r9L2ezf17JzELltIhxvvfnQvgvd9LoAT+nN9
h5/yf34rjV3PF7vVEi1/skP09hunAJw2ab0paQJhfqsv4T+GzdUFazzmUhN8w8Tn
83oNxjc1p46Cm8OWZ79DKcyU6DCPv1DvKf2thcgbhNrSa33a+tl72Xq+dxtvZYg2
BWUXmgVaWQHxAcp1oSnPyl19L+pgAUf2eAAEGueFOZ0CMei0wEywUfgdtq4R42pt
wTzH+LAHPfiHJ9DEPwN6GspN4rjUVEy0J0L5IdnYwg4oVzR8ojzIOZ5HAuC/vEuv
AlNF7wdxgXGP2Oiw/l6vpTmr/0Zs2C3pZA37P1o0og/SAOsk8rTSM5H78pDbTC68
tQVr6vibyx1k6o2nw9OJjnvIazyiopNIBTYLX3a/EpLe0yEvjSwtUFKT0AN8ny1O
XdaNcF7Kmj4Y87mQW2zBfh9paGCZXmin301oPA8vaOUXETTc4+Uhsn0Uq6VDIwKa
+4ODjaHmzCZV1fF92htFyXs7GR3VtdOadA8eT2doYNQkgqmo3W5xiVYUltQ1LxFH
6sHCwhGWKEPpkM4nBQzNe1rvInTJMYTyOmNlNeoNemV7tgSxn3T5L3L7CsgzCOG/
6lXtNgIEfPtvbiRZiOyFNBlb491p4GDdodTlUhOZuHOYFZ1Mxbv51NpIqDwYbTSR
XhqiofrR36x3bIhNuJ4USlGgKfbCXAGM2iTtuPeSB1+ErB0/zR7fqvBSrcIoxOgY
/KochU17M0S7C5w5rVsiTTVtPiX7EivZEC+HTcfcNKMkRfoxPWy8bWs0fuqCDNyJ
VzC7TpBgJl763NJwxhLfO0JuKbrJne+gbAMGW507zWHKe4PKmv0V/KJUmB0rBQrO
APetezAtAK/YO318Hn6nl280gpoMitW65q/MeL6aT43jzTQ4OS5igoNEn4IhY5eB
+PLsSyKS3klBJULHlFbb9JUls34Q9fYsgP8q1BVqvBOg1BRxtLAlgU0gUaeLz/wC
/Bb7xpgspIZ17HutCCebWej75PHKus1l6lYLkHx9XOwv20zKPsmYCZH/9O8tfTHS
ju7cVkwlTsLnT8lJMlHDTb/k7WicPyJezwjMVzUprgteKOApd716t/qAqkGV+bKI
o9mIoe4TctZCrU2/08tY+WTCrS0k1VI7mNernmHm3nTopVdzOviVTwHlzjCLIu92
h2UdRWX591zf8aycsI9ekcoBGchzIqkAP/NoeCMPKmkp16NMEDCArhYsr0nBnBns
y0wauDnoSwEJBjDKntjDk7Di0a+gdQ0NUl36AoW478jZEte20JUiDqtD4t8qSLdG
8pRhBknXV6frAMCR8GRWfJXo+xmPy21t37zz87HCisJ3/UOi7May0db7Mpl0//ON
6sq693D68mYm2Y1EHkrR20uzFAppTdz8Pv0Cl9oAZRd4c3zALofXl9RZq3nQR7hG
03QeaaAhdw/0Q7JNGS/MjZnBpaMsv8EhndlNqkK3Lh4H9p6Ec/Kb0+oQp9rrO1+u
qiMIs8afXN5e+bnkJijaArheFzENycY0cZWJpnLc70oFi5+fbkSLyZGxySXKmKlR
aqrqYgU90io+W9/reyOB5BIywdguXo8oz4QDmG2Q1uby5RboZV5+Ch3fCNytJ/48
62+58ratlS8sETOVzGlq5ZEEfEa4zLuNY0v4Wi9Vj/lw7xwkAb5ZkEOsr3wUOK0Z
9wO3AISAbAiZHpQ6JDNjjEBgNb2oBmA7I5Ieg0qUaPByb65mK+nDEfU4NjPC3Sko
tZ/Bdeu6Q06YDLURXjYRIBakN2Q6YNkBNco0TdDLCLqE5IczYZCsEqxcMwtNce28
qEbIiR8Xw4gkqehrEyw12onSa/+nnnsX5IFLwwiy21qG8+pULHhk5VdPhdye8ijO
+lVvjRP5AXkjxN7uT/OKXhTsUtFJb10hYcJPEcYChjYTKU1gHuHviGL9ft+gTNay
fvhEMwCfti9YPfeham0CPT2zZEyXPjx7GcIjqBy1C2VIWwgo+iY3hYupVSVSOa9c
1U40QYt+5XdDdjFMmWQ0hLqzmw8VwKW5W6SDp/s3r8Wi2secVDDsrOzy0sW0hNsW
23j97GkCEjRVKjol0Kap7gXMNILL3dzfA2tvWX5fvpLrhjlBpUAJaKktOQuPJ/+P
L4KumkWb1XDcckAvLYsR12Zpr6UFoT88wIAH3qcSakSs/XU8Ss+GNzVFiCrpxmbu
BdsT7yUeptjVFqKhPCtAMxNL8u6hUPqPHPcfFK8F8BZsbLkOHHsZpwcVL+rwxvFw
EofLHaisT2k14WXVcNvuxyVgng6tyKPLP5Z777lnTipROaHstomLUlvGWotI9D8A
9gWWBcJRPJfKfTJFiep/hWU3v2L+mZB3+T5RL28GZukaFd/UXQBHB2GDFa83dyG0
tIsf7vwSZlexzzCh5unwNm7Sj/ldzggeWqmuiHkzcoSD0HeMDYFn408cxHj80qus
yzjrB2do06eZgg52lhs+1M0Z4aVU/7iersOJB7FPdafokKNSSMRUYd0CVn8k09ZH
bp+tGo4NU+OQTS/8qansyHkgj/DAkvb3/n5Ii4nxsPaOuHGRLqNH3YJ/RM/K/4Cy
Nq68vXzZC6mMqWs7MbYNumDH7iNAr4SUnrrQ1xANUwGIDHfXgib+EW+0kEDY8JcV
l1h9JonmjuzhNr/uh/H6Sop4ua93mJZfFdlzdbGcJhDwAyrpa86epAEhu6fmxNNH
X97m40t6AEsitL9RABEDVC7+Sk22ZuGaVmiQogQdNkp7C9Hcv+mJZp7jWd2tYljS
JmsC6K8uH+I4dFLe25tm34CXzFXcQBsl/M2A7QC0KXRJtDoNf0CxLLRITT9BjtNu
vCscU6iJTkY03SAI1Av6mKc358EHRrOlRuosVOP6CG+egWGdS06VGDcfKQUktD3n
XqIzi1xVoCvAoaot1zYrGksPoQBmp+aUZl9k127KKv+9hD77SBmET2KBuF+8HxJN
1IuwUAq9P/omaDCjqMtRm41ZjWRCGqpf13RFTO4cg8TqYZdZQsIT5T6WNCucTSz0
leT+Tn4QH+1QDZgkyTzZ6QNQJvPR9YzD/XtRl867cQh/a2ISzolSu/Ah0wT998kY
RrIk3nepmymdc5ve65w4IqedNLsMmEQFXLjsMuaOa7ZI3y4+6Mrs+OpEq72VDF+Q
q5YJ4xqwSBQagwbQWmTpviZpChyt50Ys9zZHBVToH+CbvZlbmQGp/7zyu1WynZk8
+en3xUh7Wz6a8DcDAojvJG+jQ4kRGGXsuvZ7PsU/2Stx/zB2Lke2HgS9wXIg5mtA
WUd81x9BEA1NAYyzRKVBdtpmuW3k7LnTWweFVr+geq0kDBvRe1So/XyYCUkQ98zP
PkEmK0ghPkvAzib2E2mjQSuQUurMl7nZ3BqAyOvHPFK2osyWEK6jjzD+1pah8Q3W
iIIVeZiYcFzUhvWCSF1FC3wXfKlX+hg8usA1uQo4gKzgrNkkX/kPjp+Qf5JxS2bl
20HIV2zAeRxSTzuTg49EuzM19tqnqbZHwX2k8FuXLZyGC2iHN/RgQepfLGTuly33
B9xrTFG30W7N6RtTiP3bncUseBhe/UGg1SL2101pCNiyjFv8YueiBeIPJpnD9jc4
bNxaG198Lczw4VP6SdOyn5tfW8H/DsHOCWHfSwu7pUbM1FH6RkZYEASUx/Ge5r6X
Tn+RbutYYhz4GnnAEcCZokRZQbQZUrlMPIWBnmmy8VBqliDBRCUFYghDTMmOMnT5
wz6UScp7gLy6dDSRKOBsu1AeGP2fxk2eaGxvC083PfqPxRCibiEmOwv3nX4iged5
1hIDrzbhA/jOXsHYG67yMjBx+AljEPjRc35axnfwX1K2sgXVh2Ob1b0Q7EW0ihdj
sxURj7BTUIqnhVzvC5yRsvLFtXvJY2LITB8b2dmsSn2jc6HcFplFrp8evxLvfDUr
Su47BkkYhgi5MjOTmlMOX2cJeLW3dn6u5dPJEq2Y8bYJTQIVeE5+OmijtuHbZcxw
r+scQWbnUhQYwggSdZirUBSDX6+egsXaGRC+3ALw6VR0xHFdC+U4DQd2ZJk5fAW3
0vDTTcD/DfmJ8fAzxxs9oZhYHYaSIDQEWgiS8kQUJzJ3CTHIkuOLbqZmHqCOJ6fG
WTnQOPl4mjV9FTK3E1JnV9zPT21wg7OK5QYcyFC3zt5/20TQ1YDe7ba/OClw/Ead
TlCU1v3jurit7L2wWCr54rbjnN68bttMIo3ZbUrA+XBC3jTEfwkREOxzgS01qhPB
dSaXENFznS4dP3k1e19Q+OkFScij0vEDiaTU/g5jTbf2vgVhTQ/eWsF7zkvpRtb3
vuupLsRdlukScW4fpMwE4+pP29z1/UVlXVI02MXNqUgSi/fVK7Tx6zxT5AxgGoDg
Z+rDWgRS93dSOgWXU9RUIg49q8gXMb7DrM2fmpESKHoOlAo5WnreEJxQ8LW2z8wP
X2xg7E//UmFrPKCcyxeVR4JbhpCI4TSpSG5mRuK3FZ89RlLgsWqJKpAKKqnoDO6F
cmoO6j0RK86x36wVLV8NlLvmNUtyXD8cIrRqBw65ImBvDc4F59yGSnZfNwDgg8QS
Q1Ka+DojGMCOBe8Cf912WPBYnIJV6X3sxoNCvzb5awna+M5XrWrxLjX2EDYWCsIS
4fSJml8L6wmatk/VquuF0+Zyaxzr9xd3QaESAI6r6evpHNqstG7f9ZpLpPo4PnDo
KGuD4TAsrRSgqk1Hv8YFIr6e1lkNln74Hj31nnmkhhynrxfmm00bA0UYiGD4td/p
uvzJWBuwv588zIC3Xq6WRn2yxkXPbW094HqLtWdTxwBoYMYNK7DW+hRn+GnjojUi
SAuBKzvNgVoc/71Drl3WZ9l6OygzS3ZiUg6L21eOBa/7Opcv/S9cxnloWNECWfBE
BUR6LpC+3Z1dKwg6cJypzGU3u1L7JQvZ86PVsLHLr8DWxr6xZmv+c+bXcfykk+yz
5wZBYPFocEgj7wZUpa6mFs9LjViG2V7prvJlJb5tsETyj0bN4ylGRNWmzEPT75eE
gTcQk0QBmTLJZYhPBgPHTWWLs9Vg+2dzcyM8YHQ+Kpw1T0pHscHBbIZYXVHmAR72
qc3cBvN1g2VgnaIfmqYZ2Lo9r8+RfKYoNVPMLlVbIAenDn7XXN8qrdb3QJupk+0/
DM408a963HV/+u3aV6qTeK4DJsvdHFGQN9Q4EzWWbgYz2KouP6T/ekj3I6NgDAhw
qORW8o+nthWSCfTVzu92RilMA1goo7BIEoo05FNiS0vRgIsjQGhTDEyYroldTV+o
viaTK8vUWRDZGCooSj/HsZ92TTi42HWzRqBGOaEWPBS944vVSeQnviox4/6fa7P6
OVu3BpufoITanZ6eg6YkD06rGKJ+OR7R4wt05EolXU/CcyYNDpWEuBMC8P1j9LgY
NdYXuD8m+zs8AwYTRLg2FyznIDkOWpNRhr7i1ncJqQ9D1JPx6wrmd4zqo8nI48+O
BsWMHtYUTA/N1Zunv1dnAbzm006m3OgKhSJN/+ZE3OtssUzwRe5YSK4ht2eOC946
D2aKpAIIOZPilj6tNTrKV8xgDywkwrILBUweAEXaV7B7At5Bck631mVKK6P4i1RE
5o+hQ6atM+x/qn/kX+OkyGWiLeEbke5dKs6aCpb8GyAs/4dN5cavYBWM5X8f9pcL
9KD/PRlKy2jPJTaU9ycQHLVOMV7IqZOldG4+qTJAGeZIwPZ2f77ZLLKB1zWJS/kw
314KsGXKb2fRJkkg1eMM+hxvOrvuHOAfp3N3i1efi5xR0KfvF5lUtXPEZyc9Adyk
EYMEpFEaznNEfbowfNLb5KzWWJHq30Oiq5xxejMz4kir3MV9SecNUKeVDgZpNt3k
rrs73Pt0Cpw06VrOTOqv4E5+0xFo8UZ3pfsi8lMtk+2V90bFyG2J5ltefuImJ0NG
wOPRw4QZYMWkXRLKS2DZRrfvc+WLpIudjxQ8nVczF51tQNpwUUZctLI6GyaxtYTx
gopyxwe300MWYgPgnEBLoiuz7qc+/vXZldPNrxIyzPx7j2QNycqnm1s3gOyFKsmz
G0GCvPlzlEXcke5KF/HLJMeUWkHxFuTzI0wTWbXg5KWUJwlvKRPs0q0qSkQw594k
/AsRqdWqZCFtJDmLSAp6aMKk5wBJh+ZGDNtCv9o4L2wEvCVPk7gVLA2Oy3QoLHin
Ebi/SO7uYHdaFLdUZ0SgwicejSwOEE8Pmq1j+hDYSkqRQcTssMHMA9gf+DKlUtNh
w4v5wZ3i8ELmUbOmEXjC5rhL/UGooWTfYox9Ikh6Gu3AD9TDJ1rA+jGuQZlft9sV
ZUp5GiSPaCF+KITmKctIx4k0AsmGr6TG5zjWmMO98TV6GUd1hABBa+wA2vVGQ27z
JE5CUki73+lZNMH4vJAieKp7yJWnQcjq4CAEdyZcHwMjWXpLGlJ/6bqgFtTOJNae
cP554aYdUSiqVJfOvmyhWUyDudN6pa1+sWfFstTSqkLqOrIWvxnF5dMjWdDoHNrV
YHEr+P5hdLGEoBiCdU1o1AhdNSo0UMc5EiQpEQXrYO6hbC+vqeSn6EsiAD+XrTUr
f9R75G+JAd1FihuRp4y7ffqjwaXzIFBAIAulUcZvc/U+ImLiZujkUiO3DYnYIu3o
WuGlbhTT2ErWlqQGXWwMNCtnpW6gvNIswaHcOU6sD4ZmpGYTlJTPKA0cccoH+Tr2
9q9L/b3KWmDrn9cXENzt4emJ5AzA8B7aoNrEm0ep804qEtzncmvvgAWpR61uni7i
0BIcHleND/7P1MinLonNH0Mh7lvyX3vFm5XXg2AsIFcLOTKNfrmG/fp9W/N+yHME
G4NByV2m6Fe6WMCaDKLo8Z73zCfMdP8kazXqJgJksNx0e31sbVqNKt0y5juz5xcV
8396m2zRng8MzgOSdhPeEn6lwYcsheDJ8C5LpsHmiq5dZDs7QE8uG7zuYdlt2yql
UOj5Tm6qaLXkYacHmGuRo61Igus4w3m/h0PeHQh6Sg4a3afM0bPZanzFe1qQ1h0h
W8FbIdFuaVXheDu1VVOXxS7xxAgkiLGNwDkjWw5hBRvLXKM6b5Gfjt67QnDPaWHV
eNQHevoMv/fu1YjwNGEynuf3UE3ndlTRWmY0QBMjnmMawLuPP0Bs9PeNqQsG8FaU
M3KSwxRYbqrye2lh9GJuXt4U672XG6c8XO+46Tej01ZxfTyyCCg9NCJud11EYagN
A64GF0iYjKlPEMSannKkKQ4F3EZa1CepdLG6LYTOcjdcEKtnWWLTEyr2WMldLtaj
DHaxh79FZcBUblbAKJgI2ezZ/sDvwQL2zvOneYZTcrd8vDHKKnmgw7fb9C3TUSBZ
e6YFrm52cJZ50adKuhtVuLUZp3fIQNqM0kBmEn6eERhw/1AWsupBPbpl0toalN5Q
rGKoOvuVoKk9WvwCG+8uT6vneho08WyXEx/NgOMM6FilyTeddN85ug3+Ugt/uqUX
ct9gN/hyH3Bs10bsE2efQnkNFmk3ZJryLO5Y2VPoC3KG/28tLp4on4Rr8AuxzmAU
SJYSnm7QPa8nCCgcXl5JqOOknfR0ErY1y96M6c9Gk1tGnu48/ssFl/57jT3VYSmE
/LSg0njBCkDL+1q4RwohXAd4Jh1iCXcgTir+s/Vha66NAAq0kQETO/wsO9uJkk66
5qOyFXwRfCKrALP6dkRiJf/X5bhD5FV1/YeknA8GYl45PbX5N37mmFfyP7330eV9
lH78porqE6C9UG91oQ5386c2TTwe6Ep/Zb3pTOHTHhcpIg1exPriYUHeJgvwDj+l
fAxr7qSL9pebSlcyHRVEyX1eonnTEF7wK6XoHWO+6HHLbLoShhH5JIvVn3a/vZvt
+qu30MJ0HK29pIUEk6lZY6638amhAy0kK5GEwnJDJdJIlYR3QaDF+FE/T4DbL9/f
oZrDsciglZUcB4ZZ077t1aYZuQCyI1uMpBtA2M2aW1Ie8kBCSgl5fsYjuW+ANjOE
NIll5IbKExdt4UZaHzbYznGAQl4hxQeBXQOLKtseFewAJ3TCy3EG/XEfmNgEqmlk
IY6YoIWo01kHIk0ZZSniRdSuy2CkWhWZlZW7p5iikmGo9LLNXus9u6UHCNyu4JhY
NbQrxg5eSQL7MoElkgpa7+y6/wbQEg41J/ZAa0D3D5C0dZctJkv/h9ZZvbPXHIMB
M7GGHgCK2iwC6JqH4JTgjlvneh4kLEXVpeCYiyqesike6ufLRtz7rDy/FLmrx8XY
qPZRtBYS3aF/fdlqd2v9BAQivSFiITxqYjJ4o2omllB3o+EkN8Kq8pgazM76na3d
kh1YzHiG4AmC3nkRkLTWfGABbqWbKnAMpKxjcWzw6auWlBEmvYSPuBQGLBEY6MHb
jcHcK28UtLvU2biW6QKTt73s74KVkgll6DePmua9MvMyVbIg1KeyO5+ViFRkUSTC
bzZp39cK6i1pgULembHYwBbfQpOOn7wR5patNB/wAoeNYkbmBm+6P926lQCkC1Hp
2LfDQZ03fhqFbQ79WP0lhhaFnmfqt7QUX1+4twtZ7jHtVwhJtMLfqRKO4mgppN4J
yuU//d28s1G+USfmS2aCgZOHpX5/K4XgO1+X+JVwgc9SDXhd398GOMFPBhfd2Lkq
SzYAOklYCLPi7cCYdFOy0g0exiipke5DXjfwyv04cgZ3T7kCanjsAL2AyfMn+CG4
JvPgPWlP8axIDACPo2Lt/kwKlzf8qLBUGu/vsOP9Q8JGclVhDnbL9UpquGQvXa+O
TyqK5mMW4qe+oXBBfBZCbLJSH6kzCT9xmetw6IS95jLMKZfXKJg+1MnwS5ncUdFJ
fN3u/9Xj/IDDkJqHiFCFgXKoRt+C3asr1RVaDMecYJZPOXEg1L1tKnbbWUrWs+wY
Z2gCcUEv274Dkr/Jen4RnuPiSQqEWnIykLnhQ9Y+h6y1L8L3vLE7H3/FVfOxj4E7
9ndBD0B2njMT1z/Wdq7uS6v0xmQnQulWnyZtwcAFUGuqBaxYRhbONAWe5WUHSWJb
jOoVkn3eM4D2BiCDbsqx7ewPUnHsCWBV0aGuZgS8aPWAa17vf0d9TXOWUTaehxdR
JLKt9dV3Y4vPfS2EMUJ7qPkL1WFjnJ59J9xvFq5VmKtgcoafmri0PwYCYzwRZmB2
uwSiq2lRbhL1Gh4PF3hcSkBSUeeimzazpWy6JR8UAHu7bAKF9A869mkouiAwTTsj
cIBQQDYylzqzdZnmdChxb1Kev+S2MvZFOTtvyqDQ2CFToCbf9ZkUhC0DJFACL5mN
FtljMzVv08rsb0bbxyjPz0UjZQpvou3xh5bo4q/fYKmxW1UAOBeWE7R6qU7hZsJK
F2Rn30+qQxO11j7zW4ZEFREKSftNGbUEd7Spd6PSlgLgRXXHRsIHmqj/yIa+lGj+
0yhVry/1D8dh465Ubx7O8/JqiMDO5EOuwn7qiP2FCg5qO1ZD6CE1FWmp81RdHyFC
oY3XHz2LuzG8e8mrk90QIFL7bEUHKOVoRusmtcNQc0d4NhoW1u6LBU8GXVReorwj
JytETmQPaszC/rLnDwOJqYLKFjnyF7/5EoBz/0YOEfu5z2AzWdm5T3B3K02PSL3i
cxmQQWEthX3ijlQTqZ0ThMDTuLiyIxBVw8/FyVfV6XVJiyBTtckkGn6eaFu9Y5qY
e7jVhMfKTvGDTr+ke71XpmePsbKTvcQPRlDeViTf+umUVmrlHdLcYxA14z93giT+
wkY2W+pnCks5Dyzm5Dxl4h5LwZ0mZCwiuQii6LhqQKcF5e/9AxQYQxIRBWjpVXpI
0fpH6n/2c8F1YA0K61UQ3zqd2AwwngmM3gvw2uqejEEMBaXkZgmLjRAX+NbQ4srb
J1fLXJXfAI5ryn94EXL469CVnnCBVn601LDtvi5WyqdwhA3IHmJ1chz7y0wTDkjh
6D9PTMvETyC8aaQW8Flp3fiYmX/7susA6qjkYrEcn1mI1ELd0DcEwaMRnxRYJI5B
g1E4SfBw2ynIgpufzT5LVu/NgMiGe5IRE0iSdPqnnYu+wItw0lfQeVKIYaleFYDC
/ycgZTvcjkLmtkcNguNZYlMKRIfJIDspzmm3HKuz16oZQBamGamRFlMIMSolWsiH
Vl6at6HKDm6gtZmxe8Ecsi9oAxGrEtKc0InIzyKvT1z/x0nmFd8zIiOjzjVMW6XY
q7nzJiyfm8JazELKxfIjpFirxiwEdudKH3BI3HgbfRahfuj/U3WJ1Sa9Ha43LkjQ
tkRO99S/YsuYDk/jtfvL7mmCMnZLCTq0lo6UQBon5ZyG3bF9pciaLsTzdaHq82pP
2/UMM8kGMY8JDDeg4J/rTziP3Dmn0rE6M8g7VZAvXOiAVBMqzC8QRsoMpmVM7Q4p
v7goyz79fX+fwCoLDrpMnWjd3mJiCO3Lw4wO6Rske39ZYAsSxd524LXQzerN1MgS
/KEUjN4mw/Ot0oxmbZgdcRaX1xs1TNakEGb1bG7uChrABijBXN8HVXFviuDUpzB0
djhktQ7iCzi+XSwraazAbLKWBYZXLtGpPl8qMbsWD/B8wEQ1PrY1ZtlCJAKX9LE1
im3f1ya29LWyrT/70sRgv310PKqBK4BFzEfGmIAobZEwIpEap42xvbAyZg8JD4sW
WfuC3/s4rlY6MLjw09cQigXbF0Ft0iCtrKNPinmB+ix6r7vw7cC6h6u+l6inH5oa
sYYBAw0dkJsYmHm4ZPRI2GlEEZfMFHDaXSyX3JxOAul7Roo6eoHw0fVKXPxl3LfC
Wbdf0gyHNK+mGPBS6USZ96ZcCDvdFrHpOabr9jiz1pMvIX6ELjam7gXdPTIU9Ano
GdUvisByDImbqlY2TFNRVqcV5F1q7SGL8NI6MUDhSVPsrS6UwgaDDCo7zz2d8B2w
c9KlZawhhwNyYEunHRL1KesOs1eipnnd+fy6yBcRA11Jysz1ei+/SL7qwt2ucUXV
FYtuU5sW/IvDMs7dUiSJJwkh+KMEtqbW7Q+9esrwl57rxCjSBKCVugl+6B04WeW7
ajT8r72DDD7ivm9mra9C5ah0QyetMP12v3YG2byno7jTdhwl/QQTOHMXUePry2Tc
q7z/MASIpt/iBBnw3alw24L0NBgl2qnvs+udLT2yr7kgY3/cRVkNf5v7vA103Ev2
AZDOpAU7DTVhxpFeoXOqlPNtsiINaAiZiOgIvPuEGm/LONlrpeY/b5TgT36tOnjj
+bON+DU/T+wLdaZYCZcqUnQaizoun6o3muqDaXUPXSZIRMo0zepehRHXsgnaah5/
hQyXrDQBI05vgwq/e9AlISidVSvy82nZlV4WwhX5n1Y7ptkvzh3nCtLw/jFaR/LB
PBGJm1rt0II5OmuewOJh1DcHHolF8RbZY6mDf9MytHPTFVvxe8rT2REUGy9SexWj
HjxdM4E8cvRN+iAHfqHygqtztbYUcGShlWxSXkqOYHwuE7sGVVJ9TQG2c3w+uUQ3
7lAw+eGLiYa59F9kPwE2t0k9bla1OQrFu4Um2E8tU/Nefe9nRL8ssOybxUyuJSMq
J4g+pvEFFqe+9kSD7O5k5l4B+uABkTLO1VwzgwIQ30z3rmtZEIH4mMpHcVSTjx0Q
ASWsKXqBj8miKsEwb8v43yHA8tBrkUZFKPaNjKRfPNnNxhOgQjeYC9gIsHOvfbBl
j8T6kMpiRvTJUQRNhBCoSSVXIl3YEEyu34pYpYbpoaTiGQQMhEuoBoX06NRUL+5f
GZycPePsE2QGe/lIXrh6k2m3tEpmVla1boxwiqVMUsAcwFxufPbR29eE+uYawuE1
SVmvVr+ee5SZY1j4FNcU0PMzwC0oDzJmi6vUhhSuVb3gOSRpcdhr/TysxFRvGY3g
DFUhd+Y0j4lYDsiyy8vJeQeJDPkLqcaVRQv8vbgnc+n2JulMNslRPH65HyMPWk6P
eBDMUjpKKcqttrSnNrBUPiTYPeJDURkU39CRu1cBifX9vdEgtVNqrawFhYR5mKJ/
Aj+OQGhcYZTXVIMszAr7mFVQzJr28D8oyvlQN5YmkYbCA3MiGUQmmQuMw9xbK0G9
tArCFi2vmjF31UimRrRiMOq9OFMnKLzmUT7XjvytKjorHNzB21xopqduiwnYn5oY
toZJpHirTil+cHJnTysywS8NcsMnM7PfRjhFVRQlMnHh1jd3dK6DvSbw74dxwK5y
ncbdJzjz3ytk75FYFeom/5+IThoga4KPZGmKfGROHRL1BBhp7dVEkZ+swF37uTBI
L02SwrBnLT3R6KS845jAoxS5zbOaARLYnc7gTDRn2A6mnWOL4+eIo550KoExJfQl
MBUcjcKhhElQrkQA/ASNI+oKJs6bw8UX+zBjjOtylz2EbrBmH/yk40xChLJzZBIV
hrN3C5pg8/Mf2W4ucECniUWnygBjNUg8DI/Y6lA/GJ+vigK9FMb4w3Y4WFHfVpr/
l3+7he2QVA5CjJvYBaiilBoxzBDROQ2jrrZQIs2TcKunVFLDcKQCmcGRalaQBzkb
fxrGRkRNnBtJdvx04CIRflqUb0rqWgWoffjtDDW1PUPP9TxP24+5+FgQkyCCLauy
RtjqePRpcXL01/SM8l/U4Y4EIB7FUY+GSOyMA/hhqFIYQ7YwDDTxZr0xQ7lc9SQj
qSXjhguPJ4uiMpRgdBGjRhi8yInVbWHaQY9L4d78HtoDU4mW84TneGMdtZAkOdT7
M0Jm60xzXyY3OTkrNWJYQu1aQpo7tJz/h/PWXIg3mzGLm/GJ7TabqJbss6XJP6am
r1hMHrMgUVXiPUnp3hJ8F45QylqhivPKuf8/bE8Z9l60FeQj1RWDGvGMMDuyzBEo
3TXmrIphN8Zmzq3190ljDABCPb6rmIK5TQHG1Bm79rByhv9nu9otfVbkW4ZQ+aa5
Si7kSOjS8ap8CnK9ptvvMXCwY2/9lJswMZediCtLs9cDyI9S3Vq5Ytrnk0cZxdQ2
P1M/PkZC25OguazbCpuukAcE5lgJS+M0H9Wqem/gyRahiydq5avsUT131fPx3dDZ
0Ym/Dt9+v9K0Z0mN0jCi0xnAZOPVyAPo1NXOOdlzd5iVxkqi3kz37duhJiKjgeva
+B/J9+XwJ0zvszLu1i0sqLR7RZJPz0+oHmFy0AY5fJN1wMb9xf3aJPUbOG5qOoCv
voeLYO9VwcV6G/dx69wRQpOteCjiBqNvYAtU60OrceE2+f/HDo+T2mUWbuD5UfS1
OaaYvFiB161lfpGFrjusoU5JzTahsLPCVkJpGJt2loZO3Ltoj0BQB4U2sOwoNqEf
tVbyt+GUMNZ0utoWFDVKM8zqGBm1tC5VcCeLAZkoI50w+sf3jLpW/hx7mE/WJluZ
dj2lTJM+XDD2bcjM5dsLt6UFplvjFogjV03jhRNl6MWXBLEuiQ7LoF+XoZa0dDGJ
AmuUR8LcqWwdrNML7emIkgjk79/ENC3DZELLsBcVxRjyYdgFPdX885YQrYxIYB9O
iLrAE4K96zJr+S/c/4s6+5YXtlpRpKVGxSr5YifUjVZwqEJhPXdtcynVJgCRri7J
7YvwhKUKF5s8Yh97Hpe2S7o4ZdfjeG0UOLUHihKFoHHzapHt52cf+SmE01MaFEhn
15HmIHoOl4Rlm+SNKEzo34WAZeLVE0F0TpYmt8elrMl5BZTbJRe/p+ltFsJkNWME
n9xddYdpNr10EM/G/Q7NIZ7gFi2dzEF3bd/BWC9t5mMZR6Ny2wde3Frem0kD6EfL
z0bODKIVtaWktMWtpw9wMZMfxBiqFsNxMzKCMguhYvHcIebddZI/IZqMtbexjGEI
Ve8OX7i9z9FXlvXMJT8/0TXjXq85RqaSV6Esc3R8AWonv40/7Jy9tCTCsfocgDQh
E93gLrwmoKRXWL+4afJvrl4oWeZ/g4mMlM9COa3Xa5lZ57f0D/N5+bhrP5jZidM2
k1wPfpTyfVW0P3b1FPJ7Od+Ars+/ic6pIsWmn+CiGSkVwiIc7aqScF2dm8dvIi1/
fxM1mfdMpjDt9I1644Ki1Ivr61cQdy0WQx//WXPDNLjj+VvwS7rhzdM72Ad8E7rM
0jDPaijd/gVcfddsaRWPIc2tBOICGuBnA9nrszfwR/NZ0Q8k33lMrUU7DHRvlpaP
6Op53kZK9sTRESgO8QjOBj4hv+GNH6coo10R5C3I2L0RGXQZftCB8/WQKet18EeU
`pragma protect end_protected
