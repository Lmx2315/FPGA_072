// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:36:47 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
qGSHh3oPq5b0zd77pPGqbEjyts7Z/DUaJH7cwE8HKtk+9j7zMDtjr65LWcjwe+rH
pXzrfK1ugbh9P1q1/ZMDVqwY7611rdQsRjosUyRYAu58OfR7dOpSk965Mrvjxyly
2n/JC97b0xtfiYt9bc08YiZYG8chtwCMoRwiC6ZGhWs=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 10960)
Nz/0N7rRpFksPV95hw2bwlivaUmS/mBdcw2pCdtdC+kFbDgLAP+148VGL8C6ZZ0W
n8yNsYr/r1PwQjoeGNB0GEB16vtT9ZqtntLXLeWp40Y1o5G2PDBBrl4wZe0G+BRR
SqLIkAYzr1wasNJLTdxKOs8CYExSPKnCCL/WsJG7UFq+PH+aqpK1L5FM7D/QIxtZ
Z9cIf2U7GiXSIM/yM80WJ9aiRnFBiHJ9WvkuR+X5cydDPNitCFgYDYkTU5gBZdV+
79qVDRXRZQ5HweSs0g91NdxXsSSNmQei3DLYw+vKXvEwTJU2ii8ADbdVsqBpqgRk
PMZuyi+xuazSA+J+Ya8nOn3HYLT6KWS7SjGc5i2qvAnwlu+/3y4f3rjxUSz7Ti1m
Sh/xyrVQuJ/KS3m18WeRLlbWO9bw5D02PQNVMZg/RnjjoPbfYLl4shIzSXDb+jUZ
c8dHpcFbbL8DwEeuZjylqx+MhgknKpZv7lBoZfZiMRFUyqT6Y+p4JCyFs0ZERiQc
3e65gJLwmmN2eD90IJUhxFboVVp0xybmgRIhlnLwCHD/oLVgLCXn/uGNlD5qLFXR
BqSMVM4TVYwAYQu4e86A9fqUiQ+ms44hJYpz2hfPG+tNheNBAphsd710lr1k6Lyi
LxaejmK4KbvrFhjUepS3m1uppsPVhcqYp0gsWv65r/tthTNRoAdG8puoBstk58Dx
XhJ/J+VZ7d15bA0diIrOrwoQa/YY00EdcAbWKDvvp+AxCgmt6iVS1ytMCoHxn1MV
QVqRkjZdXZt9F8qE6869nMzr77RFM9npuZHN+vcd0krMQoGqwcMglk8h9JINTBbX
UKz+WlVeL1wgiQVgQRZiXrK7Br6MLJLtQy1Wo0edoDwqIHce1JVhBJk76eRaa+a6
MWgbMXKb37rsOeG2woHegM7OOTe4Ogmuibz4HeE49VOFTWGfquV1sXCikYoIusSC
UnMS3y5aRjcFql9wYmHFlpxIlySU0pvcU57ptHZyUhPvJwM64JDvt0JiGIPw6aS6
7Xt0NEoKsFiWqJAnG55hbbqWgRvD7yuNTP+42c3s8f43PhUamkHqdy9wWmK2NoUd
7ZfFClyEkSupHg8lmPRQi2Jy6fYQ1SH5bQA2SBOSa5RRdR8486Zvvakbjuh7yhWE
HYpiyzENFnTIFgSFZPp7x4TAwaVqO00ftNReLM7wqHulJWp+pxD3h6F7Uac4hrD7
b++HaGoq5qoYvtD1rf6AWSAAyqZwc2VhMPHSJfYpfdM60LuCk2ObRInyLpRd3f+a
YmBxYBgXutsxc1R0ncmq3OhLfcoWJlyeo+p6CNZJh48Bx9sh49zPVeG08mulB8uo
9sLkEtH7a6yj4/1NQIXuKwuWHmBupbQtmid3lXLq7Nxy1NuU01MzonM5sbgAkp6/
cVtrJg5T5R5f87LOxVWF+erq8P9bxOh66TuIe7yRumfrxW2LzI49bnPclBOsyaoN
fB5Ipm/8XXDH17jEny2KMqctXwfkOReH9ce6wBnIh/2L8LcR6Qt4PUSLysm45Gpc
lOtEnQyxYhd4ppDpOpFZRqvjGOlZK5YFRNA1pKKyZGaB7HLiCRqtB3mVIk6/8Hq9
1t9ZrhyDNTE8FhEGOGMZsLRlYUJrn6HTthHtEacsgk6xvzIYLKFGKI9+tGFp3jza
4LVSIFJibZBo5fXolsAFIbCyy4Vi/SSdwyz9XIp5HxGN2fPDiJXj4ibCMFAgi0zP
88BQv25f0GpVeOBQYVFR0NwYIHL5oUEG6KI6dLNkgShE76T81w5NSvXTm7pUDB/Y
utF9zUS584mhHIP2qGEYmpx8kRrOZqJO+2U6qOPdvIDSxReJe7z6JlN4a6BaaBmv
/9/XUGYZWhb8qIKnpFBngL5wygbo9twul8yXOCHXct3s0UeWOoN8aO0ZpNAto9n9
TQOIbKVityWtZm3ZdWY05HtBIQV3v0NtMzQ1OM98OU/85LhVD0f1yVx2TDKyF/wd
233vcmKp3r8hRbYutEuJoaET/Cv7QBbIPDfABYsPakQVg2G8wT2a2W3sckuUA9/+
2Sx/zl9V/iGe40kQclrx2/KEY5xBAOmZzs9u0me7rcYPLEzPZdudc1aL2BKBYpu5
U2myH/9HN0fKnJOWDged+tAeHWzrIa0ntkQOMIpdMvyAgIz5gSzj7ElSNgoOgezE
sY54A4Uj1+wunlMR+rQKCohAnjLOh2OCmAwQ609y3QrGWRPDBBcrukiPNuboqk4K
LqSsG+HWlpkqRCFrP9ZQHCU6276a37lct5WnUG4Xh5J1ep30QkVBmWmv9MockNk+
1gKJTDcF4mtvqOjvkj9/Ctyvs1wLYy3y/4Cv+i5ou6GseMET2N6iIAVaROPIKQsY
mSGQ9x9JLOwENMarkbxkZ+e8WBBKl/9/fiVTNbWaK7hqyalOHNypZDkUlHTIoXxn
YX7oLomz6nlpE/uMDj1bLGfTkrMgkQVnaOHX816Gaf4kF5HrJch/t8yQBRdU5EfU
etijF5o2nn838cbizM5pF3SciP4cIBEVJPXm8raBd/rkIlkvMXjhDyoWJJ6EVfjk
wZL/BViAXqNiHW4LqCRzB9/XNfIvYvA7hQrF0fD9xe2G4+l5/4lLXAhDws+FVsiu
XHyrFVOIA0IB2sHCmi7mPVlNB+v8r7QiX4rYpPag1vp/16LUZc21QlccDaeRlrDK
pmgWKUmufKlB4ZwkTJnQREQScBH9nCSmT5hqeOWLF158hALa/o/OVQmnGDp+aHvC
ldiWEvZ2F6+StkWmP9axMSoj7NDtBo2EpU4tRxs2aTNceVFTevF6iHJyjGsZvbbZ
itfsYbJWnHMFeVct1yMNeE4H0/OEZ7Fd0kcx0gNCwR8xAkEu1zLcPIRIkHOdsIDS
kQIMx7ZKdT/EwhuUM/6rSfm2HOGNJWYfl8g5yNRpMxfAV2n9eEKQOcng6uFcDnxE
oWSwPLLCsRylvE7LOZp61hmsMVdQuH0qnw2MwNom5Q3BGbOD4VEPKw1BJRlh0qG0
U1qkW92l2EP0V09eZjbhLxznug7rNqsaEQ8wGrIorS6PoQruChBl+ukmeCkrlDi0
HtcpA6hQ/IcLuQHmpW49iwkFpqpKewb/PjwZg4/VQnxge3yysfHgHTcqp7iHKOMX
ZV9zT6O3YCMc7n9d0qCzpA9EVsC7RmEFJzqvZ8vWE3pAiHbmeTkul2VcoqFsYFPL
08VYPE5+JtUrwKgISr5n7N7jVC01snaUbjnyKtpy9T2naQjWGOCv8N4afbQLyDMv
I7Tnz3Sbn5xZrOCD/jOeVvq1pa+bZ49nS+BcNOEpGrfmwMNyMQdSv4EBsor6qt5Z
tYoi1l264IUZsVwpKsw7wOnvDcGltRKyxyVP1wz6BF0MNVe+IMoH52o2Bk459C4E
+Ke1uI4r8hy0if08d3sp2MdBiL6RrfVYovaI3i3bUX87/CbP8DE6b4UM+iZV6ziv
7cEa41sCuYZ6eD2q1r+W1PMOjOHlgh3wYeLDuFF4U+a+KuFZQIfNoT+NcJtmbhq9
IyQv/3n3viGbi8G4zpeIgwD40dGBp4mLSx7SOCAt7xLK0TR9L0n8xwEmz9dYhqTT
5T73Nv2/jJhymvVjQPtlT8i+4R0tH1xaGdCG0BfEbqxEJaBGZ/bUSF2SvybYNlLZ
Skw9dOPiKFUQRBbYEbYRl9oN/PiigF9s8kXLJLglmvx5yiKjOKpgZB9B5hVcbHNh
cduQA7No8+Y7dhype8chk6P0CM0NlZKnWoBLqk3NBjORFGAy63atou5MJoyx9nrw
+nN+c8tZNuKFn8jlp7UfAvUsvD8c6WAzLdJ6cmmN2Q7YzvTNzKmWrEKD3SQ3+A/I
pj4I/vkHCrP0l64AcxItU8YyP0UEQF65hN2yFmYjrlfwL+ieDD7DVhVJkKdI0jhk
Lztw5bsP0ftX84HeLbaFhnY2Yk3h3bf2HmKW2H2Tf1M8jsA6ExHZaINgNOiTE4if
wMwAXZte2tjakOjjA/YmLkWRjqNJfsjlruHzd5z0IV0J8UznvzKpPv1F9iBs+Slq
O92O2mrGGJFP0QfZvFUQpQTtTzAUsFrNGuMMS8E72n6fNjwtQUzoz/0tW7YMTUrX
shYOiJrLDVnz64K8OCSDbK5qYx30kIWWmMbtkuQIYFyUk6gUd31gECzapecqJsX7
ZMbk+3m7DGkRobXVqNr4YJTjYO46gDSpFvIJIl/DiXVLkAFnigB7KaShIfyB9S4H
F0CCLIPgqjGqUf6F+wl9Zj5TxTYDIeuBFmZqc6Qexr59hSGPScTtTzVu0w6SHpiC
8zakaA9qMneWPvbmIoUWcloaC8oaWJsJas8mOt1aFx6ddj5qjlqIvekDiGJLSRFl
9P6QefNZYcWDzZ8IsS8aGF0hCmNbdp/Ou591+hdZYLrCnw1UYLDLfraEIazhltqb
K5AGaWGRqiNr06v84UKqvKIgV14TZ8ShE1Ap+UGSUKR9n94bTkz2ErUvMFNcqTuD
4A8ZteaF1rCp+mnQ+3T8xaeH+G4d9sSRSPHdbiO7R6K7HMANIb+4FqukXO7R3WEl
Ps/TQ98pQcmZpe9QYBzA8+5T3tFtJfdfH3leQr6167Gw3L5Rsqwo07axaUO3MdhG
Fsk2u+0j6GfmXChpQb+z17bS6Ez4MzabtDBZIfN7yzGzSTSewkn/QWJ5QSWJvO1m
ixybR5D9puuJe9Hyuwl4kfQQCQbEXC9iwe2lCgjNggYk54WCgdXF9i0vzpJC8Zrb
u4s8ciraJapT1oTFwl+hy2w8NCGk4rTN980pwMTeHTSaAgcYiRawupIl02wEx9PJ
VkmxMSoG/6i6eDfD4l2bIOJ1Vaaq4llcuxpX1wQOySvcLPIkFn2SrpmBGZbt3A2r
+OeiJXdhVGY+LxUZQf/EMdveMzNc1Zd5X7xPxMhx4VUUdo8NPM3sYUHprhNLld3w
+gN+fK8Icx7HmOe/OV21SbMePq0GcTva8wDGpUp2z/RYKz3IonEFFOCo2yU8SMFQ
xAry+jSfKBuZSTyQ7yKSLmojVZSseQZFAxc7XIsJQ4KMkJqc4FW0tV2SkrwlK+/k
jMPEGOqUBjyrXj0RL31j11bTRnuyeeYtY8h9zNmo4qlA+g2iIG6wrON39xIm0+OH
m1NABV8/oaKaO8md1VnrbIL+zyqdkMhvK3K7MFqifpi65oEy/wg3R9QvMcoF9iJ+
7gJ2hcP7vpjHrBIgeb8i4SXMaF7O3VokVS1nMgGH72sL9jt8EVQimS1cVQaMusa/
1L6HGUGETFcxPsF5mjhHuOkzE9i9Did9csC+CLf2MMV0pBZd+pI3jzlcrQ0nFIFX
RZALNBLEN7nr6iKk6vvPyicXdMYaMZr30fVO+IaN5DFaVDWZnAthwMK5QR1/q9sx
AaGIdzFFANluL+WA9+o0h9MfO6kSP0SdlkLYt7dsSTd85KdGPSmDjhqvip14M1uY
bbCiZ9SkU8OK+yO6/rsfP2WUcUOW6Y8xEM+4XV1v1K2HOL84wyyWfp0+5hxDmgdb
Y/cPlTtx2dy6yVeg6HNDXGZVRjNDpLAjwqUcCLowIeDbodUXzUJU/78vCoDqzxhQ
MRcZ6VK+DF1LGVv8RQq+CYuSblx4FfQVTfUFZ6AUpEUQOvaicGmRUQY7RcnT8eLz
rUqVE2gTqAFk3qM8ljV77cYo/WbbP3VZ/tMNdj2/C+adEv3D2pqhPiNSKFe5CdZD
l2YpkGtC/5gFphOdIFI4KPpWyjqFb9Q5/JIg8VuV4M6vtfhhAIO9mTIt4y3bsdlz
pYC510h9KBcT5mHHMaazVtVNc1G4Jon+Q1XYxzB1odwFgqec26kpLYkFVxHR79eM
nQ9cf9M2lC+UGvSQiJOjSos/rtnrYwSveIVO/aBguTUEZU0UNyEw5VkhFkylHS2f
sg0NU+JdUkR1NTCLyMd0pFXaqFho5ufWCXMbnsvX1hmGjO0aufaZPzTJYy2twM5B
F3rMQ99ZSwwzC45W9uB3d1cIsEsdVBjtYH5Yzo0Ix5Uhl1p/ibB8HEo/XzOweNll
FerDsC7Od2ie2ZtdHvIOB9AqcjapFUJ3bKoYfMVTmq2Sfl0oGn3DK4OuorxesxDv
y6v9jh6ciu+I+gIhIwI1vlHTUVtxsMxcrZg18w2czry3kKdDJxYFpznns9gvZ4+9
ybnVrF8DVGgYz58lulbJfedYeDUazTBwlGYwXcSvwiMoV+PejHG6GORo0GmuQ58F
U2VgR5GUo+8DXoA8QCtrsJeK2LB9JL0lzESEip3i57FoKMIbbJM0duAr8yJ0p3ST
ANFlvridtAvKP4MOwL9sgEm/qwaL63zoB+kldpXyCHGgKqvjzz6RYy8cwDfq6/PF
Wb1CciQ9pvaXwm4kgLalHouoTEcwJdsbryhnQwSYkKRpemcITZerHvR5jR/FdBNI
8+9EZzSo6WSfVL76xcr6icOG53765RIFRUADZwB0P3e7N/Nzq6PGXfPtHIn8rarq
pIefLPp6b+aYvw0b3LW07JnNXsKoJl8C7fz7lYkAhjBKiFB7XCVYxa6vzB6RKKid
kO6o1LNHvuL9o8LQTWdDYDk8LxWBDZdzK5Oiomlo35f9piHmvw2p+ABadJXOKsxA
CnYDKv0b9gf7nNa0eIW8A0aOA46TBO6H6HeoBIEGFPOVGjG6Uo3GICCN9AWhYL+d
sVz4zfnyKui8F1yRPQPc7xEHpNofjkkGi4SpKfLRdvQtUuMPKvRINVq3nTyZl6OB
EPmFnF++Prr9HS1nXEBSu+CGmg18YM55gV82Kg9dQ/PRdgJ5k8/f3u8ysd8QbB7k
ODpgpJyMtOWGLGLD/tUlGqHQL+KZbRy60l9TgriqIoqJrVwO5aNGptuAA0Fu5L+4
SLm9T7vvxsAKWkpYZy95saBK+8E/IrjAV/fr84SRqs31i1xwL8O7DdJicjrg4Jfa
z8IvUldgcjUL0QVRC4bCjS3xBhNMYUzT5vs1f9SzmZtSFX5Jd0nCHwveYeF6qA6m
6iJJkiTFpe64GwUCHiLqcnFnYBrlmzLtqMPM8NX7nrCRkULgJSwDeb9XfbKkPQL3
bps4pX+DqSwjXXXb6m86PmW7clUkcbz3wpCdBM0Kx0SfDLkNyhWd76p3rh9RqVtU
ZwZi208hHZ89Y9iY64cwi2IHeb5IVVkLRQc/rS9yPfoEZgsQZKBzd1rIJlehsPvR
QjJGYwFqsQwz0X8+oiFb2J8X5U/Nh9k5ml55qeYJiM3y3+5D1R2bSVwi1p/C54G1
7kbmEreyatbM+sXwxnLkTH2xuSaXQJ4rhNc3SBf98KsmIhazRFO8wrGJYPc/AU0K
0K1qFpIROM7F3ZNUaINMBK7gicqJWYFYhonZ6KeKyI3dUFRahRMeZ646HVKgNmca
qix9N3dZXgOU86hJ/I5Wwi7rb5b/vx831BujYAyYXgCyJ4nRTwVlbxQPLem9KpTO
7IRve22hfOQ1nCrzvnG9rBSeCOHcs1p4XzMJY6jtv3SuDGAHJIGhrc8QvT7iWu8P
mfHonMnlfjpMsKzABJSJFEBQ/zh/4tsHIlLTyQI1gA3oXlV7DNwzXyRw462JKyox
HWthzlj/zQ9zxEo6OMBp60fwCh8oCTRMzz6K+QBwglq7Gv1Jmi91HUY8cfm1YhQk
024wKUDdHZnKaVBFk0KBw4g/Z55kNx2xFnQ33pnMtDxQ0LkJAqxvp2lc5lddqyX8
XbWhMeXMp3v55/Q+rk+naTqg6rVsOYIP6BsOWnivxgxDAu1n1uCYXNo+BUXf2vC3
/xHQp8KnC5Wg7G17NKVUJ+hxqVb9Py3eOmxIEU0Y+Y1nc71vmpqyXThTqvVw6lse
Y2NB5sVT9OwW+jFm6fJU2nUNloU2jn/dDRhNbMNKX2asVB1xwsZUk1LiY7dSs7WP
SsKCgw2lCFO/fallNSnkZ6WKjOATU5KdvO5FFp8SaYcX6paWGvLtDwtSNKqRoA/J
408f3RFdvfXZrVwGmgbeYtdxjsxBj9iH/2gFTi7GZ/txD/1TpycqxQ5f3c/SF6m1
Zey6TPVugLORMJuz87IbYoVGtZq4YR3/7tQX0kewrKKKblv4Vhng0c3zsOvWskCq
tRrb+V/VEYoVHmWa0Zpj9076HEjllUmGBqGnYAtb4HzleodPrvDauUT52KaXss/g
LnBlpnapVm2UhO8NtxHRe2CfaOtoT9VquRwnPpcnymtIilTlAyv3l9cnJSxNBCdM
xfVH1vyyDoUzi4W4x3WtCVcn5RQDSUP+KAuJhfLdgi8cjNSAe1rxIBpoymCHmo4I
9OdZKNy164t87zgl/lRSJWAfV3r7rFLpkV8ksJDJk2M6v13Zd+paUa6xCBupSHjy
ZsBEb+HIu5N9W0MJjQTdu9P2lv+hAOI3zlnmJeuwJ7DwKVCtN79ZVTBlg5IE0NUe
ltW8A6X0UoQl6m+1lZoz1zXLhI7kZELQCJJrZpUcwBavvhR3NqIiOezQA0IXX3Bv
PS+YGgGxHEzWBrqDum2CUX8TxCZJz101QAp9gHC/18oS5RvWwFDG42vpiyK1DlP1
tIF4QNXHNkna72Fv5OQTBHJ4OYoIVc+J7FLBVGsGte6SYIl8rBF1DzxI/6UeSr00
lDDhkf1dArre5297zouMN6hDjsT2oSudUvPdzp/Zl+UlplQiT3qWGVL+JdkKYt7V
tJLiu8WSo98CH5d8dEvR1VVhEfujLb5lFyazMHOotoIh+zOWFUaRARlZtYoMWFLy
L0senik3kXLS5erNq4HoomN/olouMhanPbf2AzQALaovSOcoY6HtnCl9nPas1J+b
0z30fhkkICW5LyJdOgT6r/aT+IaluTC9bOEMQis/T/qALQUSJSRTTRnBZjnDa9Dv
GWDOsz4/MSiFIvrVSVzdYJtbufdpI828n79I8CoIMDY4gSCGyD01oq2fcfIc8ftw
JE/JmSfu8o/6c93ZRAUzdP44M3uBmDa1bzcQiTIfDlb9C3/cJu9Ey4ckEucOV+VE
/pEmNder8DnCgmh4+zqXKaDOjsW7i7kZ9jnIF1n+VrLI+Gc8yYNj2Ki2bK3ZSBe/
gy5vJV7mFb6l/c7d4wp/XOFNERWc9bK5fvxi3FychEPt1B0EK27cGx+USRdygyUD
cgxhgrHxNmWoazvO+yfcicW+AG4J+ki+v1+U3k4/CU6Z6XMFhWsAP340WBub0vO+
r5Wf5CLOhU/l5uTNZBThAn/iW28141jQ4jMmwfyUVe4EJKiq7E+kzVt+WVE2LAFf
qLsZFbqV8YzQClDFPPPfB/VhkEhIniIfG0bKdm4K4sLUKIVnP+eJeuKQEN2/hxh6
bPMqibL6ILLi4SkFpc72Ku48yc6IV+Rhhbh/W9jXoyNNQGjM2FKTPuvCUdmI+IXJ
8GjdJadsQSUQEOvsx2YRGhcY68VC8KVDMP6qeHySrZurVJVw9o8RRD9zQFYBrHGD
6IL4w6RZXd0g0laE3r4hvh4pfXYXT9f6NDsNBVHrRshp54FTVzI3/Tp9+VCicR/m
vOpHi1suap41RTctMael8afaCNZG5h3BR/K22rIq4mUDBaJr0Yvil+mqExsweEOo
QU8oL+SjNpwO4qB1COmCfj7VPuL/fXtyEUmuwP/MgAc4E1zS8KFvN9LSvn0Okv2d
U8mGg6Xhvhz71qhw8Rl0s/2rngpTFOcqWAVNZ/lRLNSoubEi7ZrOgwSBUvQQ71Bk
6A5lK6sl50Qkpgve1mtIaWjE3AA8JlNqJieQsJ/PY1ebkha7fyCITlFku0BDBVwY
+zeWQg8HYb/63EI3dBegba0Bp7LHeKXcPuG24/CM6Hso+vBkYZXnf+2ZWwph1cjU
XpGKQCodvjNOycSHiadS3gopVuzmkC0kATnd1/pNyQxAge+A9OB/MAYLtqNqAPOa
bfJ1qUw1wFQPhAyJll5Ye8/Hgv/Q0HPgpbF9gENJgkcCyd5LsWE3PuSJpl4e6LWm
GPXISSgQnNV5Z91cscq58eRkg5lZvrfq/iEPfIn0g7bOVSHg+tEOI1opPhTaKDgx
h9GqG7/Px7A7ZWUTuHl3YeBgmaRYZc44G/YddEcjTUZ0hMjb2m3txRxAf5sid1qh
GJOgIH3hJhSXrpO5KafvhLuFDvGADDOUXS6QWblLYIwNfYPkuO72ki/QLz5cJkX2
dgYjg1sU/ssgDabgrMy5UbxP0LdjUUdeVFCj1XzvYVJc0GZGhGnpjICRTuCop+6j
RgiYT2CKEGkydJ+HUyEWTg3PmbIWohCN00+3Zf7tTb9muTuZ8cb4jk1m+WrFJd0J
S32tbDc/yggcHp54lHlqe+bGMXxBWIWpOaBHOkCGwA4K6lrNi4xa+0WLie4+vq1l
UjGh8FkvLkSJIyF7z+A3yNBTORSLFJOBPhjEqQBMVKhHWA8ms+EUHnIysq4PXrQi
kkp81n3L5b8yN3dlsm/vwLLSwcLPgr8t2rEwJgxG3Tl0JuiLwTCGFpis5Q27U2Ak
WdAka56TftXdg6GbxzlPA6ZLeEl2Yfdi9xwAYwJGK+mZimndYEnZZLLkuVSZk47k
ArMsBmqVYRjZN9ZfZDCktznvshnoqjNHS35fdZZMxi0Mv3nRFS3BdhOG/7YvOTAc
ZlWB+BkF8LF1LmTW8nEDnDXB8AYVESnYSg1+f5gBYIt+94NcGoMeayy0w8Lqie3v
SnfAJGI4s9H57B91hlGomraiOlSkgohT1PVgRW7TYnurmo0ikR62N9O19Ml+7uYb
FxFlwbnmjD8b35lVoN/VBilxVeFPgFKGHoSKO956NR7zqj7FH+eNy1LiMC+Pp/iT
H05omML9O0FBq/37vD0Hq5ooNojs05NfwsMJpTYTlJT9SbH0QCd2hu4bxxowZbmy
4vN78uYkueXWHP5i4bZ+Zt3DO7YneA/NIj4AWQjLfYNAwni3ZBZR9nkZOeiBt8jl
PouHQGMXNJrirVDMDMa72jVIlvmVauQq55jlUhiySBV835APYM2fjBUTlcqPh2Gy
hXPzn4wqTcAkD1KAJAk0XgDPLzxoXV3DGrJ9iFdOssMqhz0tGe9zpU8VV9hDIB7p
UB4mLCnIeuv7aQwSDmcrRQeo4EzzY9mypqC9kfqw/f1eqaqEh7XT7LeUCxW3Jnwp
YeNBSG3pFYGjC2jwgMxl1k2wFXBDZ1veBavA6x6UXgcyKD1WH2y/L73NGhJ+rBsQ
j4D6JgCG+3t2fGTF91XZbil0cO3qGyN/KMjs4CP3raNKz9tsXm32oh5CtT0kLUVV
dP3o06+oeQBXpLEjPYMNIWXP7a7U0C1sdQgHUxF1hsSY3hLuZXbCMpGgX5tJCOAR
269SNqtcAB3LcxQpd1kiDrCdGO6nvtQXYnLAccs0T6GSJ/dCoMyMvFEoQQP0WTo2
6NysMUu2Min3FjQtqPbYIzv5N97rEKzUoW4RQyx1AO7kVH0oxgURfath+SX6fls0
1qoKmLHyq47zcnwLRwqR39RIDkhUxK7s9Jr7o4+jx2sL2iIosyM8mPWwny0vtFzL
xSs1TZTBFc8eQ98wtIHXZCYEm74mJZV/G98XeZwOOGnpE9AanjwxiwD827N7Ctm4
gerSoJUlRzot8Iw2aSzacTE6i6PMELZU3wmOrX/VjyEpQ1Ja2tmwJulAf38OHkGM
VNTFvoyPlwllgQoHugcjJKs684SirzcVDKzre5toyuSPSnnlr0hKqs3KxkkMdxFW
b6wFE4cCiZMMTDBaE7yJtSryyjkCij3bbFQ/9SfWIPBiPe+XLRtDSgKj4u5ZoY0q
nEgaAEWCOyv6C8DrRwWWEKWG1XMbqWv4vo2giNskcZmPIg7G9zRDG1N7+HhhIjg/
WlnV/duENWn5QzPG+68gwAwPqMVuTc+NkfGxCkKKBdeHHccvnBtCe6ZxfZR0ypl3
ONQBB3Asp+z6/+LrkrS0WbrfirjrhkHu036QXnWPj4CV9k2Hj9Sxz7JTTFtt1NM2
gqvqYyVCx/zJ70lNns6cfZcFn4i2oJZAlqU7j4T2PZd1qlnF8/Bd0CciDrA2dm7w
GHf/edSMTFI6TmA9J/RHAYfkpcy7nEdal0Rfc+0sFbhvjVlSB812v59GUoHbU0SB
d28BY1ur89eLHR5A/DAaQNY2QlzBICiJNlcedV2FPXj/sywzyQkvLIhsiSy+jR0Y
H5jVj1CG/N32oGl/6sH8VeHHXodS+vH5TUxH7hTZPbMR6ZnxyamqRNQP5kxDtBvT
jGpvjI70pdkUwPTio0O87tk+/uVG7PTDHiemv26YHXHFKRHkacLS31LCsPUrNRsA
r4LlJK2gicmXR1ZgoOLpVKHXKAX0XdF/fFdtRZZYbAmqPnpze9UMHP60oPQ9dkMZ
NGViiGtpMfVYvPQOkC14VMwaTo/wHrllI1WIqAIU8JUEnmyaa2TQOhU6oStbv/wD
JTXyq7S/gPVUunmzQMj/MGFgy/2LQ/vWKDbqCVr/qH4MANAS1/7nN35VWLTD7cSS
+B7q3so3Mc8rWqvRDtEZFK/6OBiC5MG/m3WiR7DsV+SBxDmDDXn9zRnpmvD8TnNV
4zBd7fuenlgTOIsCjgWWc9WiHzVydzK0rXguab+ae7NP4+ffFApE3IrZwIV2KyOv
v5HSxz5GzkCZZpAKtqEead8DUNC0+lGbF0YiBqk2Tz8G9P1ZekGcZhinorMBXvza
v+rQqf9h+LxQWBcccPExkFNIOs/oFLYW9O/UeLbKcpVyWO6fRYzn645mtJ4J8RUi
yPcmaywHjl1uPP5r+znvBl7PHsjgsZO/VITgJxJB64hoYpqBHrlr4BLKYR3q1WSM
zze1O/f4XkK+YeQ7lJ933jo+yp1Jw214hH1aw1MpGmLwXn1BeEizC3JD0AW5m4u7
lzrfWTdGTyJ2oPrKoweCKLUGDiCnz0gDylEIZmpAzDGpiNZ7Gt5jKFGWS0hL3PZj
7a/W/rA7RtubjEvYy8vdyD54r2EcbPgWUOzhcm7hXNm9wI/XlwiFPze5pF9R87m2
5g8nMGesNIpNS9gix8RQT4Pee/3MyHwcjpDZ3+wzc5hTiDIT1Ou/J4E0EbZo2tWY
RtncoHxbm/FXIx+cUt3ZUWmdwPMXVLjQbPLiXzawAjd5G7l7R/Y4RuzNKayXdSZz
sVhQdkFVkk8rFjkCjiXy8R/RdaZMURFS18TDXhGuV4EIpeDAisqfqopkM6LAdFAT
0s4hkkibzmSv9FhoqP99/QL79VU4OtfJWz0rjJE/l7gbSP4BL78mqgEZy7VQ8Mob
aV46B7yy3CJIDk9eRPmM2HiyJ+Dxc4IDIat+Gv7HzKomOuvPJXjBL8F2ajyxnW86
SJAAW/f0LyN1cut9dSvVJP+zp2F/bPsg4MMJ6Z1nnSAOd4Hi0ltqS/JSwY5CATTQ
O4+HoojrqsPBYbS7Tc1YgPegMzFmP0QzWVF+BdiBJkR/DpI+Io+rbV5tyAiVVz4o
/1RtJKTxu98H9Pyv1FMFV776HCKK4lN1iez6ZmrpFZ/WXsjzQOGIOmd9uTQpypv7
9uWxPnHaWJ7p+6BADLLaUSNjFXfZzGdH+fT80r95bO9tGg7q7PKj8orTKP0wHMv6
FwWG6pzwa69lDgqXTNlpx5pB9Ej9NRsTRqvIaCgkLNx+Mu46Cx6do8gESPByKntf
ZlWikgx8s8ybMo7V5eGoHn/zYmYzW+mekjlwlLKwJ5nzTvXc14K3WPEbdgaWW0mo
rTkCFjgAeBpzElzLf6QYdHpESChQ4mOCF7rf/gBqexPyMUXwP0hUPZX+enc8nck3
aMvotItqGCMnhGtA0MZYzWtVhWRIsGX2huWwMeHIE1oJq73Wr+tcQ5XvnrH1Vdlz
rhp8cDmIVkCW/mvYf9lRmOWamodVs5usrv17LxTXLZKAluumXbJZ495NMSB8ma8m
/eLIDE5DEVxiOTcgco0c4TA1MYGEL0jkY6WwenByAyPOTEHHd3pA2ycMUxLZSxd5
AI7bYrPba7MJ1vCKhXAP1W9gZpXdYHubmmvliTYCcOaokDLUkJPqyKz+He9yWkvv
Qyy7cbTOhuFwyakTZpD8Mzg/I2I91AKFKWw8BJA+cXdb8XsCzyJIL84TLqQnbxDe
9pAw0qSKWFbjHRfuwbuLN4I9HRXCreE9JeACCbaiwq68zbPAxQRsQDv4sFfZfxMI
UfWI2hZx3pjfVL0YWs/MX4///Jqaa5gtaICLFG875IlXEQhwipRdE5QRD8hmWg17
HG3BKlQzPYuMQWxFfi+keoChIm14LxD4ezaFTtZkISMeAlBBs+0en8F0pQ7j17f6
6cc9rCRmYuRxugaq+h4cpyWa0TupL7rI3HxynDsGHWDrzDKocKARXpzA7la2g1Mf
mwrUTQ18sb37YM0vi3AewYttIx68P3750nhl4ic9XJZg7e5sjya74MDORwgmXolm
CcA8eD+dK5DEmgW++Iy4Us2xJ2w0QJPRkg2qdOfYU0ZGmKInHzOeCGJ2LaSZOzU0
XrKA/ne/8GRx7QkW5+wVwKIqk02II/WY4bttf5smz0t2ooffQLesJl1f1igclaO9
TSriRoYTntwjsU7a62wr/G2p9eOaf2Ibsf8v8fWc7Vbyv2x5wfqAg5gpxcFvHoJm
QI8w7+JS2HfqOIeyQ1IlAG2w1DXU+c8VJMCBAOYTzEnPRIIV65qD21c5ECVeJMDL
FSmxXFuGj9r+emzdjnYduw==
`pragma protect end_protected
