// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:37:06 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
HDTa0n72WzbvocYmDpEYNLcf4OoPHts/oh3vy2wd715FhnqNU3Iqifc8H/y5QgRS
u3FNFS83MHQZuGLW5q4gIo+abES2NVkOOC8P//AjIOHgW9sopjbNaFksbfa256bk
oFDb4WdpXX2/WdN4W36QwPniZO6bDY7z+SQV60HjDW0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3104)
giJUsAmX+Z3mp03sZ42whGn/MzvLxigJEJry58cSYKl6GaDIFsc1GQaNXFiU3H6U
1Ciwi1iWpbcCwh//7r0h7kOYxf5rr9MjQUQKfksKm6AX92oNBI17Uer+OYlOD3wT
IA7J5hw0vP0QNH3qP78qvF8Wmh2qeQl5XIVLoHY/8bj5c87Y8+u/ywLBKlw4L7qq
yK8fh7V82QwNtd/wIfuTBYcxMn/G1ZwMJOKnhHtjM/zI1ifwBfEUkB1/1yxg3GhX
KfLBUBz68JGJzy8TMzOoNvBEorys174ZQ+UECWFCDnyqNs0euxL/nro669dehpq6
7G+ZRXkMJJoDbtm/S9Imvg+kKbJChj2KZdooOBiqyM/SnJ4kc+u35dD0GyFjHS+m
eRkK0TFe29Ewv17Cl6A77mkXtTiTIlZ6YaLxMhl3d5RclBwaQMSHQuq75J3ex+zt
2Opw6Y7bQuFg4yWPP44XXzSKxAtLxSALME6QUiMPsiz1tKu5Cqt5LLsPJRdkVkQB
r3T3eUZBBh6B0O36P6jx+jeOyRVUDvc1NKhcJ9ldb1zRdJgTglIkKnu9GXb4DpkF
yKATSj4bA2I6rxjUv6GrB3GOvoqwBd2kcjXCjtqdBN2Zv1E86ek4r5qlMyTuky1t
yDJyn0AiuPFPGo6yqblr6NenVVAgDn1gdHfvvbW7L+FeK2fqzJiuuV42cVgqhlmJ
1lZiaIkuCbSl6cCHvDUtqoAhbVVTPRJT6JYQaQwdHT9fZElQ1jVyN89bdnwIxn1W
xZbJwCAYZOg0Igqg7GsOzhoEhUcl8Lb8r/wmC+QKK7RmmQK/KQSf5QuAyRHgnO6V
OSBYXGR9yMfboQOhvdyg+9MqX2JTfzb+khV/rUA6ZKSBDKElzhYfODnmmKPEnplD
y/hAP/auc+dVsxBkXS/vYlNn62x9GJo3b30FIAjucdqvwVwwMAOlfHj4DK0SjiIZ
AkFcsY1crlB+vgayCPbIrNW6xGlvbValfdoq+MDIr+Wl9me9Krq+5wHfRN0/AXU8
z4uUfo1W3yg77JYUlPpLd2pV2DyTJnjVz2f21U9iYGHDCnLZ6BXpw4l15QwjWuwb
kif5syEPbxGQlvaYtUk4o8SfV29zMwYpHd7d/4EQtYNxJdPJ2lbYT3F7AFYLpsWF
hrBt7NVviEoknUOWfXMKvwBW/D+NhjJ5FumvXxbawAaKkOE2F29mwGVx6r66izm1
0OwdpAGRFvayYXXmUscWXE3c2Lfzd7XDVk1E301WNprflxaSnINQIMzNB6148drt
QitPIjxlBEKxRrLr5wGUlUs8REhDMJ+1dY94992p0awNuRCiVJ/CeoVYUijjM3RJ
o2Q/1KyAfcOJHPnbKmJX9WktHdhvSVPc5p0RdksRRWd1tNdtNGpqSyXhkRQXJJMb
k9yugaXMIHck60Egw4aJizz4W/BaJiMdkvwPXMCK9fcenvAsYwmw86OkuqVFGAs7
pjkkEDPzyezcLfMv8xpKr39gsE9B4HVIraewBOC0UWuRrefgJlg7RK7MyjHA87xb
heJMdiBz22cwyT2F+WVEvxvoFY4DuqbSw1OMPV84Bz3ZLfLRPEA3XfT0nkLVDiga
s3OUKebsPvRymf8mkZzcGHcZI0NQIWkBnWWJupPArkldb0F+TglBHUUgEjWhQsYp
z2JQ1pfB0IR/eVgSryzxE3hScbgNm9NBI7/6tlu2ZAkZtLepeZPK6T/6S2R2ARTy
GN34dLHn6iYQz5hrJ4k2IC71RoqGH1Tnb51odehihu5jwghRK5FAUVQL52NZmRYr
u04aS3YPB+SgXf+sPpM6Xb4JrAF8dEfrw5qXLY8UG93gl41Jl39FTOXF7ooXPqm/
JfL1QpXKScO8oZQS8I05LH7gsgu+UNUiBNgFAFjXf2MTUzx3+qqMhscHfWVyi7VK
Nh5nYy7aH3jOfw3psGy31urRfwLihsQVNtpIV53LYMikKsuNNdO3LdxxwRGnspY4
n5l6mCIyNGXNWPGqxGZ5Kb1+BcYW+pnuQQx3sSTBqKAzcIChZA1NlLrLZHCihbZr
IVu+QcqlRmOij6zqwV8ZXcKh1v7WXBNPrTATKp5/0qOpRHfp2mik1QTB1tM1A5h9
EavIuQUsc7PIU8fGMgZ/LuWJ/5f4E5g5FvvmA9g99lPURCTsAnH8P/hjqAZ/NqlT
S2nqI5kiFa+bSIyXQ1cJULYWoBS12gUISNbovtghZ/zFp3hhbgQWUbcKbk9YMhNO
U50lafz6g+zyokric+/e15se3JOwA5TC8ZYWOBA1tnkw35VuccsXk76IZagHWYdC
J+sJB0Jx6FfvGZAKaE87eWBsRmt9oCeepIQA9rlxASVUkBePT3ZajkjX/f0wc3wr
W/vZxe1bUUVVw+o7RHPbiHfi6Lrw5EeGz1xVY/cJRnZ5MNesfgJF5t5BhYxaN+Q/
kjBY8BEpta056QFdqhszlsOVsy7L8hf1+G8pydA/KTM2riT7OgFDAkyIXRwVgRiJ
P8fuurGUF5ECQM/BxilUqwyrY6pOUXIxQQeTqzoOzzEnc7tE1BhznzZInlf0cMNM
ZmOl052tvsCsx+Eu4TpuDFLkOhk2LO8yTJmi0Ls5Mq2kYsanB41RldRWy0C+0O1L
Ok/hfqXeEFa1VgTE1GNo5aKMrQaa2/pcOLTfu3/q3hMHmQJuFYv919FZnQqIH5Ea
2EZTwyuMETouJpGsdEh6mMSEHt+O0y/Wy55mn8VbLuUTicxzwljs0OIBZST/NyJx
nbFIVbjaQTUeAPDLvcbqTldJjhC6b691Qe7HFspRnZ/eQXtuOfcNCO/KwYB8i6aw
S4r3mi4Q5yCCRpC7XPWuFmmM8+CkK29cmTr6C7Y/UKdyDVyZHe7r300ODvRtx59Z
ag3ZS7Nr35wGyzkU2sBaqiBiRBDrMiR91VA6aPztYvyP2HUWWTbb2vdZDmA6oJBw
rlSFNHlYjEGLYdGY2x/7XuXAH7zEr2d1NZXSoruAG1HIWCoA64G9DHYJv5Amzm/+
m6YgLvibmIXUS/k2lpJDsCpIfdpz8XJehVKNJqm1tw69zzK3MduMUedhO6lK5uU8
U/XMO7sgBJ5HubcNR/m0HGJaU3reKBnp+Y38W+Su+0YChS8MBKcbmseDmdWFYW9S
XBp8BL7UZdEOJ4PpzKoRbhu1RV9P+qhGpV9xuzg88+aX+7Fi9xoRwJwVGtmOS7rV
EupSDIbe8V/wF2ooXz5lEFf7TF33C+EtYSTfz1t6tTWgz8ledWcavhFyKD7CgEHh
5E5PSPAy7O84DMkKEL1JdULvUCy3QZ2AQXFFhyBhCJsb6Xkivp5ZkxFXsIxEahC4
zPeVbKtUorDGWRAr/ejLgjxkLRQwkA8eMBfmpc97YIzZAO3Go/fjrxfCPGY+m4U7
+xWQNmD8/a7GjGDyMUxlsPMeVAd3+Ubxx5d8/+LsEPihyLhaEeAFhucc3Iwn60qk
Dklmy2xeGpFABvMm1fpJaWuwEcDj0x99DQ4oybPUN3Q4qNdNJIea0XHcGSnXmHvQ
bI2elR8ZpC/HVgxYpZVS2KwgpMyOxCTFq/ITTcmOTuoIlkXHja+CTpAseGHcZT5o
z6JYvNADKZqg/4vPgqti1uEglOQ7DqUesDRFoWEdXYPx2YMK1AM5B7Un1GGDK0e0
LkX4PBzg6sI97HmhbYzRKtjIYhOOz+TcSvPGH44Tewjnj5MQvYbrh6WGeEvGqGnm
29a/7F6JYQZz/fpQ3f16HrSdBTgPg3T78982JCsz8DdTQpHwM26or4yI/ExBiRKE
ONgV0al39v8APDimCT7aulKOwIURig6ljErfhMo1XKOl5BJG5y1vxUKK9Add4XkQ
BB+oGoNCpoMthlslWMu83JWWKA6YICR5mdmr5QiOlBNBWJ9Js4kv6QtltyMjknOz
U1uwf8JW4hW1XJmT+IC2SEPIrLCMX1/6gSyg3GszsGQVMLghOkVDVUlHAl9gBGAe
yuLRuwjzONDJyWN5DJk2PI47erRtSVE+Ah2BSRQUrxqA1WHxWt4QVFUTYysyNZsO
N7OXtb/TWUTPBkaqKwlzzzKfwusQfkuhQ3q3EL8QwZPX4NBH1XjCrqQ42Gjgd9R+
A+6phHXxVe/IFpg/Y807TnJ7C8QiQLs8HcC8GZ8Jqs4=
`pragma protect end_protected
