// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:36:46 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
DVQzAy/j0l5TTpcZ2E0dCb18GvX2eAUAXAmBhWt/3aENe1tWVBybqKFa1makmTjk
CsrEnfV6XD3oU+0KrB1d1JbSMI4OTjoFocjyDTx5J0wDNt1FX5P1+tFXcQplbhnA
XlTZU/ooN3rRW4Jz4hs3Cu8ko+sCH85M6IpAPTXFcf8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5648)
ChrGbI9wBFxiHT2wzWiFJ5zhZFvnrYfB2IfvvmdTJwoO/122XePJOZYw1eOfLNgw
Jycav577qvT91LrxSii3QYrAJIYsSXCMXCFWHbDrNtkbqtgXSsI55d5ij3xgOsY7
Ss53VQ4wkq2y7Ch5jFODeLHdhnwDSiOEBTJOcVFP2nxBKv4fCu9vGmEQiH6a/l5L
cQQ5X/N+lxElJPTeoPH5mD1iZqZj8Ki8OZweh3QPDmgbVdp4zgW1xNzAV1dgSfrs
XPwpzhd15rlPc9fLdafTIJgvFWa1xEUBWOp9iINEAe58uw2KTHdvaNJ3UMbhjZ/G
mo8mN2uK/HZysjjnUIQAGDI1oM/PlgbqUKuDtj7D6j3QPR9BjsCF5NEg305lx1u+
j3saVR9ZVYe0VPEidlJfBq8h4SWpKFS0NoAXe/GOPBH9lBVI9uFZFUdaU9F7aNAk
AO920SOUQDc2iHr1tTbp+m7WIuLUf7gNqsIKnPUpNx1ccU7v1yh4Qd4SWMYbBPZc
2A/tig+NQ/hX6tKrz30EZ9lkW7fQIiXWxutU+9+97KSG/5yEMJfAXBnDJ/Ghf/i7
saIMsy+JtDJmf8TNt60aVEQiouSbx/B4X5nLRgPwDKQfaCRS2UYUv6pa2jAc0M1t
S0Fg+WUnJxMXRoY+hiTHvWYhoaFfKbrwYKDbrUD2SJzgt8ybrQBsYxsvCN+rEp4p
KFdDMhV/hpliw+PFyOfkjOPM3nQ/B56mogNn35ZtmLFMJETBnw+ri+ysp9eMNz8g
qWwm2DpweGca6F8X4yAu2sw/i8GEO8t4kUqnRBue15EuvQa8TMs0NgHvKc/R3AEa
moHUCoaELxgGRkQhD3MK0HtWDzQF/KS6lHNoTY2y9rD0+TpZh8JFe36YKB1bmcyu
Dl9/cYZPK1Q/2FFF6E0EE4HwXy9ZH8ODrip8HahBsWdcyZ1h2SzDSUds+/kyHoyu
++9NRNasbQ4saksCrmhwQPNZPUMQimGFTTLeSJwsa1F1DhZSd2TTVsDbz5bgvzB7
kpK2eKZr/R3dO1p860Qi6USvb1P5qjumHPHvtfVt+Zw4z2FAz2GnTYEe9S+KyziU
4mXOFfC7EB36DR3DmUP+JEPPGkfBJHuUhBlOqbuXLlgvQnFsyOJoV6zIcLr9gpag
6OesNx34Qp5yOfL4TEuCr7MUKKCiBX8ybuLoXeiO38vMqdDrFExyC1I1WKNZ3/0Q
f4Yxao2O7lDt0gJytj60VPG13WzsH2a4/ORRuzjRf+l6V1ZJSasbmgDiSo3KxWsY
Zp6+u8V1WobDWkdZlXm9EsLOlqcpKIyWN6XAPC9ntlue560CSWYO3XgnOBpuSHVZ
AO60Q60LMfavy5bLeuHg3684GyMwFOTlyWcbXNh1uNgKpp3HRhHAAENjvQAAj7ZZ
vjwqpF3ErweXkQ0V7qbH3TPAO6+nPstqe6zxXZH79yjzOXaTxFpQN488XYRdKlXe
0qzhaVRCGPw6sM85/YSjUdwgZE/H7bq2uocg33ZtGr14qaqvP1AkNedvWxQSuB0o
ji6/ajP6uijGariHIPlAIGowKKVPMPzUmpnMcsVjb7JjxzDqlj8L7TcRksGVuDOp
wy5qv0OpOsHyNRq73KpZSHfsNngTmG+gUGe0AlNlazByaDaNk9Jhm/QpXcUYmKSr
gIYaNUjBSPakXkWrXh0QQfZOkH0qetrH5oH37zUf+wRH2koNNrcKKLCco6C7BfCH
qh/4VTSMmMgdHbdZ6A8zUlkdrL2ujg1/d2YbmPGJsXiY+bJgHIlHfLqi+tvCd9eu
aifbZCy3ypRQr4j8+pRRnGAxMXOOuTsV2V7Jrww1G++72T2z4KaF/54tSB3NcY0p
TdOusakAmXjxtp+pKviAOKejq7WSAxQ+poSS93jr0S2LlP1Eh4dnDs+26L80+41+
EV5l1RGtLsiHKBwp0+6rHk1j83v+ckz87k901iMtxhae1Yu2//4GsItj1nU9VqMd
kKy5g/w8UtpUWRthG9Q05QzPSCilr0vSlbbRwTBlIq68bml6rUYI27RIAM70f4+1
UIRl3vM+WvrWIX9Znv57beWpcBeNIaQiWvhu/+DjqG5QRg8gMAwDC/9yiC8iF//n
fSn+pssflwqTaOrEYv8UlZTzHLjFF2qoawe1KPe5SAf9b5vlYiBMuqgmcRejQcPr
U1gW6dUAAfzz343hW8ddqjNTY+u02s9ELnGWnHeVFTyeT2OiqAHQpLbG7Nq0ucOa
/mai4EytsjcFzKwohksSqDG61/TbtggrYmD39eV7yVb71fC7sxdXddfyvXTeKJj7
WCZuxskVHxZS328CAzNxmVbEjk3hzor9Z7s8x8PrvQqoOSFPv2s5C7UE8QeZQJ/l
GtF44i7vNJK0pkOaNKtoZaAxtx/ebh0R2aBZu+Rj+j5V4Ltie9zLpl9KDzURdwu5
O+qBPMpVWcTVdtax/hbwAGRznqc3QnKCvLRTOq/B5aj4vBJYZ4V1GCB/Fi0zoNBp
CN4ttRYoEQZoA0RNwqteyptsDew2PMhUFAc1F9IkgxJFpPwloZ7K5G1sFVDK7wjO
SJj8hYglfE0jsywX79oz4bVogSBED9cwS0a6yih1LDBnOiok1cdC+6YOUmcnQT7C
+SRo4X1FO1+UKzsIaWiIPRoZZqulGLD2glmlk7MBQpm3SYx4XEQyiQOEEOyLkjTb
/L5JqdDRhi8belo3s7JbtQRzt56sbUQ2g7MiIopNQmvTiri/7CvsAR1C0rA0HdoM
x+Wuzo1BwiweS63n+iLhhwceQWZXI7PtECdcg+Z0qPTb7hMDL9nSL1egLuJZWnfU
OYZrUzucd/ilqZTg+uauJtqPdL/7CYzXw2VdiCwl1KBYmIyyHVx7+KAbrv/Bruuv
dTf7QqfQlXGF3EUh0NEgcpJeOR8qp840eq19II/VznT+12sjAjPHouGxdxA6d6Jc
pvQCZQEmoWIUxjPtvhuv9F7lWqGo7mhvAJMjTuhQgdzee38lGn8Vv/XqVS5DFacl
gP7bUnhzWDh5FQJCZS3eCW2B6MvO5VrIunQBEFDwzBAr+zopQdxW8WWG9tsayRYZ
NxuD6hYN6AQXzZhjKiOvgRRwGo8QeQ+VHDQsa8K8hCNMSRtmGuxYXp/LAdZ2mMkr
Wa0ZmueoRRxKo9lbqjrTyE3jlxR5aEoAwbNS5A0z/VogDpsYYCpzkfSoY1/3pXsf
v7yqlefo1yd5J/0+oZP/2k7KdlcMpuWzlbeJmR0mKwK9KHnXZ8HWY4JYUW5dqati
atmDucS2wQEsU68aH0de1sWEZ/Q/ShA1o4KH8P4qKc80xqKz+m15s6+lnfuQCjqc
mOEx4cc2AaRmLKGw7asIwX87jdcGbtN7vfZf6qhNN8URf3rCnsxk6vyqLOIpiydE
DZDjsPxUW/zzap6T0w2U5WlefN5UDuphGTGrGMeHnxiRlPH+mbukQxdy+RZkyUfr
48UCyUjtIflzGyeyzEnKBXyQMEDtiEATndPzAlUnZ+sQgwl99b0eynlXBE6S6WcC
pWahrDhzp24J/scfEdi4q6NMsHxxrLiSejgxl/oeQNQtTnm6Cog2arK1EmwJ8I15
WMen840m2FFhLf58LJ2S94rIg16Kw6Wt3wSFG4051b2IdeFmt08/NBG6mjP7s14h
a0CPNCmGj3j8ZoqMFGkCJ+Jh2pUCbLxs7oafKkyXG/ND2FWUjgadFJLGtvLzRZ3a
DKtiE01tK/aRZcZMjup/z+54CmK/mpNJgdRpOHt9T2DfVrLwYGfuHyboJyDmestH
gsBZDR9co/4qlgfrRYmEF1ZpjX500sXG1V72reLAJtrxfDZpfSdoTYA5ntgzpk2b
OHStxZqEBJdpWl0Jq/ggwd7d9Df6q2PoV4YIYu1+JkonjXtR4001wnKl0hbytkoM
GztSKh9jTWC5yA9vA/XVyZRAMiiT/GITG1NbLd/ZMRHMKjvy4IyO8vz8tEVugnP4
tI+avGLKkmjezLn2pRuMVDcnNGfTpv1zrNHrAU7P5x+YDUb12MqgN994kDtn4/Kb
HcCV2pr23wOXrtFTsU+EI9aygcW9fslUV4+85H3NQ7hRRZi8JhJom0QVmbVFJzbg
4pjTFGwTAwn3iL6hDHvbZ3orO43tZxVIGBAof2AANBn9X6W2WSsAPL6MSENX3srr
yPitD49+NZ0Dzz2TOPhnMKXD/6MvC0okazbSQatiUzK+geufMPZJ10JEYJkoxapW
E9PXf4vSLYRLMI5a+vflu7IMcrvXVpqCOhyUB6mCcmBvAU2Dhz2bBQt5ImFm3j2w
kyYzFQHwStDfYyei/+hdBT1tsBtLlYXPK4UWJ14pmPFSSg54NSIxF1DHMJFP831e
+iH7FRl8o/X0ZyMQRA9pSMCiOJ2ldqOp6LrRZHpcSIcI4BqNJDMfaae23UWMvCX/
uAgufBGs2MezfQ01+dgDyf9mQ/Sbee1W4zeo1mTMQOz5h2TyiP66EKK3AojQwcZ9
ytaaVqJv0rlmd+PXOv0UL6AIAirPGOP4zfG/uNiAplZCWARmryxKp+KvMRfrz1sb
vhB9Ptg4ByCNXXa8GUBNP0iGPRwN9MEutvWUbWb/vO9m1m9bCkft15t+sIDjIoOL
fXJ/oEP4iqMTvmAiyeypEijxKTK4C19cx/W+PdBOdVRA4MghJjKq7IixBWyAXtlu
T4Y/2/SCbnEJpdhv9MiXpyzFy42da43xwZ/aFM0N2AbtVG8B2dSkqJBpgvOz7ObL
sC3oFoizcSyqK2uZH2zVAbLcmg5Xv2eIaKXuJvl8iaK5h6N6VK57qSUKAmU8TslS
3P1iXe6eQ7xi5rWKO818fS3ELI1krdtNBV/xsxh687TUuWtdzaDuC3vUHQmIU6dM
IJO5j5K+bfYcGcbsVuJkueaZEzZOPUDNn6X+VcfuuXNXWngC51mMUjIBYDr+0dOc
ZynqyCH6iD7UcvHXA+lczDRnvAcolRxGtt8UOhLwUCpn6T/4i0MIfp4GbbHXq0sN
ZjoOgZg494Cus2yus1JGu2V54pvrzWvipcQpkL8hoE2sAdG3trIgkXMjpa9Dw4m8
0HZadJcpTdSw1ixC2G3jLZc4bpxj53pGjnyT0emJ2p8XwK5Lpcbn1B7+tceGOAgr
U1CEl025vdKFH1tzk897baIFI6sw2xKspcGslfoiNjkM5Gl9PVOwyzaqxbZXmKDl
uMWXwN3J25kbuMvjNi9ZEK8QPiXhPpRTsczxucAzM1w7k/p/wyBsiSELxyC6PCji
lDifej9LXKHJeybTjPEL0xt4WjpA6TK5L450UA47cVIAnou/ECL8HKcMdzKLrkhY
rBhYlRgrs3RoaviD+d2cqPtoNQ813M7EP3qNQel5+t9NCUZ++Ee6aFneq5k+xqCk
LfmJdWZ5qml8WHhNChIWeTfuJh9wxbbYCDiCg0zO+w2Dou4e5zzfRbivi7Da6GXi
6Adg97A6NKo+D2aV8oICYhnBXWPWtgmEYFwbPqw+9CGHTpZiGj6Nvex5MF6HLXDG
ruAYTIPUFO3i4uFNMe52DdX+TVPNniTr3PCriXbV2Hg4cSrw4/zneKMeBkCQ3nJX
nu/0CDzbO9SHEOs/SOTB7DHNZfCnE1ykikhpqFtOp3hqdzu0KWU9YR2Rr07sNfvh
jkZDdMG82cPZk0kR7NVPzbrzmQ/0eeDDdGWVbZVaenEFeQyDgafZpO4Yiob4pjXk
W6ypnjW6RTMWI9yK6WASsEsNwPpvIGFYrdh19XXdF//BhCGgDPo76Ti8aBcWdB/8
4csW1i+UQtBU43dLjZ6r11fwRBWGjslS13j4dbNhFA17dOyuT3uQTGXXp1UWfkzF
P/M/FufdCzvubhtmUBSkigu1OmzF6CzQppv+1/h9mMz66oJZj3Ddu30Eqys7F+zI
6GQj2yfYrtzfPGxpTHRMp19Z/HqZjueJVOUj8U7WBY6uRYWWAqFu+S/n0pdCdApo
8bGI5rz7bfS+mL0MWhVW3aKwu1LDf9PVhi/zr2JkTMbv6T8990Z7+WAvqf4VBs4N
MpAJGhyHcaO/jjP834lYEckzMM4UEgt7isWh8kitDnDLUglF64qf42aMbWiE9IWy
pDiZJDobciG9fHBrXghY+IRI+t4+YgKwPZua7fMheYffLgc7BoekEfHgayL28+fd
rFX2nIEcvK8HkAg+mU3uzqgeG5VDJqrMoXLFh8rQaru4u0cKUkORHqZULu6KGX4D
I2/kA8R+6nD8zPJK78wcivRIM7VdH+Iy98C/aiwhNIH70bHl4TGslrlwJ2QJpdXn
AkCzSs+6X3jiL9hAvpzugtwYvZ6ONJ75Wv7+BmeEqvkCtTJ4cvTgKFNNiS9hpp5p
i9MmCVWrBb24+ecPFichObyiEc7i+aJjvJP8NwozMUQ3FtPowFkLHmgryere0i7i
fC1f39X9RBGsbjN3maEHRFPyQi7uwwe24QXONUbGdG7Bt97pNoFxHOV4e1PA0j6w
ipC1ZSnSZuNCNOO6vr+f8vBB7dlq+wJf9lmkWfa5IdKrTtf1mbI6+/IOKxajuMxh
NVXXACW8N42A1KiQa3QHQg6kj12EyxJZo3oqABMnyTsir5SzQdAvESsfrI216NuK
vHwfM32P818HM7TNa57t1fd1osyffQIsa96+hG2jCcuFsWbcM+uKjgwvpZ5BnIZ6
nrvYg5Wf305UWamO6mFM6rFbqg4uaismaHyq8GbLlttd7UeQjARhJUUVDmQFV2SC
YvqOOszGpTFyH++D6CXKWsrC/sp/YQg1Vug+LPkG2ykH4cedxULdSgaXnvO4rZdx
cYgWLZdBJBgjyhgTIeCqX4EQlx/3UBfy705LW8LtFLXqCJ8oTFT4qzdRemQpzJXr
0cu2B2ZMnG5+cWdnfuEHigG6hfHO+p0S221lWqBiQQHsq6/UfHxK7SbtdyswqFuj
hV64rEgx2MFlq8qa12gOgrJz31x85BDm2aRMZP9H1l/Ima92Z6sBg3fHrAlcX7RY
/YCS2G/3MZuYEKdZQuCSlOgGtpwTn5y8JCvxk+d0f5X16sFCJl+dfxKjWmSSJKvm
S7N0j/WRxJooT8XKGrPOxMfWJmz23B9I0GP33obXNErrGfdjowyQxKoZNP98w/78
AaRgznvS0AwgjUyXR8U2Q7YzGrIOi8KR/40kPTbB1Ko3VZw1+7DGZtW0BWUnsex1
CdDiq0mOrPDDBr10Eu+9W5HHIxcZsi0FUdlMWPFfnPPFBASx+Ml9n68HDkA08MtC
8tIEBmZEYvzKK2Ccl8Q1bEujL9V7TQ5nlhRbKqkY6pIYMqj4EwEMzxiTkdUzrDIL
cCFwTjrthMm936km0vo23iTNGKCSOKzusmE0IuhHuejqbquoMTsB6cNqhCBOTDSv
JTH4f5LmTOPyvyWbklNNB/tcYhbul5GUh/4ICJB1g+UbAmI4+zIyVRhA02Z4imNe
jflccojsBdMXCIEo9kQFJ2qIIs91FgJl82ndSBmHm5a8gLegRjTa268oMTjCaqBr
9rwhNT6YSItvZe7cG2N5m8uu0mn3+gbmtRtIhHRAYBg=
`pragma protect end_protected
