// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.0std
// ALTERA_TIMESTAMP:Wed Apr 26 13:36:51 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
kBlqFwV6LFgEHlS6vpSaCc0SgNQkzhsJ99+4aOkdINRQKk3LFl04t/ix+vBj5qzX
Z51mlNqDpiwp9vs8waCE83JERJE3ZoWDoQ5ZAjQF0eAaarYw8A3QeddUvtJmAOLY
SD4aJfGWSls5XaGJIadkbVRcZFID8xH4hi8P5BDEJEo=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 15968)
6rYz7b2HWtEcJE5bqABZmfwT6nbE7bG/yMhlJwT/AT+Y6LGhcmiphUCXQ/OAkWcH
w1SLV/7M244t/Tj1MHDFAGjPixRaNVM5PmstOcYzNw2LmfjOtxVgUbXpt+k+ycPO
rk+8VYcYpFk27CfXuzxKwewSQkjn2h5JkAFvXbgUisFI/H5zfZNI+hVO5H4SW9u+
bKVIiAAyNkYz4nGIkmbG55/N4PL5YQeg0S3ygyZHCz5y0zF8A2Y1x71TBhYleJk9
OP995gkF5dMgZu+USmLAgVCsnYJB73v0V0ORp5HiD5FqXJwsZlScHrqFfg5UYegW
EdmxBgEUKL3E3uzY9m/8sKPXiMe5N9lABiYj0eGc8ccf+zLS6Re9nbONYDfeGQj1
M2dXMNiR2TghkZKMQ6JIZfw03uqZIuS/p2hlJ/xiIPEwx6P9G0I1l3DqpyxsoBVH
4hbRzGQ911MvzwqnwKXL3o0zLjKfS6fXL+e+7IipWzx4MY7t4JKwYE6GLr/fsQTL
YN9FHOPvLvu2vmdZGVQzyUUiu0yto35qwDMUPf0e01o5EKhpYOjX3iMhYhCFQktJ
+t8ph8hU7uS/UUlO65uzU+xCSGNQlrCgQW0MU+cHhisLezBSEHqZL/bAV+cY+P0X
qcHE8rdCEjs7HvUK2KxcLrQ96IrsXWb373ajaxwNOdie4r3tMce6MFQKHEb2g1Th
6qNPFrOxS8YElaQ7zBZiZFE28prVqFa7lCQXuoQQuvEorbWmAKGrJov5L063n1Lz
ppNpZUXA8bkmSYCEZwzghnejZ97y+uwXDVFxPp1ilSpseOf3kQrmIeju05lwBt6q
EuDaGCcBXRnGn84/o8jOv+7tK45vBoRUatW2u6SZ77+AocrBOVZ8apFkEYg7Nez6
rv0970wTw6MwAK0lWVKHJRdxezwoPDFLsDPiMzTSKKTXh17IN0C/sFtcr+zPb7IJ
aYegqAY390ocBgEGbwgCDIblnqGqeSdgNQD3PyrNc/r1/h2BMYCxNNJuUf46QN6/
2Ozgu1OqKDpbhCuApxrAgmmRealE3k2SOybNXdm7SV5Oyguy3LrXIflapH7MezXv
UFcIGZKnL9pO5E4JgMWkHBZqXBo1B/wSHsMni2A+ac4Mjs92hXVe73X80PuWK6GX
FRTwIVR8s8M25sXjO+Q1fokEfAmFct9ozEB4cCtK2erZUt3eONw14v0B7DC2nUtK
YbdPX17t3Q60SB3sttXVVIo0g6dqXyGRhgsmXZrntW0ogwMzMSHGN3Ra3Zs0szSj
rM3vLV6IJUcMqXb9eHTvv3qYsbsYuCVDa2xywR+E6VemS6CXeXwrfUiqFzG6iymG
8YfZ22NhlreEe7qPJls28VTQxdXbgzw1Mca5R+fj7gfbe4+WKJe7XZgGs7EXM5dY
NjP+YzIuZlTvkDtWbQB5skiFcyrKjma86k71GZQOUhxw9qKex+O3mMnQrtCD2RrJ
xIVi2oFIOGoBoQY30Qm2Mrbuc9K5myCxa0EgFzzmASiL14TJxfu+4z96K5f35vBg
WBYsmAwy4MyrnoM7fYpPAsvQ1Jxxiwj46vc5FvvvOjr/2KWQBBWfW5o7IY4zgd/b
xsInf2AHEn++hHZOwAX1HoouM5fJyVseTqbEorDs8h0YcWsp5wqaB0OV3ZuxPfSo
ggeAtz1IhN34nZ621K+sIN4S677M85Qr58uWVNkB5gsTC/7BKfSfUkq9FdLhDmYd
FWtmHlxhzi0ab5hpRXhiuHJCr49aXSLOONK4+l5Pw9D6k5KfVbzETqOO7snu1b4H
m7ja8r9bV4ZVZR3FB5jNSQJxtos5gwqymA/SyT1O+jj2qUCXmLnDF5amoij2Fo/U
B3q/gXWtFRcMw6htGxD6VvkPaaW11xXnWVYD6qX+5RuOavhTMhI0BCu2wQHahpSO
xW4jZ9j0FxSNvxjZpy+Lbv+NminVk294GmAfkSlpceOLymeDlCQNPLkTSEV+X/B1
TOTcrTZQ2GHJBQFBJCOm+qcYJKsO3YgxkioJqQe85+/JA6C7k8o1YZd2O9XNEBF3
fE6iYx5DocKz5wXBlGfnmj+fXB3xQU1ISklmVWI41JlQlTyHRmVjgYVltCmcUafb
mkVkLMmj35DiHFu1l2Kx39MDOUbf6IHyAct125kNjo9svCKuCszhQO0gD+cHE4lq
1UmAkpqb7tS8uJn5AJHr4guFIJvPd6w+VUI23FsDXdVBaA98/b6aA9ag0er1lB7h
GDT2ikXWTqDWrb5NjX1gV6cT6mYI8Y9fbZzCIU6L5V00Dj9GlcOUpTHZMlxGAKJA
5vcoRX9Ztx5rlGaoE25S/2ntD6WqF8FRvyZSGMGYGkiHnz+FagJhcyq2VN7haMkD
me16/vY8kuzJy1PPOy1XABgTvx4EqtmcfXBVVmLJeGiOktxla2hLm4t19dveSfpa
0wXKTyBiOT114e6y4jbDpcGud890VjCdoj186xhrAtRfaeHcM+e1h9Y5AAjWCHkS
ebYZYQ9J3L3MLnxUu8FlIOt1wmrlZxWrCtocqqWb8EDY9AOu1GyjayEIH3crxyDS
xd7j0H3kn1QH/5IgKCaOwQUY29xCL5jSCWjs9cxkEgOL8abYV4Wip1y6EswWQqDt
jO36NT8vZRj4UItdhVFaI2+ArhPAnJepXAU3sK24HX9Sg+VY/TSbM6fvzBTtqp18
N0OgM1b0wP7C5XRv7huW/LwUSnqMGwSrPD5s+vrkHfB9hsl2GmtHz9t4izzPqVtD
gAtlTl2678Mb9PN8FSoP3HdfeDNtpE19fKqmbbeTjlw9D1gqSL7JD7ky8p8c/414
S59M2tVs7kn8hOMzspC8wGLLyeSFLNyLx4PhHrgVdqgF5G/qoQZO2CRocVyzr0W2
4sEvphpX+AahFK4aokjeicEyiNcimVKmt0c55MsYNfmtC1ttmsJ4OySihuxXM9qw
IddCH1t0vKB0jCvF86XUopu7vQfRcEuHpz/AzUlKaeW+Yq4Vg1mVW2CMtCBBNJEq
XAS23suBKQB9n8mj+aWn2fQ8Eo9jhPqMxkdwhhHupcLfh2AHNn7qTvDKgIIZ/1sI
L/7qrbTxDx+pi2eOpiDB/V4CiyjBJ9P4jK8JrjNr/QNYwbfifZUtJGtEOp4AKaLU
Waz8Syjr03xhdi/CMZYLI4KnPiR0FbbuPDi/OBhkozYQG/Rav0GY12lchRTv5Sra
127JKmLOxZgzr8EoUhw9++Lx92S6t+eRsV6zUszYN31fd0z+vcyBTOPGsZ8sN+Ub
k+kMIVJ2p0CqOqBhKxIn/IlKdtbShDb88YXapaXfn0llt1NmsD4ni6ze3P+mkPoh
w5sMwjMBLX0lHZfo8y1c5meP5MgyJrAXyqZrQllrV3t3N+YPv9B3AJQtzbA899ON
uaMD2Ahp7XoeFiIoqTBCZvjUT3m9dq9BLv3qZTlNZ8WhzwKpay29q2QazMsXB8O+
Pc5xXmqd0dssJqx2ZyTOTRAbgykNZFiH3mghCGvpskyTRtamzDN8hmtBRPKng2iv
wo/HwHWBuSQVq6ecLp8JWuhWFcHIn+G/VSg0j0nt+c9gYX1mVVBnRmgKBm1jByfn
IcAKhhNOxoho+MRZCuE3h0zW8Z5nFy3DwyFMJyAt9VexJQbXGSbTTFdxYKKCdDWz
/HXVBCD4MvKIeWIuojS2/ozIVWo7e+JRJUeex2vsqjGZ/ba3pk36XlA+ZW1S/0T5
t9a5xptYNrB/95M3pklx2Ndx2GIdBe2l2L9BtZAtnxvxPY4uFzOXYNcbIrtDm897
hr1iXneVWthjecexaZ6TDoc/HMPYFouAa4Iue6VhGaZ6jCeZOcFCA9qswe+Gv7fu
8AXpDXckD3weRXiUKqnKibj5w8pGg63vu2jEd7uzXYXADCSojwl61lvmF0L36jyr
JMpGOZ0S8nUVI4VvTQGyT8/rOKrUUvZq0PW/Q1YWNurd3P62gMfELWp0DxAxENmz
VdZHy8Yk2Z4lyyCXCIcDyVY8XL0mhIJGrn+Gxm/u5/MU3Xc7eG7rENOdN7lv7RnU
xT0TGTJeDTt9eAlREE9eRkNZIZq/OGgZfX9XcmoSKIN2DUrmrRLwwEo0x0d0GQZx
Ds2km9hgU7Ko+l/kAjHrxwWn/mjeqXLMNASx3PP9WiJGfXSctLs+ER6X2+ij7Ubh
bpcpdkDAG/vUg448V+6jnk9NcRMBe7MdlhFGdfcSA90nphNpZh1cAt/e1bWs9/eS
fdX6LgZBn1VHGnN1qobmYg8eXD8VuNSlCbaAEoWin4ND9fbmXkt3xkzRVsZXDB3S
Y0tUKcbnoCq6/aMJbCsDwPFLSbC48xsSzDkViN3EGrrmTqp8V/OyCdJRsvtYBl61
NLzPBPddqlpnEGQ04/+VLcXxkG+IzsmHxoilL4N3i/nMLJwOn2OLk0lkPDlbwygU
q1+SMKUy/pGOmLRcutgQAT1KRhV/0wZp4udr3pR7rnqLRbwiojvCssfJ7SnIdPiI
nDT4zjtoyQTFrMoyCjzHtQtaoO+GJd/7M6Z1Cga+5jj5khDl1OshTNLVqzJuErJe
mIqKuWPT6vxZAY/rqy+yTr7dqhWLzVzoFTE4QRhQLGXv+stdv/iv5dAm1P2bhB6q
khLczoi+/Ty7ZyACOfDgcGc8r8w1z1NnL29DxVAcucwK7pjQefl1nY44H7/erS6l
z478JIVfbQ6RJ0KsohJRl+tsjnkeATaFBrvTzBjLWXWyHeuM9XfwgAvel5FsanqV
TMjWvY1QgJzzoABMu7gSJDffof/PPpoAImQ5DXfy1soAAC7wmwp8W2xLLwxpgnuM
BIfFZsCtll7E1V+EYxr/6Ukd5jJP+A/gYfjpjvP7WmD+YGbNb9qyuNoUTm2Zoz4r
TQt04H3l0Rv8XeCCvnpu5Z/6eaTwuvmHg+mhxn8qN22dGlpemHZJXg86kZdfjsQi
fyROnch9E97ICqQK53pVAYM/aWBN0PTY/q2LtNyyH8oncLQQDtgpZUrkYq0cqAq6
NFNu+5a5ROU5iONZ5uQP8IkwI3WQXT1as9Z+YqpLRWX+F9wrBdhu77iLM+vT1Bx8
d2nm1LeA7nzV8Slh/NnrfK/EUeRp5neYITj6BQm52yG7HXBgQZbpOErAvepTU9Rr
5EsQcuaBI6o03MeDsLqFpXH8RaCuxMZe0Fl0Vp6TaT4inZW+J1pkJR+GjQU6ZD+n
JC/H0YyGdJGhW6fDVzmmu+HRMb3MRMSkbte3JevMNWx4xohgMksH4oJeJn4Mce0p
+CMH0nvf4rVjPo6iWUgW7gf1iyJe9Sk5msxulCtpcZgw5e03ISO5OVI0fbA4y4Nq
GLeHPNwdTkDrBtV1ZTJe2bRoQALmI2o7o9lOWqCFK9wC8FDL3qs/1vx4dhCj1xsJ
JIn7fbcxWm2sgyIuZOKkqqH4vsml9sJvSjWFNTZACRn4YFs/htsO/rh+zLPYO9qn
wMHCNqVh/zcXU+lutm0AYLVgvVZxFg41cwo1pmUcnl/Q+npLEBtn9smgPnKqNjLc
zf7gOoZ0gpjhHNCCgTkz3e4uDtiR+yQl8kbh9UU3xH+ReslvIIlEvTXp7Soq8p3o
AJDxJwYvwE2djxkQEZKfOZ1+SFdSpnSFXaPW0xpqnhkDodH9WnZ6nsN2EshxKbLF
E95adc46HchfX/3O4tQYv7Rz+0im/6nQvPf7al6qA5UShsFTa/Ap2AmnVQYuBTij
IiwBZ3Co1RPKxU+WX8uWJ185H7oFdjIT0/Y8Ko1Y4/p/QmtM5ak2QOhpc9uYdRwE
UZwBxwffHlHzJy9SrHar7X0gpK2TjDdTKtsbEunO3BIjVquIOTb/NPTqncxqkxAF
YJGnSXTIf8Jqw9YZeQa1953EBmQyd48hv1vVfoj83juMsHGEijIn+GdjL+p9qK9Q
o+6qZElhyulFz6c/T0hA/CCuozLKc4qcY4UoPUovElJO0XoNBh1DTeyAdFUJq0Wx
zRHU6bax+jr7dfIvUHeG9uirJwL9cXM3VIEkCi3V2FyvNEd8661bbyTvabxftEW5
8OtcSyWf2HNdA6kcBdPgRkXwMvqJo30mThfKQIVkBHtF1lBS+Bn2XDQLQi3YnRCb
g/pUOSc4zPYI1VRfnzbipca0Y5a7fpXn6tJyimtsl1h2BEy/NKiY6eMe8yRQk44m
HkjkogUfZXsl45gTn9D2MEhLfmgwz8jAoJQLp3D1lsSzmXA8YHPkbzXeRWKqxu+u
HReVe+hmv+/scKIpWZsf3b5Dv2W85E6iw68JWLCkjXJFslo2yY2LPTu9EeFewAc3
85lAyGYXqgz3sq9FfvQQK05JE16TYe4DUveOh4JFO64EADmeAhPYZH9EUtsnmXb8
ZHUtQomuWflYDVpfExOrZCBkuwjOSfZzoNhxWWMoRm2THax4YEuZQcFNMi9Erx+3
DJEniThdumIeTTlveYcwalb4bvA3bYb4ai6HrkvUyh5X3q7Vd39GOATULX+dAdA1
aBiMGPk/n6Ofwtb8j9wJvGiO1z912qNx0Cg2dDF/8899JtdG+P9+L9TRW5RlfbRX
1gvcgsztKUGI0j4azFu1wSdiSO6Ky7FDTJtdOyOHZ8QvwaId1jYjbnNTcKIJXJJ7
QxFP/6Oeg3DtI/79VynLBN1Y64iz0ukgsYNboiKLPEgdEJYjl9fQfsMj9yg8NVIR
obkLQgaFyCodkjOS0UgF7JGnVGEeFGPDtZZLRKQoGE1/hcEE/avKm1HYTf5MhnVm
re5PdrVf/qR7yKRKPiQ1XmGRcJI/wMacFwN061b0FQh0qLpgAl+hwLR4fWu7j5WF
PTPBi9HY8uiWkB8q6JX+ncKR9FYPDG+v0f3KlgpRFU+F1SeozUkStRR5DoYXxcWo
Am5/otdvT4MYeUvOYUa7YcX64Z5/mnNuwCzGsauEePmixyajFM+PxNxEbf3salVs
+olvl9uMAmnV6RA0Uh3tYfoZMOlteNGLC0e5m0WM9LQJQ1p0HirVqu/o9bYdN81Q
Lb3awLnX2/aRbLdl3fDQGoIlMsLpk4XRzxLcCEbYHIxoJ8uA6+HZt9qojomxuedl
Cb7Mye4eGT/EmuaGi8l9yg4roDPmKmAQ6zoIMdRmP0mk0ICrA8cmfMHqOJJrbOOc
2wYRfqJ65dkhNag8CGOOJrRHUuG6fmeREQGCVB0QOMcOTz5WZpMABWq0SuMMqGLe
IuJ3kF68bNQDipczsLTQFFv4Nz4RbrrxAq9Ks0N2WNpOikGDL5zuyRXmC3AfyLrI
9QjS1KGyVOM3m9YM4KqVMi/k0KNxZEyIWqG+HIge4a8DW/UfIpyEqTflyaj12Rc6
Zj/i8LqddvFPZOjLcLeXbqYRmmfs7C65c4HCc2trjgolMNa4RDiBaKEZM6oDncD5
x+7RDyc+D+XbehFmHeqxpHARU8jWf+kzTL5mMY4bo+vPDIXt5AkLlNZwPv57lV3x
/748TuEVnHR1LQ2WpdgbELUc/pb1lXt3li1UTdzkvvGbUTOvjSz+ttJ2Ugsq8UiO
VFTiWR1VArBuStqRFLbfKR2aV96TNyISDaxv9YCiIPUI/Y3PoIkHsDZqnO2RTQ3C
vLe4oZIWQkfehD/31HoKNHuhlHeuEUeXnvKHp2uDwM29RcspasxAo05JJAuro2dz
sOFal8/KzNqQa+HDfMEIpWsC56UrIaEhEQOEuL/rCUCv4tdFtQNIO1Gles23sO1s
ASGuHWf7hHUpAySj5qOQNSlzVSE8tHGk6VoEP4ZeNQqJKdowhV2dyrZWuqBafPiI
g977kn29TtgzpzhoZeCNY9yQ9ZSJrWO9rW5wkcyk4SLdwQUbnUASx0MubN1R3+DQ
4Yh6xq/slUzrb2O3/ySiuADkvmfrIh4bUIqLkYVuAaUPECXv4dRYOg8dKpuPOFSA
85aaXP8pBdJ7fgU5mDTJbAza1akK7SheVei8pZtXRv9aFZW7vIiwA0UEIy8WP6pm
oV15m8MtrgORw6Tinwm4bauuSVBsgkSEeed0L0WFg3Z3Y9spZS6G32oEYt2m3DXk
s/qWtDZ4FPIOYr29gSKEdj+LjJBxLiRZdSGINxjZz8HicVS3JWZ7banaaL7Umxbe
XmUgh73lS0fahKrZtkyj2AFiMmEcL9ASKnQPGWt/fyBcMt7goL7wMwyZPcmvMyt8
G5lYgBzCJbTztXZU1NcikXsQum4onhhEjC9XTZrsbYqMmj8cUvCI4e8720iQznpA
53PMq0U9M1arF84rllQ9kErtEsnYWvuguC/7ET4pdM1szz51OpZJFnehLCX1KNj0
69fxQUIrGYdZyAPSq5/x21y1JbABAb9Fh65xoBoiaqBR0ucTmLMcFVsilKbR/mwS
+9l0JxQfBAqeQS7sj+FYvQj+ygqqM2nHMa24zbVJkpiNrHH88I2Z/JvStcbx9iVV
gTw8N8JLLnh7FVfEeHjvNHsEag2F9oWeYimzHIGvr9KDmBSx2S2urE6EQ/MJVfMD
lfHO3do+TZ2wsbJ/900N8nqsINQ0jcnXE+1xO5X/npdXYRnaZF7iI/vfrwyulLIp
vXy6XgytZCUaJT9wXRwNn/14nGqlH3ejLm1Jg7zA14ou8h64IezWvQffye3ZjpEj
SFN7IIvir70zzM7kQ0HceVOC3C6OWWITvrRj7jVCselz8B8kD3Cv2vOLj12odQB8
UASb8YR3NujjMEwqYQvNiPkfa0g2Or9Pl+kTuRBZatN61qkzIs6Dh9CbCBZDdJ7E
9POvoSbTCmGtHuIfq73BYOCtFwW4WBg8j0AldA8z7LgPPTPYe4ifyrk1rwGmL5EU
/0VNJcyN0hCZ4i9BZS0NogO/HOg4CHclPjqHlTkJ9W1seOQC65jNpFCAuohInwx+
LiiPXC0X2agMkcs4/zHEvIeHoWmX7tJNJhdsi4XtAkI0sX30+Kt0TnlGVylshzpw
dAAeCe21i//cwqw9xqrsFZhatX+h842s67IkKb/a5Mi57xTMYqPdlMGViaKXK96B
z870MsmHoIsJUuOlUIqQWWVKcysWmK+u3+1puvNQw1F3400dqnJ9mwW9IyBWrFYi
tuIAbV7j/1JJ8m5F55IItixivRTMVVIEW7F6mAyIKEhNK8GO6jQx/RsHRn1iwZhB
I/ydAokDfX35x4Ib6F4Q3cv37BU9Br2K6UwDqjffXNL2eOuG8J2RrTNjDR9ajWe8
NNgPQDjMANaid08tCb7SLjbWW18w+Ub/S7A0/IV9rUFDk2xvPpov4Yt2TgEfnYbC
W9IiHDUx9E1gg9m9/8FtzPsQ0NVoenRR+INOL1qnSf9t3AR93JgvpjSrsX7cKFci
OqgJgKUKW9Q/ueqg8wMIbkxtLavleBsAAx/gbkc+9yKaCbViTa8qrHCXzv3fdpHS
j5fGUI7tyoV6evhhheJ6ZGKbNAJ9Lg6M1W6ZKKPXOM6JXOqsO5/31GQyLmCN7rLT
l0rx8ueP2L+2vqbazNv/8y7b4L6eMPqgTZ+04A9+q6z5MhRdewLgwPudmKztnfF3
JwcoAm4aukM5eXz1DZ93xjAckKexxbC3PCFROS1b3aN2kw0uFV0HBbRXfK0edG5v
1JejngUH4Eue3bTOrM/yujlfnjyRvv+5GyFesOv41IqTUblqMjEuEHU9gV1Q/FDQ
ErGONKINjjdp85Mp8l+morraaHgrRlcwjTadntmos7HZIncruByXJ3w1jEHU2JVh
vf4DlNjNkHHOKtHTyU3n1w9keciAethP/3+vbfbjdynMeelvYsDYTd5Mn+JE3/Hl
P1uGCReZeBJhvKy80ZYicHe9JDNkp2cp8gyjch8CIS2hmebCTADwViSCMFHljO2W
rA7pPE6NTPrAZ57vrhgE8CCZZqsjMC9PVpKeN+MfYJ+xmTXgtyj+TUdHwob+b+NO
wnXE8qStvPl0mlzQ3U5hd78H998N9XzndMyBaXfGo8n+egRb6yEeV2IS3BmR7o0Y
z9vB5Jo/zUkToDza86LEronkWTQx2zrX6drX+5vAIB6iRxhee2SyRj8X7IyUcsgK
kf+edaqZNX2xsJFtYKJT6jZk1D2zhh4/cHlZajwNdHvgU/Elb1UZAuZDlZMcgRIR
zGK9aVca16NL+5RfuXOKcFZGJAg4XO9WVxAnsSSOWLRF1gqp6CXLfdGClqLEFlPK
z313H/ZwK+Vv+DjLt833anzGC/0eTB7QGgzTkqr+kKc7bdJp+kp9QbxF/HNHb6DA
Sx0asy6svBwgvdZvx0m+Ai36h9EzN3v2gqULd4/+KWndf+Ctwlir4xzE6QGB4mgl
UdjtlVHgDtR4UDXRXhG0HxeEj3Z/mw1e3obgOZC9ShOLIiWCnbv/b8rSf7vhr3RN
hsTOCQtP0RQukjY9LAQie1CXXjrflHxoilUkqSQJJ57wCW7B/trCxxeUa70W90Vg
R6LR/PQ7PxZS/HfjE2rRBMfmYM4pX2LlDbJwcOPTMS+KtD/PzPtkCphhUATfnRxx
52z6yqhqWf+StAVIB7rzaslYuSKsXjSJGPUbCP0pX9bqA/HqF0GegxqBrlO8qExk
Ow9Ngcq4Ng47C9ASX7A15WIxOwctirm7YtsdEj5DDeLZhbgLr8PIC2vNLzhlV2+o
OHF1l1ITjHC9AvOYzSoM6gHY3iz5F7nXCtOxXGMkbO9U/aZUfKV/NzVjq8HqShQR
seUekT0fLK0mG/QuoaTlHnqE8nYn9uq5jwEq2k3cLVJ+lb9mkUneLK58PXr7xr4/
JCCaQrKrqajDRIHaqypBJWU0gH70iQhig8qTCKRyDSuZgN82BFO5haHRRsng1yLD
ckQAhUDU+MkRF1n4x9KbpTrJ7MGf/LDQ7erYtunPt+ozNxXa/HUniBrWWKxGavkB
HydwHKW2rypXT0t4Pu9yII6tVw1eBrWPMkWr/oYMmSw8pR2ES7E9vaIrYYzNl9/h
DZBmos8qTCNHbsPM2SRRyrItRHdS74nT2CkSUdlSdNK/Zeq5WzDU3A4lmUj3fBk2
rfEjOEmHqbmDB3J+l63rBl4oe3JYg/Xs6adnjiXLsA7JUsUAnRCI7+LZUTRVP54j
r0seEdZsMnHU+7t867XM3aqHaAIAwTKFN945gxOOXu+ermK+YIKkjsEUOOApifPQ
F9BM6/msxp9VEV/5j66P1ybQVIIZo6HPIuT/S/5YcGVkK57pY5f403YYH116Mdd3
XqoZR4QH+ZMbZYTYOIijXQvFKgRqyWVVume4bqoyaAECnhjx5La32xaXa56eqoLa
/uLIi1arDp2ABmzZ1GQ8aURwUWs7axvcx8Ez79UvXiB7WXEg9cRX7BRLx/GiPLQp
yuq310DVeWDK2nsK422P3fYAvYGhgKYdfBzaf0fX07Y8XAoJNgfMP2GpBE8SuWuu
gKdMeVhAYPoCmJ4ks4bBnHGLR0nLqd98S8DLYZZKCFkOsNOZcrKEDY55JASdXzy3
L3oqxji1Ofxhy2bbeIHCJSphGjW7boXxxjULaYf3Opuass75D8c990SgTa8SDr4N
2hCkj3hxGuMziJiki/Q0TP2CZIGNBqI7iVkh2pj1sKQ7drQOzE9+EW7DJyUNdd24
JycSpvmoplTElkyteb3h4zVjdwZmPngckVyHMbHSLK4jjndODlZjSYyiwVR7xEPL
G+aMbn2VsWiCge+NIFqbjL/09iOxUsuw4EXbbES41uUKU8KLm3O2krySv1vhWHtJ
BbpVQHJag0mwMaLjW8zvxstBkoqg3gBiuIlWudGorF9pLBxkgTkZCqzoXUysmyjV
N+h/PBolVGFpAZeGNmIB9i8KhmJLj6N7DOd6M/3aljTC2mPedr8kt0HD/pty2NAD
EfQMdL0H315Hl8Sd2+6GquVehnb6t2c9u+cJhY4jd4LrFBVmIusTBilBm780pzhY
6+r1Jb3dPAQL7x8kn1gojtbh0HJRSN+fapmey0zCsg2WmhHDZ1uiEHLhHRis2Oxu
9UAUtO0NC9NE9jM2p94fhf63dyYeK6L5jG/b5rOT26iGRUNY2xAz/FXBrZQkN739
eOmU4UoSUNwXg+Z7kHoSZ6QJnYZz30Vg5ino1K3ZfIc+ZygVA8BYnJRE0nhXHAbN
gT51DFweORD3tc0GLs0uofP/yDzZ7YMtOFeeeUcVqCRfP2y7KwNhKNgFbUStL4K2
zYyue64HkFoS4MhmhkLiR2aBfzEaZ+6A0J7Q3uXjXE0KBdL27HwEQnTR4UQ35zJb
P5SnmPfCiKD0P6+mwdgc6NzfJS6SOXXUigHpcsZArUFhxp6C6I7nWVZcBdBt8vVB
X0zxkjzTh63c5xuddq4dWWbIC6IVoJSpe7haXbc5CpTIenEjX1tEEEm+SC6HsCfq
Sy69qEaIawE7DNurCzTUZYATgBRn8CDRrb0IgK/zoRXvjU+zTAIf1P+I07ouU0x1
0xy2yzi1ICMtWsjs6BfQciFQAlAp2FoTgc7Gl2jQnEftN8fc/2s5lv9vDh4l+J7M
CR9i5tihmLcpYhtPIxIdKtpT5i7hLKobczhOgxhLRYrSOdJhHRaEk4YZ01bSbKzP
KfFFT1YMkOsOu49h2v4QB5uTmn20LeRoKeRBW7T7ag/G51l1BNxggK23y/GF3hey
RVntLcBypUQjeIsV1n5iB+vZMNSHWozjjca4dkQlRqvPXlgK0xoPfzwBompO8V7H
6dc/yZg6i8AC3DeFBw9ztm+UyDwx23sDhZu9I5zcI21M0SR4D/7TP8Xz/iaZ7YBr
9C+/UhUEvmY+lksg00nv3C9+F4rBLGZWRyRNMVXR1q07Hwh8lL2jpH75kmK5M1oN
WIJOf0qg3An7x7zT7vaQIhti0WrQSvly2X1oqkf5RY5iP0xlndHhI5ofDYuE2vUM
zyx8ELjkdM3jLshykLqu+Xjd3oWvz+2g9GhAFXp6cEBayYPXtb/Rz5PgkSXdPomY
Ai26gX6vKvO7OBuDfQqgBsL2PFzKbJJbzppQjMU9sdveH1hZCn1c6wixoZu+qwLv
wTzVlggHQ3y48/nLZGyWK4+ud/XImXlVMWHS4N83ZKMip1YJhEtQNa6h7qubx9Gc
nIfb6BJekPNLkHinn45rwRUkcxMPespWkw1VJFLrmNwoFbocmBn/yhLFr4Lwln1d
JhGgpoJxXfTEwlcmkwWE6I+BFQz2QxF9S5+QZ9eEEQFT4Vqf8p5rGUwvs+9Nzd/z
KgSu9x6rzdlyG+4bH9GiP8H+DiSQMfqbg1juLQoX8hAg6ARFp4qyUCWNV5e/BQwr
5wwPhd8NDD8w4d+HnEgGmcQ5+U5j2h13nHRKEJ/s+qke7O5/bracwOsRNiXN2k50
bGmJMYB1nDftQQlMwaeJSrRiWwgJX+F11ldGVh/XfG/AW3mclQ6efMNVETXfGjmm
QJgSrSOges2ntMTERSrms99LkUd3N1Rc/xg1C15uiyyip1Ne7PRlXMb1odbFdR1e
e3RD0K5tKzCmZ2qjWMhGP0iHU0T4pUft9J+3c+sPFn/V/ZMy8F71YsFqAEiYyeqM
pCtkNpjA4N5P4PHJZ6u9alHXBzCJorsbNrkgKoS+Th2T9PPnlJy5JpmAJy6VRyp+
ry8Q7B5HAQQ/asSd2YFw9j7kYv8Ur5dB737GfZUtnWGjY1PMeFglvcp6UTKSw1lH
bvb5JFz8K/meJJ4X+fdy7WmHfLjmJpL9KTkdFcwH0ACtcbwe81glEq3/vYapjMju
mKBUjMmp/4bZDRqnWfRQYSRAqMCgp2168HGq4uZaSNE4rVD6HvoXfolKtqN+/56S
q/NN5oApsH2IQjKqZ/y1vobPTLWxWffnPd/ks9qMW6pr2gLl1N3TB3dg8H8OCUWe
SYNWs6E2zxTOTKIikGx021G1zx9+B2MAB5ZFMHt/giljURhu01ZWPZHTDgSua348
gdd4IRlLNqSLJ6b5i10pwea2Fkm+/VZel6HQUIHdnYTVWP0qLGXlxm2awWbuEiap
4yrXOFV7mhbkPFHfJL0hVDf6G2BgHMMX6+O+7SCQ3mJr/M1jDTerD0NJgx4D+xxh
NdBctx6aDGN94Ea9G+h5B4G564LPRIsCBauTKCeOXuw9ZefmixVpZnUGxcBf83w2
/Sl2rmOIWgKBnDuUZV0BtJhQam+wTUEEjXbeaa91nJSBFXoByrRE6HOIjacUkRw2
dFDk8OmsI2ZyWwRfweoUTjUl1UnVqaSuVZDy1Jnwh/Br+B8XBVc2wGTAUjk2LWmS
7nc0eNi1nQG9pYB1g8LocNItnMeledMqQOoQys0AL2zEwL2vg5K33uzkPfvgGP4B
tYVFZFw4EY/1og0ITFRc7RLa7DpFA7Qp9NTuzOVPPL6BDc3jXNzmeyTyYjxJaVvX
UsR+HEziBwhdMd0W2E3IAjfW/lcKUs9iC4QYHPsuH3dubMeYy3O5ejWPu581sFg6
Nuj2tZ6yJPR4gZs+oGHw1v49nlf9/OqF3084dw7Fe6OXs5EniCVpAARifhws7ZpA
gN8cQdkFdiiR3stfQULCUI9/KnNqKqNHbkWC4PldK/onpJdE7ceV/YNkRXLp/4/s
pZb9p4V/9lDNXFg38TOXkjZvOvQx1z/QWA6MPnyS27Cev2IIEugoYGlc6PQYKp7X
6GbW43BgfWIiW3GNAFvVd40+079BldorhJkPcRkhBgymj4/8IvP3hrbcTjV9fPr8
HxiHh7zgoR0tVRp+znyD6eB8Ur1Ls66laRun/++VvcWghC5ckBHLyInqXdmCvC7H
27AyyFHa6f+3UkUDCUSCPrWO5grD3gvZke/9WoYo4qjbtBjdkSuMaQzigWk9YFue
hznadeUueXCqFYOBoFZLvPHG7FduwOlD5HeSmmqO5qoupi6VAwgNru8m93jV9yKq
m2GYQ86yZ+VlqkEdVJ2nmS3X8bstUcoFa2ycPCFVmA2ZzkAM82aC/t/ieepDbt/1
I0IuQbNqIPE5E4KTDw73tt8crje2loVjnqKhQgy0Pc3IsHYUArQEvXM02SlWkkI1
yYdweSEBeN+LpTLT/m023QWHPram/R7qJslazpaTTmEZbwuIjfOi00dpb948RsRB
t4llCuTePo3LmwPANnzUfYPJo7CT3vpeTyrNl0fFU6Lg+YiL+wsZJxFovfLArITt
5Q8vLzObzjuTsPh5UL4Fv1pem+57AtonjNac0I0DMNWzG24PpzUeOjE8LLm0QI/W
44czTVl/neqZtg5VfWKTf0rtGcsvMtSz1AlyxcqosIyozxPk/0h89lpdweHSFdJI
u6t7sguRtDSyzJWhD9ufl8C70kaeWMCirv1dOu8H8oxbxR9Bu0P3q8lnewsCJVL7
sOuyY2Gu7Q6m41oDCiSXOMzn9O3+zfQuoh2iO/iy6ya4ZtgTLxGGrIcrYCwVpIve
mXRhWfEiGjzkxOVmXa7TFA2EB4BQwrk3WU1FBdWbJ72XqqfjDT7cpbOLhSKJylCT
Ufo5i/TPIuNOplXQQCJ6yQUWqZEsjRTG/lzCxKhIW7N2p7/384Ttsu5cu3/4rMF5
BdzLYqgBSLO7s3lUqIAlPosAV3Thz3KkA0VfKOkFAya/42ZdNsIq+gOGfsnCU4H6
KhVhPcmxQhkZKC5s1wKU98W0c2Roko6FzBKYyheW6GDqilVO67iXFhdvKAgLVlDA
JPhokIGYJ0J0ZR8yrtJAm72EfK5ORcBu2a9Axc2OR+KunjFPNin3U3JjKmUDQGXa
yCUrXgPhqElQ9tgsCaKNWmY4+JrnT1QNCEd2pqSOwlrVJkXCs+YlBlo7t9O2kPkP
GgZ3GSRRE7QJF8khuqf83ffDWHtkqsNGsyvCX563VB8HPmrE8IG1WN4mGzxBGAoZ
pNlxLHDgDTp4hn565c8ocReZSynbCDJ79fel2tPWV4DaV5Wqi6xg4xtMQOVGpbQC
4wDaxFt8KimbZ+kvDdKIsd4SZjYtbnc1WvamQ3ic1cy0/QbcTS+kBQiD6LLDcx/1
Oazn1fGkBPW7KTtoJX537KZ8XT2C8uSCFYz1Fi8o9i0XrqlGLKi1fmN1NIZxTY+W
ySMep0K1pjNcjYXUeBWdlOqK0SXQ38ci73lFeFGz4jiRgBGLh4ZmKDhuxIAZYPEN
WAlHvcNYXr3Dqpvl9Ux1dvfq1HyEclg3n3OudoENzLucRUV1Vf6zfq79Fy62Gyea
dYPq5fmWHCH+K4uRaBOV6N2sbBxf4UTysK0Fjwft/xpwoddpTv8J85PsMR32MEU2
LiY9oxi3zF3gEAT1CtdM3D+OuAFFxS12S9xS1+lpnLvSVg39M59LSKQPwHfCyyeZ
qvLimTWxIW1ZTKWYQIWbfPefWhGfqzVo58EUNFxE8bx3NyGJF2cv7YD4fUNW896w
MLtmxQsxJDv1pJsISOGr8h54wrr48A/2xYjcio1D7alHmf+sW12RrlAlGoPb9yMo
O+tKi9gVkG6FIZ3tLq9FmOnNVcsvQ7qiDRncn7vW3tVCLdLwqkmbpLvnynZEYFUq
6uYH1d2xFQ6rCJ+f7V0h5XK5/gkBsYDMGPXEb3GC3ZLtboTsSeZhBWh0uiptmqJ1
2LIlsAqC1v0EXMRVTf5sQRf1cnyZuhs+8pF2ALgk6bM4FDquT5Z/C9LUhqkF0853
rxS5rhh/6Eatyj6/pvW2/crnjdMP5bjtpcvzt6WoWBGM+YfbX23GV4Wy5uD9gVh9
edZ++eJd3/wkPnrBltmgbLKe8qb1hLDlTcpBpA2gL/AmUerSWA7m4zO4eU9Uq4+1
A9LvNAJPg9eTWEgKrKFJfNh8EsXN92QS9lxu0td9cRuQFErFMLZwBciXIArOz/vf
t6jy5DDKijIL6Ppn9lMNMjbnjacYLfYPEaborDOOP7cxlwRgVbizZMfQ11mZuEUl
wZOvwaat1FxPBql4c6S0TU5e9trY5fu9pyL7hu+HQ04ms5qzrQmsBYHrIpZmMme+
xcCg9MYHeKfMiVCWvXu52qPvgv5jZECMsrjSEXSsQLgdDlCsbP4VIVpY62EB/jVH
ErTIX33YrpeTwlsY03hT2ouYUwm6BA3+liqJ8N62jydos5UERsrFvblf8iXz9A4o
1QwBI2HTNMfmo3IWe6lx+ZRBsGxuWOvTu7xKre49Hz0UQbyi7g3gG1lf7Qb6RrI0
gz/8TKRQCQTb5aKvZeS16A5V2MWwxNXfJYZ2brHQtPw79rA/uafZvmpFIU6fwSyK
LPr1RNqIUrJPw31Rsqc8zaRqcQAaXtI6RmnDdUPRMnQPY5lrnzAwvWR3qqJY1S4f
hULdWWvMnSziCXJfRzLm0b3vGGM4DJBplhHQVZdyXjJUMtArCkEsQAFoSwfT8kF6
0+u5gg9efpguJAwYFHLfHJ4QJeosknIwFDPs1E7KKHC5oKbX1rmkh8Kh3OZDvqwX
aIpJwBsDk0D+KxEAf+04n2Eyduh8SRgVD3yQTqOPVM1D12s1DswuvjryViZ3odlH
+Cj3gbFH3P60QrkHVzKiML3djiHi1OBGbCCNlzrBKhlLggAjGKSH0uzsh6NyAaoq
GCQ5k5TQ2vz+//kC43gcvrKiQqjQhaZUEelTdOZ2Fvfx4RjQ8pezXtaniE8lMESS
t1ZlTv0JbITmG3wTCpaGCjLSEPu1Wnsu9oyGwd32yShrACPRTRu9ArWlz9wyzOZd
qS9ydTN6PHuCWZVLeJxM8JthLOHq2jEFpZTsUJNrrfkQ4HQL4wmxHqJ91kDN7Y1Q
a8CJFSjFnqsDkwaQ0bFFqMmnvIrAhUbh/zWEYWo8TZT4VBX6aI3H3fVyY+v5HfG1
xoblJXBYAwmUfXWie+H/pjQRBr9Ie/hldnRc1OCEImrKPWxgcSLJpwWQX5f7fB2E
ziSPCHZr5sTwe2bRmxMc8Nw90IAxkRb6tZawqMf7ad3D59yKxtAxg9sMnaaHDHc6
gjsjkB8+xNqrlRJOmhpVYEoXIudRgt5/PWEUZXmWewdd89MqJAoCrCnzJuPSQFb5
942jpu4N0je+5769HM8M/dujp5muNt7YZp7rnHeoYN6j6LLDSmcKsnQFtkkccS0R
kYjGVvTlMVYb7uqBkQKKltihuMuSfuNUuyOEFaYHl1TmzR7xnHqjw6zscX4JtLle
bY/UVY/36tejJjGkpQkWuMuDO6IMOyoM6WM+VrBx9TDCJEFk9zv1Nmhmo1wf9F/r
4C1JariI4Oi4FhRMrhm9q7bq9myvUAUnFGb9GveG82DfX62G6AHFX7m3cGS0yG0w
+4wjO0V/CuEkMlP/zjnlF6sPxp9JX9HUJixKHAlgd1bTM0mvvJIGhjkw+ccjpnk0
CJ2M9FIRHAG+KDUQhIv845DgLIb2P59jaQPMuCAJ6az7xVnxqKrkJOonqlsYLiNL
M1eQBt/koNR0YOTGzgFLEN2ORhNoAaPiJqClBOTbJ65vWAayipj/ZCMs96ZBYczN
SWK0dMAjdQ1+7Rmm9D7vsD8X+VPGppNLRTUSPNIHqLI+gQNPkUeuOPsKXD8rQdrS
6ZF4QZqgxIfnHbYJQsmGXApmkSmsTEarTZcHbqJHWsmgaaaZGF5abEFe+KdiR7SF
XHgvHIUQUPL/ZmtedxNyooRnRmpe7W4Thl5rj8+wLKTPhuOluNtJvBlIkA0LKPS7
Sw5yLcU6tSiZlwyq0z1KrYi6hzejPEO476GlM662yt07ZYPQKP8mw36W7NQCviYT
FfELpOH3kdB+cUsgDZPw49lJZcmdiORMvUwCGxxLAdv67xeNwO2+R6y6ROTNBsU3
xHpTD+oESrzVkd18yaochMw6q52Sz52s7ynv0YaERBJOiO3+zKEW27pcxIclNqII
zMMPj/pq4Y8SzhzIJtcvKac2kfvQ/ivAjpwEL1BLwzgjJkLwsCKI0E+kR3e4DJp1
Ph3OZtsKnwbrhcR3ZVuPjSqVUXPzYYAgmp9CyBsBcTED/Q+/b3xiZu4RfS7OEaYB
vEABijG2CpkotYE/+v22h83zv4ji/sxAEOUecw/a8e5GXZDJQ8yTxzom7/uvVC1P
ouioLAPtvcqxtRVVG7AVjKi4ciSz+FQ1sPk5qkG4nlA08MBndP2rDaENSMmxY3u3
M9X9ev499IgIbUfLasITbHQswM6F48+oLeAU8YNQ9k+FR56GrIeBptW4whTxoLtL
GVDQiZqFUYUU8rk2nDC0ifNVeuPvHcC18S55emRvwJjHIdRRHeSCLYduGZH4UAeT
yPnnrBPF/CRSykwbm9ofeD4BSICDpvM8nV6P1rt7go2QFhHG3e42MiM8u8KZ1qV1
1QnDdAjo712CbWdNsSjaB4cuIq80mdHFmLrbSfbV6FEAzsrzLHz3cZR4l7OsvgMN
9do5fQoUQkbcoXihEBnnbu74Iw3/P8l4083goMcFJ8POVgUOD9UJ8Q5+mdXgmxNt
oXETEaboyDasDyujcdffHd+SeE/FfAOzaIrDPBhzOPcmFsAmoSz4WZ67s5YjnhoF
JkL560VQIi/qcCRmAtkDzmhKPrkJjNtxgdyTfgmiUej/yjLiIVsEJKgoN1bUiUwK
RxNdVocqL+NCjFmJXYZ8TBr+6hOVdvv478jLMB989awYRl6aATHcCf4qV1bRZTBW
xx9hjaxPyPjPdBuzN6Tk2BcGxWEJ7Tti9MgvvpFwXnDiqXwFAIy6HB24V8XI9XVZ
QcZr8lCTepqlmxHI9lPpLZHhdyrUxiKITxE8wVJkIqHknSb5sXZZh3ncZHlTgCoh
fCh/seFHw/op6gUePTFCKB1VoD0cXwtatu26sj7gh5n1T5dt6lTbffZ6fInVrJPt
OEz2v8cZ5KkOfnMewRXQl7YP5iCdtpPE7raLRCqFJ6RFFp1FjL5izOKEAD046PWR
jdX47yuTDVbCnZ3nduxBO3MVYGTJ7gLI0a5S6xvYVhVeloXHDRjr/YHs++V0Hj2Q
uqbikLV5jahJCbcDv63uTuehsBuf1M6IMFuNYic4jeHT++qWJNaivlf5nWFvju7G
FT89Nl0Njy7yEqWXmkL4JusbExDe7fE5N7+fUK8mhp0KvLxoe0a8vIbY44Q4idJW
Qdou5ItRZU/SD0RWGkWbdF69b6QnqJQBQoHZoVW7732emELRRUkqHQ/+7weMjdyo
A2BI1BskCgz2pIIDds/CFSGpeY2jLmMh+Shp+xn2KJmaGuG44KXWdeUKx/+fQz87
RnfPhaYuL21JqfuWPwkypN+coY4IV1uaTxk1eK3XSBn+U39dLWQs1F8m+7U2mBLU
ANSt6py+7aKbt+jYp83RbMokS2zqp+NZO4CmQod8h3FYfc2qux/3G8vl1h/TTrKC
k5Ov8wkw/F/4gJkmjrkkVN6PnpfY0LiRrae1R+1InYW+TippKAeLHqR2en/MJ8yN
sUznoU9ctEbkcMVNJZj3F92Qe5qPvf3sr+JYGP9o6KQSYURsARg7w56leeDHRkyk
IuQHS6EOtU8R0go6kXtb6FIczQsjFKeggOp+/Jbddm8onm8JnDq3dsND1cGxXMTA
IH1hqZ2jBXs66cE6ul+ehvRuVURj6J2qICm6D0SmdTFvtVOiCUYSm54SCB3YHkxr
+uJRjRnyZCspKfm4TbZLd6zznx+YnjeqdF59UyNaS2OPW93RqRrYB1RdZfQpXxrG
LyUi0Xg0Lf5UoSC4QZ7OMAxY5u3/BVN83gjo05XdbIIz+PGsI1Ix86x7Qjs0DVgO
vjqaLm+03tdavpzX+EXnTZpeZPfz5LkzlZ4aEpJPKpJqiByM3KTtmerPbPIa8cIs
LAqimIHBABNL92RxZq3D7C1H7BctK4xQZMldB2ryhUX4rCTkL0e3vCLpX+iqx0Py
NdOXbXUrZ03PhU4TINzkziCJncFMXPCfwcap3bxUTiE1p6gkZ6DwNeEzp1MYmcG2
ErtwA0t9F3hk2HUxRVSBmPh78Y6/6iu8q4PIiPmCAgYHG9/6LihJbH/RW8scUfvE
kewcToI1UuaA2kS4gb/8bJYji6cZ3LmWswkGMDBRkYSx/p2FyRVXSbRGqysWlUzv
Ww9GL2v3HnF39zXyAdcC8u5CmAsfFnNG1+a1oZq1gF/bAvEo2PVghC9ON1hEc5Pz
nVmLOTTVjLIQb9iPJRGiVDpXfPgdluWCJlfffNUeEtrYLHK8jVSXAzH06g44nq27
dyOXZwGI6aK3iz1bqTmBi1DrC2uDMf3u3VnJpznf4bTTh1Tb/hucyEBOa1ehshYq
X7bIVOB5ewIsq1VjBEi8s6I4RUWR6+bWUYp40e73Y089gEsxvcUkgDJ6tmf5YRIM
w6Gc16I1Vida+CMLnyUs/g4esBGRnImFsULbOPzUYWB8RlYWiKIKAk4q894HMUu4
ZVXD/NG+AvlTdrmlLlkNU/b8c0Sl+w3vufxXnLizjVd7WjGzIPaO6MhZ0Yzi4HWu
eSMqt/MVfYw+yGUFW6m0L75W9tKHJY52KZl8OtkrQy8=
`pragma protect end_protected
