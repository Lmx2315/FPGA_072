// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:37:06 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
VYlTTMksI7U7Sj4mVa1GYc4ATPIOph/SM6pVe5wufpspvE3uh2ZSyrXjaDxxfXaH
DCQEFiPH3dS3LIEOuiF5mvFi8r06INTHEfB/Sj/iIXOUBWRKUOU86fgwcSkZ9QY9
THWuQ9XUIHNXEfH83k3/Q0WUDQTGOWW/sjBAYUeON5Q=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3040)
fGHGNxBik6vUvjeTYVoHhincSEBV4yTuu+aNq53TlDvlGvgyASVPf34qAdvuYYjN
6iyL7Iq6GUrhBKuc6F1ipSwSXLeOhGO7SmFuEfAJOYjVDoiatsI6PRXwZ7Km1ZIg
qAshMdSo2bMfkT87M5b2h3e9lC6P/L9HZp0gXDbYqDrkmDh72lMpDcjdoKZt7vz1
EyZsjiv+RUWtEPwV7I3cOfMfI+TbSpVilGBuhmVOmy1GqKth2xo3sdTVZAXZQliz
9duwW+gotF1fMrIi/GB7QL+OwEPbt8QNk9uU3KVe+fPFJqx1SuZzUQimj2iDMhGO
nKIdknvvWu8KEW7vfaZLiVF9mFKeRBadj4nAwF+SkVtW3LYLdRlgFZkh9XpKKw2p
Lfl8idmP1NXKFVzkTnHcb5V1cdiyIu46Nq42ndlZ+RB0WDQlJLN0ZGHbr2URZGA4
jxyJ9SC1GpIqt8gpOeZew0p4RgYMdEgYyJnybVtd58po/7ZaDiNuQ2yj9w7k8i/8
Q/BAb7qx6z3SnRXJpCiWQJgvTEMZO+q/9SNlvSDe2JVtg/FPwdl7v4U2T+KoUV70
gE3vvAWV3JUXOXunuOoswaw4M4dpxrWAMYEigIkGLh7EIty+qNcJ4vF9sgvN/sZi
HYvtdSSMJUFi0Q6880KcpdXiR30QxUhNBiJVauNA6McxnQLX3qb11c1trK2WM7P/
NzCeVrpSWwaVVRK9OHZxNlrPuPa6or24agcyNBAN5NE/8jbGpGnnypvHUJmvzcEx
TxTSQCSx+r6qe6M3YzsntVEFbnLIRa1FvTI7gVmUnUIDEPTux4+uddn8PuAaS22x
JeV494LdcnxUIMm9+EsaHnjMlM4UsWznWxdNAJ47e9p82Jr9/Q0wNXQdUOYnw9e/
Nlu2TganSqC9wvdP24Xw7qsbxLVlB1N9tXAbPMpq9mmzlmgM1JF1/iCwirHlGZmY
dNLJ+LSLjecdNXaGn5xSMVPbq2tNGoMv0EMHUQ1mfvUTdtabXHj9W4rzdonnqGeH
egbOfzhQ5aPJBdCjXN22QlkTpIQbCqZO0EwzF06bzysLNjBMKEIUIzGGq8O6/0x2
xstfw1p4/sC/i0D9exln+jw134fZue4gxZp7Xe4bgRHMuM+CfqnvWmcYd6sVY2XQ
FOOXP/8tw/jkM8peCpW0e+PnQ+naKOVNGp50oTp9hnTMt+lmjuK0DcD70Ioazpgu
r0AbASL/rNPQCzS1YJqygPt8WdGea6EZTgfIC+wVvFw209PXI/nWdNLOg+06CSHf
X9mkC4SF8LZ1bB2ngnWK4W62mpcfbepWzaBt1bmXZIcIu/esJRNjqB3aexpy9A7X
upo68KDIVJjXRZpsKuS5KOhIHnllxGqZeU0TGPMIHKPZTfcF5tg+OO2+e+aNWIU1
7SWF6ezPvb6WOQyhqIGBvoOcL7jqaCdWYIhXopQwc39b7keZKpbFhfQRopf8rnel
37HfnIhqfa9N8xbQTZZQ+JWZikxmbcXX2LlA6b87MIdlzcaP5aQSurjVj78eDt2g
g11Du3xOZVtu7wR3/PdHATAVekA0sghfuJb7HPnMb+i7gf0+LZpk0qH+UW2AzV+k
7T6xXNpLVKjJp6c6cbbY89A9NKe3g37tWRZQQHaPnNle+5yOaTOCR8fMvqa28cE7
BsCeVCO+6s2cSA0d4vjkRah2vRYa7sihz4eu+IYHD+M1UUeqB7yHtOJlZm4+bcyT
ZFWAPr9Q5UPjBYZQVnooL0C8wje0P/tBdVL8X5PfWpewOeIy7rhSem/GPcULb5Uk
LwDN9PG13b19+P+cG+stsjrX7kB2zVbhMbP/O58jOrekZTbazzMk1OMNL5itEuGW
f95tX9E7pHxLh07abf0b7QxRTvzWSCPl5aeyii+4qRCrQCvGVuIwCZZL5oJQICI5
x3OYmbVJrZ7cUX2mXFXAtbviM5ZFYFDzG+OqctQ5S7FkVFYYeH4FOjzTg9Mz9sLb
0IG6gYhd79GxDMFUNXAaF3RKTvXkOeEVDoc9uMeLva0rCCkuTE375ZI7tyM8cFxa
Mm3i0AizvADRbhb3Mkc/5I3pIPS0Eqg06MWbE5ShqFISzQ06mO4Mk5Sd2fA2CSSO
b3qbiAlunR0l+jcB8sY+u3sGU7mupYuu2S/u4oLdaa9N1stcE/82YY9N7hljl3XW
8CiD+1nypO1O67AHP+Njim1kGtx3C0p1PjRo40RctcBs7D0UrwUL8t3EyLaXMzAl
dqiq2ADg+gRg4v5BqGxi5Nb0UBDNblSY9xu802kIKaYsiSMQj4LSr9lR5crXOsdA
KmEaQjJIPq9qV6hsKNho8AE8zXvkGmCDgXGh1Fo7bSeh2mQ+91HI+nYj9ha4Z4wj
OYKxQtI6UjwDeLEVaUQ3HRmS7BU4KugP1nawF9IDpB0nEBae3+P4+rtecksHY9+H
LW1hXGgndiSbkboV3LKtApjpQhlK2SqHQy1CIz7ct5YOJB6l0Zz2d+7Z8g/Qc1i4
9xY8OjC0A0RpgSknluT+SPUuRvoxNTGASFjRw7s6JFU17d7NqFfovzDufyA4DCdb
j7YkFy7OoUs+2sIUFM5F9eQ2047JqU7XtXQH6pri0PXSFwEsx+smN3Y7ZAfoCUNy
DTod+qsJcdpfA5rVblO8GDmFpZk5/6khA7mcY/8C/5lKeeH+Nql0r7/373w5udiH
58dW//5NYu242b1Xw/QR2kkxVCf0/xd+/ZcTdwJQFvKakpNp75u2zjx/CPjPni/7
quUB0RQjSPuQHbQLv86mm2eawa1Vcge9QCebWBEgvnXkQH5cJ84jslw1wQ2F+Rjc
tc4j6Pq/FFLLLp5jDaf8YDy0Q8Id/MiShY62EVyjyqYYNJiFnW/MD7+9X0sCCgAz
3P1BsGdP7AnmWNViWGJog7bylFgPzgO56eI7OnERR8yuFDzhbEK/9q5OpUc9p++b
rown2eNvNmOJrRkG4rgSS7aw9Llmpl/shvPAuUiZGl7bdQLJo3gyOG/KcxDlsK/3
9o8R0pPzItVgEcswdvq0sqQWHBLCNuKTYhAx/gsUrib6SkwIMACNkDREcKZifWZN
xr0HqrioH6vOYQGTySczqP26h9oe9wrR3ZE3ClvMLzUyxsbaCsxYEtlZPoHy3/p6
j7NSiTqnTmo4LkRguQ6GsQq8C4PtDvmciQ3ejQbJIaDpiB8DKf4ezl46MsOFN2WO
kHLDSkPYthnsAZ5nngcazYH7BBaIS61etvRRxJLi01XB/J+vY0xYJAvEqonbjlW8
bJyM+fR2e0hBi59uDchUE1HMWXwhbYcPDqc+SV9NbUVLqQSUmmXqAi8eAhGU7Z9o
kBICbCjV/M+HKlPeLJaGNAcHJyg+eYeEtTiJfMTi63tbvBQVb31C60ZvnkWJfnHO
lqH+qT3PtK6Y7zUUX9g3XaSoskEaf6GWMveZFNZ8kJTcUYsKp+zagB3N56tcTG5g
Kn5CGARV7W959UvHUZAsjYlZ1w6akmQXVVY8kiAVuu2EO6NngYgLL1wb0QWpbrCZ
Rmzf8h4CAxlhV4hUVqipiK4VJtNBHzsBdXKAMpDKKw48chNI/55mH+2r95Buv3AO
+puMaBV1LoNGBPa98ckt778ZNN8NfdhK3f6estKqd5SU00XaRMLfQrKYTcyLyztN
ClTGsy2YfADC3Hna0OcdzFcldb92kYk2PQNLxPVywtEIIONaei5dwPIx0gkmb9W5
9ZZC29EziB9OfhMbX+Tzf3tHEpiqGTBM/+q1bjgmWN+9z/j1DFHoqSvVaRRg1nl2
0Sgm6QNSfZw5c72rEwsrnbteVVhdoAiDe+SXE+h+22PQ5Pd10EMIsSlPCAO3qcIL
hITy/ZE9qC0tX1vL3ZNhgHxB1XVF7Biav6Ev0Gq5QBPfeHDUfwjHqjnDlFxzurZS
s6EaJW7zYU0ViLQjFw1yJLtNo0XM/avZbpXZf9BX/IdtxZqbQD3jPCapCAVF9sHY
AuNOFKVF7ZDgiO29R6v/5pjaEOfS3O1x7AWdXRTid7tZsUqScO71fZ9Lp5Hjsa73
h5mpYtkoogYSCBOc9NBhkg==
`pragma protect end_protected
