// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:32:31 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
F5h9A85IdnB5lz9co8ayMjkQ3xgJTWeedy6Q/BxrEwA2KAhuUH5uP3HPI5J95oSn
4PWCXBXcSW0LZTWwXdkJARCYIZLQSqBoVjv9KWDUwuLXsNHdIyCzT/MhmakiVyrK
kt4GlyLby4rp7o5iQdRCWGIbZo6YbOno2NoN/j+fzoQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 28160)
g0PtGM2O344xF9oy/3OatxwclG+xOT3rET0ceP6Gw6/j/0NEi3/C0e4lLTVA1hJI
VPOiO7cDn244VSTlozmJM9TjrR102jWHBb/wb0+JTutfn3mAIQv+ON74kLwGtQaO
0VZIm/kqcEIBAtznfLf8yw52uUlIqtHALXygfXVlO8aSQ3wjK/RFT6LhtuyzfNpa
2jp+MyVbQeQ6AIlXiC2EnN5LFfrXSonyT0Li76pGDhYMY48AzE7uuGuUIZ8zWu/G
9kqChWaAhZvUpJTT3ag0dTgTIUBCutwpZGEIlr2KNbaWutH4Z6S5+CbxL1hkoIvV
1PdvivjHP4jjqJLxYkSQPWZBG+wT3h+dFa9Wt8NSowO9g8ydB1HtZiCSCeAiMLjt
4+9KlsRGCHa0J1OVNluMzkeXrz0jb5CIRTGJVMhpUdiwFC1Qp6odCgun8z9UQYBs
mgUWuz1aVTxiilJ0L5uezHcpcANIY+yXm4Hn8g14vdGcqBmyfBsenskRZduTCGvK
94xynnBtdfsQBx6iqCyCjtyd1BxpkhMQNjKFTmplNHFsz/C9ph5AV0Ae4AAz/k22
BwBZkHRhGNWzySgV9eej5N7qEmvwOZp1IobKrUBpP0Y1ixtaqJFYvgbncYS8Y0Bi
a537e4u1ypepWekAo2YjhnoDSMP70IzvPLEhVox5T4CJhu7AXL6ZRxV8vPvkd5of
6L7Zl8nKQotEHFzfl1TKZfo+oNDRcWxiYG/1Kmp9WK303+2t0skXVb0R0sxdjqaq
jnkA0EMChOoewSEaa0GDjkew7XH4rgOUsjqJBMoWhwJxX+ptJxiDAGmT9k7rndGj
y7gT/j/SUVQNK+SQ8Su9m5k98mmhgN8xT0NDzSpULQFNzVN5r1mfTMo+6XrzHrMO
wjIKfkg4PBqCMklPEysUXOR92UPslDmvFOzca+F9AXuf/Q3U7zkZwdnP0p8vISZi
JetAgupco/6Eprk86UN5USFWJJF7lN8mD0qMHsP7lWEJOUftFqVWtsr8ULbRZ2GP
tqAkfyuMetVKdFgUH5Ujl0wE801puopBlhCe4gSicnxXiWhAYEmve5TOgKkyDIGO
1CcxeVavDkgt+J6TYTjV1Eiznh4yb/y1G9h3y7OttpbBqADrl6yWOk/NnaxRN74I
OmXLT0FFitHAqRxiVs7yrnYb8XcMvTtTIDKZ9oqZDTrIvAVgGocoOyOs4lm88dSg
MgAY2K5GRfMG8fIJpRJg0l8Y/2hNpz2gjWlIVHx6sIpZiOGkmcn0ATJmhxCqqmnr
rsoSBn39OMMtd6UhL2Iu6Be/MfkHZBLOWjUujuVi7WT82q1WOnAqYDVhlVyvOGad
eTGkAIgU2rYe1QqxvDOHGoxOdxB6XVw6eBwEh3DDzcCKX9MtLXliwFUPVw1G313F
W6ux/DV3NAjBPumLFHjwt9yf3tCIdW+9NFJAYA8e815goERZede3QESr4eWisACE
kjjx4MTRNUV9TOaixOqLU3XUgntOwREBwkCZZY/YCLjA/i+j9naljdq9cNZVsdCX
NeCxPSGVT4HMg9FtTZ2HA0T3RBTGVvn6HxpVA1NHQpnFL6mUcD+gpGe/UPuwvgNZ
0C+KWv5LtBtYZCpierARrtleZSzxgZumMXhu92ZxZpEy2YbIU5bozgNTTGVu8E3C
UcjXMhSIZWQbFAjK7n4l/UkmkxVm5fN8izKPW8sthzZiGzPNcQr8v14JnUnuSJxV
Khpv3rcN9cZSfUpfHVyVN/TrOiphDaVA/hto9FG+TNFap8WNfgOZ1HNae05aKE9U
A8O1Ql9OJBCujjP1pVM7+K7v0EcfQTej4KJ98wfhKH4R5Es8KHfZ8kEDIF8Khb4s
NWbkGnxHddhWAszLYZJFPMrIBJ0T3tToylsRpTPn0PDp9aQP2fyy1M2Bt5BYI46n
igz2w2LSV2j33i5AyCxvNc4F56sa0rzocnl22RyUobVGWBMrfRYxkfZAR3sWEmOo
RHlrXbnK7mMKM9iSY6qWHl9V/5XLvPRVU2lX8tvNdS1XLE2Kl39qtQwUx3lgGc7B
i2EiZ8cL4h6LwA3KDKwJpft4pCm4XC1xo9ybx//tjTOQwtwy0OE34O6NoLCfZD3e
xyuXHjUfF7kGTpPe+DNoHqiDFfTUuOdIySWLjXrCpjpdshn8+Yr+PIn65dHcjkr8
xQm+lQ463pETr4BwBDmMRr3F2OJt4kCN83KDruavfqaN1eZ4hXdMIvVf/mDGr4sT
5aDlAe0eKyc+vxhtnUwmmyJ6IgV1czjs6aX7iUU0XiSkcl0Sv2SxOt6UCdIJvr/t
0ulv4t0M4Ff59zhhablgHgJ+Z3pLGlmsNVyp6DmSRRFHnjjnbb5eqmCJs2Qhgs4y
Z1nMcJplbX5oIUXiOVmQQvad72uejfAIgLrAsB7T84fDAE9uFakx4ZgfvOlIkfi2
70eoPZEZ+FTucKudZ2Uznwf1Q2YXb43hbZJFeAG4LxFNg6+LEBTcSpKy2grwuFbj
P/Xg7mIHtBLM2u9HMl6+LNffqXMEW50k6GHemXdMTsBUF1YRQkTSY0iMvXy2aQx4
YMJhLA/0dasrp+F0O7dJrDbT1shhO9KyZ8NhBz3wdNJBZ8MeSxvfsnukdd9YQMNx
+RDmtfr2nwMK2PhLkgcMRqWesGatMHBofURZq60cNIlnxRRqOm8fa6qx3feZzOc6
j0qdWE69LGcSwKqHrGja3x2ary72qrXbkoI0ifad0zwzMxq3hKQ6NX/VvyVb+2UC
6jL2Rl0Lktm0kWRK+h82AfV19GW2U2BVTZnw5mlujkIMiAyuy92DJbYxsKTWrZA3
Xc3/duvf/q/64Gu2xxNiafq07t8Cbh4ph3QKMAtaT1Q0VnMl0dtTMDfhlSKYEYhv
sWyihIcHjuce5JBo85c503q8yWjb80XsKw8CymwDVPkRZTgI6gI8b7F9VvnAsSDi
iJUzpr518+ZET36IfW/6CVxDnwffcPeFjMfGe6ZuOF3PIe67kKF0Z71Kkw7EcoW4
5kStJR5BeJW/A1l4DWNLNUn+h9EHl2I2z84dLDD8hZIifxXzytBMXZW0p9/Pj++m
Ey/gBM5wL+uwIhdr/ZJ6woaHVAbeJhDCkrCvbCtCuxnFqNpv2Urg3mFQNqP/oeug
+go9S2PshLIlZjLDaBVfTmvII2pvITXnVk/YwDb+nxRLavZx2LqoL+kpiqp+QGOP
9sly7pqvf+84oahgO5+6Gom709PpQYfsMa33EzKTMt07qfa6+fyvXR67EF8LNAhO
IphAMqwf4cPWEERxM36Y9/h6WHi1tY/FSbO9HIs/+pWJ1oGDuHRG9Zg5jCv0CjgQ
NwTEWO7oYolK2Q96kdwVofO0orpElUuzv0BqSeenDobc50vHSrYPmT9aC4KdRyqT
LTE8yZpcY9VCSroZp8Sxq7DgQYuqbvkjO7cM6lf5ebuOf9ps5awSn+fVAKWgUIG2
lt3FvSAGM9RlJ97yFlaZzalFLVSvww/kiHspypIljEuoxVtUQIFpIltrOtmZUpUp
UPtntd/g1Qy45U7KctrtxUwIbVhBCqBMXG1N7PX4SNn7do9M+TRnI7IuAmjz98US
ZaPiRupGmgFh3sLnapj2QNi72PirrfNHY6uBoUksF4USOjz/Df7LZXhBuZraczTd
tywlaaAiiwIXQzfxa58lATwCXDtmUdzvaDUVPoGZdGsFKAp0Kl7TYo0eKN4Z7SjP
18nxHzMfRKEy6E7Z/VnwBYDLoiLYYdUjtPd+PiM/zSCdxWTIEiXGeKkxZsHtLEbr
UV+xFNVhB6MR6JGPBfVEN0FtMc1CDrbddsn3xDy6KRWO4e7llsF4TvZ5hDGZwGIA
lcvrYGIEC7z854OyTzaAXWbrGbhek3L2gJLPUYayMIAh2N93fJ6+W9aeSN3PaAbL
KDrpU7VGuztmBCtqT5eMqEM/XS1QsqGqnSWOZ76Enq3yyS731qt9rmeluXHepcAY
LF8DR0A5kF/mmNFRPV/75trdXeNryESnXiVPAM7IJjI2NPpkjeL39laZ9ZDoPOau
Hs5VbiGfa/HIJQ8JMeCbbvrV4ep+wKgUikl+pfgyi+FG5EmFRQFBiFZzZv8pMktr
JNsgvlp0Fd1/ZCx0iGk/6hh0uMRWyopwPUpclAoWyduh/zQji0LSkw262R0440LA
fIItfSATwPOZZhM5VVCWVB9oS2q8RBTfKKxJFNWr+/tfu2VQKQracTlfNvt/znaD
sDsGK6fYf+Y+VZVIp9EOtV09OMISwGvExyfYoOgi8YEe7J1tr6DUKehhVSrfk/3y
ukQHefPXa+ydfGuHsuplMmE8/QbHyjzU5x2GMWIUI61XitasB1rVENMJ1ToszNkz
OD+6eAaO3+6b7RYN1a10acijxqaw8PGmeTaayQxN4vzIXVevTaHt+HEcH/r5A3XW
DMBTQvMYV8FEGpRWHJvMGS44dQRdQ4U6PGGaZBfwo4na6ja/3vVtxVXmo9OPRXEI
JsRNzaslSFcAe/JUIhyi80KBcLsWXyqpAfj4TCd4BvIJjw7aw9jdcPbB9EIY3GNV
BW82VxVFx12d4OCBhI/cUiqJakzevg8uDS3BB6ReIDrxAhGwG6Cx+IaNKs6iXTfl
bcOPrxS243NqtC/N6C+/cnmfqXpD9EuQGadSTuXExFDR9KtPkCxUJ3gNj172aoCu
BsjUlXjxKjXRzsDQokCWdus5Eqa1rx+SRBWpZYVwda5JrjEZL/4B4k/7ftvnStb8
2o4tK+I6sVLbGudWKKH4iINAOTlX2u/s4R1+G3d/759qLb+NBsAZ5e2OT6ds0RRO
xurzDxDanHSPx4kDLoRH8fSc4cydJeoZAuDa6BSGMVnzB8/tZPAFtyUzhsaCINgc
fdRDvdW0zUGaH48P3m0NJ/5viFaBB1Xlj4tHVuWm1jU2WdXKpJ9QUMHkrUixGdZo
cIsFx5dl9o7W/B3EXKHEJUqmE7uRKctgqU95sRM0RSiQGQfk/mKGPeOOEFweq5HK
aUM9TeHugs8yaNIQbDJBaYGuV3ZLI+kRkt/lDIYz1MHSLgR/1iFPf3rMbeFD4JnF
zoFDT6JBA2FXAKWME8+dSK+MUNWNNQYdvLnGLV9gL5OP/5iCXvhhiQnftW6IScnE
du4Y7YfQXpJ4soC0T4niBOSGQhdmNUwfzb/d1GZUWxAneX9rBRmZISniYpHWyrfX
NcCN/PwILuIY6Pz2VpiMJAExynzSfuukMUQTP60aJvW3V9rTLAxpY5uBQ4x8Gj6k
WkSeiNsN+ZguyOw1XEA1tZVQfuQFcRUajC9O+lrJD5OvS62LesQdjEC1o7MZAJFb
dgUnyM/NVO+EBwYgRYkMDQbnMqIUS6RAXRvb1dRUvbMR2N71Ab+N5U0ydmBJPrgN
LG5yGycIt5D9q5cpQPOGGFFdD8RAMfEEQin9kpIDyyFBZowhZHdRskgzac9VAKSd
G4hW832TBA+q8h2DmzGFHHmfVx2BQs6wvnKuSEvhrL3xgErN/IH/6kRJh3cUEMQD
nuS2yvPJ5OqeNG4faRGnMinU9dY7OdMztkVqzy97nQbbWqzw4/aUWGB6xSHwPZK5
aAS7SJyQd8PUNL1ty3+wMyD95Oh28u7fl/BZbEE9NRIKr6JrU1aa7Cuc/TTjkHNE
DyYpjcHzwO6CLJxdfm8eMsq/PxoFP2wpnmzpMqQXESZOumBVPUt+YSj8JxZC122C
4b0RUeqc+BpQjdEG1gUOqzB93HkuQtiADbTSSbxZeYPNxwOFO9sjUQYkL8UjEU1B
EXCdYJvBPC0rpEFgRUQV/91IlCQnEk0hnpe4MlY8H2OWrmdFIRGQdyj1fukiX/YF
Q8RaPxXyLP69B4E3DxMEfp+emkqC2gpYPNbGnWgLkYzrHLpP62DpZPMJAskFMiAO
Fn6wjA+ItliIsts5ygEnduUdl5bcTHPHBZtYfT1BW8fyxUVkFNqAZI27PxyQ6fm4
dV7IRY45F76YClpW8g6gIcoU+abbfdguKLFBnzES4/6RGWZ0c0DS8Dwtbsce8GKU
jAvMXugkaf9K7wVkGZ8KUyg3ZMkpbAZUaDVUYRDsR7PdMF/TnlF5dkteDAhy+H6C
fs0guneXs/ItBvLTA/rgf1Ke8Qt4gsbX2qx33fdNOUI/+zQU3eBHQo+LC3Q2l3bA
aodu9SrAM7i8bgZ5Mwc9SNzrp3IjPVA321UI+K45+1AtW1fYZp4iK6au+GsTGwlv
ZY0RNCjw4iNXuEYp59pXv31tdAX8YJobc08SsPXGhLaixj8Fdk8tk56BIG3pFTfC
pqnmuoQDGYv9Za4JldTWOkyDgY+O7jyc0ZD4JzrUvqqglwdoD1FvGh03lGXUd3N8
4C2PVdZJVtxdmJf21kzGRf7kJHgqG+mvaaBkrXuo/UoTw59ILQvLTk+WHdroyB+W
SHusCIJz3wegET3k8hsrwG4B1s0wIU3sLatzoK5Hhd1S6gZSO2FsN1NwjiSOvykq
s0D8fh2Q3705UiJKIOFqmGg1MGvcvacnd4glIXO6R+BlE4SXptqu7wZj/dNKOwKp
r0aqyd9c0Dfthxr2itugrce92kriS6TJPrHhDG0OopblDmzMWdwySDQdbP7yD5bc
5LZKFkPzEELkLMN3Uk1ky5gIIhzMxE/qmUET40UJAsA0jtF/oTw8OQ31aCKudskj
1QSsliny6WJNLzJ6vlYaoLhpIVECinY9pEKL3qlcUn3tW8Un3CWzvOLxT/DJD3d5
DLGRXDCILsc02cheVibUq9FyXC7rJnTZPvs5dvMUap1i6D2f7d/I5gwXoLAjuCKa
kl1g+6K8d3XJmvJ6VD0okRtPE7ggpuL316/CoYLpVIHqb51ibbPLR+L978zIcG75
suQOINYc4M2SEIpSCcqZzuge+pXtTfmDFghyiSNI+4z6NrSsY1bXFDALcN2l8b/a
TCN8q9ZKr17P/6+QxasVX9Zmon+6SiyVijBm7RX6LiKi5Xwnwde84fmy7XWR2rDP
J75ljuJCx6DSHOviFgsp09lis42wSelO2zBXvOJiAs2NEGJ+hOS3Xijzp69YUXN+
fUZXHaxYzrOyVrZKDUm9onYIBM8gnIljClH32rZ3PTMho1F0f19l+Ws/xB0x7vS9
rs2d5ouRyQsbbbvXksvmwjFp0GQdQZ+1N9J4snoy98oG/d8gPZun8lcg7/YmiJ4G
atipxxy0blaTASvM98OC6YL5KkxZPy9uACfZkvkqYbh7e4C4nNjFH2c+eD9szz8Q
UlpjAvusatWNVWv4M82KVHzZ12EGBc2F+l7WlPHvr12SFOdTKzKDfvuOI+vvl8aF
FOnKG2b1kZK1BrYRhLYJEPyMWpDQeJwLUQyIzJAK6DxMPfrLTD02BPcSrohXMuAk
MQowAwhEVghuUQPTSf62YEv7Tjx+jnKmtAsyraBF2cYTSNaXZ1bBzCZWuJFHgFMi
JZodu29RBsfApTGouNCYKPzaif34pBkw/Yg3mwePYF5Dza9ulJfR0Bo7ktwF8915
vde++/zd/BwsdkggD82naeyIk7xqwZKA9YYkmRg3HhxtTVP5i/LWIIKNie34O1Uy
8nx2FJebFRe3rUjjD9woy7Z9XiL1P8EexiElLgpk7Syoauf72g5DTxNLk4CpiDEh
dvSuIlVjfigA4qNy+7dxaCLNh4w4GkhIknjNm/ozE2231wh2kv1X4BCKHMoqs63f
NXwcG+zN2eDneloe1Efsy6u63OZAvNdMWQdLceOYvePqMtkthkAx+bmO4SbFqDV/
hHy8KkHQEJv+aCEEeoeabFicMeoEQHPj+ZZw7LhU0GyxIhWK6YO5fuOdpYGpXt9R
FjsZu5tBhrR9AteUCmbygknbxZSVafpjqx4nLP4GB0DkbIY466eOc+dj+ljthA50
IBcQC86nrdyzfvC2BBjgqqgrElEIUAQBf0lp6/wxRtLYcs6cuHDTjNKiHYuMDN+g
bHJDWmDz3xukax1TbAjYCxkpdow+7qgK8P/GK3DNQBUHy0YkM0Lkj+8UrMfLhse2
xVq1KDeXCtacY+nmitXlg+S5jSVukSxMrjSzRF5eNqbrLdasK2e9azS1PNTpHJF4
ruQIIV2t+8XU+c3Ejy01OAYeRDMm3QrzWZTQeR3e9GNg2RnKAnrl+3nupUNUfxgK
ZJclnC8v3hZoLHA621x0PnTsBf2EdmbBrKZ26MzxQC9LVgsroq9NMjBp+h+wt8ij
DGi0n7N6GKPf5oIAgVKWl/FWMnPUybU68MFrtly9cuU+MZc2rRpVl+IdoI4ELBZ+
6t8ust430DdGFOcR3m3mEZtp7Z9HGRm2g4eLoXVrVXZLNqmyOEqtwNwYZw4k7m/q
i/n2zmcZCwnocG0p8U3u2ps6bGiZleFo6S4/GTzsqe6rGObaZsuKyp+urRMQ9qsK
uiiddatL448pQcFYPWl9Eq+9k+4DEzRh87UZ7MdX2nxuGCD3aduOtbXcbnmFKwvZ
ZZ8DGFHy4Wo6lr5feyYVe+BtWqvH6gUon7cJ4o+bQAHLdtbqr9WOp9LPRnQNJK1h
Ewevs+4t//fSO/5OM2gv8OuiW1w3wYSmEh61Zi0ZSCZtodNvM2vH7mzS66wIpjPn
EB6VyI0s2EVIkN24hq7d4BhdE/X5UPLSj1fSfsBAWpkQJ6pUsb6w37D1l+/rjPpp
EbaN7LC9kz3NsE4MOQJSqPod5H5f8SNGri215J19EIC/oCr46Z/sXkH9XLUVuclb
mjwdYv0XYKe7/nfWjVSvrZy0YguBluOw9kJlYeXcPNsXrXE1NLd6TrUFqJ6HzyPF
SWEeH4B45dYwZtEjQHo7HgiCTRrD2hnBq/JppFnzxl+TfCZATarEVAb6xrwF79jR
eTQcQjXK+FN+ItknMvBSFox0qXRTPhSDwecVdfc3892AseAVwl/egiHeUiDi810P
vnpJx5SXCNmC3siAzavZBLQ273jdE9u0hhEJ8jJYMH9KMQJ6KM7jOxagFGMamsRM
6qR+uVLTjCn3AGPurfztPvNFWbLxif+NjxS6MY+aarQ5DVymLy/QI9eDYrTZPUx2
166oyGha75ds3VYfPC9V6C8vlwQLBHPqKMp8mrL2XUcYNrmUW1QbEwhAPYXhN5Fu
kEJIYGEjOHFhz/y5JFKVNT/PnxvOTIXnbD8hyr8zN8ADXzlLi9rLlLrDjFQRbj0b
ZRxB3mG0L2KETinaTOTTas8P2lsuvVFcrkr+5SNoxEiuWS+E6UjrnCvoN0nzOm01
AHr2P86m8ZTS8uP6JQL8RsAkbtICFFgUnRsJguIEYwbSUktaQiE49CWjSDod8VJZ
kkbvlRNMM5IjKv6T5KqhiKBvbLnoadJ07aMNJI07ONTcVEeTcNdIv4gDI1obK3CH
SxXZHBLB7lsmPG2P0MEGISaICAMWmnD+wLls+RWJ/RC180MxJ6QvqPBOl4XTIPlR
ZYLpo/FuaZhYYS1u90wvJxWRLEEEX0ikXRYDYUfDbVOaDQZZ86I2A2KjRq899ez1
77no8rggO1S+tpVuJRlnQVegv1jnxfFtOcnGZ9Fq+af6lu4f+M8qDgdqjxIH7zCn
6A/bfyIFow1O8K1Lk/kISiwp9tTSgukhS5l/x2A1Ke18Rk4ft9Z5Tg3tIA6HajOP
yj5Dw9VfZ0PoXyAEkeHL56dvBBx1Od12FZOLMx9hCPnEsVV2fSDUnquaJf7q74aQ
FD3zysMW+oKBdyTLhEvD1bpO1E7NPPPlnWZ5/ZSLp1KKwKTPdeDJikipvHURzrHl
I0paJpI999WiyPDc1RTsTFsBvwoCUXB11qTtikqe9z6/EpZsPSiy6QE9LyHzDgpf
HCDYyaJ2gkS1nsneFoj3UEO6tWj+MT+Ny57GSeRaDzr/Vaf2ljJGApHQr6IxS/rH
xCeMaI99fKifFc+nU4iGA3J3O6yHjA1CRaqhcDnw1yFzf8msZH1GPzpc9Ybx1N+C
pje0s1TxOM/3tso+caFup5UebwCiHQS9lHtIxeClfwY2ORYqgB9Ue/hqDkxJnclM
pkQ80EEZPzW2xmU17Ce2fd9JfeibgsLkp+fckiiCVKVo/oP3+E/CkCpQC6SlNRL3
MVktrtyfpC8+2ERoaZYil2Rn00ncdESwJwyu1ZJ+cD5FGl1r/GJQEFT5koEw4hOl
3e8bTSGp+yFU35alpCc19ypiBROAQQjzFIctFCVXOxZd3LdH1XAJZ6VmbO51UZXo
G6teeBVh8Z3P/VqvrUDgqHUSOd+/8ekQksYTIW1O2EhWBc80jwYDXWtwiJTLuawz
FnS0BShL61hfFafraIWbnx0fs6Pr18IMcruci+oOrPHgx+mrhUPKefp55GzkC8oe
q0KsDolXC5oN5isWTpGyF9Wt1215vuYnrIKcQJKDii4DSuqXNiq3NLhR2v53QTAR
ChHPYioYkORSAUiYC27wRnsj/UXER0nx1y29Y5dgAOY8msc+HDwD3be32IOD91ot
KneVRIgK0FvVSwD3ii4sb1l9ssXdF/ABmyPrdH5FamI2U+H3DinjW0ENfknwCk39
Ipr2zITpDzwl5QYJxuK+co/xn+d+yy5d2pZx5gd39mJl0mOrxfZBGsCZQ04YRZbz
5oAF1orKaHHDQnjP2JJxDbC3FnIcB1b1Zen6h3gE2gdHfsY+OcHSzDNWBNGU2h/e
g2WkBkrk9zjijXpGJNAp2VFo6mKRdk9xyZiSF7/3or2zP4MkWzyKMQcA++CaLt2E
IGb95XrVXwagl4uwu0d7x4u+Mh6tDXdsbhps2FKzTUvUhri8a1ux6Q13cJdoy7uV
DOIWShFnwjUtRHdRGtsRmqa5Qt9tu/m7RULLnfor0/1sahK3UX88w2K05wNJXlvz
a9rzcK2PrEOVkehNuXYTXhon/97XWN7cTAU3a6bJlc03e1TOzTuxkAUlS/SdPG+e
gOgjVaFRsrX47Us9iCH/HvcfK9/WEdFUXZE7HbO4pgUOuvM1a66XJq52iV5JoE6X
0G0kh0p3oGoLkgVMYI7kdgZsStaKQlgXtuuHa2VF6OIkC7CE0vWPPAh96Aj/gQ1a
gf9KmMIXyNPlpIYi4qT3w8QxnepnFeGcx8ECAm62fzpoFMUH1/ml5IJXpO+3EKyT
LXKm/bmp8Xt+NYVcVc1FOwFY4JXQSvcHbTCNJYqGW08AW4shCrKzTOtzwPZrcbdX
4qk8K0U3zc/0z2dZiDyftWKQwN6YDVZF6Wv2dCwZk0nhaU4EO19iBYM+DGOQS4Hf
iKyoTFrIUMMhk1fEO2psyFlNUpQ7sZsIap93UX/pHPHqtqIN09RrnNkihfDGRXr2
vz5B+CHEu72JRU9WGcZkXhhGae8+hprERnM5bCyEUc8ohqCknytVq8Fw0lCUg60O
2dsF80a6xNaZrWDBpC3ldANK/OQz/3B1Leuqd/95zr5c0+ZNdk5W/87a5NUpyayS
HmzhwUWvmNVlQXXekBQ3J9WxFUs9RNHZsjVrIWfnoNXI86nSDczoWFL8xIlECUsR
IWi3EtDycfBp+lDoyKTGEZRQHslKUTBo9avhmrAi9TmRdl5EWsTUdOsuV28GOPwz
bSkcvHUe3dysaeg5rle/dOi0FWbjUIdOGZX0Ahd9jqh1Bohzy8bBz+kdSn/cZgxE
K/eekVSoIfj/eXKSOCjzgFDibOjMRmVVW3jrrETdqMak40KzYI8WaOTBX8lmo8CN
PxM3gLH/sOxQto/hpgpzx2f3S2/1mxsjZMgEDw//nZywCVtgjKYDzcIToi5QKr0p
MuHFVAfYoMrQ+aczj5p6G/Ok0itRaHX8i4kaX2I/Tf9wtThw6DeKKThJjGT/WSq8
JDQaRQEZoHgpi0wBUerJNLK74imq0auqlvQm7Rlfb+lFltIRYQmje0YC+YVaVxnW
VUAHZ+7wNjBSc4Ia8BI8Q2LVv3cuPlZCFxDZuyfwq6b8k3vngREyvcCMuxH+r9gk
GdH9ZOZcX/emTDygOyWTpCpdrFI4eMuPsq497K5nh+g+3yjTrmuQ8lxeYqzSz7tA
oUudEqzO+8bgJ9Vt3fZZ2GoBXCn4Ut8JXbLDz4cso89Ql54NFk8LEWVGYV9pGm/3
ZQknELFg7UeddQ1AjjkUG2HtCDWddCPKu95H5AwWHnnk8GPMYBKvky3rehWbgK2g
zA8Y8a5qzCpf2v8Al0cTnauQUIkZMqqm9vmkscdx5jjq3T6i/4Epwex39khXpJzX
QhxhyLIEMyqorED2Vd9XqZvZCjYMryDMVUXi0XFJwOBsnchTPdeIc0SPHd2UTzJ7
UcPmwCWajeIXGNLiIdCucWuSyLozo6Gv/H1Bn98a+hw1k1dQeX60WJ2/dGY3alnk
QrONbo9bVELGzI6MwDao4zuvWX+tFtmSyMtUJ6pG+0gCxwq/PVVomoObZrP5RDic
kBZTmRaB2fk/3vaAH6nH4gj6hgmMRd6zMSg3fjcQyS5dpvClnt726CNq5Mg+DQHY
uLzWtHFDCYrO1iIVsUdICEn++6oG3nsHOO8BK64YXhBI2d3ioc22s7plgWIE+9Vq
3rdPCGWdsntzA5qm1cP44ZelnbF0ZIkiV6oWHV03Wv4C876w42lWFURvNbP41tNu
HXIZnRN662A7s7uxLD9yyuYWr1+Seq3KgJetq364yjxrCvISDinE/E0SI8oEew7O
Ar/n8MnK2+TnspDKZLD8OQ6ky2lpphDCSj4axYwsEBZRuU7FqCdIyzShvN8FaE0X
OGHnZ5stwm8SeOC1eXtmQws8+J5cbpc+yVDJefR2NRaagabGuTzxbaYn576NtxxC
WeF0S0GMWt+UBaPF2P9NWzIUVxe29OJrx1p4GxF2hMcBMvGzHhBNrUDNDpxK0crF
HGueQUwwiMMAX5JLuXDctWPG45B/A0XEAkDZHehZoVqd0U3avejkK8c68TkqDTw9
gbO6wLFN1NwUNXKFxBHKzlTuE1rpknTpHd55a0JRKorIjdYw76Bcixq3bFhKZ4ji
e1mTmaR4XmEIjkW0KTJA5/SFkZcDZIx5Loa5mpC8wV88FBtcNY1qtOanB06O7ghV
ZWWX0xqiH8t42D/ocTvU9j9OfyjzFWRz03CnFrv4tOFvsHxkZeAO6eQlB2t2WXvW
N2DnCPsihEapngAwcMjY2XzPNTOjzCxLFNomzBCyOuS3DD1bxcI/ybdO3itqmXYA
CsXg/6bG+LW63eZ/kn4lDp/5cemk2nDPhmWs1MoHhRFQOodl56H5jFi6ELinhrZV
yum+P6eXt1B0rC9WXXzMKkTdIyx9CqG3W1eueBdtXjtDk+gBNGljmfTAV4fcvtGk
ODFjcyyC5nLSFEPdQbs+0Cp/fqNnO+5w2lrMicSM8K3FhapYtLE19iLINMPq4MRP
d+/nsdtWADFDF1HJu2e0sPDLeQb6LfeBgpxJiUl1YuDy3RWaTXKdTt1coEU5HGQj
nlGu0ZroXEuLDSshN9/mJDVqCxmUXSsrw+hhofJQWoF2b+JG1I/RmzzcptJQrohd
cloazpOd4dg4s530l4YTimjBETPaYHZ8vfCr3wbJBXuBS+dzuSxvFHnw+T6e7zDD
UBueuSTgiNdKH69CAHyiLSq/J2/y4AKTzFr4Ickg45jM3GXTUnAuXicjRR7VqgeW
xlXp4BtRqL0IxDr5DhmQBCQTZtwDVzJDzIMU5ZMLNFY+bMk3DKQ3Kw2YKdzs2Rmn
w14g8qfOZjnPavk8ZmVXOgzSrhpwuzfz+F2t4fPKI7AIBLWWUPdOWZRYTFKLczqR
+5031/i/eQxPTnjchhTbpDJjHIQ8sGrDufcWa+kTS/03lw7TSJjnO5epQa2xYXRP
jEisiFpbw7AVmlyEpiHXTM2J9mOh9bT9tghnAJ/XkJwLXw0ZLu5479kwUv7SiBHi
h1dXGZuquqvddYbfITb8nm8QqfjmS1PlJSwqptN2U6+KR5MENSsgZQ6k4wZtiXcJ
aIJ8NggQ95RdZIu5LlKenrP4651sSWDv1r2qyN7UqnRxfZfbp5KcGm7MTT7xoI3j
N4jw4a0cgqJQguVr+7jWIXr8UB5gQcsjvTuV3rZdNLcObfZmUKRsYLcGmDglMLmW
umlvhDrHsZQoPf+OdEAhwvuVSJlQ5yXHulJLIM1zPn06DQmkDg9d5w773m0m4Xiy
IQS4zZdlK4GCL1VW9uTZl1Ld20j9/MBiw3i4bXks17rs7bAtODnoF2Yf1BaZPVqc
JT5EhfFh8Vn/ade+TRBQNTF1T28D0gMk6Hp+O81bl1rwvwqAjKo7w0TiWNbsWHHW
WRJHdBUiQRFeLc1qPGenyhjK7AjxEtqUWcZ1ayMGs4WU7d8R49tVxj/efsNGFOzX
pnl/Nlw6Glh08nAKvOS39HFbBXgrMppp+G/ZvUD9WrX4BgNm3NLxxpub6ZmfkhGi
WiXuc0poJDg3WUF4wtR13ErYvfd2lDMyRkx8SXJ6Qmg/i0t6ZU/RCx+kh1CzV1gZ
KezIbsehygQSoVpDVzHkMcGanTzeXYt0Hd2GvYiaL6Rg/FTC51WSb1QVJ+TevXp4
bEgIa3biR33DCQvHz07PuWNVUYcATRjmSKY6jLE4x1zex+ZK3QnDAfxpJOhfs9Hw
6mcI92GtFkFWKiVP6xKkrqS8Cj3HVH5ReRZ1uiYa5cSE/proCyWklVL3jLIzQfQ0
uD4cJ960MlBrDlOkpHEia22x1pRDeVO+YHlmQYvj/z0U8so+5HRHH/Qd6EgNFyNE
hZEz5N/WKOmhiIQVx5Yd6WEShe25ow2VhYZ7zcQzYaSWwP42JhZq2oUehN9zQkqj
4PdTLpujt891rLD7MsCfCBPOeFuoDSDvP5E7VhHLbF/eteMkwbe7chpewFueI4Nq
iOPG/60owsJOssDc9QhyyFaAEOVX86bFa6dp44HETUsSRAuphLK7gI76o5YhkFkI
eCTwy2sZA32YoX/PujN7xD9Lt1VzYw6nuXS3H22Iqb8Kc3QQyWfjKqzqft17BFCo
xkPHhvWAOLl9eCnuL7QmLf4HzSBwo/0zNfuSUhXYhFs3PIZcsLitVK8izY4ELAql
BAiu3utsq7T7lFbzHoSy4Sl+JGjZovDkcD+PwT+IN/gAB/GPn07igdijiy5jYrgx
a2+sVr6+pi12f48zqlbhVIBhHo6zZ0+CtqhURDwhUmIU1TxEzmR6xVyKOesTI5DJ
BT07bfg3baUP8EvGCrim31vLJtwXIPD4l4gjs8F3kA7cCJd9bvDd95IWuG2tnYoG
+J2eyBfpixwPoRWSonwd14mOpU7I7UGqoPAUiQh5ujvs4svt9xTlhZB5MK3OcBwb
jDzB/4yrzBoSa/rXskJ9FSHkYqr0JKZeY/ZlDPpuyGR68nXRj0mkZdBZtZNV52Of
9qii1MuZLFaLSU+uRY8kYglDYCmnozIHQ/syeTaZGdHnBtRRMUCIOCluNQUZNb5l
DUndhFONdEOwQmjn3RD8wze1GZhR19TsDLjR6ad7t5VHDA+Co9HXTMqN6yzPHewH
9Aoovm0W8uvIrE1nRh/5CYsqI9sgcha3D96uPTTdGOfHskxy9qobuRKAzRYTTq2M
7GKQcGEDN9yRDNuxdjapLZ9bSnvw6AUpVFmxsBIHftfM3FG1GGG0c5Rhhe3Ujrew
N3H4BtQuw/e3DfGFj03WPPBDniXYRXSO54sFyyvRwvpvorkYhGOIGz6cBrQ2fg3g
WX0Hq1ZlCLN06shjXml4s9k4eOjBy4/CjEFVhrEKSN2QQ/l01wGWdWSHJswZpImu
UmuOOA70wUeE08unHCr9HjN8YgIpOu0FYJIMy7n21dWMo1P8m2iBTH2SZPAKn5yF
zumqZqb/URv2mdhccYWe8/48I72nnjdzTGFYPrFi1YCe89MH3aaZgoFooe2z1j2i
5EVY3uzwlE9cf0rYyvo1Ikz24VetGvCuTDBrJ66xQpn3c9qZ6eJl2wIJNdSmw8dq
kPD0f8DUFKC5N2i4qdxe/76BOIzaU/mvSxblsC9aZIf292vzLqi+pU5j798+W/Qh
uT4rY0paju2POTqhNoi3umk6kfRMbmYiKEnYtG4AZBUT6iqcSD7iJ/nP9zqgJ+5w
fpi5QdkHd1Jj6MPTw4UVerFyK+y85CYaHV86FkuSKogxk0KCcxto7WySQmXVdQZb
vJTYUFJZdRAAyx+CAHD2JeuwPvXrOzdGxThyAYU5TzOS5SNJt/um9Q7cmWk9vRXz
YgQJ+hvcJPWWDrs5KByUVisqM+T6JHx6gV6Jd0L+DFixp0tLvy2oHN77Jeh8QIHa
sqvoqLPlhZWS7LTHsUH+/17PNMwkbgEoU7bP2mBW7yxpzZdk6ecOVcCYfbICaeMH
02bL4cv+z3CYrUOacQew1xy9XCVDME6hI4G//nfTFHhQEw9vvnLrydYotyrYBeo8
as1yME2kpWlk0tByCdRWCZhytztVlA35jOG4d6OoUIlDt2hmvcldzlezzrpOWjYu
K8/Wrb+yRx0uYfw29pdfDKmn0iM3of01ii8Kpj3TXViNF1tqFC16sd9pl+LmjH+2
1JpZZQeo2FbVcVTcr7FcFzRYeRy+EpCgKsv3yO8PvU6fjnycUQbw6nTm+gi+psBo
sNnkWX5CoKthqQmZ1JBcZhJJcUfWIkIUAUdCBSYO4BvU/MOwsJraXCt0o/6GBiSj
0K8sVEnP16BskN8s3CIXp92Eh6YPdEEJ+6UdkVfeo/Mvh8GP64EZatfeD/92MiO9
2djhRMaX8Xj3EpBggDFyHiJJ5IlZcIVCyOSCygTy83b0VCPei4zLoiga3PBVCas5
SN5NDOZxqi7rvH9zHttVz+hW7Ql8xY0c2laoSDLxC/L0scdXcVRhY5dYK1m8AoOG
a1+k7nQqBcFpue+KF2fEkvFUhurF9GBvqDhCQimviUutB692kIRMPYhuk3hlXf6x
8xDDdFH2dwANlvALm7THxd5hBNiibumZFF9ai9cgy8CcjPNxDEsCVjg08ghbkaz8
zj5PcTbf+p7Aa1HztuJlgqP3l5qwb3g6GvRrhOJaVWa6ZY91DUaPVitdCFHwKO71
OGrgjsPxl9pxW7quy/LCDjzeipJDqaOnUZXg43QGnCSSWJfeHuPD3Lg9wsp52W/i
bH5LEhA128L+zB2eLmfOmWHOP+6EwUmV1Nxf9GaIfgs6K8G3bVizaH2n2rS8i2pO
C0GxVBuzhqYk3svZ3gnWfl526cqAjsdlrJJzj6yfuq06as+Emj1YjuCxH1tUEYXz
PLg34TYs58hEuqM4/I5kVFCx6p3wo2OIbg63pPoDCpFjzs+97D6RAb24/Y1zhCoy
8t6XNneus/+nXyArXHic95/2s7lKOy5gUqyHYAjfw+gyS80JbCmpoNhM4LjOYJQy
WHLKuS5CRtKAsW1oZQx9YMMWk3b8c1euD5cwoTb9v36c92xovoMCfGcfDHbA3pQp
KDO/EzBvibKMpopCpAndxKinTy6NadJ3BUrjwShUGt252csHRQorgtUZVdHe32tb
DINOScPZ+Z/d+HdqT9fp5s94iE7KKRSTAC/Oo5ZiilKuVbcJqkm05epf+6gB2v8X
sVTZLaSwy5n354PfmdBawTMM+/t6Tq+giSWfCU51zKiQ7owlOHNXvfXcjSgNKfgP
j2YJlW+bDdtL+auQdjOvGQV9fhqk9+JZqH3Fq0Pfyjldy9L9KMVKxTgmErtIAHEQ
BfS6iZVtYD11tmW/uXnHU8xqnqleyUalPPljW39rRP76qkV9fn5sL0lrt3I4IYs+
brugwWi7Yw2t9PFKO6a5wYrNxsKAPhgRWERFReW0JWKXWhBqhcYJ/Eo+SfvWXe35
g4BkLKIenZ9N7Dy32fm+y+3tAYuDcOAHZDAEz5w0nbAoZTh/6JBP0o5q+WuLKewX
BIvDkRuPdY3TK1Ej83k4kofqA3FsblPD0fpXwf0t7MqOBcxY3UkkJK4J1/2BHcFN
68QSYYrYKeNjZDnQc4rv/roQuLBbY/5kM1KB+b/KGCEqiamV0RdC+sAdcyaKQkNg
/1WqSBoewlpPJ2Dv/XdguOZGYztlLAGgzGHempH81nQOpo1xTSY08MCRhk7WMKPU
7TQg/6Ntrtcvxp6YDkLYUTMNQF99b2Srse+DMog6xaV6HgeFHkmPdCerFql/ISGN
s9DQ4gwaJo+y3OYAE4FFlErI87kdwzczJn9VuRzuekJPgjk+WImW/apnGNWEmZIi
YwGtaPrAtv8K7tMj95XcAvWLnvB5E9QcuCgN62lp8qo4dZn1+QiFdzA7fbyISnmI
PSgdrtxpFzHIEFlx52kojfmQtdSJWSLKtOpkO8Eyo3FE+XkM+lp0Vt9h7kMYeqMt
IbOlXmKwvQmmjEo/cjFTc/Ee6CDYlOz0OogcMp6JxhrZRl97deghNcFjrSRDvJQR
EoCVKqVd06/pxbpMGnRX3GrGidbsopAKq8z2cvK5IGf4BiC5tL74jrpruiUl/4ux
J+8shVkkkLoSfxZUljhZUdRwv5NI9YoXVLvx1CLlg+5liOX6oNWXiw5OTmFxE2gj
89A5hgiAv0wMfC5j+G/Yx3cGJdBSdlSntDjZBfYx+7Ja7eo3WOwlOf1hy7kL/ZlL
zVTFgOQu6RE/l6oqQFicteW1p7xeVRnTNjFBtW/EY1aGtC+E2sIQyXr6nnntrny7
cY6Bn52p3cJBabcjz7CZGykcBQTYMX36TEIFZYxqcU5Lcau5Bx4A96t/dSp2OlM9
Djz4wNF3VcEMQgVXjaNFAFY8yU9LxkSsq7izGdejCUsllUzXiSMJYGJs//cZxVdg
W/x7Vd0INiMCo7A3L3zHI7b233gSm3DP8noB1L8ojlJtEbghO7RRuNbA/JbM8Y6h
kOTRrNtWq5Ajxf2SNOkTxQGejhj5SaRG/fsmOsiiZIV6j3Y1mBbJqKSbY6xWiGgX
l1Umz0DNMdDdw8ffeKefE7eE7Wtd3rmnqHJBSrupA8w0SzTrlQdAGYPAWQVpkNOa
Uuc+TDhl/uf4KG9bbVRRownrsPoXsYeh7AhVKRvR8Z7GoF9VY1QNFn/BYgdnms1w
j+TVRjXPD0zd5TK/ZE3d8+lEwVXrkA6D9mRP7hRaSH7ym249AengHuX130bNztwr
zhi4fCXUGyyXxTiRIs8TS97nHQSILpwCHyV6IhhcXPzWa7f7Oys0dfVXexluIzgp
yNyvI4UxFhOaw27Pd4+ByMLkWm40QMnY23J3eqYrKwFLbatEyefLKQAEfbb7to01
+9WWFOQnezY62MUDK90Sad9aWaI1COXYvrib2uYvxil99TkCAzZ6JWlmFljraAOR
CdunQZzbYrDiWctNXcJ0hvMsJM+nM/JFYPhxcSv5690l05vQxWX2dW+DJabExcha
IVEBr8m+Yml+P25ynXX0RKgqh79kCJoknO/RZUVnCiP2eXSWlyceJaz8IGvkzrql
Bq0q6IKTapPkFdugBiy2t3Mx5xJaGzoKRe77fYhBDFzUhv0muBehosYYq8Jkm5pL
+s4CwkpJtHRIMftVGWYYk1XLZCQ4swGXK/+sgenlgmoa8aXy6zvxl6UTxvU/swF5
0DRkOCFANzyeEthVT6FIJEtA0W0kD3gWSqLtjXdFT5ewABy0TI8OHQO5c4NWzYlR
BxQT8LMo0sxhZ6Rr0LqWfhslbnZw2hARwwzifRkgQDX+ALz0Bi09NJZ2wUD+YBPy
9oNOUNsd4Cb2GEB1eMEs6PQ/qiX4nzrL5ReG5ld2dAu28CGdFvqjrbgVaMIpmmPW
Tb7gsKdUms0omoTBYtve4tacrIgfKEHJE4Tn/ZYc5IBXGiGs9dNB6pzG5SV+rtnI
iXIdRerBOeuKeAber7fgLvzqvPfW6JzmCjU/Sr+/3BUz4ou4iPH/wVrWD5HSSSEx
eB/xvFYm3QdDNJQheqYlkyNiCpgk7yD1sH0JkUPEaF1t6AaKMjVip8dnnzdq8H1V
52WdIzKZCfjSbtfqQ/vS/dclVi1nklFhZ7DhC+QdDLxObqjXTrcOYvhHlthloqDO
xrB1Yxw8obS0+v57Lqw2tMx20Ng28Yzars2CAJL5veGkwHnJC5bHT10FpD4Yj3yk
YEX/ewXf7D9w9L3oCIhxq9XRg8jS7Xd4GkWA3VxJexYW84WYJ6AZYTwsVHLuNJhZ
1zJAQoOwSH0RShtJ6ehz09dgDb+C19WCYRmWx2Lb9fGCbH6QUjmq4lERSLowU+9D
1me4jxct6ZEhPO8jziikpQdx2HF7ozpWsezvq/MZMdtcwCzAHlOhJ01fOehSgGDl
JfbqaWlH6/uZVCXDvJjjDgROd6RHg/DT7OmFb8UpPxhczrggF7uWfsRj+GthanPC
CtA/POfejMs6yStDcSUaaRvXx65jOBIEAvnpbR/RFYOl2AcefJobrGmwUPl/AGNz
BVUPn5yLoiXoIRRKT/3e+BIVgxTfG7bLzW21He7Ue73L6j73uPjjXRM1/zyiMdfM
C6f8b0eGyE4WVYnIEE5GyHcpFK4THRBdSnQxgJE81AwEB87NpzwkSWtKqieyLs6o
3X8XpbCBHhdpZED2qdYVtEbWV9zn+udq7NeJmsbiZQVknKOzEf93QAvYMtolVnNc
gAg1PNk+h/X1mS5junsK8sKZyl1x1j9siie1qFrdUoPvRXyDjhaZQYbr69A9GmQF
uKRwVjKkh1o9aDFFQwcsMTuoDikLCwvOlMrMjVRfvTkOf26RxZI7boEIPonoqPkI
6UIoaoMDXGhg5BP3HfBHckIXlfQqJCpRIq/VjwKky8GP9DRWEygRngF9i7OvG8Df
zQIZXiCupCYYVk4lqPfCwOql82ao4eo/Xatemquwjs7hFZohUZve8fwFCqteU2+a
fjTYzFuqWX6eiNLgTD6yfIp046aELkLhWgd5na0wbuVIvqW8GvV12seDAEjJKIrR
mAI/yMpuP83XiwobCLsE0ultaqwJKUCEv+9kBEv2P0Fv9VbMA/7Vt7M442HHVNS1
AjT4SqMF6Pf+3mGP/6oS6074PfiGoMFJP1nR6sTBgl6L5KpWK5E2TgNle41gn2yb
ZtW/K1/zd6Nu9Zy5I0dRgAaIixwLlch8f7ejm8WD+ERnJntwYR461mHj2kEcbeG7
L4m+RYBJXBDtTqqVFy/slvk3pcEMYhaz9B/oJvFk7hy/lCkvoDCjWKAA0kQYWvCB
OkWZnsnqk4Ll0UYxgPZ3oc8o7sHzL3SYhoQxvXdtbk4ZHUDjw5vCE2ZFHkaD5J6+
9eL6J3/SI7Q3EEXlD2PDLFvuQaWe4UCvjmYyiU5Rm20Z+1mCPyM1pfYhIVrE/52e
ZI4skqiJUCGi4FRAVeSdF+YxooR7f4MJSIM7LeMN/vSbmmhZDqu5xgMAYMfP5gmI
KSxJkMt+JCDpKQAStevY4flJPEg3euDlqCmgw5Bzb1GELLDwPLyP4XM+p3tVBIq8
2QZYr/gE4y9ZF0cVaCL9v2Hq7o7orAr7CxQUMuT0cvlnL58xAm+rvciOKmQjJz0X
l34p6dgsw0e+gQBAr7rcq4DND8s4MvSd0v3n5ptKmejECq4vxVns9FaeJUbeoJP9
AahwvbAxEv3J8QP25+8ZvDMvrZT9QFrckCGGIntmWdjGlI2L59U8YUnVgU5RGrqn
8mpVr62mAH9MeQDl6UY7eOmr6NFaz0WSlQAwpjgPVaKpsXFdU1uJFZOdqQ6LkG4I
i7BaB2ZEWSPsjv2ggosNct7X6grwIHFS9lO2RUGBqSmzF7Fy3D+RmVAeC08w/SpE
pa1Nzv8ec/B0s2e22syzOT/sdaoBF9NcIJIRaTrR9MQcyJb5Z1OqzcDG5SkBvXWA
oJvlu+1JzajYuowFmIQ3bfU7uckCfZzw4u+Xr1wRGJUiInW6aoyB+6eOLyZ72i3t
zMVjt7KDpln1ULMWMAJecEp6xedUGCWta52JGJbRfHSGEjCmxVx5wVptgnmAJvoB
XSICnMuZxjMs7IGKu7PVzBkOSZaMduS8KLPSAuq5KAYV9qXcSDm2+8Ug4fsFnL4o
aCp/HSoBOorcgrnk1knNkKByJ6Fhk7TC6I1fkPm1/NJqYIrjF84hvenceD/VTJ8M
PXi/T6Ii2omPjMW2pvahFXmfPaFZ97LHNtT7rWHqO4AeWnOxISV7+wFrPZ1raG5Z
VP+Jd42z027928M7I/YB5/h7+kggC8PsN27/HPo3YrdtZWvRZuTiBRAePT5it2+L
aWhC8vlTyJAI6bQtORgrEJEgn7qjWKkelA+Yhta5p27fYsBTsvuyWN2vU4Ip08Lz
UBXnEo9j8xeUzohFHsoY663OPs1J3W0xJ0+9qhc1HeOG8yTao/R06azA8GumhVLw
zTltAgUdvNN3/G6Pl67wun7XH4SUaO55UdqRi4nK1Qau2HVfzPzpkD32v5p5Cb3z
2bmJwN97GX+Ptj+9z//nk06zdH4YZFvMtGwhkDTb+DjJ+iNZEnYIuOqb7oZjl6rd
R0D0WPbJdO47CVYNVZVHy5jekzZLE1euwmmpYABPa99b2VyMMBdvD3PXvu7nZp/A
Oowk2skNBI5QEhTVjmZi5YS84ifpVSviQPdBWioi5h9iaPfDeiEY5Y7Rmas41VJP
AZuc0TJ81lob/4LD7FU9I3kqn/ibfZcBQHKHZtvA0aONRDes4W0VLCgz4d1es2Wj
Vjj+7+Ri2t1CqrrJBMZvZqR07jN55NFCYZkIKjR3a5Y1TwsRP0lteSwynUsZbyK0
118hRO+4llyhbuCP8+Y6yqNuFBRJMv7kx8eUFn50r/zeQNGMdJlI+xLeF63O+aKu
wwpuTPrvduJp+fKGeFFZyahSBhrhwnArfByERQaoklG7F1F2v/v+iyGRxtlzTHKm
9ieJo+DHjnmC9ztbkuP90ro/vp3cxYh11ZwFiWUQjULkvJXNBR3vUHnA6CEB2BBv
VBEmdYwUtsoGer8pNtVvfxvJuhOCkFFnzfCs/OUTFIC9UEUcBoMkn1Xm9GUkxICf
ZlGTodLfW054J/JoXp0RuDNy6eoJYkUY82NMGVGIgnNVjSWiqm+vUSrQhMuEL/sn
yJjXfnYbBbvEIXxVzT8tv/RglAyFBSto0dkpLSvHR7Bt36d3a6/qTKUJVinndAGr
eyFeoHCsNkIqDY6Z07FtMS96p/lk3jcP3TUEBQ5K7d9tQQIs4o6lKU3AMcu/cT7e
2bqjRwyxYSW6gNtwv4NBp92HAxNJri0UP3nPIgVF1+OI5ZUez+7DRNGptWOQZ561
FzMe70beOAo9vZIVBl3FGZj01aB8oQRdE3cCsOz+65oKYHphzG8vRWJkoRnzAYV0
aEUZOf+4xWZxqBv9PTXijqs10dYDTxqnRF5zJUbGU4J8RdqtV1EFOfjY6gsgOt3V
W/pBWqQTROy9z9spuHDOjJz6wsv+/UXkQ9KsJIDgBSluLyhVxGiJFT640RD7AeoB
fsWgT4B5MmKRn30Zwv3htk8gAYZpRaebJy7XNiqXQIA+18ktNz6a6pM/4SHAdH6v
Og/aR9lYrkmCKtkjqzaUYUM+OZXVUl98ANXOi3fk3AAtHkv22ahmPzkyxFceWoOA
kBomZtGjxz0WzaBuSzIphvvj7aafSlRIT8+9AdL53DfLixEPD5A4MhTlV7DM8lZx
us8ikqmK/5jm4oKXz+9SJTh8NYZ+B3cdv/dDbjYBRf/lL1TQq2LT3Z8w6vdOdCey
o1Hm+63Ui5wi37kW8yz+D8gcatxca2No71r+mzTnqRNaYitxHZrYBp1jLRXxo1V+
xNGO5/pljPti2EB15cdEl1fCuKss8i5Icov5a06/ClfilAQTmEco/deyLnM8OSme
YnbtsfNMl7HMgC/NTKaxZ0uFVWp0gnKmkEjTx3FFezhb+5EP54Vkik9IMyWF5AaE
+kIflV6cUhx3F2ulgKsubPHGs7NV7y05f/DKlIemwW1zSQWi7lVQEl5s6ZXeyfYH
7xfZFx4WyjIwqB89cLvLsY4n9q8FsL8XNBHhj9qwYJw3EmHvw8TQEEiq5qAZ81Ir
8uJoGA8i2OFdF2DMJwG/EmTtIQxfFNqC0a5Ges+pTvAwZAcbABBM7fB7xkVkIv9V
bA51chFJwJvY76SAnA/RAeaeYIH0QDiBj3e/SOhDgvAVgDMDjdjXIPl7XL1T+D8z
I4rtcV9EoTXqP9R29xB1V92cAc3k9QEIoA4DGhyrXfPw/1LbNLLkeyzw0I65Y9sk
esWRprdx1QfhFrUf1L7txcPa03X6xKCfT12lVnhILrueam4rQDgUXtliW5zQWKl1
jeGvJ9LJrvNTHEIUg+EkgUAncmIjmEyd+b9aRU6t7SL/4xjXX6bmAPAA2PtazWTa
N6ZeyfKyK7IgdcWZgC/fvJAHu01bBC21hi4hge8kwFMu7nAZoyW9xeEnQVLhmcNG
D7dSTmCHZCswwE/fgHV+KzLWanG0hkeYG4xRs/rgMAl8EtzIz2LL4r9IgV/byzsX
/LaXoBLcf5WlC/DmxtZfzauHguOSRFl5BRGVOyIRgstY1h57m1AS5vqDqtTLtrd6
uguqzVOHWVtS4aVMBsYu2shbBAU51AVYRcneGt42FTPKMzGQRtFcRLX+1+Rt9hns
xuDut1XOHIPQlrSxILq7wcmVECIBm/KBdNl8YbUPvW+LVBD4h5Z7+2lO7HoCHpm/
8vYPS2xsmCDiAmRH2CGAgN9+Kn/T/NUG2/9zuJEFfVzJiY30ULQHgS/8Jp82I9Wo
3dr7EPZpQihWE/Yr0Y7kWzEUJ9OPetKD63/ViGCURwIWHq6Jv+MiCZfLQ3YEJIpp
gZv0XFMtsCruOMwJ7UR0KjLAlc2DuQ9VM9NfMx3i6SktVwEHVYPZJJb6K/UuhdCl
95ZyxkHVckfYFiE0RORZ9Uv+Gx+HTX9GvVtM3Ljx9ih54VsCecWB9X7/15mPEaYT
reifD0B0NgcTxpT1q/VovjyU5KvhX/nm6vY04MAsLLS6RerqP4EGSZMJycuO5p2+
rs0v/6Lb4WzQa2tPbzoLzdXjTVCbPrvynI8CQQUUm3vZUJ4xpEv/pToZCsK0Ew97
NT5q0iRNazreWBNe+FztSfw0fthpwTsYWA8SiOnbnS+NwcSCRoBQOyiquRVSQCn7
9KnnqaGSJgMYrj0GaE14j6o1jxVGXxiWigBoT4dHtqggfBm9TCbiIECjN/iK6WUG
GsRbxwsVJdYvwnf3HtXPEBkL93G2u+//PWhZWb1WcgS140fG9nHQypFhWVZ2arFf
g1NYT5MMwokIJKa49joo1bqzp0qsZ1UKDkA4q/q4t60WkfZ9FzZIUuh7PZEiMoAA
f3GUrm5z54W81MxiCQFP3noX3Z8DArnZzVkDmwrH19m9Zjlh4hMLeW3jZD2xmkK/
npRMEHGkX5ujg3Et5B1ex1uD1OgZm4CDQgnVSGhNBYvZboUSWgz5aiHjJryQ2R+M
7SC7uANPn2s/wQLFX9WdsT4OOOAKYH9cKB3WLcjD9hjS6G+7KYk7Akgvd4qmFFIS
Ia2jQT8G5OP280xdQcS10hh4mXlbQnZpHAJPpKe/KELGnEBBzAKULJ12LNymufiK
CTnzEjtQos0WI3qxLmQA+XnWRaIEAI/An5DxmdCRO/6Lh/HzgF7lGsyHy7cUkiiS
bGutvCTDiYix0UzxGqX71eizILu0yDVmSj0HlE/9ZxPVEPdnk97G01THUMJ8T0RC
eRt2w3m+VMSTttW5pNdJgjUx7hngGD9ZWmld01oSwD95DnCmyt50nX8C0e/tMQnR
mxMX47EZlZASbqZi5sGQirjQ/zZ2kfgD1QKBvqk1O90b+R5z6/uRMIUASkD0U115
rErER2z73o9zc08eR8cRdX2Rc/LClmfkNBSE8skCZ+pZae8eBrXV5U/vr67hTquG
CB6iX4QRkFsn6/kOg71mWabjrY/c4KtIryE1vxMm6vQuCB5TeyAHjojUP3JYK8SD
luFXeBlqtkPhSfi75Ecr6hTXEM1Alf1QJiAjS5MBOvF4eF/iEcl36uRv+4fcgP1+
GuV3J84zOOdu3HqS0AYCooGV0UQHUOWS85WQlddG1iPy0QzA+wL63F1uOooLfB8W
Ay3ksnlq2Xp+3QeN3OBu9J7LOS0Yun6XcvD7A6QCdyM/TB4FS5b1u2NBetuYSzCZ
Lxm8veqlxW9q49QGf/1C2DnsnrDMTmxyGLHxTP1e58g5y6WDSCKZjBckwjmPR9VA
53nOfN0nlxBdvowPxWwlCfg5OKVpSZJfYjldtewMeWgbfjRBRlGZBIwwjz5eTBQ6
anNnI6TG6bngE6Gq++5wHp2HUYlNR6Df5uFeEALDOzr5rwwehECTig05qeJrAUY0
yvJUef/7PsLS7h41KWc0juOV0fl4MEH59U6kqeb/DoRCOdhnFrXDTRiEZJAPI7eO
sB+GpsztHrqqzjAY5FgkXSuMNN11yJmhjANJ5dHK2qq5ZBYmc2Hi5CB31dJfcCej
CZISKcXMOQaY3qNKwsbeGalYVTdUaVbo36xJBq4CpG+otMAgW3xZnlB0l2mx4JYU
lnEACaNI/IqN7xA31NuFnPjo2EGwn9D2DR8hiQwWZ+aK23VSF+r4+eozSsVcmS9F
nd/sJkCJc46UEvg37f3EBUtESqlJGaFlmQr0xAFS+zEuTswmBITH+nprgi/E1kQi
RmLQBmgCMKYfZadZRBT2tcFD2PnThpmMoqF+d8i/CifLE2O7W22js0yKekVly7Xp
EBstVGF2B4DSiiTAji8MaU+VrW1EgiYOxZqU4dG4QH1tq/xRox3GxLE3rI6aU6V6
fkSujvt7RXMgI6FW1y4nWCfBK+XhSHGPAuYTHV7WVs4/q/5XPeh/A65I/zuEfqJO
yq8bwsPfzDSdXToUS33wqhjvtWvgpeFlENE2SF2orTKL+/XfRdU4RGmcpLWY2I2h
SEd6bD+ylmvcSeO3B8tlQDr5ycXP9s0Ed1/KsS7zsRF5IpvF9r5+RL6NLaVgR7WX
7qRjcvsqpaybuoYP5M5c3f24WdAWK2V63SKoOzhesro2b2cAQC0Jf6z8jhjyOIG8
wovMfo1kXBj/pTojg/sMv7NwFX8oCXJ+iVCnCXmWV2Jw23Kqoql/MWk7k0iAcmOS
obqtuh382tXo8w0X8E7/mtv2JRUg0Y3SG9ECUn358Sdw66qR48yYQUcJj4EyMG4W
9BfYrVNj/iArtYms57NOPyO+OcpnPOdkHdZ97qVf9tna6EVlz3NajzA49eIMkt3K
vdNFpPLdAGrse3PE5+/29QQ0XVhIJJcnML65etZ+dajFlg4p+QWmvd2eM0HgoSJR
2hVF48UBUU65QoYqwrwaDr0hYT54SAYq2Iu7q6dJg5xifxYx3x4veg7APVlhNyB0
ybB9zxojxfAPYv/XDeQAUu+k3N39SHrqCTy42+lcvw9ORh3k7dJeESItsdcneUW0
Vc+rVDjlQ8NpWuJaAeEpmr7Aovx7LkZSDOvcSzg0ePbIxQIg14avPruuL30OYAxV
KIazMCXjVzwExRW/ozM/9t4XBoZHjg4LjbxQdW7P+IS0Ferr3ZL865QkcoF/tSwn
vQAz2wD03l12ktVNoGcVo2lBROiehNFLCzjP2lW+cXrWT1W6PGWWuUZJuGPKpTDL
W5ZBBxVKHsHHNDwehMBbe3Q7H3FIK2yNaDoAc9/JpsfZZxAJOjY5aJiCtKaOEVBv
KTwtncAUji0guisgGqT5bnmBS6UpqmkcWkCv7wctcTeZHsCsgNFFAmlPNzuB2mfd
WrSIe/I2bsIGTLj1wnRJeypMsFQ2PaLaLLYTJKIZraDFYNgIlcjU+bKXHsabb3P4
PwyjYQlqmwbX1yFlWAyi6jzvxb6dX08fAaoKhG/oe2InsWfMrnFz7n3sWKgkYIRv
TVRK3SpKAHM7j4a6OuD/g6A21RauTocznQBY6bwqjp+gi25GysUgaeLH0mcCyxEp
j+xo5U6IBts7hgzpp5V8TANPJ8qmIgZije0Nqk+70NQAtMtHGC0GSSKrLEpVpNen
YJzZLf+tiZsKTNtQQJtjVwtcPt1SwQ2jWyE01Dm3ehXqZO5JDKpXPBR20kCpDKqH
Vqa95SanY99i6pPAM3rCvhk9t1YPjxRGtW7gOUcZQvFuAyxJ8g7/VVCyW48Gp579
EgQra/3KsU8DORSIqmSDtmIyEFiT1Wd5i96d2pfyZLDEOg4LiTJiJ0HTxOh4B1Jy
OMulfnSrvHVwWCCXvNq1mJd3gnYv7rMk1c4V5gZOZfSBjIL1DsGAV7wRmYiy0cMI
V+6qzxbyKsJUq1a3hJF3XMXsFTUEhbp1+Vt50Mq+AOYN5eAQtQes2EJ0KoRWnYjt
HElRYR6ieF00ucomsGI/+ksrG8H0DFBvbEygrltvnyUKIaEDYZYFznAVUuZ61GLi
OeAgkgFjZt/Tw57S4YMCdpaz7voZY9RzhfVyIB2J1LoK9vYJRRNaqbglGodvkMLO
vnurkS8rKNycj8TO4/LzBM6lCmTeqEmcNtOw+ihzx42kFKDs2NZtejziO8vS2VtM
OBzISQS5zhdM5oJZ0lpbHKDkTXmiUpKJ5c+hQPbbVdq20abFXhFKg6iptDc+jhji
eoqCzdeJaJc6PFAA8hJh7ZB+eRyckpNc+eYeX+uirAVvGFZS/SVRomvYRSZjICN8
nEsHpV8aAMrz+yM/iOQY66g4LvNwsqMbuZjt05peST1M88yqhA+rjjMPkXthi/Ev
N568XCIwkqZlhkbnAl4w0ptctrvNSIH34jNQuEWf/3jmJ9B07QpbuoJ2D3qrKRn5
v6JDBXDaTPZDv11/A+Id3Lv8oaWGIwr5GJjzRvtKSAktAad+zlhCkSWsA/uROFRH
fIlm9iT6wskEntEhczZ/tDPA3q33tC/CYj/2f/TRgzlkk4oHv4QL6L4nmdIQ64nw
cHhWAaDk7IjGl39rzxb28OhLN6QizHZv7HWed/n86C4/XaxlWmJhP8PNOFk9351P
7TJQWIvW8hk5rUDGd4juhF5DuVfYn+mHREBy21s+lXNDbcyudcbDxT76exqHrMCS
/TRsANreVp2msukOa7vG9wsxGZtU5UMQig39S/9IEpsrjepWUOniMaBXNKY4VxvH
lG35aS0Gzikb4/zFtyDKEvB21xvB1JsVo1EiYB9N9HSia30+Ofiv0LCzLzgJAOw6
/dAmRfOqtREEaBodxwr6vzNca7umNDpPxxDMU0y5Nq532pXCv7nS0If0xwKdje7y
NvAcfgXgU07eIxqF34LkyQ45HEHSsrWxckDg18TdVUFfdWIyV7257NhXyXBHi6AT
Yok1FQYMMDIQqMOJuCUEqi8sGnYjUTiPdFR2ScIbJiVE5WjfcsxCVgO0/URhPjD7
nhT6plKB1LMemkQqBSBkOi7aHlcL+unqtACI6JkWjMEy9REFxbYoxMbVlrKGip4l
JD4AVEEh1ZzISfiKSgN/UX/KdeR77iJoi3HPaX1BStu/iSXumARxoMFlx6JVySg1
rNZALWF814KQGpkqLruRgGVnvCCsWfUze+ZcTCkVvY3eeNlASEZ1COLFjFyNkZvJ
bcYFnxZbLmguKqG2i9neGrtmI2knjV1m3cDSxa2P6um+TP7n1nLbfQUMTljUxHL7
QfX/YcdHRqFruyxp1qFPMpDSFrnMtvswKJjWseWFU5hph+0FG3cg3ViVcl3J9OT/
MIm0qac+Y3exWJ0Z3P9tIzswC8C9NKKS3Q0TpTyJOzjzhmnRkgUJRhl+eCGoRwe2
JJtaHG1K5vwBHChzUq05oKwuVa80oKCQOSE+35kfmjX+K/kX6qkqVg7DCFxAFkpb
7HmOBC9jxTIehWHMWCc0arwbLZZnoiSU/gt192GNA4bMjCuGyp96St+MsYSimk1+
sSCCNm0QWBTmM8A6ExXQLzftV7DDxmc61apWN/sE6/2YpmUjy0U3Pe8e5ER8943m
b4MV9DIIcp80JqMjNTqBzHZGyp53Px68dRaP+4Y0pmOvUik1DBwfujzDYnhP8LvW
1zoTVrtqQT2WCDTZp1pPKdoZSqAuZvRFNfIgQ5DuXwwPtA2Deg+kgbrZwRrlnlr6
fddLe+O4lhhnnr8GAeed1kyIY+5WaH2vcPig0OS4ASP+QnS/QGLgMgb8q2oDQTFv
Fk3cvW2ryoBGnkr2n0QJYt1xN2u9jwV0ggK1Hmcaf7OtWZYr4pNGkmGOXcOEvbPs
pGeyGgPLs8/KXyTO1wk5T42j+MEvQw3zpszWq9ZCiaMPZJz1SK2ci5m1GCnzwp/I
/U8oMI2sf8BF2tXtju5xq7CFhfxyXkTI0MzEXh4IlnFEAb3tl7Ekx/eFRbcyXFIR
RLfi8U2mkJt2b+y3V9NFO2bjDrd7Mg7hcuuI++QD6vxqkKENDOW2AZ6hHqeEyMIG
2wDoouQcmoFjvEXbnTPGU6lcMHoBUJb9bf6tCJmKyheE0kluo8ohvQ82dBHQgQ2B
g2jSGGm3hdFIIotYBnQqLwJa7a/cdIKFfeGjkZL9dwKA+4hGjiCo/pgPux8QPYvS
aGXrFnvm/ItXDDoeQywZW5A7A+cjQB48a3QCVSXx3AaTHBSX/H0oKL7Ymt17FmeP
5xFmynN5GjtGc3zFs5UHNiBkwGUreMlt7SOYVC0E06iXePw0QLp3Vd3bbaYeC8qR
yVsu6TtDiVCb9pSCg/kpQWZCkdNJ2/JOtL/cRUHbzAFGZ7JjzRZsteDOcZee+Pd1
U2DyfFH8J7OLVCNGS2sGqM8LEr0RWdbFDUCk7w7eRfQLldOB/VvyAdKWkaKRiJnU
KJBUtHKhIzwErluLy45n4DHjN4zjMmpns6z8kSEVljHreR3ZfSiexAlIgln6BxFN
mZ1HADkLPrvhvYLsf2Vkt5YV7oMKLzW5+hXax8uAOeFk7GjdHiix2uJmLMhSr9bz
hfNpeR3LV7+Jjsxk8dx63rWBs6spRqs58KZtknT0GgHysTm8QaL6Yp8kK3e9dRhR
97/y3bN39OwCT85SrlRT8rWekrrZEVNQjAteqGmSEjjtxSVl7u4hF+GRwHoMDjNw
NiFwLS84z5/y49TBrD8ztS1rkivlkiqq37bwMcRIITaurY61F81zgHh2UvFyAalV
5nzxhEgVYIE1eNkCdyHTogwUyMyV5WUrbfNHmgOiiMyxsveE6g4ajzuu3ZXU8eeY
j40P+VBl0Y7q3FlfskKgvqt7vKmiKX251cdIZjkm96EV9sRyWiQVbObJ6oFbJGFK
oeTbJcxM+CSfWm1wAl1/bmBXh5QQMRQpGjlmGOHtFbDsLRiwaYKuxFG3y4EzETNP
LAmpBKvQs11WcV33e/Gff+yiyMScx/xOGnI/AKH45FGrNS9b5uu7oQ9JcgVQf5zE
n0SUk+j06TgMpmYuuKDTkQs56WbweK8uBGUWIfkuu/oXRDzDjFF/0yUR8quzMiRj
VKETeQ9wl+jjEXhPvGKDxCgJCAg2iHHdj2aPWAzZuBffBrPzPujM3uMV1lbOfCM6
sDCWgeZImfMAqNko9Mbmm6NcbT8QWD6hO7ZtIq8DLEKZd7cwAlrlmULZoSRQ+2rt
KeI7tgn8UHCrjHg0KZG5YLFSTl1Xp5OFiuktAaJITztUOeqFtSRdxNXdpK8zyA7j
/w3h3kBUfulbaiUNwduzo0s7g0EDgEJCk4r+PmYgUkvt1E9szfja/QuOgULhnA72
VuPtpnrg9z8fN8lRXI4t8UuCbmewIrvN+XXl4PSoRDb298CK80vHf+4N+mKEEm5X
+ufkAQr45/Kz7PszPOme3Q+q6Xy13V0sfkX68iiE/n3tkqoqKVeC99yZxRwv/BWv
diyL6oVuoix7nEBoVs4EatHbKqUvQNTpWg+cguMnXenFVF1HTfghSytAqTH56XQY
E93Ug8YYr+jxSTzEB8EE1qrXF8jo5cq6PtfT+q6jfjUABDCa5cOmtWG6ArCTVLsq
tbaYIOEqCpgmIsLsT2RRbkinr532YnM4xgL/RYUb8JYbJ9/rBIg748touPwsih5x
NDHJ6W/oHyRzNWxhm2NNpBsxIFbKq9bpmQXab7uQ+gDVfIgfp9omXweINng+jq4X
9dsTsJYOC9tKmlqWailvZvkS1xysB/DIdL9OZswCAvmDqQs1ESAW2zksZoyB/Lqo
8c1L7ybB3x/X4w5e23Sl5i+1V7fnjiCjWsd62jogmkC4GrXt3ZgYBIY53cIGsK1h
zkqztbeOP1/sAq/l1IK6SF9jS38s6NsjQzSEZX+ioYv/moF3H5jW9oYytUE6Ss0p
Kip3FynH/C+ul5RlLHmWI4vzWMl/Ql3528kmGPa4g9Uj950ruRDex/40jNsYfOix
kjgGa8rfNnM/3jRRFgF9iHu88V7BdSlxm01ensM7HzlahlPmvZ2iaQdWTN2FQ/hD
UZK/rKZilwsBkVSYpzr4Bnyuo0L/cFQONfq7lg55bRsNBfq74gXVatW0o8g8Oj+D
qW5scYsK2aRWfUkR0gza9NcsZhX4jH0OrMEBEKfHMp0IHXBY+KiXYAeyXNyH+6bk
acCHI4O8gvsubSiteJFxS59F7jPF9RDoZnXEcxIHYJQ6v7ZjLYb8vxn8SuzQn6mY
htKyde92pXpw+qWhefBceYHEqs48mXqP3U56ALeC1EThDIrZ6g9I6F2ZODQZNM1H
QuTd37VwtY62bOSwtfXXDHzXcRqR03CzhthJcxzUIF+7HBznnXXb1ByihYz9ryGR
t0U/K+VKTYSgPPNhj1U1EN8iU63iIXxeoSg39YVvE3a4+tgi+/a8195O1sIX94KO
/2D/0EgDJrv2K6aaRh1rjpoHIshLFMnw65D7C3KeNv76skYpkN9hVL4RdNAl9jJL
pLJPAMbqFiV2f3BDN819TNY1LDfkzxDp/G9Dxz1+pBEBJgZ1/PpNLSRP+MZLowHp
sHq5BjYRRsW+RJff5xt3XsuPJRVjw0kR0EC9Lo0J2SsyXLjXpXK1h1Y/Z/Q1fXkv
2+bBos1AkgXQ0wMKeJ8Gy+6/u10ubBTMiZYEX48A80ADghPpWz2NBTu49jiNzWE9
5CXUmkCjfmR54/GqETSxVcRk4m/s5DOyqY0dwehMUrm+u0UFKsK9Czxk+9QGmT8p
m/9zl5zvOYI+JR28VtS1VN2RfKDEIptQk0+gbP1dmEpxdySS7o1znPwWkSITnB64
zXL5bDPPM9W7TyTXAzZCynvzAolWhBf01GeJECYv5wa7C+5O7KxoJzZrlwND4dmE
bJwykA8CaQL+KRH64E84cAEI6m2le1gK/obYEmngoMObnHFlacNzOOprG8CGc2ob
xfPSSNNu8e8pZ4ZP9i6uLll8xcEl7vGVbg7YwVe4ff+N/OaJBX/Hk1bSHZZIC0KI
WBC29PmoI4WBLaPSQcM8jAgnKswXmVBjUcddFkU4c+tDx/Zg50nQLtGqqavR/JvM
JaZOxPGFpLNuAZskBhtPWEge1V+Rvd1ADILeHK/jaWpMxq8QEVhWm7zmVA5oAagA
ULFrbt/aex5UPU/Rem1HBTk+bGef3YA4pasIAjDwrPyTzrO2vvYkMyqDGEf8BY97
1xwSPpMi1zgjiE4MVu5bDJOn8+cTwhBpQY/gAxHXK33gE4gCnFbxQZwOvHXbZsEB
E4c+/doUQUzkDhIVNE5qPXat8wpojoNntqwfw0q5/yBkE2bykm9p6UQS4Q1Dl/XT
ryxEsRdZPcaHn1B5TAgkgvGWDEmQ66Vr6j9YGhCgyx5JlIJeT6Rq/Pgc5wglefJX
h9WLsQxOJZIVcfMMbGX0R2OyySrJvRGVF2rtjO/rTjvsSSNf8I2teDeX/KdxYpB5
vf4SbfKRySztUNocjA+FZRFkhx6mObPg2/ca11vieb2Z7IUy9Z3rTXZVFAFb4Bd5
p4W2eyIAq3VmKjlnwYRESgdXGjIoeYe7kNHj0G9G0rl5X1p0eNQVrNJyatX9UVvP
Y0L/kFQur+BklE28HoXIzgwpsxs+NJzZLciVq+TULpdwLagHFYFl2VqKQrZrZrpn
xu80vS+Hj//SyShxZiNqybHPXWRvUIxm6voSaejO8y/F0GOwjHHdOz/QUV0HxdCp
H2Cv1Nsxoq0I/13im4ObGc1pzInr7VH+SRmu/vMH9zSZw4kmIc1s2Uqq5Xg3Hy9t
keKMSJNNnoaUOTpP3L6cVe7tAQs9kotqmR6ZBui0vMzcTTGKJZIouO9be1ILCVG0
+G9y2kJDEsiO96SBZCqgO/faTsRJRxqnDIoL9YTtjzFznEdgQnoJMQLfMJWZ5zus
Y/pVAMmCtO7r0ZbPdPdPXUWvTMXHlSjmM+X0lZv8dwb+0xHRjZnYy+288PEbJok+
/F8BVL3dioVTyWRGQDnDRCLs+5n75COswd/s6CxJVQ+W4dqDUtjMtXfadrgVsa/m
suPi9bop6MCWa80sOdQOaLSiTXjImo1PdB2okyBZCzGfzDYF9QXQN/dcM0Y+NmRl
bEh93++VX30DDrLxs0j9KUHbBxm8M+1CK+o7dzynhPS1PDOM39Xg2L2fwSsd76xU
1qH2u7I9RCjfZhr9kwYdPSehAHnt2JwG57C5/MoJy6WC5Xd5sfzXfbNjOZzuAT9a
keIjGv8yUcGhpsl0HcVRa1kOlIhku3UWmHiwV4fLu2SS3f2B1FBG931P5zmtcQ1z
17nr5SjkuBW5srnmbptqukfEbqn+I0W6ZgWL6vMZO+vnsQ2nr2beuOqXqK199Jql
O7PcwrTHwX15zfG7KkFPo1yW9T/HQp5QKh8woWE5b31iyI08LfLga66CJmSt8DjL
hqDWMYbLaCrQnWP9puSAeuY6I5TkRD4hPTD3T8tEeVpEOXew9069iqnJCT6KA7vq
lp3RngUkKxn3d7ohIbjBCeL+6DuIDan78W4CCUHweHGFoOhZDfqIxRQm5pVbO7E3
6de2HMSFJRKOBuaOIolEociMOz0+yyJSyXh5s0vREe8331N4m8gLBe9OwA9ph7aG
KztxK2McQOgZbuQRnycxABwDZk/BSiNbsTjxJrER//0dw1FmWtLuEmGlpao0Nvkz
oWaTXJGqoAXpMKbNliM1xOc517yoaiICI9ufsiCQ/twuC37B70r2JMSXuGsnv12E
w8oYiyKRWXXYvQPMkY8JcSaKHgeX0ApGxilAY8Jd8dSFUSw3jWetNBR1V4f1SCPa
KDfEByj74Io1gbKtHp8BY9OmQUlUcQ7zQ4Rc3iqwNi+OTJmO+tnd0aKcQMyUA9Ua
Fe5fcJpVBYTDd9zZ4ZzWMzUqvGZbF2bSGpSQhzHEzshGRNtHUR42CtLyLclEIK6L
C6VYsl3btqoDfI+lzkTLTi+DIVKnFtVljyjo8GVbq6aletWzhA7d2+1A9OG5EfJC
Jz+rTCbCMSpMF1XEZV7AG1sVOoiJu7OVh5d5OFBRaRJ7JYjEOfjMnGUrSQHEcP+t
c1F6sCn5kyw15lT6L5RbYlGwxqA7S87n5x4UGEO74ITWfqkXRvixZweHdNvhgYEf
wM2lkP9apvwLL5Eb7X0k3t9y7hWN4mIYMZL0bSx+sHQuH7EwBqm11YSO4Vej313W
8Vzeq5YGFD2GOfIN6BUgm5m330xNAdEhdeQ8kisbSLO0eyYEfTRQmQPdAbeokmGK
iqUHDGNEMEM1az29q3iW+D1zGuttxwkn836YqWDkE9g9w6cBVe4V4h2YBeKgTsex
b8VnrMZS4qrZwtDDWsEvBWHC+izqYBeTkc5a+blNFI1CiIDCFtrK4sj+lnHlRTDY
62UP8vaZX0RX6FsnxrDxCUGZcQDVQNbSuns74vqD7umkvhVdoydpc3r0Y5J4ZwrB
2rCyRYT4O2B4AXhHsn/OpQma/2+T+J0uPVGIR4eiD0abdusjrMefl+NtHg/oQysz
5B/M5OxWd/tHqdzABm21hA5mKO8lUGftCDPlUZwcXUa5W+GGrcv3ho+A1Krqyp8G
ZAOFF+bQPDgfkQB9+3zfziHbqAKHd4cX2zyAt0un6Nnvy40oqbPHNp1IDsUzpw1j
lRuPeEdI8+34Z5A13L8PU72LzhbtU9v3Tlm8/Ctjd6YbDga4g/sw10VXfM+A6pY3
jMdJIbT7+SgxycLSfCsHuq9jiuCqMmivB+6ArB1Hgi6ZANSvUoCR6ML9FBjMMGhZ
PKFGj3dBeLl6mYzo/S68csbn4TneEza+xJdeG8Q4hgq/FHcBUuVsgRF84myUp9Qa
pkHaxeLEGGDbi4clsyMxmDttf3x5jWJ9bJxAXQpvLRkPtQc6XGTJNiSM04R92ZHO
9DEJl6yCqX4Nwtl9bWOZvUIEcq8bIpp2OqB8rDHjXXP/MpjVi44+ieqK6J9UOU1y
tpwkm8NybTItyRmM8lNelNS7fqpLy69AYq/T1anY62D0BvMWRHgZkxZDqTKncIHj
CO74LoByM2m9CX/iWNQVA8M96OK8R/uSdXSQ2JWR9YzVcEiNxrzcRIH9wTuvG2hX
LHs9/8fJVLlor5PpOVczooSh79i2PJQYRNFMh6QLcsXvCj3gREY1/xi+blvtoDD2
ziZjjwoE7zo4pft6rBJ79ia3+RXWxKeYMlYYyiCJMUvCyIfYtjaKbG2bG7CWcrpg
1s3RzBKV6IueTx9QQ6zfQSgfVZPAR6HK/yGkqew/pKK3nm4lSDNduVzj1SnyiykO
nWYmserU1j+lB/sIneu6NJS+RfiazjaxhNoNViKgw/slSHC9oYhkRjAdthtVJs0c
5Daxx7aoFktvQmRKOtW6N2l40z+adPr84nnjEy0Zn/W/xXfwx9SB8lmpxzP+ZKAX
dIRTGt8INaIAixsnuQnQh6R5/PxFQPSSztxu94jxAFD/3E2CAIdNZN8P4N4BEo8N
wbEo/RyBrW0DW841Geti+LfQFWathv8A7TaiLm0x23uoe+7qlDhP38NnpdUBARUZ
r3rDjJSznUZk/lMQRhKlhrLwGNUtmfRYuQCHjmzIOF7unff+lt7wZhCL+ES7jbIL
XNmQPAEP4EYJordR1Bi7/yJg2nKqri+AHr3Q0FGa/ylVF6JWBdCtGL05TkeDDg+U
zVebzD4CZgr3lCC5LTZDy9KLzAprM/C19LvXlypwsFKNRStuCGoamybUegNb1Ezs
utxql5X3U33S/zWp8wxAmGrkjjLvGaBb8kf790WhxJpJ9ZMTai98wMV/NadtMvJN
DY4l7jyonfZyUM6saylNBGgQWCVnEZS9Ns/9+oy1DACj9Z0Vca8wVIwCBRmOkUpx
FYs5cdHzrgJ3PtUeIz6VfwdKhO/4hCgTP5lJhvdWQ83npcpNUN+yAX8zUQZqO/ab
M0cs/I5N10eG0+ooOX5N1oXAyYT2oYTjEuh4TZ3S1KAb3RapEJLTLcptg6kF7RqF
77IxVrfnzi+1t3n7dFRu2z7d9P1O1uvlhsGUmdHn2NZ73w7lVS0rtygW7vk0ZW6+
FpHUU16i+ZdQOf0xApmigzxrIAyM23upUUj+/3z/cW+jtt/emUNu1i3q2YWL5L6s
ZJGkk65xJwBYannx8Jc3Hujwv4ZESzBftv9nMfLMYQL+UoN/oFETmUYtJKnPN11w
wHegDDsZevfX+yv/hM9Umi3EFeXNpXiFmdXVXJQNMFiANfAjlo4ugoP/kvZ3LSo6
GrD4kxuRA7rVu53+Ht6N+ECrjff7ReXeigM5RJiBwkvy836YaaJrln1Ni1B08yUI
trnI4sTklWpB1pw0xs2aaJQvCch3YWGKIMQcqG5t89jI+uFNlLK7RsYmNlH1G+xL
wqNAIm6eWbSahSe0OsbpLJdKR9ykGgsd7i/NQtvA2Fo=
`pragma protect end_protected
