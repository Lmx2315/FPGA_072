-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
aVk8JXkHN2v5qb6e89SgtrUwcZYesXFgxkxYIGRFATMCJpMuUJtR0k8uYynWSeKXTc4iPAvUw2zC
xqmDPESehpENjFnte1wLbX2irr1YMvTqn5WwIiFoFaoJP2SQLMf72sNBbLQ+PoorhN30PzxNYbdp
qk261M7nl5dibOm3qctCPBjOAzr81y26kGTcMKAK08WHkQPNx5dOMHEdNt+i7+f1T5cCPlPSQoP9
1cTg+vX29dLTUlpACzf19EgutBuHFNOhNiGY9xKmdZSXh3wMvuYKXYeuBXJ7fg1jclpFO8NxRW5o
fdYO8nB6zBoIFt5Tu7z8IM/BaPSHnkxDe5T/Mw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 5264)
`protect data_block
MkSbtyVheHIo8dD/Z7W03IoOh/nft/JhUX0dK+RYpQgOb/GDR5zVaI/29CULnzv5DzHZO47l0v3I
TC5C/s7rJ9F8NSibJSsQ37qFLnUP6zWu7SBknAuzmaK/8dM/FMoR6/1mglFILiX/mB547RMC9ZLZ
N6hD44G3MV+6snZ92CnnZ0PLztLypnEgyqpru5DhjJp7Nk1UgcCnNQf+CrdAuDNwrKtFN0FM1FlC
/kWbPeeCCHxlOr6c3XEcyE0d/VN7v2KOcksOYyUd8T7A7t90dL1P4QokXuMGWVKDh4xHdKp3QCKe
rnWutXSXawAYxRNo8ZAHl8/suhQImCyfcxipWDm19CnTxzfwrbZq60aAPjishpG7k/ZfKPc0WGZG
eAjBWyFvELQBQyhLLlzklJjLxm2BLNVQoQI9uXslsVhQszrLpjkFQ4T7TW30Nr6BCDjWiyP2sdtA
I+3VZjS7aIaLHAXfuvvkeG/ZIArk7okOPpFbyV8cf/ZB7at2IMOluWCCH+uZXq1PhwYvKynZvrIb
EoTsEUzPuI94BB71gfuKNuu6Od0u0io5Dz+XfGaEHld6BE8zKcexzdJKSEaqrli5Okooo27CFypS
COcQszJsoYYUYgCY7nDn5M/h8zWXBuyBb2dbmWs+fJ0vGXfxGIk6Qe6KxY6G4vHetXebOHd1d3XP
YLFbFsm5Wafaaz+2vwRsVPIGlwqLQOlDBLQjMPYTme+XTmTft/Dj6eGnKh3HpZumGQ3ML1irOC2k
G86ju0GngIFdfMWu1EVwu+sitGB2klJfUAhFvPsqjNWCnE+isZtmDa+GFFm78X73e8JuHk8fsPV6
rgO86K4jcmy38Ko2zj76iPBPZNFS3pnisrPaLHxELh5ixJmG00z7/qUKNmpih8ZaMa5SfzHMF84q
pJlkgVFFNPETOnZKF/WkA+jfWiTFvJoBfFG4T5VmVIdfzqVxCNg4vRRNqapPsiF0V26OLDJBxdGQ
zFf0flXrWlUNZnaaqNajoAuoj9zN3s6UsRR+/kaYRm13KrtCSPW2UI26jnn+0Vb7xu9477axDIoY
l/q9tshMnjtT+Z36jZ20AyVS+V/A0zwc5QdyruyokcLcpSbEoUKKdyBqc6fsO7n24m0J/F7BOop0
Azpz/LL/7fEzjkTz7Fjq+OJTvVUbv9Lo7i6OSo7MPF+N7CxnImh2P7c2EqZHhpfyc5iKNA/qEbID
9KdqByjtzEGleLh8Vh5JB3srscP4raXPmGeFVk4nbqnFzuKGaQ4xLVHKnGo06jnoYMyqOQhmemGJ
905u4Taxy+QMrt6S7zXN8v7VT0xpmn0Y1X97VKaKzZIT2V440LmUEZeHKNXtqUxbAl4x7x3v/xnY
26g17dlP4fPjY4yH93r2VkY/E/pB2TrQrjEkYH96faZWYAnL64V9EaIhXxns+mttPN4x5jzYeY3f
IPoUCch7IJnQramVk/jbbqJq5Vync1ueABcWmgOJsOHYoTLczSwhy8qcYKjphx0FhDDqCYZDwknw
dpyW7eF0htteApoPdor3hujqIo2Kr58xCTJROr6oqYkqQor9O5axpqCU6ge/ISozl+Y6NNMdKE2T
FoVIpL8akmWvF6KCf/eybAkxlGM+mS+fD++IKBZa/3ak4d9jt4CYbdSzkIFkxCa8bfnijWhjDaFZ
igJxXQEi3IOOvJDBWsXtdE4u+ZWPfRNGBYyNs2qUA3q1tWCgy4duuM5mDO1Ke034fsMNAewmayE4
1azgaOAGqz14ckZo9RHWM8KFznGAdbRUT9Z8PR2iPcrMtBaeQUD6prVqSA4kT/YiqvR5CYalFOIg
goN7Q/svP7kK6/8jiQ1GyAh+mMlTktImPUFsiaS0wCbaiJPNcIdhAbSWGojLjI3movLZB7l9G06L
zZY+k2dwEK8CW7R/GomF/c8Y6uiY8WIxfSZmhe8AjLvdUUS4oB8zEh0yvPGu49jnqsZ6Vmxu/RJ3
OtEk/2XI/MMDMzoLwU64SJQT3AkxfYATOh0mOpYvSablwp7EW29B0MSzzA7nm3GUccksS0Ajt7w2
myelXGvJctXcHOErA8zfWL80c5KCmv8lyVY+J7RNipXUWNvgLvdT+XLqESlE+SmeJFheREEAQhqu
52oM5k0r0ahe5m19pHcsh4iCgmMbiBIVjPtCg1165M/0zRQUTeOH0Bajo9R2348P6yH8cfk5rRoc
d0N4p5srEalMyTaWLp+ai5yWuvjTqyjyOE/VwwTX9eWxrZUBnZAtZSNCMxg7k00W+m46CTzv/Qwf
brtJpe51wIVtZz6KeQIZP1iaIPjQtyJNWv5+k/2Ym7q/lAqj8spRg9BjwIlRN//1nH50eIheooqj
GyenCq+n30+z9o7FyzUOqbbMWQmlQE1XNyfORdpYrBPfSx1PRdu7j/L3FpqE0vrS5t5TfT27dcrA
W9BNmMMZrv719CkaZKbCOyLOuTANE2jCacLA5q87oWhJZQwFH8gIofGXW/HVa+YZMipDB1pzhwzL
k4ScrFxX5JFJs98V03ufUmDQosO8oojv3KnJH7p3F0qMjadk9VZAkUWgJkP0ObmZBMOXjZpWuiv5
Kj/73beqxm0GTv8gkeRlbEs6wgfL8A/V5Aj/zqI1ZQWyB900Z/377vZAC161nigsOYiLwDzpn7LR
041yl+zcVRFr/fgYoKy9ZbP1wZAuHbhiY+x++Z+FKabrsQbukU8vgbVnF26gu++ozeze0CINpsOG
qzn5lxOGEFa7dixtUv4QhAogk/rc8dg74WAaC3hrjxRSgpHXW3ogC0HgzW+fv+OUCOuGmIHfe+yW
JojwLHr/TeIy5154OyL2/iJsADv6MYOfSnUirEVZ75aSasJjZC968uInm+xrNZaVVLdA9/dI6kCs
fBTF8rQyoTdsg3KixI1lXM83QZeJxYSD64L9obTRd18shHUyLc/byksy5C1ZcU+9Pcjsi9f4cG6f
uiYboselYivjs/NA4gaoEXSWr5N9WUxX9S/KHxXIwgMLYZEgcm9U4REtyrqfVDvT4EGAJK8RSQIH
udKr7xLM/6Ig9YM4YXy9iUDfAVjLEfjxH5a91HcYlnd8uyDnyEBVEfmhnVgPqBDerlWdAMED8sTO
ckIyU/gFvy9rBD/uZYDlEO/GQG7j13dUkCu/Mng1Og58Hx7sm1oKpjDOqHsWRgVrry9W6b3BjQ+2
/8p89AzWanMtwSomSLlUlFhjTmTgyGLWqOIvCW85W3pYsXxGaOToeNgfgmWXdwVU/zYhNqXfencF
ZcY5biKlZHOwJ6BurBYUu0Ys4xYyGViIz/16VENZHPi2+U9KKDofCqTY5r+UOKk6NTt0UZmA0oEj
47sqTb4/jAyNmILL9hGn8M3Ud2/GHWkbkRxMlxPRchXCqHbrPzlYgEUjx8g52aPZ7iE/cO6pVM74
Z8QH3YrZ+jGtrjLU/iBCrhfewXhxwnOQtcP+wMbWTnEjde58u7DNTshNeA33YVLdC40Ib7eVteO4
yL2PnqQOMqGIY0h2wYUeyB+cpoLCr1LrCIt/K/uE6CVHZ9VGe+MNdLHRCDVrcGTfpsr1BWDyjhUI
/bq5CRo9l0RtiZ/QcopEmBfrriEH/F1pvwzTYTk9Ay/m3iPCDkE6tx8f3jcKSZST7ptYdJ/DgxtE
AxdF36TLx+WbTXGSVGh1eD/wsbdbqKRxF4jcfMgD4sGqt+8Mzs0eFlBkxfVWHu7wa3YumwI72hLK
Lg6NDoDgXLCxrEfAAZHK4LO96lyK9GBEBzcUf02nKauIO31jjvmgT1oQ92xmIgjmHPQbeq3Whxwv
1+XR/72aOm+jV0VvpBtAdDni4SiDOImSgzzzIb8NW0oioy8WTujN5N8GQUFSevcy4QiLXBdIt5W1
6Kv2YTR5IXndG6j6XtWiIW1Ddgskerz0LScKCFK9hu9yj9pBS5C4jd5F7Nvhxwsq1CR4Jayt109i
Ir4K//NK7LgxXheVu6vHt2tFgxMgNzeJItOd5+2erXLESjvk4q9GwHBJVF92wsdg+t8WKyBkLMOn
68y3AMdcii8LV9xscIWu6XTfhbMbHIq+k0TOzdxwJYjsSfPbNRWyVwXh33r9t9aG99TIwDVOg4aq
E6gFj6x0ETbTI/zuUdFj96gs7QyRiXotWI6pjCKjCxIXM2qv482TzGSRGrqYxUybi6MzRrRZErUF
hDCL5gOvsJJxZ7qHGFtjz5b/b7jsCJ67+SlTnpoG5SXD3OianjYyYBoB+iK3tpvbyGAWbeMmjqSU
R26QUZEzwIb1owhoEm1k68kenGKyB7HbDvp+fE6+XqDovX0zN0OciOyWWW4rtwRJVTgNZvBrKGzH
mIte+QN+N1EuxbZsQLscQlO9uYJfh3OjuGGNSPcMfQRanSZMKN6LYPY4KrFcvK7eBTmlQI6c5IBJ
NnPVs1uAGlaYW1MvYcTpHATkp2OLAIy3nwDaJ4on0ka9V/n43yy3MHAiB6A7sPV2xjcf4blJonU+
op/jXbPR7EhVIgcgz86DifDJbI9hGdf+36HE65xQb8BvSVS+IXXAYKcDnI7rTlB/xzKcUQP58+H9
E7n1HqTC3E5i4yBnUJIcuiAFlCraviAyZmuNW0Rb8GkRVh6tilAUq91dOucaQf5b3zk98HhxfYiJ
fzxi+XL6/tMPXGfXq43g5Wc4Aeev9o0C4gTesSavnijUEMepTQ3KdD4KcY2sjIwD7DIIyuEh907o
ovMmJ4v6wxX8JDMu1nRAY8qUj/2j1WORKJBhs5YzMYGv+Iubw7HQq19CN5v+bwTb7AOLfIK/TGFV
2aAwnfFunT0fgv9lZWdmX6H6l3yi+Ix8zKoUuS1hVWhtWZej/t6woRi4nQuMi4m3P/Ch7ZVkkeCC
RTKatDSPPcGov0X8wV9Mff7Ii5e6X7VUNQnQA0kGhGEFaMON0k3C8fbwOiRrrXtmZwtoB0UuRbqy
jrjND4+e/9QrZ9rTpMeZnhmfJ+0jSBzNDRea0UDatM2NkUmGMQ9mV1QvjjA5XWwkjnsdb9ybQegx
nQX40VXno6ZihtQ9/henRHEBiqS8uiftBBrJ1P1YfaVZjrlUkj4CPzecN/ITaqoCzl2ukc5TgUQj
eryv0S2YRibWdiSp8LXGFaQgsdqqll5ASf9eRZs1y3nvQigkozIpq64s4HcWzG2oxAl7IaKIyRh6
gnPyLVZEnIYac+xIg1fKwEujVqLeLQvY+LX+uzVQuDIGuVlERL0+rAGMU8+p2S98ncaFCEBBnwD3
AdVoji1Wh7iHYfO7OMKxOViXAu6FHAG+8Y5NLr6yHE4RBMTmB04+mZ+wd+LYHILeUUmox1TPquiJ
+TEgjGGb4RrTOpy5BiFQj11Ld+fM5oxLnHxIGF/1HcZA87CWEHMSJIBU0huoeljF8YEDByyYjy+/
5kjRxXJQY+uOr5k0BjEMsLRUjiI7k0uI4wjF2LbnisGRCBhYUN29DlXFfjkRgJfDajMEt950JIky
BM2c31MDkyDCNIgdM8tHPHlR+wDp0+n076uZRz1MeA9AjvbWhlvSorsYLfaLIaK0ROxG9bRdmpbl
zxpI3J0B2TUPT3vux46bcESWQ8t5q2fpOCIy5JAtbi15hRdmf99//P+pNJbVPtdBLomhaeLxLko5
CCSlY++yzPByqMnQZsV57Gsw2jAmISKAUFKvbJgP3E1wff5tpJNl1lL2gXDfthtYr/stZc1RuRNS
u0uI3fcSroXSQUyhZq7fT//6nTk4A5EbVAWq/QXDKC2104kvqNRTkC5kjhchiqPKH/3nkNXYETxN
IU0Gj1fIzP9N0f+W2LeycEnFQkDX1GBIBU5byb+py4eIOW77ZklWxJfFQdAThmTXrbRI6Q7vYbKK
PeCGrjeDIJjwuLT8Kh3LluPCRna5o/KpPdtRFYYllAN/+NGwbkHy2FgYs9Ilw9NL9ccuEs7KyN2j
mhG1IpicMGW0zPRQKwS03FFk3FoRrXcACP0baQI25wNRzJPFoFA17+hgtsUytjE77QRt0V17/Qme
kY/yoxjIK2yW0PkILRK0KmtUfU/6rC3lE9CsNX6Vsfj1cMGKmoYAOd1302TLCePgVZuTZ1uqOd8v
KRzwmLvcbd25a6qYTH+ujwYyYOY5E1w6AwVfWOspUm3k8jwkdvTYx/kC8LFNPpQZVbygs3O5yRkD
AWEKU5T5jNMyJaHMfXATqFpYK+cotmqaMX8JPL79E3LsiqK9aoj37AwF4QfmtYIBOh2Vs5c3AZX+
KP4wJbzuP+NgbvlSCiJm/vKqh2Zubu5soaDQn2tai7ny9CDFzA+UQq1Nnk2q3Wdmt34/6+69fwhw
2eueoPdvSjvm2iVPnG9yH/4rrj328zM0JRpDchOIqUu71HlywdsdM5DArtSYpDB+ZLolKD76nMDO
S3RVQTx9EI9xihDzIAAFYoR7207elRvp+0kweZrk3dBHbgn4Ulxz5wqBwRZatoMi1BGv2K++5j4C
MMoy1SvOojHM18BmIoE2c1k6DG4A68Px7AO5N5L0jd/4RaJsgr5tr54i3hhdNXvmwMZMLMdY4tWM
V31Nj6uDY+jVBNaIt3MWfo+svbyToA0wWDIBGwqWpT2aZJfgrMIOpBsXv+OwmR9V3LVo84t61XtW
hktUAK7UFNVSub0DCObwpF6C1jQ56k4QlPPshv57YCe3BWonqsuG1b4QgRrIoCkC6uLs/qT2p0GG
BKyQskDqDxgESk2GBMXKDAaieQBaJmP0YQCuhH01BcJE6smqgH9dzKlL7VsqrYoEUOm8fidwKqfP
5nXz9EpluvlGnzwBXHbITH5PNvMjgJB7GavPi7IiVx9ERJTIqc5GCxOZETXinoRdstQD0ggVYNrs
j+4B5LzLYe2KF0xBlTbHDsQWOPQ1ug1zZd8qdGTIBBRFS14M6JbQuF3onTPgEyZVsDFVvY+UH20R
wjk5A0eyPHaVmwlClidbRFn1tFRjGkPieUcxUU0jlLYi/T1J9lzfN2vVYM/1bw6YPAGGq24C+OWM
h7NB62u9J8neScoaXB9+kELbcMk=
`protect end_protected
