// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:36:51 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
UB4Xk5XygF76qaY6aybRpOx/tB/lCN1H5ImADe2XR8eNntlovcYOt5rVwFFF5Die
t+rfvrrEH+kpMjleE22gI1vqLGcBl9Dl8+LwxNb5d3tgDXTCT+vqiFjL4r0Lno4i
S6nwSQX1fOlF+VCmV91iAGmWI5DXNYDri7IwNeZ3I34=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5184)
4Uq66sIfZbV7YQOEvmw053Fl/nnmcruon0uyXdHQPLZ4hNmq68BHSqq0YdvyGpUc
vcVfK4aZ/bKGA+0QMOxUna5WKhDYevYeLDrDFPYHJDg0L47SklbHVDhaIH4k7zd5
RiwKINfb8McZBebvV6wLe+JFDGCmwpfxkw+z1WYYNKaNDhqjwaVouZO9LIykbuFD
GjhvWndiwX4RDs/aJa4h7edr8ZhRA8NxKybT8/w6rWSTom1a5v8xLm6FEPpph4U+
MK6/umxPiZitMDUGuHgcf4zspT3x7ORqmGgtk+BflQLQF8jg347755IO3UV9jHZa
ATXfik6Gs4D/rTwD9Fmv5LV+dxfxTHCSouQI/udO666qQE1HCoAg1ILbGWThiay/
0RPlDtwvcWwflV49oa1cuOawZmS24Oliu0CN3mV7whJQrpqXpqrEGeDrqNIQfvYB
6LJuaWHHdkaC22z7wlOaVuNKT+y+y2YtyrHw/Bp0fUr1v8vU7kM2MqK2DCFh3w5E
ICS0xjtxmrG5g0Vyf0YqmHsO/GI+U93aWjtJtncAeThRXInqoCUVDTdm+uvcS3NG
lFzraoZgk26FqELLqxCFXkBR2TTWJVH1UOuGCZcilDdKYbfLwYHrRi4M6FUu+xrF
1jgDo9w6AG4y7Z0RrS1lLHIno05pydcfPS3Bvi0YsrD+iXRK/yvCORvINLrqKLjK
HFOn7r7M8WP9M76Q/DACzwucXUDDPVLJjLOKr6DNuj8j8kfH7F8t+6UD1EcIn/SO
bBWCgvr20gkNZo+w+sTKlvxnzJJF5pSZpCYFP/EE/dn5PmGtwWMuGKwaKQLIntaP
QvpbNthdmFDzumHWMKv9pGDbLudXQPRWXTYA90GHYuNg8yQ16K010v12y1mjWvID
o/jZ5obql7wzPU3RJ1K9jMElByMoJzKhWzD3N1KzUMXIgF/QQQIAb3M0oB8oZqtW
NKHQzLej368YiZHcyTUSexp19aCkUmdPZGW77onmnyPM3pZWem5HicPYIaP+5/On
cijRfMzXZ8e/QXeFEj/y8pSxr6Z1O5POxWjSCCddvUXxon0hUX6R4vJx/SGHQ8cg
Z3mQKDNY01ugy26YUosYUbeIeqMLGiTsKFB//ujgJBFbIWb6wGizUcIDv5iHFy/J
noydUh6P7ub49oLXEH64njg9NZ8tkiEmzkoh7IqzE43fJ63p/Hn3oOuLZxNCHCTp
KHq1s1vLZ6Shu0aJ2DxvCq190XauLkMYhGMnSudn5dwz3fRTyX2rM0Xz7lXPbSUk
MdA33XD25HHkzLvalOzmh2OrCoJSJL+F4rwdHQdjgVSyBslwYDlaIg+dTdgbUWTw
r65rvWEs4eMOunSiz5GzhH9x9st8TNT/n2jBpC6oaqgBxc8xHIQb7TUbqY22yItr
pPRRs5uRH8Fk3S9o0MvU0yfSVkFkzsJHXxa+mpnKDCTByDuXopEe946I70bQQLYr
5TGJ+xZK/eDKVIPlpD8UiZXeU1EE09jmmPpCgAytVJ6OaYapQoBbnVhosY9prGIf
3UOWTTJaL9SFIHCFIJO7KhhC2zquOn+CDDKm8sAX09PanIEOWod3LtIfRn+oIKZC
ZNQY5p8ftjc2efhWVqUah9YLIe1PHwIEsaYeKy246HIvmN4y7H9Kpo+F/J+Xd8L3
r9HKIdXEY46xBuGzSAPSNbavlShMIWSJote4JUNGRUK/sriqFGk3th4qY7vr+oHF
YCpCqcqJO1b9ODDi/5OQQ/505oHEBfanUnivxd485NJaPyo5bnCQFUEqu+USwP7r
/iIQph7QefaNPtHqPaFu13B1NoN2jnGNuhjsGHbiaZ+yjZ3P4NbY+1Cd+tFy5Jh8
a03IPcKVeuIzP5nvDA1h1SDBf0Ie68qTfqu0m6qtobZciy4XoNrJEFiexSbuE7dd
fc9EyhwX+03mjBGyeoz8eRupIZ62lmSypozNMNR0qvd2aHjv3SfDqKosDRjdb5+d
GXeQt6YCYkVP92JzjSOrtpL/PWCAV7WJ1FjJuN0BW82wrPTuNqT/htLw3zQd/FiC
cYcWPZGLsE26lGFWt3g7HqsHf/HZg9/7aJrMkz6YsdCpwD1exY/M1EIhbKB7JgEu
yZfYHpwPr/WS3W2rXq+NVW/4lJ+YWRGt0jk1mU+rI9dy7PavEwQHZ4jqUvOvv8Ih
z7+ZW24obCVdO3Tam0e6EtStXxR5JHE1eXO3rxwDByW+fSbxkP0lw/2Lc7lv8No8
4O/1IGJN6XmfnwkF1Fe/43eGVNtFEofq+6S3eU7eFvxffIM+nGX7kHyBJN65NFzd
4ylW7Va94RRdPzdIzn74Yaj/NEhbft0k7oVErjDSo7QC+tpFDifNJKW3vVweyK/b
680y2e8rUiRC0fQH+rRq5Gcp5+qeYEq11ygtVZ11dNE4DAID69BEhUpJyltwVj1h
aYLxxVrz2s9+RopH9Uw0NT6PqpeW+xlZzyAfx55YFqt36+dtXxlgkRCgAeTAqbkr
moOAoSOjrFtYLvx3gq6X0WtOV5+j6gfXfT1OhhSKOi5PAQ1ew6wdpVshb/QJsClZ
B1OaenPbsFfsKO7h3KGs0QIEEFAls8iRvxs4slpHyWW+kYjl6q/F0IM8VfxlE74v
cXkSrJo/+dbrkemUY2dACb3f1mF1WNUbybq9bZqM4/ZFINx+kN9MUpV50MErLDYf
TMkz4SAoVnACc1J0aW9vvU6aNlPulwmWBx/JAyn/E4KKmXHdf5eQqnxE/LB7Ct78
XmX8fnWBrG8O9D7DsjiZZbbUCzI30U/tAIFvDgtQFQQJ+VNS63eLx7uTcVTloZq8
peNqWsC4ILLiVtAtEeQR+f5tWK2aVANkUxabwM2a/X8f2aeYoEA0Vd3v54XTef1G
STWZ05M3xmDzQj/CNpdQ+e2xgyA8zLLKAcLzdb+BtFkJTmjMRXJ209O6v/NMvjCJ
+k/oD3Ku4CD9JojhdIvL4tCLL+OJEp8YpT7e4oBq2nUYHszrOCYywhVQ3gIV+bjD
QaS4JEo719NUohG6XLz5MBGi+oq1nFolo4Q2LMggAmMy96wNis4Y1ZqHEsXtlzbD
FW+whpDGWU1QFipe4s9D2IBpu8NouId1Y3EU/XU/TlMKoxmy8cnd+GHylrhy6fXs
zj/rX2pBDluptCkd171hspGrlYvfP/V/p9OhZ5eQJicEHistce2NdN9KAc1rSsNJ
JtzFYYSov7+xWRgVx8UCd4Mzm/54V833qNSEJqDqA2fexdPdclmJXAxuPFYb1PVJ
gfKnCfSyaDe6qSOpC416h+oaOh4SLRuPsHymTukkF6oyBHaW7roHzPTbjQs8MYg9
sNw+wbJ7fy6sz+KS7RSblO8nGrE5GhBMo8CSVyunQLwBYqHWQkz+iM2vE685qdKw
Q7AuKFoGUfP7MXlg7//aD5Wisau9gTT7erCluqPNy2Xx++XPdJAYKbfVEqcPuHO7
m5Jf18fNwY9i3wU8Gw7QIR3cgDzycBrXWgJBezbhP/ihhfUpfuWwqETtdo3PpWcW
l4rVURoRe+kRnNgFyfGINKGI0Fll9259gJxsQ0COMv9LS6m2CmDsxg/ro6PE+9lH
MFdafn97b1Hcra0ytCzZ4R17ecFPQKa/hlysiWRlx7Mq78FhmVXvZM0nrc4FVdp1
3DC6uKz/rLkL4Ki/HaVJnbuCnZcHO5DCBAUWU/vNs9RA9REQO8vy5Ab7t4taL86X
q/5WTzCd1q7lh9m/wXEQLlO/CF9kiBTaUtkLxxCdDuuJXV7Z6iGgXTNIio+Csflj
D/taHi0HLD51/aDb+0ICoUuPlxKVBvrVzaCK7D9O8dcPFtEdzNUxB6hc9FKvYSrV
bF74vOp4CxOtF5KImzdO8Cpv2XwBearp0OOzaYDBrQPWP/p+ZQtpKIkKNJDvIpFw
QIBswvXgvdlRICG18+kVbObNBy3/x3qiwN92UAwJ7ZBM5szEk1pDllZSiitl0oJt
s1FE4rDAE3lfQhiDVJO7EcPru+1kzDX1utT/xDDyoQmWrr5AeTmznsJpDJ2zKu8I
8hNu+dOXZgcU5naqh5D2JJj79G6I994arH4pfl/1u0u2CM31+rTQIR5xWlG8RM7y
ri9fr7auvsSBXReJMBSheYfmBV/BI9yVSvYn/KJe0DZDfNKOUx2kEcUON9o4njbl
sjXcT/HrHvbpMmLW4vyWJIseHOhmbynrepbjckWAK1Tlw+yCmNVGJ15wiFyzZnfI
kUoTis1gmDRmUJzF+Ew+PUstA0pqrj2RpiG++OR9QeJ0OmHInhQff3DFHUWrz/gt
Io2diAATWU/1MOiiIBEb4ZjQHmF4K0NzFLGOq9qNduM2WQ5t0FyRh+0s0zlDbtzF
9NlKHHgC+JVY8bJ+qDjhOw/+iz8OnT1tNQFdmnFj9AX8Kr1AotCJj1eKrrDi9uce
IF79el/3gPlRebLq34z0QGXfQNFLsiLHL7mpRq3ZfogBSXSJs+2GndKnJShYxXL2
ytYc82v7X9EdhJApBi2Q27I1AfD/XkrIjj1OkVQsl2F/fIj/4QIv9o3ohBnhu6QG
WynAF/p6zWdufsTcrrk6AByNhNI1z2lcBErTnRPoDFNgi7ezByb2Cnf5lkfHDHCw
4usooO4WdSO7k8oRGEJCavrzgKNktxLbqNWTmg076qKuRNkCaTAsiPqx4GRSZt6L
4rwOZKvwroVGb2Fvj7AD3RoLaeha8LNs/4waGrO/vN7fxxKvZCdk9aVz9fA9jPvE
NkLMT14kpxELTa2FQwMcezJoSRPcXcQ+NZWNDLq5SoCsESB8CY54g3KeVXQIBIfX
xDSncRoBb5LDdOoixMtGNXo9IGwVt+hZqYZ01u/p0/YyoxP9Of7FffwsyrnZVNox
W6GKL4GPqMJdzxreNNyxGLskS4i820oPYWwdwaU3avUjlps+ex9gfGEYD001hVqz
UbsmCKcYfUd+OCtV9lVIT4yiVnWxloYM3zipycy1qbTkjMvSDE4h0FV+OmbfHfDf
+dWbjO0GoLS4A6dwbLaeFePvqfjDPRs5d3ut2W0fD96bJbr6yOajCWVsyDyxKQCt
iytLfdiP2R2lTqJWGWXbPGnAcoYaps92BYmwKv0HllwT51VF44f06LrRjv9rgEYT
qoPcBN1dnpcFHV4jL89gwEf4te09hraXE4pCxQmDvYKi8+3zjTPlreGSwsUJ4YFo
jDPUbrKKkO3zGWCiTjI/oDRt2pNxFlHvuN1x/gK65SJkxV2g6iLRDpgYDgVwUXiE
mAaqjQ2zz/LcP4iwHVdt3IefoZofsbjXP6NYvb9JEo28zoE5CTP7rv2b+RMdtrVY
fspDkVDjafG8YZRuSbw6R9hpopElYuLbF0oYrrtDN9h62CXFgavs9k5BR8ENqpsI
2xjSuZzGtvvj33jVE1K5HeZlaDAQ2K2lVupJww4stmqyTpL86fkYVrfzJ8vlFMWE
3TTSxmWE5MbpYlbXblYpjtf1FJASpkohj4Aee0kZ+Y8Q5GnJ7Wc/A6NPTMDMpqYK
fDzXwa5TJihBEDDqGTBZHP995S7zEyBE5LymhMeXpARYzxxUcddxLIxg9PtlkO3f
/ap479ewft2I5sJ3MGI6RGBHm3om4XgSkQTDldec9B2Ct8WB6mK+caUn4HgYT7t8
E73G4YcCuz/+iAkVt/Rd+3v6FNqJolySFj5F9GXH24mfh5BqR56u/3tDhyuxvOwD
fcGyNa66A/mc+WbwTL/D7LG00cX25FRw7UemEZkzqPLbac7WfE1XWq0Cu697Pwpl
sGtufP/HI3XCFh3j79TBFd2pEbFjdLNCDI0CmdaFVRmkr75oWQSsSfARa5O5LFGC
bY9CuPdYlOKqG0Tz7syeLPcOtCMSs/S/yLu9NWt8AMPEauxI8IkXcUaI6qCpgTuP
1tSraRu2DCkM0xw1RrsQz6AGscsRtAq+YQzjx/HdHP1ximaYv9uatGuOpr5mXYYm
VUh7MjBbRRz5sHF7iItE3Y3kZPNfV92XT3WysHUGZuZ2+bnnTt0l0uULMyhFRrt1
Vop9agmGlgvZ/+QgEg/1HWcaSpmNcfbEuFHIr3EUJf/LoKaJ5OkcZVliqN7nM2dl
lZL0E1cRx9AzKTQVmAD10dnxhlVkrHInhImhd+nOk8hc8cQE2Huo7SSEcdzYxAIr
rVJywUuxCEoXvpkPZcDlE1QaFW7gR2TevN7MT/Emg1SkC6+eyexv09nBXgVBchj1
oahb9eEaGmC4by401c7ZMu0c/iBSfh8X2ZkvdYEv8IFlGRg6NSsM4rhaAM3rT06A
hR3ePUx7Z82M4tDvRmEo0uLuZP8tUvAJUBX0aLtx96EPYSTlojUojxvQRXOmfK/d
VEVTPrvUIzZvxluMeGIvxcwUuJoZKotsUBWnggCBrMMe6L2qerOTVRGgfOI4YcK4
FDbtFxJ+Q5PTgQJ18GPKWeu5WFKxiiJVQJyjdNMowUO9VOhBsDS6D5XMoBitvMQS
W81NplDm4Z7rcdLqgVE+RS8FYGNR5uMYzChY58GyF32VnLlZF3ZGFq33Y/Ud7MEr
5p8oCCkKpyCxbVixlgysjCSp/JXks7mzZ1Ll+7nK1WIYQ+inEIuk+dvm4tKhw5nc
imaiKO6wTOg1JrHmQTTZig+jX8707zuJ0i/rbTaqpP+olRf/DGN/8r0VepjpjL5s
ZtrMpgqr1RFftGDd+Dq1LZ4T7VY/8DWDJPnKMOp9vo25GOuoZtUVYaK8muzN/3Z4
y9o39hZWj9wbY0qYrHf7x2C3u+PcwoCw5WVEPMHVuFO4Q0G+IUpfPIZHvv8RYhS1
HJn5xBLgoaf6PGg56ptOV/DXdfLLjHIk3gzH5KObygJ0WDh1YFaNHHFqVj4KviO7
tEfoSP8LZD81T9RX6lHwqQI1rauNGGVNchFBJj6MP6JbNsek3ogdci+SqTcf4Xsy
`pragma protect end_protected
