// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.0std
// ALTERA_TIMESTAMP:Wed Apr 26 13:33:39 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Vdh0qfjgKmGuDrgoeXB+DJ9wG5VFQhK3/r+j16OMnFKPLddRUGlK1g9wehi638r1
UxgRshHWeFj08V0XbJBz7y5zxdiMAk/ogUbzW3iP4OliungOEXPW6Ez1XU0hWFRw
RSSwPfVDp+OLcZiqp21Q4hEJCvolOhJPHJNxvvtdcgQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 10256)
KEweqbd1eg9OcqaHnlo5oAMaEAvMCLkVpBEjqqv9l9se10B3OpJ2eqaWxSRqAsCX
sGrWvYnIftxxTsKEaJHkcugJOB/ci+Kca1Hoja2pU1EoIqoLp4To55u4Vly/Q2j0
NgB1G83DiJprO5EpAneFrxs/vFcBj96OWwgSRdYOFLmisV1qaEG0CWFsrtCG7bfD
EH2grbizzLGXhc98KPE2DksidBViXbhcZRUDnOOlwUZWOpGx5wHHcnAdNimThYEW
c7pafOhQCrKqdr0RnzVKHAAtSw6ruNRE8DOpg/xT7NPUs0hVM+a8MJooInfq6FnW
nn1BMJMYD3JfbTvPYEI1T6XUYONFAjYm4Uk/Y0yajKCB4ydtgUfHnhg+pQ3zC9Ls
WpuwMbDRtY52W6vq/PQtyfDxonmi+inbPl8EcCLRDlCFoon4He5tHwucfhvwKgXx
o31V63UhUODD/PB/ktt4qRfS9NaNrfSNWIufJ3ngWQaXl1mEr9s2aRGH2IfIyIGS
4H9Ew4cSPZ9910esjpwfkpsr+mInW2Y9HVZV5OCtu9g37Ju+OAUfElKUSCc8GfuO
zV/NFK4FnG97bG9VlGX0qCE7xJx17HgBXidPU/vLEThBKW+U/uIzyMBmo1Zn+bce
tbMPsYqsagpQrIL9Ev313cA5XwQ5AQzFgBG77kWzeqy9OS1+gmM3DyCc7JcQj1ya
U31CA+8wq0T+ipqEvICCYCs1+gCTofiPC4hC/fc+1nhrVlql/VT8/irShC9QBEWt
S813dAlZKOTWqpgDbArw8de6Lmh13Qh6bMrm6GkyCn6rxbJzwynWnQkqaD7VyT+J
5c4RcxLFKWk1cLQmkF+FXymW+AMVO0N5c1Iag5aocE1wIa00U4Hzp87Azhrtu8cJ
BMY2JCnaXOmR+yc3DnK7Q7n5+eXvfSryTEQmyDHp/kB/ATn+NIRoZPO/aaAQvHld
fEX1Pkt6rYUEOdjuEtMoKMkM7GMbFvB5aMHyOD4kmq6+iETLTnudTDmu5eOfpwfW
KZBK1jpKNsr5qF7nTnI0vIbo6gh9e285efyROf9Ts5ErgqpMWJjTAErdLtkPi/iY
VB+LCIiKoowRCHlZLcjK/YwaHllVWisWRkHx0zPr2iWmJ35ELGYe6WEKRdADmtSI
6UZfi0uJLxHhec34iDdALsG1CkFhF/fH3fSnBxPjmmJtsRHO/AkPgCN2VWQsCBMm
qj0ocSFHJg483oXLmj1o3QcS2WsBvK+XFU1mvZe9KnohVAZaknqLcLSVW5w7XwA8
r8/swchWeX1u65elZhZWeAX7tm99PyakguUEh5FZNpGiyi0B3LAAkOFRF1Kj03/r
emgkeaGKhiV+dJITdGRcVpO9dpkfpJJ5LQP/f2rOzVF7WmdY2Ifl8XzOzjGlZ/Kn
rQq7mhmzBVCuA53Eg/pToWCg8RFyASF8S7CmgLVGWG4GxWRn8K7mnCqRmfGCxA9s
XEMR0uY7fQ8CGYGOX8xhiWb2Kis+EHGZ1lXnLAt7v6bb420rj06eha2MVuwEMG6u
G3/GVmiS4fsxT6S9pPKzEwLhyHRbwpIbnEqHdXZOc1jKsPJBcqVz/GcLRi86jdY7
sP8BipBz6jtgLPUx8/AVY51IXTdYL3jhCBenz4JokmnJbDgBu86qw2FeXAZfmd/8
MhO27/qnkpR9QEtertocNq0iq9chXPCkCDQWGsGzaOwmVGgXLLaeRTinZw1vCKpw
VULF4PAkgg6dF5gqohEFVqGDp36BFA1+nj/fiDVTefEm5T9VqYgcksOUCriH/CwV
CznECH9aDTVwlcvnlC2cu4DnF6eDe3BGKNdckoURlbj1eqfBEWyGOKiQ9hmQkHLE
/t2C9B5/OVUuNwvNTxPvdKB13FwGilGZ9kHTkGxjs0xqWwWWzaxQT860D+9MyL9V
D1GAbXBQ7UpFx2YXDD8W7pMQdPIJ8+AV7MKeKqaaA3jxf68e5dD9ZXhHjbV/2PcG
8yfVMUfK3TOoP94E6qoxWk1kH9Bh07VJiKL3sW60IV16daM6Q7gSRvQuLx/h1gB2
FmzKco73xEMXIaTksQls3RFnbONjGSgK1UJ5AtCLf5MWkfQoDr8DCC1uWbzYKkKM
+iWfhUQh5Hrzxw9xqMuTn0r2EwXDChFdYHrESq+Gm9f02F9Ctsz5QatcURGrpwYG
wle6FMtqLPhj4NC4EP/JLiMUFpgfw86DqlZfT/bUzOVoht+NcDMP+UBeHg29pKiN
Wq5GepqLOXmg4qW7rAV24MB57xU0/2UrMi9CsYfoWtvlVYTeh9nbA5u5wpKiyUww
+N+rJBKojVdx98Q0n8ZOCLX5KILCO//WT4TrNfmzro7Z1aGZ1oMzMez26TsFZUtc
FykolxNDoz83I/Jt0p8E0Jy6iW/u6t546sLvTQKy83NP+cLcC+JjSdGPeu34YqbR
DrrwGn+2SXxariCtFeYavydtThBw9mGOr0jJP+96AlVPqiIm/ZjOj2IeGG9P64FS
0gLrYKQigO63vPfN9lLwJ6yuVKYF9fkdU6D5xQcm/o54sTlQRsjBfY2v8+ELVL4S
i1ZaOPX7aQIWiLfXCGk4aQJrXh0iKPoYyAkji+E0SnxuAfOWkf8ftejmJfSLDCBZ
1C4CDIT+FeHo8QI+QtjFBOEFNF22YQ7Mr40IXin/aQPr/KN6pWX9NPiZBJQjEgUb
SgPw07pH3B604VSfGPoMbSyOY55JlXPXC1eAvE9b58eIxCM3WmmBXXLdG98Nz+rz
uSUgKJTIgcAizb22sj1zj6fDqh1MYOh+7DRh2WVmQrtNr6+QJA4rvpq1QVMZKrIy
HZ+M7RcO6MbA1c2Vo5lgA8znTzOWRNxyNVyjMPLDWmL4cDPm5cy3B2eQrrWGBqfp
cU7q6efkZDpaCqESaOeTK6hvKAHTOovZ2znDlkYlvvhrr5SV11HTyLazgHp2NWqS
J8/yGkRuOeqvIeeHwcwFa07prliuBpySNKOq+oiJkiMREgiWTRtQFvL6nAoK2hSM
HoFNOoo7HOkO/5y/TkNYy01BsIkf8KVHX8Xr7gwgqsq1DjE56blOYnmkM3gqagR8
NEt/tNyFss2BElGxB+ftz5kOovDzD1lLkGlGtcP57z+T80PbP6Fkbnzk3rZ2WAKL
ZutXpowlAjFx3It3AyIbvEe+jTZH/IwYa6pSCIQ8NqQO8e0L1iyoNn6EEi/K4+za
dO51JhFvyTm0dWm396qvhg0ErYW5JdZ6OSIweb6Mshp/KP/0CeaOPhvi5ab61y9E
053MSXLzFzhPh6WuQOJoRmF8vYwenMa8ibiNCUL+/MEnJEOHUECwMMjgDe8wwaNi
7uCW4uJdCH6lmIDO9U1OkcpSTyn92MmK/mcCWS26n3evhTZzEGwIr0Iun8ppyvXj
rI+ER/u2LAn5de/k7mYPqJEhjLDEifMWa+a1h3viMfcy4D61IK/6/UA3/lPxvlai
y2ewpdF0knM2pvSIov1op8qorOD4x3lLP1wTCLiJC573KNqMnr/s6qsO25MNWn5+
mdPLzDSV77UDHUChEk2wz62JGuX7NQvS9XQvUDy/8TLK0dse51yz12p526bABWXG
u1QZCR/QRZISObEBh2v7kxFplbyZMCIxYICdZyD5ukt9aHcdy9ztE7/CPt8wAiJA
CqYuwnqpt6eIvv45nm/XIjyi+p9b9HMqG+YGYUyB0p+8RhwR26SaM/51S1VMV9Hh
Gq8lYdknMVz0iaBQD/CEAZW63vy4VNm1KOCeXwT67WYA04Sk7lWpsSKGomx/y3sK
tV4PvFEZLMrMH+mBVcEwQjOb0rrHiNPPlNdEyNCh0cAa/rwUiy1eeYqnl/MWgKF5
n472xWxdPUHDch5AGfaEfV2xv94p5Eoy1tpezyTCqJFZYKOphGWipwEgoHhOZcwT
5YhomARPP8K6NMN4AYIq+ZUTPfSiqUlhYREorlLuqWNbFu/n7Y5cTAf1Mi8x7F6c
fzCIBqV7iyti6hNbxVhUNFGW5EOtTHnYwP5N9Xjd2XaSgNaRInAYstAFxwJchnG0
qF0TwsS3aMZj8zhA85R7zgUV//KbenUDEcFiM8jLxUylS7LKk//w7ncSN42UeA87
7WO1NyaEihGv4XjIPnVuUNGSqtoV7gJzhnvO0LivutemMVeaH4O2P8KKjZitEJhR
p0cShjc6t3hnrafTA1Nl/PZ+F91sgLaHbOs4+xMYfm6FwtxJPUJwpLoWTqfGwphG
9izQ+RGikgVEgtSkQMG9EOJZ6jctAfdu1L7Sx/G6GQWBEcdhZAnjKbgbU5HeVfBl
t86/+DXYWIOl4UsJAo+Y8975RoNPCDeZM3xbXRLMuI3MytGgwYZl7b5izgYaIBm+
jg5EAJ2EQhnuOfi7OMhaiYP7pe9xVPHG4SBhGf4AT1swfQbqf5PO4+cKhgjMTJGF
6cFTQ1Bdl67Kuk2thhYSTcMPB25VprfvF0S/pttz5elqx8f1dBiPH8bLL1SfKyUt
p2+cGczbwS3/9knRakRkDF6//OzTP9w5Pbjsb2N7p5lha7rA8GF6M+iKnpLpj6vF
cRyxHfEgDyBs57K+iZWiLziuj1DsKUTWLSguM6RPTFd+4MRgUZJJoyr2MhQnHd5v
jz7w2jPVQ5/85XaZLSMhEDfoSjsw0DI8sql6GQcQuJVh3W824uwJaj5ZI1nF+NIv
XY/eaN4VpI+JPx/TyhG+qQ0oYtLjpTWL5M6YTszkSHGk/t2vTCeHE5Yy521GV7cK
O7cD0W6Gk4iIomj4vs+sy1ew4fBEveV5eK++Ull3h6cc3VDIx3vzUzisMYbEYtAk
PvsJ/dA2bkYjXxQfbgoVnsJRodflxOh5mH9oNPE1SpEcbHFGVND3krGCRmhPUvts
rggAMikLV63PuV3FAN4A20KZktVxXmau0ChwBiy31DxbscVLfwQ2LCLecDBYLNiz
U33PFTKTSNqxp3Uk+7yyqoBWj9wRCIx56wL5SWl1NNgbulyKJR8Cy8novm5sa41f
lIb0uUaX67SlMR1gFO9qoHxlbBOWmPh0tJB/pidD6i+wbN6680qHGQZtvh8Ffv77
1lECkL8G+eLnLKrl3z9AlnlvP3N9SkJkmCXekcunTNxr11+K5OhG2esp9kqhfMr4
rfhfNtF2UYkjer0RlNLtCxOPa5wzs2IFzkXDQWvuBJLDWFrw6mzrl5IUaOZkGU3J
Ddvb1C64GBnkQrwKaFItk2OQm01IVXg3vTjTW+cnAor3pd645hSlTFjur06s85Hi
xfEcOYnPhejZi+CARZMzOZ9of0nH5OpM8DQl3aceDqJVvIpK9WXrgSIQlHTGKsfD
7n6SJawxAy+EKSPPRCqNDYnDhp8vOB72rOLEQ03DNSnrFhszLhG5GpdgWVppflH6
18039oaIEtkH7612oKkhjGOgllVHkp5+RjjKWrqszrDddNdYBdA9GNAfeqEPDQN/
ic/fBKGQEh23DkMYNVm25jkdPNjsB/n7ikejne19lu9L6k4yaq+Wj1zkQcrK8OKt
ENcoOt0/9lrybp+zX9VYxPaIhhNlqKaiQa8yBoDzJhY0w5SuUoSn7Qi9YBWv3F+v
q7JusaJasxLrBdnmwHRdt/As41FZrW3hnveVPU4xb/TAnfnkZaAbt+2CtCr6dy/Q
1tE8dGXZQmpPPZPmjFSZhHHcoTFrIBx9OMGKhHqpJy89Jg1zWBd5/OlzjF/SfMi2
JenHn5Ox7GRl4PwACZvDJzUuPk68jTEg0JcBFPXOylCP9pWSnXFhF9hLetLUSabr
qyMX0Ykos/ayqxdCDl6qmdB9arYkGy799DzrXGow8Sgg/AzoXLMdGMcYs4JgSJWM
i+PuFr/spcmn3WXC6AEKU0R4E1bYWerkfH5pH12qrZngi1KpkE+RERIRdI99kxZ6
0wEkEhr1uixuzaHiL5qsyB5Whx39hWqLL0Pm8+7iSbswQ/OVBxtITQxfE6zenJXS
XigYaz55jqRbh2P8ui1f3Hm+2L3Gie2GdR+NFlPDvXKQxl1YIfJdiDi/br9pKjdk
NV0m+/sx+VA/Upg7C7rF2AmG/TrlsDunTDEUiG9t3DaS4NyX2feOQl9gn5OuJ2BE
YyySF3+JN2C1U4z1F/mAeA0d/jnOgkT9stPRiJc7asld3/OWiz8pwUJ0qxCOGD5A
UbFETjrCNZQknmGnaLnAC822kXFX9dtOvlhy10UvFlyJK1MH6RfnI76mf7tyQiJq
rmRtUSfJwCE/PEdB3uEntdbftkTNYV96yYLNPMMqzTjuyLI4JbsRLpEjpTmIyE6d
zpNp7nINLafjS3CXArxCs/g7i0UUDJUR0W2uANCceuJw9SWcQhMxgUy+zJXdop7W
gwGvtSjqZ+EaL86aWBsQ+tVfLzeyXT73vnwc42H4EzEdz00Kuh9pdz4fwLe0r8zX
7OuxOsTv2tgYNZn7sXJKouqFM1zzHiplC9dh203uFH906NDtJcNgKfxfkJwjaYun
s4zMXsIMO3VFkeOv8dIZnd/l0eemcovpoYlE3ykT4Xdd4GE96MntX1UzsTnsH4Ic
boXI0anqizf6PfYJwp7UXs9ehFLgOg2+SR1qx+AltKW8aWMrOcVBW2yHIFrrc3w9
bsP6txI9RmEcv57+LI6nJVzRCDPdxqIhbPktwwXmWsV3L642IHlRlv8guNBnZxe2
GzyNLuxzY4s6zQjtWMDQpTyuFwpzwFYXIUkP7Ip/b/dwnJ7NCNOs3Ky68zQrgjp3
g06DJeS+DrMwidEDGMlW20KZpZtggJno+hHFJQoMD09pDdnOCa3MsSRyZXwGNNlC
OJJVr0E7TMmmtrHF8Dznh7iSqGQwGc7axc3eE9d/7V+XyEdr31LKZ/LmZWm0wYd6
fYododhCPCvdGg/hzB5yUE0bX5uYkQav7NX9bX+BWN4xm0NxMcUm9kDKnyx2v4UT
tR4z8SDi4ksVnrZ2tVNfZUytWNSz/qrMbES1UkfNrkyPR677B0TuXHRudNE6BaKm
udqfOKda1wfvS2WitfLdQv0qTurDwh9fsIqg6c8lSLrIUbvoCOwlt5Kl7lLui+s1
1XSB448cNvgwudOVdlEbC8PAxrWTnW7Gkn9S+DtjaXn0foDDhFwyR/koWvVgatY7
RKEUEHBhSoAMWRxcfGY582CNHItaq+ZU43VSUPLiXsIVY0c+je+SXJO1tjhaQUiH
qzEyi0wcxgVVg41WB44SiTKdFTSDQGFb+Jb82L491U0KqBNMlD1pnUnChrCtKefM
6rlZFGQQqK1LQ4ttvsanNoP95SzWZ90PQBGomH6PCoCMf9XkZx548zDGSRYs+8T0
MydBYLSsbvOyVJqJIwG7+ZqzHz5mFzc2oTDV2c8mxmjS37u7RKEC0fU0V7z9ibuF
hFJioE1SsJARrBdQzlqJwSzsRfnD8mtBABMZ7OKtsPh80OsmJ5WiESlGWzMBNHD9
dRfgGWRWfuiVbJCng1f8eNojyeHZkPdetWG73mHoAv4MvB1LZpbf6ekXDwKJIsH5
5/5VoKT+d1fe96+MnLPbgszXvbVO6Jipm83CJru4iW87MGkmNoDrC1SWiAay18CC
vpCsHMLF5NshuhZx1/bKnX2vD4NcxQ9O5Cfsrsa8kdYYE4Hm06/2hKs60R0xhafu
Idnbo3XtsWuvY4rEv3+7JvkxbEozBX+f+lfCf8wlRI59AD3ynkva6Ozi1vFL+XSJ
jkd3cTOWBS/e8SoE+979A0XWkpOawnDErnrdsQQME+BwTr1mdSMvpOochBIaYBgw
N0IsqQE6j7AIPmEdUN88c2A4luyCm+ljXuQYC80vBDwldRf8cak+XVMlmr4+e7ot
x4LMGXzRiUNnVV4mKtQXOFjRryEG8M436Q7F7UOKPrW2GA4aAWsqgfn4gFYIbx1t
xWYyuIAXfJ5TDISDRAmUFZ4F4FlEzCDUysKEloXkl7nyIbDoKLsUBurQ5SdwymJz
Qcv/Z4CNokvEQtBgej+QrGVJ8wV0QbBoY2IxZydcFCZEyqXrJ7Lcss5tfPfAT6Tr
9cpXVculZj7UglrrfIjnvf7VPaxdS9DhDYHWAantR/vLkto7FHEKD/PkPF0cXNBy
0j4kimQBuobxv36d57JZ8mJ82ulMl0qg+lTrwEP76kLtRSwHYPBvuCf8i6WoN3my
ab1iWflv+xa3Kzm0s9bRddSmFKqgHqUg0XmCTtBUXnWdcrd1N6ji9EnFU8G0ovzD
GBK3I8yKpM5g2cnjTS4dDlYMogpEOxIIcvmSapD1DUivrAsV0kgEyeSS0oUoD+PB
eR5MagOK2PPkuvBy8FFSb4+nPwhE8GlYu6gmjsajKrey2rJTditYphQJ2p+4l9Tr
EQBTtKmTia97bKzlZi4i96KEr7jB7IDlp9yN6kDZhVgA0n2Ft2ZtSsQzL9vLFJc7
PdzRPwmmto8hRef1t0iXHq8wrqNu5tcsXBq8WrBKGvf43eHUvS2ber8mkLnK3wM/
yvQ1xLkRLNL9bP9rZAFpuci+dZJB90yCd3P/9KSIyX7r6GRvK7rODm2lnkj+1bMY
HIlv+JKiUrFXjgLkpQEogNrsC5eu6n7c1S6PMFGCCS+Uu+WPtJD1qvF8M3vQdjfu
1a+AAp+x1yjDaUwJRSS8hH2PYtBBuszWoP6gZyvjSGcbakFLGAN4KVw/qCfJo9VS
unPqVTugJqRxZIx76jQhB3F2NEMU4f3RzDyYtnjw6l27fHba0K18PLZ4g+WE0LAc
3LokkTPJLTphATDnmWVdknpwCesGPm90XRwbKJe2lXrRCX0bHBEaMVMJPU14IvpJ
6fht0md99NELH7Wp7pj3WhB4zR1zMCTvHU+PxhSZP9ukr2tJeGDUAWK7QzIp7lNf
HIO1EYyJNrJ2vubR2o4Y5s/CFe/+JSALMVpvU5lX5lPMTYAhc9Kf2WXEInC3Ko8o
783I7uwPoZkHTNbqpmNFNaJbJcCKN0Ydq9I5VxEpYmd1BNBWIDq1gCmYFwJL0T0D
mZ0QPxUHcnq3DLe2TmS7kjT3I9WPOxteJ2vpcWLa/xYuiu2B1IZxHf0sfN/lCaYM
PSPd7nBOWHLw8XYwtJG4ch0wL6CAPNe7UlBmMA0fxBTOSS8WT4oLxuGvE0zTViXF
QGTtxPT8legRMaEsA08YkgQ53Syp17wXqfxNiG43BCfEaYmk69c1WZIUW22fy3yN
TimoBKRkdtgzl5O/Um4XZivQhvDMYQ8wdP9mpBwRi7xjC49+FVd2SOWocdK/V69z
w+tN7g7vp8y65KEuCuo2D0c6GeIMi3Xv/t6VpS1na1PpzPI/LmzaCDD5Ae7eKqBH
8U8HefyqJFSNLqK3UugrHQpGMFmOqKFSW9P/LnYhp+jKPeivcb8QcHLtZw3BxSW3
0RUpN0CGsukZSkUVuqpjxGXno82doOi77p7xFJL5Th+ZMEFgwgshbs3CzSlYaVGT
3vUvqxIG+3I3TKnUi75/kKCOSwv+Ifh5iaLdvewZjAs0W4T92h/23UvxBhHn7N85
F8ni5LcKNcF6GgeIndo8ASPPMZSOZxLAbpemPEfwV83EhXhyn5HkTNKeTIxgZ9kx
dxT4tmLmF8LIpX3plxX1Cd5D1lOc7oKNtL6QVXN7rLFaf4fWMutNfVcHyJ1Zj23h
EvozXWmC7YxPUuN4SboXRelHTha+BuTz3Ljjz0d6zmig6ZiSFZqIlzs77NMIont4
J06iTnTFYhKDobCx/s9x0sOO+4xFmi04OCkdCeRg15zFZTTMuYtniT2RZ37iedq/
a5gOSpmCA2V/jF10AYLq4mgCdJeNOolSfd8OFClVPdhQ4v7Z8gqzyBhtXkoXkS5R
YK1GSN15FCSRkkGMzhUGznJJUKqNJoSVvEDlfWb6CKCCb+4TV2yzLSdqVWDKAZuy
Fkzua/r9e73DCFYOX0HvXXBBlEsaO/s6IDdYbsIv4nYV3E7nbIIJ8FAKv3IDba16
2yPYybktBXpbDY6qOeQJ38ithJ/xx60g5CssDunb0Z5Za3A83uUznSmC+EIIq3hN
WWJC3bztEyrRhq3ADCLr1IfMaXh1SNp9LMC0gQdDbmcS7UmqkjXS0+s5VWKiDqQb
vZZxe7EsRKrDNYyESTYFu+BADEiJgtfwDWJdwTJS4vlRy8f22coXHK0WySEQDWHN
b/xUSW7hYaXChhgPNSEmPDBDML4KoJlwMhRL/LuNmn3JvRNH6D2abMZKHJEYtrBE
ImnwW8/vLaVWQZIwoTMCERgCTlGl7POFaMmBUrFC0OXliYHED4I73bWBBvMCtefB
VV1qQabUj8SUoKxxvXJYJLGgRBacYVV3JkzEs+j46SzJ9/690LwSNQpDQMOClJEZ
jrFpGYmG50MNbAnGRJQdegL3UYVbS6qCODVCPKdlW9LnrQ7WYg3axC8CDBW4PHGq
Ggd1e1/8eh7M1fOCs1p4paVkYAI1SAfJVYEJmGlIfAck3QZ8IJAr3MshBklybS17
ENqA2ozKRQLxr/UgCnuQcEu8/6eCxqT2Z3pzaudBXAird65Wb+2gYWcbrtOiEt0Y
Ee+IQ3AOqg7X7/r81yYJQ2w7CPxHsvDybJJBn7rPdY3evxuCD+zgcmg1NBtyz3W9
h3Wwmpsj5Em0s3w7Uu6BosWyYG6JQd63kGG78+3qKVnteGny35BxAQ9P4euHZZPh
djD/FsxPDPdVsLD6lSkSbqhRntp3boQ/JOOqMQuDpgA+hs0a3+xdMFpvwiZDInBi
w913HcMbqfiEmTTojkzce91KbO9E/g2N+ZQhPzpyoUoidZd/yVdw83nPWps8IjFl
OaxEpeDnqSg2Hhnpw+dLZRzlF4fWDonVF3OkAv9+GpirDlZEg0X/YUAaAWocRtdG
iHE+uO1t5cQOaPqo7CqoW6HUTB56esoHlGnfsFcyagw1o7ti7rhcbvmc6Uz2iejN
RTOLny5ti0UYpGdVBsPk5OU3NYSJMyQTF8Y4fSw/srzaVG9vlyyMeCZWBTXQnYxY
+1EIQ5HqKbscHPwF0GUm0UokwvO5Pi95vvzR9SlBtT+AOZa7xkDE9CHfd0ACAzk8
HdnS6NRkRJj28b+apPB4zXW/3eFZcXqTkwItyGvQPhsEEQwmVJHsMEKMnUyEuOEV
DdPE4hj74ZZfQRnzRe8G2LvrsAkwht/SUcn8Sf+IVzg8U68r2DkP2ij3GQ2kE58K
2/65an74bhjHsYG3dxAlLTwkC0//Llzo9hDGo9BC1RF+ooIfykEI9UVLa8Q1+chD
7kPDe4meASxAK23ai4+8TDkl0q6qSedL0DZlxlQ4N7mu6BvoceFqruFzKbH3eNDs
k7DMLUg9SgJMoYJ3NO4kBgDk2kY3cOManvQDOd64sh+lqn7J+2VwgoqruWiDREl9
sFsnTOd7MiIRHt4JwIoR5noVRrmqBAaytPcbn+z6CD2nbGYPK4+NdGIvFgSKDxeM
6Ve2MjHisenaEED0sKT62fwsJyL3zOAMgBfnyYfUYngJBkK4FqnmoGtSbO9C7VzH
exajQQWtYKrrEd8Rz8L9tUO3Fkr5ZYBjfsCABL2wuqu35XVa+UC/ojm4RFzcWC4q
A/JZ5+Dmn3RlOeFZ99JbPR/KqHGOmZyEuJ9USmGo5W7WIp3cgdU54c6ud23hvj9q
oTtX19ilI5bSEO8l/QLP6196bOS4syPafqBNYaphetvE+1Rq0odCXnlOTqhL+O0f
bpV7VVrRn4EWbIM0WDPy6n1ALylcmm/eGJUjIZviTZjTl0Qi7LZvZz6td1Gm8IYX
MFKGmyCcgI9zl3Ds4VDkTrnSJhJc8DZZhRNrR+EdMLkaJW2swo5/Ecj+yryisCZs
o4UsU99FNMYHIq6G0Xoclex2/ezTQZnPx973Z+fjUoNJVl0AdBZFblo4DAnxWsy/
6JmTsG6iGig81aMTqIj02/E150iGqO9gDhrWVI3+a0MgH0UWognR9g79G4BxsRRI
JFFFB2puNmGNlbGDEc/QQy5i8hl/QkF9wTm7LmDvD/f1co+/RkQQGhZdSIzFZHYf
zW5y4R/8+Xr1J63JLK2rqFWGNmfj2pyMHH6YEwL/DoxrnHvUZBwkiAdtsXj/1UAD
15pQsVzCvxOCwWEicWIc53cR7jvWXL06hmEM7H+dudWTKFpXjy1FuqxVJXvQHjga
4/SAtfKggLkurTwmF2LZ9G+0XeLK0+1Ry8CTkgBvq7Rr9Fc4KLgLR7iUVRj0YDPq
178JGYA3wZONMWk3UKkbxDI1PbThQ18FbQA4LbO22fE3TAtwOPvsAiIc1nPFCVl9
pzYF+E5ojDpY+xG9b3sJiX2SRVqE574VcYJCd0vWVG3WF3BezrgdFHhd6CNyyTyg
9Uusx6uCrnWpzxJ0x5fwlgQx0k4bkeIF2NowvSaaWQdabrPKC/ME3OLuKIPIrpDm
JF+ROqnzxQDw5eC1aceDj0POfrF+f4W6Bg4vYSx6t6yjpLbSIhV/7hu6vvV1ked+
rcyXlg6JMVmdTorozIdk+4sU/lIy78ZIiGgXflMDMhESbpTriXtYN65dUg9fFmZ2
SOAFUWHSaP2aeMq2fzNsyEvmMa8KVCEW+Fc5JcgGBWUm5sJ5Mb776jO0WAueXJGP
YCedHpvFfyPiRpa56JQIlWcqmmvWKxbrM11iA7oSuYJaYosTK5cHiWQYXRLWFSak
vSY8DVCH8RfFf/IUnU2MQNIKJiOVXCGMozzOBoh3VJP1DKfJMrayz9D6TrLmcYrw
fKTJuDLHXSkyIotLTp/YDDMU/aZ+0n8QFkFRP67cccuAm1w6NtuI0TBO4WuvsB5+
SsjgQkf9LZE9SHNwAdPCv0o37YECaWz/XqiTZ3t0zdetzm9K6M1FLUpQXnJdUN3W
z1hcSyhVOpsyWCwideskEoimEDIDLHwArMjkhIGt0+z5jnPPREGUnzVmk7xc3Zo4
YWP5tUPxuhid+aJt3cpk9nq+ts5x3vKzMCaI2g31JHfOs7CVJG5w8jAVXvqUrHSf
kRS4v9nCMfcsg/qHKkymnOt6UlBqo+4sNBppVGiBP0HxOh7EhYG2RBy23jkQZJEw
qyKCf9PD2KEW8NaKi/PYebyiXmEMApVYy+UoIzOjZJFHo4Ih+pfcbJztqqEkj2aK
jgzwbvxW1KmopwAbAmz5txCenrhnqPCeGk/e6oLWqypNcHRYBc7xvXqvJADNkzOl
VoXkHOp3NzPJl42I431/mo7X0OMTdo76fioMm7RdEGeRTG6VNjWPkHyiTL2CMW96
7DkSFaWGKF93OCvk5Kjj0CWvDFkrjtYH/3bL/FvulzCWt0iYgVpSVullNPytpQS/
WKLkSQgk49tq3aMnWTFhZkAYNWGySKDi8PRM/eQMDCiMhItqOrCwdJNgsyDlDK5L
9kwiS3sWbUyswbKKSpev9gnztF28taz01tRLTlo3RHmUACkPDQtJjE7s0SPvlqQC
CMBZI4xW6yThGnpgcTkdHN6wXjnnb0R+JT8likiUCMxDbbbDZjtVwpSKaMuSzeev
YmLTOlCjjKgsm3Y3+oAp3kbVir6u2tzUv5rPa71zs7HjF/miJdh5Q80JqKDVEO/l
m0CogSlb6BLXjZYNiStpI/exAiR6Ay8ozrDQ4eZWiYwfEkGVes2pB5DCOm0Ze4su
DTkU91a6auspQG/PdlrR0neiZr8LAboBuf/dTSpQwdBsLQ+CHTUi9Vf+4YjYLZR1
9cg5KYXOTPd15HsiNRTeEGhpgxhuIWwtDrypnoxyXzA=
`pragma protect end_protected
