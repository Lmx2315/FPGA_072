// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:32:41 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
p0rylxAvM5gyWh4uKHCHB0fA+32M0u3StJhkkSoOy3PhvaEDpKad+lfW6BUtR2a6
9Lc2hf/Au7lOJfvc/ENmFT9Nt/2ENj58dwn6tiiG+1A65Zo2EaijS/rQkGaUSvEk
qlDb+VUPyk6/zuoSxZq92ZaxjYnIuT62lsKQOCPSUCg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2352)
QT9y7a93AhGm9rT+p/G5DnpkbPUCDdAYOFXs00nUs6ey03lFr9yp180enRhWMUsk
VTmrV+g3qG2M8/jS4374ktNTZuV1aSbkueO0J6l0Z0J87u5JZS9x+Dd3atzd5ab3
JarypFgWviw+w5RDUEf1dtyl3an8kUgoLKz+iRTb6LDv2GD+IM8GralzXUH6glCx
eu1nG/znirV3qk7wYzPeYeWL8Dqt8PxUskeVad5mVrYJaqmZ5aaBV7mtB38nVHrA
BBtjIDNwWyKVKm9yuy+XEpk2cjWgYP8Si7b6jw5vWF6tgR5fqIo2cYcVXv0nbK/E
9LLMfKdV9Yt1tJFBNusYBPu6IpVqitYx3aXyDH3RMoPmLbUtHJPc5IsoxV7VgtuE
+Y5f7UShpaCg6VKbrX3ZaK4wNmxmz5NnbiVOghXrux1SZNLAF5kA5pUfRbHMjOeV
TdLuzpiVZzkUoqf6AZuk5m2SB97btAs322/S4qwtTv9793aSG3UBKkjhXWckdhIC
FBMGQCrDfH3M4XrcKXCIJPGh9uEMeP18dVETHlJeV0llcyjXMjQtzrIxg1RBsp8z
xvQCg+mEmkG9CREmQ1WWl3jidbh6DofmkLZHkuApXewK9UrZcwrMbjIttGAjJcy8
mpnN9jTjSw/+PwaJAFrCsbxE5G5xU5D55Ad6oztw7az1Y3mH43QK7cVFzryS/gGH
NAoeGJuibHt7lInSuyV4A2Vxcz1YVDX/jWMk8USuE0ekPx7HyyDuj8FHWy6KNa90
SNN/KnrFUfHgwKUy7uB5+yYS4FJpaq4ZR9q7ry6yiYMjy5qlsvOLd8DdvxpfPbSJ
ywvRCwLSRPQFpGnjvKtzXmCvE94FTknpZqdmSF2Mikw5/juJtml0pfFjMyR+9fg9
7n3DqG0aocrq2vek0EEZOBVdLRcVPBW27ESY7wGrvKLXUcbX5ALwdHu5KciRrGBS
SPlbW8VbEi0LmVfVjjEtJ7LHl2FORSEXvn+31qpquQYoytaeSahhb2y1hOf45EeZ
ZP+g7rQQzNdIpL7hVKd3qP+gqIzutVscP4fFrXyEzKbzXYSJZIz2LR2mj6xdFTjG
LsTD6I6wkl4/vtayp1Sg8roJ3BXXrkaLkzCC9hqpcgQ19cQGrSjSRRDw6qQ+qF5T
bY374Kb2nrY6SJkq8KeaaWajv4xXxzwOwZM5NpgguPUc/TcElC9EmO+vjlqcFREA
pnY6BkwHg5JPmPTGl9xtNqXMDc263DnjnxOyopRJXyd3z1G4R0oxWYK9AHd9k49L
FVo5SGJKaZp/N7TNPA1Ftm18KkXXVTuSeCzNyezyitAEoV3UfeDq70ZtPS6bfdgM
bXlb3KdXzBGwNkOVxR8yN27nApQeWyFjtIjm5xMxz5MgjKYxQGjLC/sp7rZWaO/k
KdgFOfzI27IkHXP2bwS/2dZVtUofMIsZsdNolS9+dGa8t8OGQkoNDGyPnoMIEbXS
8p7r63rR2QviWlq5O8g4jjyCYhlFl/KnrkMxeIqgkqzYrncHq0Avhc6ixZbT2EhJ
HD8pVVDC1y8O2YmaQXN7W9StZ3Zmt+ruOkarllBfV0j68j2szsb5YgBDt0P1NATi
iF8GqDyQPAwARDqsQeUWU4oGA0EDJgEHxtIate/3oMXG55zmBAIcKO0jK0goblIk
d9F2Rp7swbJJuBG3WO9OsBwJ1L3nrbk5eBl+ri4V3J80xq265mCC40TzbeeS6XBb
EyGZk2uXEvjUuTW74vYHrJXrseYOtfQJ4tY9DEcb7IkoZgtFmqygxL7fhzSNuQB0
6/+QsSAySfGN+6lXuyjc7RV+jBS3mAGP6pbxoRG2avr6C0KMvVOfIeXKNIidKZcE
RrUBxcNBYdlImzJWnlqYWnfu9w3e77L7C/X47Lt9VYRZ1EYfzPr7qbIAZjBymd0E
4AwnL0D5Cjjj90Oj+2myX9429wZHjvzZB7ekuLnIyrcBypMDbejBDoQKBnVvQ8zy
WYfDIODvTTspPP0pfJmaw8sjs4OUkDjWSmuQ8NuSPU5XqRAl7N5732su/6wEeIaH
qnGDXxK/+X28i1qUd8swpFVhxTooORRb2XcKEYuvzldxg/I8MIwSyDPuJbOmMkQS
gerMzeqvXogM5/B8qxG/r8mD+fD0spM2YZGs4JwRVGy3ZBu6eXDv1C8SYnYjl6q4
iJPMjpV5hYG7gzyAp+Kft34X1DVYvbAYd1RMz2Tf5xKtehNiET3n8ICMcVBFML0Z
qEVztaC/JEdgSmG8bVz/xzPm2BdT80NrMh/zDBvoB25bcvkqtYhAX/ItovhQfJ6y
HjkB0XwLPGXxZwYOEzKjS5ZSZTfkFABaq+L9submG0YyrDAE8pnhzJYtNjUcrEaY
Jl485+m0D4o8AmzpJY/MrzsUk6ClErda4YMtj6aB8w5vC3WXxNdVELcxtIAysY0+
n8ycILEN0zzM6u4YdNmHADsU0+s5L88mspUUQcCZhy/zSmTGD4Z/pvzmOk1jbFkI
li8yjKew3pfmKmlVveSr8qZ5FYPjBzAPeXJnWiadKcFAmrjBOtGKF0Nqw5jBRIh+
qcbfC/WMV0qkiZ6Y7aNe8m/Tuxf5/4jnnXVS3q1NqAVxP25PUfX3siDv/H/d/J4B
EgdN7fvS6xSvw2FYVz9VNv1a7ryvwCvz2H/1lT2yWVDkb5IrlN7rOgB07fOxE7Dx
SgUPuWpvb4y6mU+fmVOPp1GidUFVG5ZZosEuzHfOlPcValPJE4Pw7v705y0hj0ym
m6llQJTfNVCn0rrTSMJvwdkGTz4k/A0cBiEOTW6v8c8c787CM4KewYKmuTJoMhMm
Q1zHu49PFaQyBC7n9g6eQ4FbM/AuUqANA/1Cf86am4u100FCdu9tDliboYFB6ZRu
vUaGkZf/twe+KYeRJHN9lnuaroxM7C1Os7j1vl/e0cmNIrayszpWXAb5rtU57xu5
9bjIsUu45nv2bBB4LcDMUXUdz7hPF+/L3OevOVe30iANqdScWcawynRr55I8WpVq
1EGRpKuvt6Q4v8U28yuYewNrJlOaNq3/huTZaGOtiIkHRRm2G23wS3mhqj8qmZm9
pQ6eW/hA6/x5DjKuY+uHHe21IxKEK4mHcRQxtB1MZXjKEAbbjTIuccUMSBNXKuiq
`pragma protect end_protected
