// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:36:51 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
fLUEKY9LnEygYj8+IsiLLHgJMP7VbpFbS0mnGi+VDMDJxdq1MkUl7KrMwdX5upOE
NHbB/If/tQ4xd7Nbsh6ndXDfUm1sSRyxo26lMd3Q2LX015V65GQvM0TvKYygjVTW
snlPH6I36iYtolkljZ7N96KYKoTExuusX60UVJ5UGto=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 22608)
HA9MD29e/8pBM+adF1HIRZl2LwEiqYTFYHzA6nv20iiXZF9xcxo1iUQ05k2VZHfC
huU21V+j4iv5vrD8WSeV8zewZYOi5vWMhIVR2JaWYpbSffDg4Y9FbJM64jsnNrGD
wcp3JUc6Kg+THKIJi7txQCmNeYGczU1lcizfEXNOdiHmwohyvGBhd/rL1ExHTdrB
wb9pCru1JBNw64eaBHwmaPSBEZgKUx25jg/9M/lgEIP1fRfUYNOA4XiQqiRoVfQf
Hm5F+ayGaSzYjbZ/O34UOnsvUVJgJ7ekAxn69joYdJgnIN+7chE0LlSv1UGEMViC
JpWxaKA3yGu85jwoyeU5wQYV+vK8vrJNaZRoG9o01PvC+2FT9SUbnGkz2DdPMoAA
SKZhvMKcNHEsdNUrRDXGzUI3R70ekplMAr3Smicg+ePwGWx0R62NbIAIrCnYIbNH
Z7jL8P18MqmMMqZ0Ejv+uwCsbcszNU1rCZ1M5urxVNHasTq68N19cCZpp/EP5o1s
hJhjh9GhDDPu10toDyNPf0qgdkGfgS0ht1AVdoCqg6AALtaJ7azFBa5bM9oR5E7N
OOUniPciBA939GSc5QWYEjcUOYU32zvVWeFK+uIhMol+plhi5T2CEIofyKD0CVEN
x+JvAW7yIsq8/fnFID142BO84rK4YD35dpyo07HndvzfU8vPnjpHLF1fWXt+TyLf
gnbFJ5pYXqO7NtJ6H5mRnjaXo+L3g/2w/wBk6MW76hdduXxFtw/s1DopezdQvX+F
kLQnD0CFrGbwjwZVt/qkfN9F2BpncreAu9pvSawjwx8MDTHweyG2rhoLgfvSz4W6
lFmRnxFkV9TgiN4ixyDHjgsXLLANe+qvhDGGQcjXSqu6BWvuJexDEwWK/GqbN0V1
FMWDnSE1tA+sYgLRSdFB/6Xlji++3ILfe1PGL/GrdGJEgjSAGKXDl04pWQKI+0se
hhvA2gCyyVJsQG0vTUxG2am8ddY/HJFp+/9147p6GnPEQBgYt1mLG23RmGByYHxu
585ZERtuv25pNqVhsd6/XPb9goInW6NkGWETtjzS04IkBOItrPoAo5quaG0cIpUe
20Wy5etis9QghjzrXOmSSGimPSgSLJuBUv309nT13xHg253hVSnDMS6cs1NQCXDv
EnU2WfERDDddHOOe5e1dhK+daoMGjm5foBQCj8+Cd/49aMU+I5cbcOSrQGBes0el
gH/V/Stw9RmSSzpVncDLR4X4+eIR+5dPKq4DWI1dbGrB6Fk694nztxA/708jf55E
OJhGn2a0LwocynANDKcqjtNEvlrPhKhQgkvum9aQm7EOUCN9VPq+pF0WcQfzT6qc
sOSN8t3Ciuy05p1uI4ZxXxwKT5kdTCEUBrCw0RLI5Ic4lhqd0QeGeafn/vNtH22x
wKh7kwe10v7U40nld26yAp8nZcS7+cjxPcDkDe5Ky8OsR+kyYUTKRdLPH+Majftl
1vWZZQxw0SNGD28P/b9lwd61knwngexQldZc7v/MefFnFKchJOrIGsA24D0CAJ2A
4+hftSM9fY2tZmiEqHCD76GSrzEeTVJim32+mYNcy9vXAADeosM0xd/h16dBdvJy
OOVO1I+DRllzyOSiZTsWGzqJK0JQuKXdXBIYX1Uw7PZUSyQ9uPnHIM+w+8OFO/bt
VrAJ0sZILG67ge7YrjVZHSWT+2oRQMto3XEHYkOZhr/nuNjHwwWiEFKo14uNHmcS
6UQwrtcz75kNuwQWIyqQOeLCzioP6C/wQgoiGVGHdFIpC1P5BKYh9fZJVS1Reck0
PaqzhZ6qLGEl7Z6k8tmdNs5LiI7MaZjLRc6saxLeHPFZDf4QBUTfwQYoEHPvFKL/
NQm2lkZPeMItfjyXGj5nUhPFvcDcWY9kAf2al31RckblHDTvar+Ot6Czb/TJlpBv
yhO7nOghopbg0oQ4hgEM/u5wQtCrrqJMkTREvh295mEMfTdnhAwL9L/lMq6XnGYz
vhHBTawqEr17U9rEzZwET8tLojCkSOMTyyovfnSkhBkVSmz9xcOAfbvuHpyGwi4k
GekZxt5If2/aalvG6k2ADXMcfhUf/15EcJoYMxQq0COCdt3A+lw1qdpkRSfXVt0j
pfi11AcBstsNiSA3kFdJkk59Al7FO/Kaay6g80GQ4Za8PuEqCxgL7cJxmk+0Z3Vr
RaULEEA+FIgUL3/A+KtEyM82FdBYCYyNRgkJLriJvAYmrWPd+JAnh1DGBY5TJvpb
UJmlTqOTH4/3gPCLcO6ajx9HFG/hs8G35KjQuAeckcalL3CYccCv5F3dgFa9Lzwl
mcaoGCvNyXaagNuuO5ScRYjC3ec9H4JLkXI9lADhVI3N/d2ZM4BtfRXjbEYhLZnZ
7ewQMgbimMpP83Bqso8+HM72EMdvNOmgI91RWar+O4lfe4QWvo4KD6s5npJtF58B
pL99G97x5qQQ22T6IDm0rhy3eGnQbYm322uuMUE93tOF5zLedwnB4g4Fb0WcxNe5
LttFNZJdOuAVwc9LjcCn+Pg+TgUoMBLLVVWWEOHulfVXX0PZzfM2dd2H5pZlqFHd
KUQzcrYwV1f+k+BzrLN0NkZdWNUT0crt8fO67o8LVTo2BQIrykda8HxKkyUTb2sf
xws+bfG2xYvvWkUCfVp2u2zWwAJZCCvnaT2noURSPK9PkKCDSvhi/R9FDWUI+uQR
mm8FkNoBU576MG/do5AzoYgImidd34GLwXqMzlxOLb0SfmnwrsFc5rE1nWMNdujG
F6bQMrFx5X8BhGcHZuIVNloQjW1T86moYnqVl/gZZPb6bDF3l973hLytnVisn2zg
op1+MdmPoVfQbD7gtA/m5tPjUxbn+gYteZufLURBKKpCWTiL/fUw9bBaA9oHocto
BKFEToaCgGLX4blzt63qM8q2EEEBIakgNOGtFkmYbwq+C3WwW7mB4CqG7g4QdvL7
/jY3d/gHw8FWgO/82rtUiHiZYsVkkLKqHsq8vST7w/Yo370qVvEZl4hMkCOLSTqH
JXHkVPybtZdruprx3mbbOkAHLbL3n/Wew7XsAIwNx7OiIQ5wZRk0UNDBypkm5c7/
8urlsAhOZ5mbL6PSP0AwclQgOohyoe78xafeizwU6F73dXQgKAywRZt2l/XPL3bt
mrYRiSNVdHrZkckBldUGOb15FMvuKGq3h3CSub6Tz0A00mh+B2O9XD6N+TvPqVTg
IiE9KsO/OkmEO/2PibVifQnURwsOivEwNzKqkm/mRXBmuBj1dt+/2eOMMD9glG22
GdUBMfrH4D6no30couMs8eMYg37Z6BWOhcLvcSoPj8ZhxnFKqQc3tRoe6KvxdaOc
0y9lSjJxd37f5NbOCTsGq+YzVl/meR2oeVtn6VNiyUf+CnbXa16/fGn3NU/gfUOM
fawxMSa1Jh/GSZde+zAl/DRPxXMLfAbLG4kh6UTnSwcRIcpdk0YgnJkrkzEdkq9q
zVzEJgnYCd8oB9mBl1vUBF1Y0AMHZ+JvYkaX9mJPV0NdStUCtxXjo+9LoNPYmzBH
0zMjfZjpFdMfJlJLUaHOpKNY+54g3P/LifiKhhdzaJGhHzprS9TM2HA6XTdAazOM
qYxRtCgQxjkzLswDrjJnxb5vv2XW43yTDUw/P+LcOLbTOQUriLaUnqG+ps4iaMc8
yRZUvJTN4U8bBDQz+cA+pAPzPM96K6Ek8vM+4XjR/m2ETdO73wVKmq5lKvkD4Xf/
G4jrB2RruMG5t+3ULIqgJXeO1z2i8pG3VWZMbsGVmY0z5rzhEholAqNqCUXqjpR5
LzD2MObkRBgfxngzyI4eYSNH2GbsGQNg9gHH7e/FILjyfJkP6FOy3ah49+hUOq0b
vb2zJafgo098MbUxPaHz7WTTWcfDn/Z94KklokNFICoazs6u47ghXVOLSvDhCvTL
a8GedSYJAMJZwW/Iui00dNNaLLy4/O3K55owxdOh5YUjrxHFBu+goMv94X4UHbXy
6TRkK35iBh8ywXEy0aECS9MOgqstzjd+nV66HVsB/8gYlQMIELcXsar6z6s3bPlD
lqchuT+ryrFb7A+IvWrHepElEaR/hHLkN9DLQWk+9MM7tEZNtxM4q0Atar2AzAYz
4oVPqoBvnpLDYjGJloYFP/veNoR2zqTb7AWxlDFwRsu90VRVaXj5YifUlJO5c4Qa
1old04XPp8AnNfzZkdSo775k8xRYyNmv5FvJpNeRDFdp2S4iMhDBlo79z4tHCISr
07yqrIi+jb3BmUNAheL10dGezq36GSKbQ6dAeULN1cvINxwr2C7J31if5xwLVeAd
k4w9wFvzqA+YlpXLZVbHX3sXVXFXL/w65deOrXfdG3cLYi8OjhN93lf8yenlDyi6
BrGRccowUN3NivgbYBMuIQ07ppRyjPw8eTY4CvHA7OfqOk77q/Gt6gEQdNAyX2Dg
dakpO9PoPnZzMQ2CdQ2t/erTEsag1wXIE/vzLO8gedCPpV2kpAc8Db9dEM9bYJMz
vZEgTzwUmzH//q4e1fro0TtXIzyajGGOuy2NHuySpWNKd/M4ILwn6IVyLpjrRZTp
gJOGI6oPyF1chkgHm95qt22SuFQQBvcubJnCtIAhaNUvehpkZ/w17df+mkvx+SaR
hX+x8+CI/s9Vct1znMIzM+Tb+aBH5gb6oa3qMRmwlW1E7K3bn09Q1Y4nepkg+GPe
Lte0v+NGfN8QQOvR/1zWFRz2hiisTSc+9fAkx7m7RgoBNlQic+JeLlmM5T8KSY3i
b2J087K7oFqzqknboItOncXxLAFaX5X1aKPwDXMP3mEUbE1ZGMvxTx2yKjO8ijKq
g1qeJuMjZ6Zr/mDr+zbl6lADc9Qkzyxws78/gXNn33tDG0K6NB7P1O3DUCFDIK3s
BuX/oPBjb7qboTXLm3ARo15uykD786iO9a/ZN9ibHdkBFxlyXv/ciJPG9zAglvqE
+QnF5bs/JXmptcW0faOZJ/7PRLobT+n4biWUAUBSfT7OEBvy+b7W5Qb5iaLIvekA
ZbNw7qF00ejSNfoeDv4UKveNEjfAB7uAtBT2FXzqZmWfSwHc864Way1Lsl73gvsX
XkIAgpfeoKjhgmi6l8jUcg96RfsqFuQAZ4k2fWzRqXGqhjEXcbbq9J14S286B7tS
bkXBPdUhKPHCPGmeC30h0V6kFPTrhXkkIXWTjpZCgip+p+8OcVnsMoMmwEjvDNTc
51c4opB6TZN3f1rvRHfeDEf28GSfUskASODdT2Kw5u/5pl85mhnDoslzlHcG0ZGl
XCQHB9FD/tGKTW/8mEkeSXL1Hgl1zF2zlaUqBn/88vpNRaQg+vqFb/3p8NdrmGy/
nS/33G4OUzKJ0DFbnwCQlDS4FohMx71OZV6TT/zv4v6w73SmKm9DnqO+eksKL1zk
ftlXKyw1dW5Q+YhBzj+bz5PLeCTvZttBXQw9SBJ9V7eM3dQCGlSkH800xXgjNt8O
o3UXFYq4EwaJtogwkrKH09qvoC7ccF6ETjxv2FLTYIgcP1sSqMFSNsLXaFKpyZwk
SHeuTjNRZJ0Q2jTKFtTd1pP0qvs0loqacp/NwnX4BxMymufNc1Trx2ToY+PzVxSZ
zylbY+xR9P2pY0NvFI23VnI5bkUzZSS7b1FKfIcoVoHFP0ZcRl3gEqivOCxPmBZS
MJpieBDD9lPQwf7fJ5SXQokMHs+MJZ6dzb4r5Tsg9tXeqUY0b3d3mq8b3Id1AOwI
BUk+bFt3qgUsLMKkpE+2lODVVbZDy8lwEFoSgZGOncwWsHBwuvf0m5kGwfQ2qVql
zE2ROqVW5zJCDUCUjzGJfriAHB0U6rbwEOehrea+3iAHi2lzNSbtZaxyJ3XYZqxo
W8vtrmpfp5UgVuxEQQOFGuxSMMvlYnZD5XR3bZLrmPjeuIpdeZvm43d6gjThhKzI
1YLoTJKXT77xR5sMXxFxB8E/M6x2NNnxWySkDQZc3j3ei2Ja/1vB4sxiUAuCUHLF
Op7JeIzMbsPm7h6pNORATohdGFO96VIHfO99OZODgZ6LiEuTQ4m86/wdxBNtXAiT
oCChWsXk0rH01kQQJRHjjS52sn4actQL36E4F6GKbugfEsyU+DRyQ1wTCUOlb8/z
Szh2IFCw2B12rI+a8SvPo2xAkGN5xf3d9+xDoOCz140OffpXMNj/YSaQzB6KcdVY
wqd+TW6NJwlh3anDFeRK3mPwmmVMjPertO/CiAT7ikLf9qjj5ZDHnN4qQWXXjeIF
szSqLf2GBugRzkFq+ZjNWkEPX0+S+GLB260VZwIpGfzyoSEHhchp6yiChW0tJzO6
avHOC7xXyieK0k6+cB6LgTHp8Xoit6c3GezQ8elGZgV2JuzrXzOuO272M2KxIyBy
kFgtKd3cdgx3/v8KcaQQriZXhJgs4GkJUn1KnNipm99fIYm0R3liCWOHCpd+g7kT
WA43GyM1qar8Lp1hOqb3IyhTQi2GRMEzBxYOk7VB9cFjXPP/iEa0vkSHIKAwgpjB
LofEBsLVTn47D7GOs6xOBb1IYUULajkiDglbEG3KJY4yeiGzdH4/fjMft1fKsZmt
53prOJ18rh/QA0j5CeM5UoiJfHkqiD92jvgceLtgLZrhck1A54b6saCjNkHo3uYS
4aL/DwApuBDgxREs1LCk/meYyGMlI6uEvNjfIowaeWMtNdkLw4r6sUZPFAmzQxKf
v9s/ZM/p3qLongyYwaNxD04B6fYNxWPdjCuiyvkE0St+L+82WSjuv6dY5ANoKkQa
dvwMWdZuNa5OcMXx+LJaLlsS13s+sDDD4qMBewdT/SRhjeMY2GnJ35kXXUOlciqU
OG/Q5lDFM6o3+9gQtpqgvEihMz6aTGjDLdbEr60JfANkiFFxeQmRI7bO+lQJr8TJ
VMPVwQE8qYcKOH+i4hXn8dpCqUX8Tp07er8IaFBCNg1l9FjCWwWFuSBtbPcDC7rn
kXWA4Bb2fn7U6sE38uJI/uRJYvKyjQYV5pawl1tUpBsuCYlHVX9wSDSvnCIxrYcI
Q3DdavK1e3CtCuuZ3vefkcYt6d7xit3D/Z4As1b7aHBorNiW6L/8M9EJ8Y4JM+ru
oKaS+pbrQhmx2TvHTwc3fvMrrPJKYN3CcAyXvDKPdG1fDmVCf7rS0Eh8cYqBxl4M
NrMJo1QHCHdsotYrI/TWcp3GTElcw26nH9u8JXHPgzDaM/SNQLItvnhgoiBUjqz0
77PM/6m71FeYoziPOEpKV6rxxjjnEuRm3pWA/lhlhqeew9K9jfZCFauqs0KWy1+Z
+PZp6ecmRwY+TLxSLXjCMluKYjODJIegL4s7+wWkYM6Xgxby6PwWap1Tx1/8ABhs
rtc+SLwPlc0fzlzktSQHbUMttl3PILqWjqvW0qiDdmSwEs+kO9RCocbvBQJwjbZ3
WIznfbN9IxBnRDTN9M/yADvcoS9YhMU8n43FS+7+Gjh0+v2ZdgxJ3Dv7ZLg9lk48
2hWnbDO+oKNLyH7xEVprzT1KraOm/km86I9kJh42E7DFux4TzfIz+sEHRKY7CXsl
Mnx8SdaN/LANMX9ghg8JtAkgWAGjDRipul+TK/TycZGfCJi30udbQcASxtwEJY1k
zdBl4eXy/YUQuHJf1rW/QGaSqeEjJp6l6GWDU7nwPMPpJIdzq1MdMqUBJJ195R72
+SX++S2ixmYgJm/t+VUg2ntXDvZkU57HabV0L5LzLspaXDmkA2DfxYJRynfs20/f
fcCEoqiYP2XAtmdkAUuVMyHRPAQ4yRm8fYB1A0J8ubLySOdwMNLGr9VtGtWtDT1p
hIjy3K+31u1M6MefZFcdvYYfkHYp+D0lBt53SE06dC7CW9a0hGwoRjVwY6CUGvRi
DJ9cbJDUm8UhJLCv+9c3+qXPNQU40f23s7InPa6b7BvX5g3ifvjrprkXyEtPkj/D
HLvqeRe+ZHRiCOSll8EIrl4l/mG/cvp7lmHs3EK/1zRsrAnmPVoWYG8dvFPvjQk1
1FjWs1MPp4rpqpv2Pj7WE1Ds9Ko7N3oX0qWM/wJd0ZhSgul00pfPrcPRD9xM9+PS
8qyTvi+v9/IZLMg0dH1MgtGw7vLqu9F59LEn1Gf7s8ZHfy/02We5ewhJvqv3MHoe
IXO/pI+0ilQvlYtwgnPTaizj2WnlYSaDeI0gzYt5pX4AnzLqOatVX6sgnerUyDu1
I5lcZGy8562gOrSYI1t8DiTL8Scmi4K9W/YwacbeQoa4n4eswgYerctr2IHVQISo
lb/BjPGZOO2gJcGHej6itOq7m5nc6ZlAHSczcI/CiVwyO/Sixq1Hdth8dU99txlS
v+Eu9yi0JvES+VqvPb4OnswjPXB0xu6oVjMLj3cWxbq8znwYQNRxtIW/kQ7Gfk2q
zQhvUq/yI7AH7WcoKKXbZ7HA8ism8OU0pE8N2TS+/yooryzN5leERVOKIw6/9sgA
ebGeGymbOux5Pa3Pey17zdKxfGszWR8zAhXImEmlSSDVMOIYGJMiqoVWzVtnyEfA
cuI2CHK7Py3soAZi8RKrVWfUCxEeybySAHkVo7kCu6n/Lu/haixWF5KW0twEeGeg
EjyT6sRSePTYz/rx3gNJRQ8TbCDRa076huPHkFpxHvoxRJMsIJ7QTlRoUMqAY5ft
HzN+qYkLNgUs2rsz++fWpxxFCyikIu9gqClTys0ibCVdcwQG3yu3OAFdl7vP5IpF
CFKD/Ul1MNSX/mOAxYdRcVihuJTPVAvGpv0SKMvJ9vyyZvqW9EiuD25vt5zPsDI3
9LpYSHrC2wMU+tQ/gPr35YzwH/5ZrnuInyKRBn7RbqR5vYBpAsS643HWvRbAqCRI
Dv4eEA8eCagCHHV0PkfTPG+S6bRdBgSKU6yVYHRzVKuWOTn331xxN2IkZQrvhqnD
QBDNAZqVxpAsF3czMoOps7bStcQSTHnTcFalOH17H68O6dDQOqkyEC22NN6Hzse1
YWHNUzUqQJXAtWMWr0orUWoWoUM8+SiDhrOt16TEI8+9qMAYmHHRBaoxOYI62Sk+
tqOdYz8M6GONOgyQRuGdJZEv3QZrNMeyzK7smG8lolhclUW1+rUWBrYbmhcHfT7V
bkCA3pI+DmQ3e8v2GGMMyjEKe6Hag2StEZOw5P2M21GRtUOu/Y1kYqRZlaLbJtzv
7o9pIMAtB8D/14Q0QT6hggDaEdQWTVkaMU7KqggIl3wXYwXzxAtGY1Vvz4h6U6eC
yc1njkr0L3MorzSAWHzYNiq9QjBPB93GhNTwpSNa/sWNqYLjdy7Gembeh1MdnIH3
31pDWOVRL1I7Ci0zl5qg8TQA3zt5eDpo7cuAhRJwVerT4okjUXpzEJmpYOfD0NCv
dSUuz02oXaRH3YAMK2O0DPKxhhgQ+TYW55ehCFTSSPyPllvRByLGpfL04Mo4tT+M
ZJUrdd7vRNLnARKLM+hJvWOC99kFaY+EP9g9MjTfq0UfQaTPmfySpHFq4NzNdf2p
Vngxc1d1SW6G3o3Hd++tUcgpUOo/HU9mmWG9aDUmJAv08HK8aH7g3U5ppXryfdcM
QeNnbZjgJfiBy3EAg5+oHk3KPSFkgHPkcBhaloBK63B0vXzLUFn2QYfwAmhl+B/6
Q/t017O4zmT8GlWEElqSBtW7VmpJUB4KTISEdiuq8xSDtYuf7PDEECubK6TcuNmq
BB/DQClDk0i7VokVsiu3BvMdUZ8ySkmWWjvSN8zg14Bs+TGUR5K3UIGCvqB6Gpfh
IM+ULLmnf/AGe+uG47wwgSvKx5AuNc1B4MjwSjfznLFQf8LZipRLbJEIDtFlksY2
RWyyNbvWfxNHeatyCh3QbDAMK0jU8FrjtIwulD4h6OA14yv7ePkVngFtj6xs0ukO
PnFo0Orm/2yzfKrnyrhajnrVf1whtpFXJS1FPjvqqmTYmRQwnFyHtOKyzJOpuda1
1L34G6kkGLHf/MJgB+gAgoe+gU/yCVPshUjGDBF4yAdkyHXCCWX+qItKpqKo4azo
D2tcydOLmcOl7KJ+nOuEMZ/CB3g30Fuckq2Wfbq4vypTbX2sI/Lm+6ioibIp9lmT
CnDgMNeAzDFgBEF6T8PH+kfThKPXaoqcDME+313d6DmvkzPRuJ04E9vnRtRFrO9S
dCyRhImrfQnaVRxpV2Gsozo7x4TKEQpB1ZxMkjR2wibzoR+CPgOSlUjPcZpMVfdk
9wvJlIKQUL1a+NfqorL6yhepteqXzDEYzTs1LXFGd16UVeGhRc1UonDSiVt/1Eia
j0SzzTdK2GirhtkIFXt9BBxBHjkusgssJHMZ8cqdPERuETyUXJMgzzOsU276n+od
Z6vAdpfSPbq9ETecVO1q118FAfYDS7kQtwqaoLLdR0VmbVFopSHG0H+YzQ0Kon6z
NkdhWLJXUZ+L8qCRgCtCijbDGJ1MQ6Av6rrVCuSFUzp0+Wmp4zsifsvypnRpmAhD
SzxUXC7rx+AAAKp0SUiUQmhs3zx71GrbxK8W0MDu+kiq6gSZqJVfCh/orwljn3PE
DFKK5UpfgIkCSclDBbGPHIQ2j4qV59eDCYKxo1qLTcwJPfD/iTjRKccQ7LJA8vK9
e3JDPfDqWav7kzibSnbr5+kd7j/k+g38g1IYcR/6GliY9+rHYx3Mus8iQHlhG+yJ
Ty4Ma6yXUzukl1qo4DCh5vVAC5+3oF7T51O3+jTKZSpTRfx3o8qrXbtQ3maJtiaW
Jff+B2mHHTz9C3UrEl+l31VrNlUk5HCp4gCNT8y+ylM7Hv4QPmH4q0TKKsj+cotj
B9o5mGrPgp8hezeeiFqmJKgzf6X5RPcUNBm314qmtrdMReFUvBrMYGpSbSxF3vqy
B1ojp830eHH/r378XRd3k0spCrKkW2zumXcdnnbMzLPs+WDkB53iGHn6YS+YVa8Z
qjzCUD+UXXgHRJCwGmilJN6CabaCjr+4qC77R9G+QHMQZRrxz5+GKZuzFd4UOQS8
/y7ERkEod/Uw1F8m+1/HLmWVJHyWvhLQxvJ5OSZ7gjym4eIdnQnORbiPsUoNyMZ6
SjaDw6DGnafhzfo2LOOV1lv2E94SIhsffYFqPACZ8iwcVVIq0lkBMKKxUb06hJ3m
HAqpcSB1b0SKsPZZZPMgnPWhOoGcI8vI4t9r5kPrFKs/4dgp48pN+wgzckhbfsDR
J+v0DkWFlN0h/gwE+ZbH+Cg0I7EHLrc0voXoqpaTTNwQt3tFVthRclrbb9Xl/Jxl
bdt/kgTOjuPncAoRVuqGuMy7fAHqzlVjQrd9wzxZ2fsumiOVBzrU27SaDMZ6aDNz
4WjjOnLPE+UmPuC+69jExOzjoib5iokbDKHxlkRTIChmUZUP9FqSNstPsNNGgshv
0RV2UbPfk9dTyO1GxOJrTRuG7o+Z/LE7VFpyudhGDCyozZ32kGXYMKbA/p4rGG3u
eioUP3vLAs9OeXSGlw/UquIYYaoH5XInXGMYV/FHYOR8KGz8BQprt+mB2v23e9KO
hH+CKmMLgSDnTquh2KnzcbpPSSFcpCNHOiE2x9kLFgnivbgDi3qUApmBcFP3AcFh
PUE5p2Nhv4KSxSZS385YP1v1kXVwssRG1OnmnjsKu9RQpyqDu1zC4jvryGRLxjbF
lflJe0F9aekYzfmQQqDhgM/x60qsOBjpV5nVg31N9xLKCMflAfTB08C6oowWVytL
Xii3Z4idpRtoXEXY8SuGl49ZzUwdOBdF5viBIJ+9aXw7pDQARBy9FeGRpDTc6fHa
6pJQvLtGVhnIRj/Pr8+gYzpnEHXWyJZRhDj8O8ZIzPHei2VFlYtMQf7ve6iq3ngp
sdE3d3/tuov+vi+Oc+kJ6ZDFevul51dN1x57FAb/I27QaESpwI1g+nq7DpCmuZQW
Wk9TcFGHiWy6kXrdr/7+PiN9xpxweoNuSuncETY05MPyG8NYNlFDZ23XCOwJ/dsM
RTgx00LhJQyzb9FZrNA58gww5kuDiwP5De9kYguIyf7odFEAxjlhq3DuY7JlyesX
Hp+KAJsItcBOjhyVc12mCj2asbEQYnf7wgUKxyWRuYiL64WKAEkiPXuhRoX/iqc6
vE8UqYhVinrakpqnd12lrLvq5lSmfpuClL+In2AHrnTYQ6DEEtRUoLaseNwn0tHL
ptV6xkjGfv0GP7UWZDWLfK31ZxFR0XOYFq0RgSxMvFAqdsyfJIK7Y5Jxol21/pFn
3MfVRYR4He2JgHlda7XDsCNl0qMWJFFl5sq8zD1pU/C+cXhR4aPZ+Ra/V64VOdbl
4d4oLYiE4bUH+D5Bml6XBr9VeADgI3Ycxw2imeJL37ExiZ1tXILFwXULslMpa2BZ
3DhJqtfVA3wKBCLdhovDnQ3DNd2eBd7SaZG9irunDG4+MQbPVKsWjA59sixBFVK5
wgPgk4phszdigeWI/HutIJ3enqFsY602m3eOUeFT51PJchuoHYP411kMScGkFltP
7fMt9UHZaQzsMnqmhALnEChpwEnOeWoI8WAGQ7ggEQqabe81JkE/UXEEktJuw5xx
3sApgTLqNUdaL8iOFI2ZZB9vDEfUX2qZJaiUx4hf9pnUHdGDcu+2NBPAJBBflp7O
28IClPpRgl86Urmp5ghkiI3hfhlL5giACWhwR7ljaf6QcRuNOsZ3D/aOmVJP3w56
5cDP9Qo997bIC1DIPPd/wkpQ4To/uqfVM+uN4MW5TCR9vzh4qPwM3tN4CjJ83Ifu
/vZjiKv8O8YxRx9ROHY5BlKVAC+ALuQ/IfvUi4OxIgXQlqd4hmQ0FVlOiw2btgIY
f4lfeDbTOqmNQFO7I9T8V0UqwwFNDMOgIVBLLJlM+Sj/zVkfN8LaJGi72r04XQsr
SFQDJA+bcbHHDSqfosgzFdpEaER1ep9e8ll0gb+7gl6AgomeyqSivalWKK4Ij2rk
RIxJ1MWgedP0XQWzcy1SmADd+e3EWlyP8OsKC6uppQMh4Bu8wY4QdCtf6Cjqgrso
32ei8GZUWu5jDjY+aRgS2Kg8LeiPOLuqJO3TWWm7MAogU/FfL9NVigrEE7ndur+S
mrCQ31VRp2bf9hPI+OMgcbS3GMDQlX+jA+r5FAA2BFqaciMVj5aXDmwY7+9NZx4j
RKnHqgCWv+zza/GvH/6ao0QCIDSK3GPA8veA2Sp03byVei5uDGNbW8/skn91U43s
5ExbbfGXwy6bdedrpIKE97BwjfaauKByB8XRlpnbP6qTuteudN/+kG3Tky25pStK
DSJmEp+rnX0ZnHSRmhV35jElzrzI2NUQ8LPTlVDrkTqjJSpezGJxeHLx4uNqScDZ
+Ve/Y2uEAm8m0mKHQ+ltZqtz1rkkIY5t95dawf1iytGUNquqy/lg00OVbp4Qj/+V
5II2XfL/i6goVPehwZBgxM6SUnhrjL4Gjn5sL+cLLPmRvj8S2FwEUmfbsZ0DLRCM
qL2Q26XVrDhLKuoUyN/wFI/E+NQJL14/vhb1uxwFZYHxune/EGL558QljzjVpF0G
oEFzgJzhdW31aVchOs7FenyqLGADVCB2MedhMbB2Rdi3GceuRXUYLzm0P5g86DJj
BmRQqJcSIDTvrZcobOmTgWWWE8tC6WYujl/sn5fMImc/VAuqLj2MnvFbZj9GZZTO
ne1mBWTnRpwzpmyY4mWv7yPECCrkazm4SaTIklSb5BrlM33F/K2SNa4QxadzH1Xa
x/OFRTlFKIjQonxtHKhY4tHPbwz1t6wcTo3RaG+XIYuvHPZ4n41TfhcpuOzw6NSh
x5R18kQ5CHgAQd260Dhz0jOCbd5ZFPfX3kXOnj/ST+pkIPxuIkzdXX9nAUyfsIp5
5+QDOgG3QkZabnjwRaeaAosJrsdLQ2jyOTqUeNq0ugaTJqzJsXUpwxMy+5KPDbmR
hjGmo21zGzPUnTt3XyeZUm2hSDkHwLYr/V5iMHUyjIF3/P72IL7ZaQx/LXzf81fX
qmrBjBZrwK2IFUX+37xLGVoQbtfgQQcmOSYq9ghEdxtYJ6zTi5lLS4sfMSxbIWny
2IqupjNpeRZh5DZfvhCCGswClL+xRkJgVemKpCttSS4Ajpt3K3As9I1aCxQspsN4
CgiL/7D3abkUK4C7gOjJXZptY7rMe/dZYseVINK6I689V7Ie9KGI+1JJ++oAw+dH
tnZIvlIvm2pTlIyVS435AeafhRA1hvqjxydYfSwHkQa2EeTuEf9WqbR129uLtIf2
EHYQ5jeVwnXewQeF5EGT/yHfLoqgcV/LO0sh6uI3ALACYmpV6E8WiG4g9D3m/IAq
L6dAMjg7n637ZYAr5du2+oliApuba9kNYGfQhcLpKgjaw3IzsuR63C3Anpxnsbj1
eP6coD/LiZVI6UL1HfZkJ4J9pyBWfxy6tkdLQ44CEUEQKLR6Bo36rAJys07z7ebO
CW/VWp7gyyuxj5hUCEioXwj2mi0S4vFfBy8fpt4bF0q+/Mh+8825YQl+LQGqbpXP
SOdHP2+6vdSJJmujMEM82k4YODO2+G3J1MuFh8LiGCDjeCg3LHVZqv66OsQqmwDI
XuXyTIcZt1LRGFntfo9swC/TSN7pE0N5olMJhH5vzjKnsF1C0Zhmyjwk33qOK3ld
XviONgE89dxJSXCUZVdlwT7ryuK19zzDiTJm/zaChPr290Vm8/80qxBI90082mAY
svopL6bEbu5XaPaH5H7cpntTVkA6YXTf10rwRFVaEy+4ohXjY53kz3AiVsI4IGAR
L7faRuZ0N9UYCBqM0mLF55s29QrZBE19+vOLgD0RVf4xoNCZiRmJ8IHLNNJuq3AN
yWVG1VnYPhq5IE9taHH6dtJKJLLMtxKrC1p4rQ4qbvLjtOHJf9yLNUiPlSPr+dCY
3zkSCj0BEuq5v3sYBFaO20DrwEtRCL9b9IlGzY/E4fjYdxFCSR2rnkozSkb3kzrm
pxdYhRQoJ4YBfB/7Nrk/+JdhrgS7DyVh2b3N9GESGdNXWcN9x854srvrU4iIxMzL
d05lz7gpGCLwH0hFDLrMFyTqhGpNw0txOD5oHa8tK1Qq0uQDjD6lRXoCd+oBtCyf
yt1apOD/S+uX4Ssa72T4syAh4j6GxhJgP9kqGoQ+gU8BxwGB5fHKpUYn+ZkglMOl
8JghsZ+tuZ+0pYFaEDgEZ3WfwGKbvY+iES1XHCZ9srLLlK/oKDbK8+hrOnztfU07
7VL/ma5QeYQmUPxToH8Bh5mz62kmFCaddJJdZM8NE2FL2LSCUGiXqSsAjiEgBP/f
Q7RDidv8CQiJ3CPL/w//ODScJTv4CiRA+mYSjRNKajTIB43ZiQm37Zk3AhR5mxUj
eYzYX41O343BU+QimXMYC/TkimFi75fZdgBCN5hp19dmQYB6bSXAZ8MzurwtSOwv
BfF2vc/bvtS5D0rQYCdJ1GPJxpVBqk428gnDWL3MeBSa5ZdqAucL0nfRZiS7ntJt
mxamopZl/W5mrgPcxdzG0gMc9F4OV35o4qLAanofEx4Dn6RlJic1RxOYKEn+4n2i
uyVRoLsLdERVCjDO8FMGSfxhTTt4uTM02meoc7PC0vMQInRHwvcPbeGb6S+LKFr5
ghMVYokK272D6loU7NkMP4X0TJE0znFUfHuCrMfBJh+HpRVh5lwchBpj2zlTuL+i
eRlSTbfs0bpwOfCFYaUAsnHprz+utB6/molaMMVM3JFUp44vfnL+yXRfwadQDev5
IUAunRNHy/JiIMqci2yK+7/5CIvr+ncrDGo5N9r5nwzZe8m3zpiKwecKb7gNwZc0
9EoPWKlTnIepAhikErv9Yw7Qb2CBIffJCDI56FPnlz+vWjgAUhoahcZ7ofXnhl/s
wo4++3AcBswlasnQUi69XI7qjyOBJ2ncuKs1kO4RBibbbeLAYUQo9kvqOIhDOHtN
4NtFvqUWdDvzcU2jgq6j3Ryxk6xkQ+YrP/jz/dR/eSy65pMTEuxPyYWjp+CNtemA
fAwGksG+cH5kCad52f1HaB2dvWKVdYeraXnC5Ixoh1DyOoZwqegTPBcMn+w7WHti
NWQax8bQNlzQVDAY/V6f3Q7bjS1KbhaNByXDKpoWWfr/h+eWOMGmdWao+XLODK4s
Tl0N3hRZBTwaez17IYMHEQ1s5b31dzM/5T++ynAPpBgm5f6e5YbYHGbsgFSmPKHc
qavbjqnQflRLtzzkbrbMnENl/5x3yA0d/tMJBmk5PAFPaFBhdP4d4eFbbg0AaT1i
JzkOYbMEqzie9DOWP+GF5jlpqeKMlOoNUdH5bvFz5Tho7tGgxpq07kJ4HYBzazl2
CCBpZV63ycaEYWawvZcA2ZfQlm7xiVZCw1q8jhs08wuGACXToWE1cKU3X4XkJbuv
tPKZC1XiUiWvIDGDt8lDwXjkl1MVX/yMNy1NLfx6JeBeQALr+m527L+MquZj2pTl
L1e8vWcBpEp2mQ+QvHvG2NrkrFM5dbKU4Ua0Aql60jR6MqMkfrAuJ3RlCM23fe/V
mPuKOzBhC+W+S9vnw387HxVLRv+aaGkGH6CKIkUBNQYbdc4LfONa7DEnsNNNEK6/
EJ3xRCvzQlWV9Uck/VZAymPOBQhLDuq82itT9eoNnSYzezWr7r3yiNapFqWREQp3
RTO2ODSDUVCfiA9T/hLYhJvjHMyDQr6mP97XGCiAo3tjzS1sUepT6XOGgPMoa0oo
ZOfH5jALXdq36xjMj+DdeDXxDWYADdn2bpHrRnjWMg5odr/AmqBaWFLmyBMJGon1
Y/L/j2ikKsiwkKCfuYshcKRsc2Vq/cIfF4AFNCB17CZr3LXwFci6bOe63MVJU6/V
TKFRqW6C/Axl1YFLxEIVcJS/SOnK+cJ2WkckSD8QSlSZnlKQnI70uac8JpE0AHfA
JI5rdEX4/qdogf28JuiiL5WFfTADIDj88/2IByGp0du8DRtK5WeEdg6QEA8qPK0m
PNE2bJkzyV+DfbNcR0i2dvqmcBWGMFPoEtYzRonz5h5LBJJwghad+RyQVeb5VS5w
XYbWWNysRfh9e6ztlbvkSHV4OnF8u3XIiXNpkuWCenjPtO4ToaBt5SauloNbmJMO
F6UBfRsS1mQxkVpZMHjV7k1kOmgwRjKkM6UdSgM4P7VurmvUW7dLblnKgmuoz60G
6cnnKoD2JtCS/fMjwNCKmx9UE8ZX9mvSwu93Jw1qkENPj+8hQl0wYTQCRXmZpQKO
xJAn+gmCn4GAWBsdlTLSyivZFd8VCPu57DK3l4csOOwJKLrUZ4D3/vCOepiBGW0w
OMsnn/wIuJj2VAzLxpWZjVqMhgo5MzUSvC1DjtiNE1dMiuCOK/ka7sI/ag3GRVaC
3HqUFJDV7tTsERIfRRo2TUV4tv9unhh2I3nZmGHb7EEXtYbIt2vTmGL4Woax08lT
pgZrxQF0ZfpoUxlKLnJub/uG8ADpGlJxClv1Zj6q6Lsbylhz4SQwoS4JM9eMqIsG
+jiiVQIZuvKyxOO9wub51jAdQWRSeTQTZQ5utZjdEfBhx6khJSj2mb2QyRvKkD5e
XESqA/erTWqlocTDRCQCWSi6O+W4iIL+D0Z2CD9IEvk11KxBelLmeDOLFFismajA
kFshIectlc/or5jedoG/+SVCcq8epIyZN90qIoMQ3aDHOzvINWCWoapxRSdO1QCZ
qgxwZLgoKtDT4yMt5KdqdqqidDdiBv733ryvdR85OB9xk5J/m1vJ5b0aVLwsph4x
+dexRmE7fqVXl0HP5hP1JmrVnLMIljW4OeYKGrHav9yO6i3iTOChJZddWYHT3Fa2
EEKdva3mtT05eB7U4VzyNc7ji/boWwAQX8vsvkiu9mWmbTZkyUa3tBqavnmKxdLQ
sT0YBUaE5fTrMobLJODJVdRa8vWXga2Kk3UAJGwcbkKYudZ5mUL8t+JloFyCQcls
EMsZ+1FBtUvMB7xoZEuk4NIfh1QfvfDGMfVxxrjtTORYR4JQM+fiAFrMdIby9Zfy
qfY0twsAjlQyyjm/roko8aILsPnJBo1WnE/Rib1S0w9AWipV9EVkN0XCJjsV3vyY
jzGJbJXu2tHZmXJecpQjFSg6lC+jouUpoYKjCAA3L/nP4vwt7L18Mrkoge4TmJQV
ghdF5WKgPO27/kx2eHfwF0wM9Fuf3pqNB6BaylQNwxWLDRAYmre92EvhvW8c2G6n
7ufxGVz3M4ErdQdTmiWndp7HMNVZwfts/Ub0x6DsUoxKP2vHJDR4042NFh/iO3QR
NZOc+r/4jXQ3kZBbI82873s0LQr+kYaSvZ3Jh54dfAOqva8dlz2EBIBH0kooQ91Q
k8rZw9A1xvR4MZFjAwORFc/CClme6P0SbBzWeaWicHJn2LutiGqB6qBD/Mq9udU3
CzGQlqAxRae7KsOAqa6JM3+eyBgs0LVByBcAtn58FbuZQs1iZqcVqEBc8is0tx64
RUC2567lCMPQzuA9O4pxSxUnkNTPFLYRFNo+UCE2HNzOj64NaHky6G5znC6EYvcG
0srF7weU7nU2XieaMn+oXt33Pmz0eMfwQtC79TvV4b1krbOiMihiSTslUDMUifcE
GS8SPTwUHuN8FKer6vdG0XNIhE2L+T2H+A11+j4mrh/EF2ZZp+SOSuFU9sqcXzab
Rtbdb23L7MzWLEF8Hf52gJhtPCmX3hzUUjoLwJliIPF53zXJ/ayGLBTdkeWsLQis
iaofQ4ZrU9vY7eTT72KlmCuT2xsIf2AwQQxMo3ju6mhfm+MUpJPaMc1jHYw0G476
nzT9/vg9D+CR2pXE2Nj4w2mnFKhxODdgN3qOXI0LVCphz4wsiSFRgAF2+IbAcs56
dIDVIHF4KhsKo7l1WsFjldHYWcHw9pwEFcPdrgCfaCsNQ+nMTUjGqIGpaYIknMzu
XktzcgFXOdZ7Q8b2cMTE+kxztPdUP/MJzH2W5ycKigCYBPpHpkefvuvDAhAesABq
HlZrelN76Hcrt0DxfBeKM9WarSt+3GSVKDdzL+CSqSfR8M/CyUIdM/8BSeUxEBzT
NO9fYzX9ASOMvMBatl1JFprOhlZaEvxSXR80KOquHDZmNo4TkOR5oAK+UfpwqRlf
53npZGm/SJ/rS/wfchoYG9CfcB0cfO7AxfEtG5CTqKOLcWyBb+k9aOXp85Yt7oQ/
i3UGzahuPdtELos2cbnn0yQKQMR8u5WL7duANzLlXIqAtyrndUH5OdmR+TDgN7Ua
rTSVqNRr27bvkDQsknrmT7utf3P4Oe0ZqIHsuTUXt9WBZyVc78WKsreWGLXXH+gq
WlGN8F6yRQnpdqRuHW3Ob5Jfx0PZT348e4FXbEtArJKzrj3dLUDwFAgrKNGjSq3Z
//n8oVEcKFV/HIXdCsGFu2+djEYEox3mryaNqNnlsnYU/heq6oJHIEmKeEsKrhhd
GJHEiIJg6Pi5upx9XTb4x9GFxC2G5oV0rwH68n0y118moT/pd4rqiVzVV0DSi8u9
qonFTmdoJno/f501XKuOTgQAlrblkiWroyOdaeF8A6+xNVZFE1H/vbOyKGloku6/
L0yZXjEpk1Htytdk26skWeiDfViXzOnAZjLF0RDw1kng0BARk+S9uJXK/ZtNzH8g
hQDWIZzHRdztX8284hjSZEJGGf5Q1MrzMwUhxWtmhbnFy+s5oQQKUCwux4S2diRD
ykYG6BXs7NBpNQ1FZGDMuesVso7+HFzl3Dsg4VgwIPvWB2ZomsPrLeq36wLAyKlc
kLcP8KNw5qhbJDGtRcBHlUT7GRuoQZM5k6Wwu04LxxBIVoJImCafn8J1Pf+/78eO
t3BMkLXvaWF1v+i27vb7dtzp+x03h3hHl3k/FhMDSdBcQ82mJQZh+LBv9tiH6fTh
k5gXtyz6G8LUD3VAmczGoMeqYZRxkTnrF2rUgPTR4mVzUVHDBELKpwngKyZlOe5w
boqeoWyUqNOxd8DcB55HZVxE1raZJThH3kkrrl9xzXXrCzwPS/vF0fjS2LPTTGTA
MOUI3zIsds+vBN4wC2kChspDwUgYTBP+zg3qE6/IfE4jXgq4wYE3VaqELj6qx49B
4r2Z8S8gb7PgQzsIQeOsgaZ6fmXwSuLn0imi9IgYYKLBHT/dJbsxugFaTtWEyb5A
mHenmV/Iq/r7SDB7QhJY6eFtZ9kVCpcbBH/lhOmsgDdh8PyLZrCpYR4ANlqMrImb
AUgswHuJbBjuYVUBNo4KSwQheT3op+a6cWXXxn7JW92BBjsFrT0r69+lf4+ZCS4V
fMGD3VE1H+aq4+FtKUTgh5baiwVX4p5ES8afwPSnwpqMfB1uti4qskSDZxPvLjQp
TCEmvYpBYlMK2YrsoGZ5v2gwaCaKKQeEOCcjoH6lA0w6g2S/uG7XfB/gEYKorCZM
nYAdRKp3dIFab3b2h643Wl5KYUG1Awn0DbAVpVyLZj6QJEbeqC+eiMajZXdMmZqJ
/nBOVXW6lkM6QLyZRWrJ6D9W3eiE78zaYQGKHZdxN4+TuChf6Ckp3vI0D4LGwUEF
9r4MuwTKN2orsXxPKAIx6cOtxVASYichECakTETzlRJLUxlQEJs0otWePwIu+kne
FYKaj4Z1b8tDnYSpWfXwSZq3dOAByjplAxBcWmh3PpaC0zxNUdljYVFYoWhGjbsZ
AJZ2v9rwvzbED4jTjJGxglMbAjjf3LE+3xFWU0426i5fz3zjOQuBMxGCBzJgYjv9
fcP5emEr2A/POh22gC6GjFwqncI7ueW3opNt+Dxd5A+2EZ+17NzWlBiliDXq/zQz
IWVYSuR53QgCDd+U2+eAho6II6Cv+4xLat7GDhJ4uhP29Liope5pV+CnSx8KNiBi
F1hbVF5PAfBcZJFZqXOZsyNkpbU+eR/KKS0bBL5FOxU47KA3ph4OV5SO+36FQY+N
+OS6wcgbH+NSquuP9u+0oWWGCJt3x7Qvu1Jih7/uQn8+M4VRcWnNsJ8/2vm7BGAl
Z/013G8vlWUGrqaPASMFiMdqrE4WnNat5CZYA8sYoTPVST0hbVlup6ZzDCGqI8h0
s+A4WDtcUfkAR77VBfVeQ5vP/yRL+Y9WPCoSHroZrKmxBWQjURNZjlFuuhioCSWw
XmB5Uj8MuYQfJYggBN7ZOSr/Zcux789TafXEddYhXnnuWGtU6JNrTi9VVFs+oxkg
DgTOLokl9JtHszQGYVwUxgOLfkDL6+65XJ2XWTzfZ2NBpHopeWkymOjURrD4Awcb
7Lp9bgx0vlIj5ouE+2oUekQzB7gXYeN4HhYDcXrOJx+hzbPhI5rd/4YsJ3CjdRNa
zwkrcl5h//z+/BhvpP69mdfuuAuMVmGICx/nK74FODmxeadhKSHwtq47mmffw89s
kWOhRzBSCYPBOYwq7oH2CybEj+8h+PKA7OLLNLenU4xsAzoIbve5wQu++n/s20/U
12PGqADKyS0mWPqbDbs6I8F5ZrEfMm5+zU2s1LYls1G6+2iKT01VF67M4pA/Fstv
wiOkmKQmdDIkYJzh1SXMRmfxxpV/dVDTOdw0bNz719P7U5+wgelBo4fIDfY4KAAE
CXfc1dHqfueIVyUcMPETQBdJr6DjThALYmwCn9ohAuIpxZy6ia0TwE9tzHhJeRzI
oFN6fQVq9fLSWyAguLvkA27dosfyWe+oH5psatP/fIP3IR3YUrDZbjQlzS7buRJX
WLWsb+ZPQ1Jgm4KRGyRvn6iX8MRs51pP6EbMVnrXhS8L6oriH0Bb3c5MQ1efd1Ol
XhSuIcK5W5PC4uMZ8mM+N3NhYv8L4BksluPdm8eR9wah46v/SeYhyWintQXiYulw
QiczCqkQaYLT4wwnlLWxktJwKdE5MLiNBuFZNUhWpLjoQv5ay6i1SOdmuH8afwCz
G0rCF5JrDbmFv/aG7l6yCX3fCvtCockrbPf9S4VYMXtTFJCG+AeJPGh4qzR3TbAy
8AX5owtNnf+NpC2GZ1CI+P1mGAYT1gHr36tMBDRmptfy22aXAFP6A9Lnsf8v3neE
S8x7PejOWJ8cKP+nCCdcuwv8zeHj8525uN4k78aCRAHQd3tx3dNi4f0ePk/NtwyW
oN3zb8FoRTYELv6xlmXdhHh/mWl5VW6+z5q+pB6fR7FAOLTUUNHMdy700UAeozqu
LvZB3evYC4Vv6HEch6LM0zq7TJcKS9k2kjAviNs1/S93Jgs2Ma5x98MgN77eWijq
AIUYS6Fh7KEwo8XFqH+LT0jzXVGgjTgGhn6U7JKqV5fuR5lfMAeSFxIxJn4ct/zk
jR7jVgn2DyQEPYm/MG5LT2lruGtZkUpQOsvAqctSBkWsvwEgp1XTwnCOByOTf19t
CF9hkKSBY/V/GYGhneV8GNFD0BhfluDtPSB6QCrhbHb13w25lD77h8YAkj5elfNG
yl6YHB9kbNX6TNbP9x1As/QismQOv8pm6OhJS8eZ5pfErRhB20F9+MXUD0WdNQXX
T46Jgxwa4NCkinBv1iDM2pe0sXuh0AujlA7mCp9ukCL1z+frQtbI589gLit8cl9Z
pJ3/6Dl+gTkow0l7UhdCzPi0fUWe6XvQ4xqg4Lrm5MWUJJDls0eWapJduW06IDAI
kjlfDRXBJS66dWrB6ZUhgOUC15sqvXF5w0yo6zlWLByPZkAYFx/U2Gl9rj1AilC5
4hGvSU0zsDCzqAz96X0kzygDZlYFbvOltQvzvHOyL6Gvlrg+SPQwWWco9JG7M9pT
sqeAySK2Ad32IP/Qgf/ycOFY5jjYE9AcZNOgXoaKGUS+yl6HgMcPfO83WqPEakns
IuYi3+pf7zQwf7jDSgll9y+ArN0/5YL/sM8mzbN8+vgyWmfdyNcJPXIKe3DG+5xp
g0PAEXyBzVtNmSYGTWsWHDYtKkXWhl/7AwjyDYVpjzYBsHJ+jCPhKb6Tq7ThCecb
slzvsC86GJlO3qWLhQ4W3PgrZFD0DOPiwBaGgxpGHiAQdUGvc0E/NsyBLew2oIGO
4cbMwsbXyrEWypA3VOsCjKgZTHNBY/Ay8GqSL6F3scBgsaOvcg8T1FL2I4iLvhVV
b6FvHcumeL04NCQiaYP7lWZe+tqicC7U8W27iqOmpU9Yctu9U+4D+UvQv8h4+4bX
2p/1kBrJXchueUVTuzjqTGfpyQXNJp39H5YGVfQ2CSOFpIRFHFBeHDZ/lDf2taHz
oOUqcRM+fpmHOuszf8rmdS4XTethsn8ePnlXc1/k2KVUGru1aaW+jYOVm0u4Owat
Br8fuiTtAjSZvYH1TCMVLzpyZdmPUP849mZM9kQO5wjOBll8VI8a5Dr5W0iMQd5k
gXp1lemHsNVdDuI8XnnvvBEUHYCOMC+dNir9Q4eB1KHpQQxqOZ++8hfmT2y46Y2z
LqL/SDlp6aDiYxq7rcz6FGlgKHwJiFWjGVWpBpvnbzP+e2sITwf8vHAYJBGrL/j3
yDuTHxynf1VRPQc2O29R2OTtH2Yww0i0+UH6MQtOSQaZ7jRfMq/KIAEoN4nxc6Xd
2T+HV6n0rYcPJG11+El80fpU6kg9O4TTTYH62qmrSVcoungWhW3ZovsDrPOeyevQ
lIHFQQE/k3hAEk2rw0Fn3duxd9uuBRFkURUCPz3lJmTurK8y0hW1VkXuiH7lMPcW
gGLhy211lTu0HHeoyCrEs0/Hjp3hhSwl7GsMH3etBUvTxIkxwB9VuokN9l/VUnEd
chn45sSC8UMDjOus/St46sU4ekADNG5enNWza2Mv/2QCDlGDvcKCuma531yXf0R/
g+JrlfSacXbra5467uUvzOsnZj8eUiIbOAgpTjB97qMwCiUoypKHmahZslP8q5YH
Wa3G9Izgt4ijrjcOjIIidy/cxoETJWYfdWxH8eQhZwKnSROPil8Yay1vuonMvpcz
LUctyiouDr+DCLG7pg2o7Y5Do7dRxbaZGnjcnJLZciKYLCeYw1PzOXYlEbIDnqHq
o1iHN3HtO4p89QWbMH+DB5y3Zc5HusjIglWYF/UjpBVjGzb9Q+8P8ClynQ13EZxC
DKlstSuKjtduNnqBsdOtV6ZaMIViwSuMDXcJ3A5zK9TooiG4SdfKtWUlAPNoYQbq
Cd7dDYSTUe3SsdRfaoqF7h8njMZXdKjqwJDzt1MVI8DJjGmDVRDl4gSiTmf77dSr
weqO8bgc/m33OEbYgXolKD+2oE3LVXobvXmZWDW5/gI+tYhE/dSBim9jCrioI14f
UntDQauPpqlrIwzOkvm7cgyNVQCraUb+LwYGmWGhKvPpHfxfNYOyxlqatxi1xQbx
PDE6oSmzOzcZBbzGLW2BMeB4EhTKnMmPesx8b+lCGaWIMNAzSIT1ZgagtMy0z9ou
qYUY06YHofj9UV4BMYk6ph0o+spp5eKx28RHWUhZyxzVjjVzHCkqoww/VMc9OKY7
5Nngqg7F5Ttzzm4XMQGcm+2JZfRZ2LJkLQiEVM4RGZWT3KtvBPbuwezZCQ9fXqe8
wdCdyAJzpG+CNP97NeVFprs2k/MvAgCaazazCeuAsk+eduf2wCQS0pvjCfjsfkcT
0muxPCkWKzDY+RS5q9WWL2w6J4QRI6sruzRd6gNDhe/A/8MQWrclITiDroHmjTs1
kLwMwxsG8WTx1gz3c61J7Ma0OgWN7oXgaymSsnWWtUpxoRWhp7G/WGNSEheZFujX
mY05sXZGcfFVUFxR32ZsHgZKv3mrZKhzK2MO8WPH+w8fYA+BVHM+y/gA6Jq9Kc9l
2ybKR00F/iwEpCjzOmkqbRDqcj3mC+HaXaq1oLCjCLYECMB1EchpSt1rGull1DFO
3/+6kMC5N5Hl2PxPdI9TfcQAb5LPNsC2SEqzPUmpdeyNbUweBC4IQrOailffdJvB
TMTZOdZH0m3XWbqC/ltXmT00JUko0nbxnoEeIdaURdlJ1C71rtoWA9OQDkyY+5ME
XWMSiHLSsRdsLdomjYbuoiRGy5l4wmBAYmsmr7qwQCRECsLaqUzx+NsJNUu7OzPB
fE7xE16DOFwW3+4ZO6KDiiNu4fROeeXKdF98wW5+WBo+rev7+2Kv1WXpd5hGSAL9
GOmCdiyBGGV1/reHi0SUo/bW3aSv1AzurQXcEF2LMFfep55rTmJ1px7JlSVQkvCB
6H4qtrLI6oFu3zB9h3jJ1omz5nUcAlAinEZobvP33b05yKNQ2XXZHf1b1hKmFoir
R+7zlf99zxR2yyLqpL0td09nvPHsqlz5DzpT4umr8Siw3vsUevN7pPX0hiQVOJta
gKS+CK6Edepa6K2nVblWeVl6l4WUbzRjGvvgQM5DmF6Iwz1CEJAjSHYfBkY1wP0x
tWD0pZe2y8dG3ty3PvsSDTRK+xVh/XGj0sSKCGZjsw8rm4P4YTvAS/snYeEfCSKO
mLC0HpDeosHwRlC1FjN0WQvBy6JTiKj++i0RazoTbbA0eMU9D9nuDYDQfOBR7lFG
ZxlzoPapFokXU4mzSNbOhFa/2uHWQoGBMkAX8bWbghmPp2yyBpO6SXUvLx8Nkdxt
jG+V4cE6XO69mkAgb5bNF22VNBJTBnWVpVL5PidNxArnlQKtlqqp1ZXZlg+1X9hZ
Ds8EJ48O8zlNp7TxJPdKPfokcz+Td8Wfc2T5DHJNqmmVtMMQO1HGDlYE98a1dUSw
rdE4o/DTsASGUB+bLH9RNir5X20XtnSqFEE07/PPe4o1x0Te/xFI24lT3cez49Dh
YX7CAlXxLrMU+b+uCUEscR3Xeak5q/7um4+PPIq6HxZc2FGZHHXLBIpY6REh9xGA
tCbho+R0LQlj+HcGVEWdvpX1nVeiEBuw7W2sS/aMlOseuO5HzKCbY5v8/E3IWNg2
YH0xJLMflHiwnCgGt17raCA/FN+BlBv4m48OOyWGj+OJCQv30Mg6kTyBGRVWYmqf
bNu8ltFapAEOhC2A89NDZ61IbWuxLK09SUjyQ0cQ39rPpsh4LD53PBaOCRntJfga
pJ0K39g9uJR7BXOOwwUefg1I4Cz1BEmmE8vFWoxN8Q41D2yAL2i0dZMltGgRHWo+
8aVh9mv8mafwf0lrrJB3Zm82E3QmAS5Lz5mGTDLgOJ5OT+MzKc3l+sBEmdnjgasH
LM/bsbFBYFLYtNNIycXErX5/z7hHFu8G0PqjoaSqu6uNl0Zkb24DX3eU6oc2mT8d
oMaovFjjNB0zIOCicpDAWxDaoV/DjzWTdFA1HGAIkQRPrgBBahcV5cPkN7qIYjR/
nOF0eRXjR+9I7Mr3ffnFKSXenuT+DCW7C0fyRIr+oQCOCgJj91pfytR3EG+xmUeo
NLqEyYGUlGh9J8tutIt3iiPTrmM5OoMLSRtkz8aSeWgCvT9zMqTXp6PyV+YfhAd0
u4JsqNC0tEHw4NNbyEMCm5S5ZCF3JSpm3ZhtL0oLS0juCBMMsif9k0Sa5jJlDg4A
rMZxClOWlhFS2GVE1R7iDnv+m5o/OAPNmlUa79ZJzaexYzXhUQlmtzl2UnkrL4dK
T4eLQXqwnA4jSvxCW3CLgHUamT/qVN4v40wohPJUDPW2c0IK0WswpK9mHLoOO3vL
BTjk2PckWtMieMVWkWe0GRDJFT+AlF3hC9w6TvlMFPjD3B1a8LgZ3zZaq9Im+USv
s5cnlYpXuXbYavrgM0RGxlSaB3enueReGEmYZPA5JGVnfq6+pPKH3IKSAX69KNpS
/8xvZBAKKNAWR7If7xlInwkWaBbm4Cw1lPpbkEBu1QkQNeFCymHdP1r7WIkZdclB
E4G2RdnpMh20Ukn3ui4XhRcb6VjRaBU6RK8QcYlpmkZiq87E4QB6uRs1mY/HWekw
uQz1dMcRq5ratuMwpvBaOJP8/X+j2vurRzEFq7RrfczXRnfcTls86SFSqWDC4EjT
8Y+VqM7whRMG5aCLOXu0WV1259MSFEAVCM520AEynJUsI5OJvuBztMzBSr1ySeGW
/vz+sUFx++nGwBhF8hWoUH0JybYby6Znyqh8W0XU3ABzhRxETSR+ruWokoGn6cdf
sCJ0Qz5NIu4MqIgLAgmTS66zzqBdZsbY+OS+KB7uC1p9YZianFCNpMA+Jy5L+dex
Xpt1HlqJH8edjc2CUu87R8OhbUO/BOS1patWwtAHx1FiiHdWnfNkDfqaOVVvsonA
RwOdzsGmk8uKDPTWliNjJYyblgvoIt5ZLmyL5FHqjUnYxMtSPGktMyjlwPuDNZbp
CXPfAQCGiK/1Q1xatGpkcoNhQVBJBAZo8xftfNJD3zwp6pmiJdcU56yccRQ1Vm1h
mSwPaa/iVFWQHoVTPc0ifBg0I3FGciR/AdPIOGSPs/RangNaDIrem3qJiHya+vRq
tgeJO4oaD/dmXXUKIEq5RceNooBTE+A4nS9/HH2fMxcsXvKmvwCsZ+F9iVwF/lGS
MiHhqWDped8oZ2kd7BL9a8SWuVFTCkInWTj60Aa4hx6ic1y1ypVkMfJzufOlMRVH
AR7PUBeBNN0nu0mMHJaXwxPgmQamQ4zya1BVcfoeM2GTOUX9y2s5Zu9aq+qsv3cp
5mu1/0HPMRwJA57UpsfZdBhg/KI1hTAjUtgBfOwl+0VYD+I08OuF4fUfptw3lrqW
l1hOwSBEDDU1B6UNUQ3NtxMJ8+GIx+5WwZ8ilqaqmgEdCAibZEX3249ZscYRnkrN
T7Mgxl2Noa5FVRpihzR5rrZG1HXoxg3UFpvpMm9yooHmC9ZxegPyviZpSusk89+R
RmJT6Z8/HMVkCfP2tn6trCdBojX/Gg4f+QGbsj2EXLs7b2Dl/q8cNZLk2byqFxzy
YJ1kdBjqG6CWooYk4AERAWTijRYpvkR39Q+EuIEZJcdBQ1DrB/hvgI6S8pXHCiAn
Ie3+8vl4HpFIGNO+LxPT/eGC1PZZU0cXf7h+7l70sEU42BAERffs2DGzd+V+gmdW
+Z5HpotjB5PDEzp2gtOVg5n0GDzOlOwY/I6CP8nMGaT+r0cNvu+7bu+vM+TVPNaI
J/lwmvYtUzzJmdbm2I47Dk/Wd5pPyx6lQyWpz+sq8lR/INx0tVKNdl/5cpR7xopQ
ypSa6RiZ0ybrDudBS17X08HOuyVKKmurghov+/JX12YyhaOC+dVuK8oGFy8NGlq7
+V/Nvm4OhzPoUYMqTRMX1LxAd6jBuIbk/P1IsJRc/Z0awXgA8ShnONurXfofOtj6
zwMoPAkkiQfV3Y3NML8ooN7rFJunEQOlENt4uvMl0d08T7QHNOmYIPQtRWbvpcVa
pRROsZH+PUuUxNHh3UIxW7LdF8ojl1yg1WXx6bUBu4D8R6NpLhiDYmVFWeB3khan
5xTf06lMaQriQPERKQFcOwl6RYyrQ+EgRZhJ/EVONtOJ7/1HO1CAcX9bgOygS3Rm
kLVkdUWFpXGdKWsBmiRd+sInZxWLbgjizQG6mVh+e1NaVEukw3qqvjtC/5hHiLeA
M3oVV/YSG+SwzHOTk9AJCuQsboraNlgTdyYVatRILjWfIB6tiO6Eo7SVQProOy18
82UrYLtFIHCD7oSAhiKyS3mgMf5AoGayWGlNXCIqW0fJMUe9jm3JuaDyFwfmv/wK
3J0MUk30in55kyHiEUWmm1PkRtzxZdFQ5gKb/7TLBQayXCT5LXS8IF6ZzseBwOM/
5m0IkFDQCNrvjsvHTdouuemu/H1Ufbw2k3DHaxwlY4HGphdQJxapE6gwHhcqb9C5
D3IMeRCGdTB6ibuUndBA8IT4rYxYWF96PlUitEOIvHVqjk5B6qZDME0wPe/k7FK3
LkDKJkTZCLV/D/2aa5DsehmvP2IW41SkIaGbKlthDjEl4v7/IrmL+UoUeYrGVsLB
fBIdNQin4H02frZCkMjwoDyNyCu/AT0oFGkaii35KUSmsepxzLMj0o5ZVy8wn8YR
jaNfm+pdm68LYR2qn85a3IpcgoTc7isWz7VgW8i9DsfiMUR0V8NkWKSFXk/4DqpZ
hmpHHJyEcx6jsFFHV4Y0Lu0Z3w8ADlZi/oju7EwzKq1D9hnekv/8MiViMjtTo2sR
iscI2Hcr8J4pxCips54HpXY7aOGkhNNSaai41NNKoJq7jZWsvCXbIex0QrUgTDjW
9irAvvy7pvtW7lDZN526sQtTbaQdmRWWT0Tv7ipPFqlPPpBhx0Zf4DDyobIrqkja
RHXWByk0NAQLgE2baDQyFymEF43C8Kwe/PN66ZL8sNQLID+0eUiOtt16TPCUwJme
SMS9NbeJtQ6zz7DTSQDq7kpoTWe3Jc3Zm2yMq+umDxarsZORJfbe6c7/SkDNIP2i
jnolsepx/mCQUYUKZRXnxzvgo3/45hjvrS4RULqx5NLOr1FW1guseEay0GYk5lw/
HhIqdU+T9aO+ywY3i9zvt0saXSAsPW76s67+rvfZGUoMOSO71a7rZZqW3GlqByQ/
F+cmo6RvNwdsfxzIzSbMmwZLoXzHhBf7aSQ9XgbEoyQvJ6DN92tXl4LXGhTHd176
nRzj9piKpFXbedcQTekfNbF+tINuP5eYu8kySZa1yG5UqCrcsS3qb/DQgrVp5HMe
lXiO+ICx7c5KzhFriFWKELzuc1ggaI/szv+5B3GAlvrJC5jxO2Rndn0ohK5wZui1
X5KDN+5kBO0wyXvllzEH/T2BRMLVQCn9btHTX1KZp8w4hPJHNVdK47iJsiiGkELv
j2Rivd0KrJ8gUCGWQvfz6SgGx0IIoNzMsfr8IgnMVRPSJkqtXlna2gTXxIZUhp5U
wepX0adI9KHenYIMfZRVVchpitUOXrkdN3yUNg5WV4ahfFosh7lOmGR7lixLuKqP
n1IBrNwTIvvrAekhUr948s9XrdUZR1ft1LtvpIsmyLX4CNpI2DEQD5YH7JQe+tmI
n8C2y2+pmfTgEQ/efqixa5J4dx7jIeZo5BxVArkYpuglHLSSWPhbhsj4lhK7/A1m
wqBlnYVyTE/dHNuZzllbQAlAXaSFarndmQ0BVCbqqv6Ac/Ol+bVuAhRhE5ilIOQA
OZU30/8f32AM8gadiKnf24vqsVHu242FhN21T5ZAhzvNIh4L2cjXuOXfiU8ceMW7
xG8HfJCZw3LHsp3xiWnsf6X8kWMkm7BzmawfTsubE4oMjCqyZGGvD9BHl2eEW1wK
EemEGwYkNMtwqeYVk6LmCOIw9EcfzKKTODYNJFelmd+w3ftGV6xfeD9Lj7JasQk6
sLlSEZ028y2MHjcO/xWHThaax+7TTa1LUbCZl/QWyHR9jmphC3DdBUCiEz0YSEpv
uYZ6m08zUwPDJF58mOe7d2IX+w2oGwBdD800oUCJVhhOac1Mq+ViIbRkbZc/YXEu
52qwgoSoaNpzUMj5Eb4OLOhQDXOuhAMamXsvih1hqgtLc2zZ15crbHKdLd1ZU1Vc
I+h4Vhb1eqaXTX3rojKFbab0zLjZxaivzj7ABm1qanmoz3FxTujdtjEPYAjbuO9r
GFUf9uYjsinMiSjDg2NGTjIQgHJPng4blV3iYMMyVJdaI4hLbO1BpzEiBzG0P9l9
`pragma protect end_protected
