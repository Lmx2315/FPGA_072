// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.0std
// ALTERA_TIMESTAMP:Wed Apr 26 13:33:38 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
QukQRBz0S0W6z0fg8+LKZmZGYPWVdLSICPwH+5xTiHsPlMAzrE6DhEDfHVc3YX94
qgXQtoBHoJPVX1VvOuM+tx9ZPwcbceL1WBIb0uH2tJ80MUn6jQedtrIW1is71cHe
3NV6p8o7lacgBqCQqR+2n36cI3hs5D/iI2tEI7FGlAo=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 104704)
exWsiEv6xfGY2u/5GlUZiaqM3WK2lVbO7wcyYG3RH/iE8oCiIwjKK4ybIFv3MEvc
ZUMMQYYdZyv+8VbOmQI4DET2Z+h9aXqHYJnX0QbW1tONiciahwejKIS0wx5eqtdh
hnwRnRPaLc2596DHhMmbN+j1O0RsNHT4gpH7+Bk8kA76ZXI5vSVTUapCqc7ZmfRs
hgNao9n9/aQXAvdwMs1qBqPcJDVhfYcbUGFC5i0KGI00Hd78fCIpcNlzycr6tHwa
F3hFi88JwXMYjTvzWKhhCI6zFwtpMmSFqwGir+rtmx7CPunsgntRzkkU8nE4XwJd
ObTDf4wNMf4tu3fg0mz958XmHwQh4hKEaHxzrIUaYlBqjNeE75YD/AZgweUCmp8r
GuIH9N5Ka+bhIXbM2WcPn+WmZY+eVYO+ccvLw4mNNPzLFmD8aAmgDuXQfp1f7vR2
Rbrhr1dXQjJrdWi+7Uve4EIEAq4k1uO+pNqJ4WE/ByKVWhwSoH56M/CbYyERmHNR
l0m6p4JSUNXhvHR6CHYwrW6xzoLmsqRqaaKYHZJSkiniWlBsyPNq5gn7OUQKcoR8
S+yPf6qIfI3LwOp1giw7ZSy3O3AMJmOfU00c8GRfj8ll9yz0MmtIiEgzAbjFhoFn
1lqdPAkB10DjYMXo4NS0scojc/QTwtr2HrYWAtEvE1N3lx6zUzQpSrEMwh8qJxBv
hUCs/Jv+XmyhQUsoe2JQogEfSpxQa451KZCuQ0t+SYKiNSB8LEY0v3WRd5rr7isp
h2zvNfRvg3VbVDHQ7jMfSgn3/UUoQaWdmHrgbz49RRkcwlNWtfmqgd4xHdXe+kMp
cSsiV10yx0TxaDu7ci1a9xdssE0n3K4v8L5v4ZQMy+/c5Rq2XH6W1KaNKx2izDKi
/QtUqWDZwzBCRZ6ArQ7T4kPimS9u5Za2GcqmwDAww1uiuYF6nvwmvIxB2YiK4XJp
ms+QlCPLP96kQ24erQehkMimqWH2/zdvRizrRMFQFC01yOYWW8XDLcOMA0fDQ+cO
cSDM8aprEbuT2dx91VQDVGcI9wbQYTkkqSbJiu4ALRo/d4jGjvcyJE6fRimZnxcu
x/X0zLEKLhUK3zAshIAby5X6jc5qNUlVFicoQJzXo6hUkKqoZc9chPoA6O+/1bdl
qUDqYNwk4oKnhHgHNMiV0GqgzbFldh7qM7oK5F6cRomeFVx8gLQ7N3fw+zb/rzhj
SGAkI64XESR7j4fYxgl+fKFlqNr8R9CL90zxlnOL1+XoRFAyd/yHx2OOKrxHOYAO
whQqyksUuWVL5GiiKOavU2dOo+GOjtui9V/FC843up/E9PBktCDHwfVg/uUa5DGT
Hz0QNin+0Ju0REq4mjRCq8Zyk3j2s5HQjMcT0XI2RF+u1rgQfIZR2omd7Jvpojhf
m4bNpwTE6YNUMKhIG885/431nBRWOUcGDIxl2uIn2+BbEm9pv0MFmVNoEpCDlRL7
sX5nUNokQn7MG+wB83Fl2YXff1fPsDDRevlIhLN+xsA4LSlGThXvwQidRtpfyc7J
zupV3w53mb1sM9YVAnNqAtceL+2+qZ/XyIRi6Ri19p+0hDP+rx+zYMh/HVGxSCp5
3ui/RQVVeUBo8Uxy0olAjWfnK2hbIUTCLQSXeKinSglcRqkkZEp5rKpvkjIRE/Yb
rF3J+ltNIep3b9wqO9ZVXTf439da2iuWQplIKQnZcJrNDK1MQu7g9Con/36Nd6sf
VQbS7bGsA0VlKChBxJfSbO80s3sMl9lEu8+uC4wNXgDIA8aLzfnAAIROw0bjZi1R
iSGq0DFW4EkQbL93PMqZsS/9vwYtZCaQFspmICDwm8O+VQOcJ78MLTcBxHq4P7nQ
4pRpUtK7LXm9chAxtIHzHEk0Y7CleYQcn1wmOH3u02o0r461gHMDm/5NBHYO7gmF
viM4It31BLfJS3sfEKBj3GAmftygXSHJoDLq6rbPDlPBTF0KDz5YaVaklMdwAPYn
KCljOTATwn+3EVvmIv9A3Hx4+LUtKpzcvy8ynmr5pKG6Br0NVIyz0oL8jGvdagZ2
dy5FHygN3040sQnx4GwgtPQXjlSUqumds7yEGjqpYFGvUub67jHHHc7fyh5CGnDo
We/VZSf9v8b2wGCYvUaODXt4DJkhJaj15Y5K2kVigRnLfq9eJzclDYT6sWjJSdR8
DUmhY5qFJLeSCTanhOlytZLiwxB3q2n6467t5fflLahmHEYwDwStu1jPOPR31TvG
MGM5SyWso0JEeCRKKlmvYxI1f79gTuqU3B+vE8d0GuB8Mxn22Fv9LGfaVzjtX24p
GKjw+X38Tchx/tf+hj+/FzzsE2yQHZFcsxS4SEp90pogVGklm9ZoIJJy5/CDRxVW
xpb13nB2be+/pctQ7upzxofCPbDFGLqcptJDSJ7E31YFk6CC2cqELlsB93uTRFin
hYJunzwU/2+qduv5H3K2pb3eNdSYtTq9oqFWW0BHu7KRhERwtHEF+JnXOB/WZQP+
TH0+16sIbFwailCKgN4NJyPSyhvFcc/Rt04zoOVHboBb34i+md1sBirTOCKx/gGy
XbLyIDj6cDAtVO/BseZZnBZbdAGnFFIepaL/jP6azUaziYQOe2oKMtQRBfGnvCZQ
ZxVBhqACqcVOnRMQV+cZHvMH5i7UazzUJo1YR9M5GTMGyA4iAskdgos5jZmaKhLe
Fk5WNU9nJIe6vCcWmgZ8Ys9Q7/1P8ADkOy5yPzeMr1fAng/ee5Ml/WUZFr8hoAb2
z483diZvfrtchepl6N/RMDZB1JDoFPUytVCYUppkuYY9bzWTN3niU/Pj0zJvLC+7
VVUBbClTsOtcbHGnScQ4g+1uLfvL2OvoyoOmcblFxCmxq7LpD4pC8phvHL/hn+Ki
LWMR8YZRk2L3m6o1dY6P4nQhDBmdtklglu1gg4y+xejp77C5nIMByWWcHG9jJIZS
xI+r+KTmk/BPUgT3sUM+c3JPc/VLK8fUOK9nMIGGgbvjPPfTAym8joroYRs8mMab
p91RDKy6SIv/NGCOpjzW/HIQi8eSTXCk8+As7zQbjdUaC+7s46a/cPoVG7UgK/Pd
ieDjj4HpIyvtU/TAx1Y2ZgL2Z8qr3A2LMEZQnIlTDfFTdZYyqJs9E+B7dCW7TFDx
KiBy5cM4nBSqPjNqP69LnwUNodqltFx23s9906xG4YXMu5qldjxTqWDmktg/GJDx
et7oKwOpVVEqaMOXEDs/XpCP5jS1LZ8v8noDN6ZduJSZ2BF9kRpCytPDCtj13H5q
zeutkWx45x/r6bF8/ZUaiieclwuLKIu1jup0Hz8KooRMlLQ27fbshTtigzY05iDa
zOjr9QoLnbiafLV7sqqz4AlIu/qCCxQQCqcJUQK17dXj/ktITrPA/m5u/YJKjcd4
8g5gbI2bOYZ/PNl+6toJBvJyjQuzNMfYNolqrxAwj66bLwoH0EYHm0asu9yAsUdW
HEsMGUc1xHrHgXtMddAyXuXWTol6kDFnCRUO43TMDzVJ+jlmxNiHUa0YuBVShUb9
7mfzHTHWcdu5Ii2kQS658JHUlRPEnDyCoKkoGFwyFxsMrBzAvj2ATckoWm+yVmyQ
YZhZ4GcVLVzWbuIcV+iqAwZFy5lGeESFAOG32ZyhzfTvuQckuxeslBfgoBjnWjFD
b3CTHvaKLZX8d/2H3ihLj2wIDAtwDscwTuVuYGE1WgGw9ZCJ6VxbQ2V/PlLT07v0
YHlB6aHgtKVLjOnnta04suWIBE2EjYrnKI2AXOGkqKO7HWNvJYOLqEBszuJu7zPL
75sgnf9+gYw+fcfwwlPryHKo9s3Aevk4Zq53xwrYwXqfzyuuJRXAiHrZt+3T2/yf
hO/u45w4lCn7vXx7nJCZ/+hgYyAZAlsUnKB70r4Z97EpkxMzMfCViZ3wII3BH9jU
v3PjnQdtk3/+8i9OzeK7G5ThnLYDgeh4Iu/As9h3cdfxOUnBu1ty6dIflqli1eyz
y0ghUcgpeRHRzyEuhDM3CMQqWflvtYmacwCzDNDvKGcuxyeiQkEQbH4EFHvYZPX7
DztCON1vcN1/Q77xY/0mn0PrNRMg/HmUMyuuAB5wkoyQR9iM5yc1umPVM69k3LiS
VafwMr4S0Wi5U6pngbGoTdNZJ4Gkl5BI+QtYfXdfGbryEcVmtK6zEXqaKGje9OFW
Br95NzpexBIBORy//AQX02A1fFPdeNFNBwKqsDjiWmbo/eXKd+MsgsKW0+ufatyY
fBvTUxe5hptaZfbdMwFqhaWIaRLNDQfiH69ZL6d0jcmBJ8ZAoDf22BifcvKYxvnR
/Ao7xw4jRvKcmt2J3xPkg/aSYFLPt3PxX0U5KWHxz1Wh318JZNYaxQwmiqPZt5gu
uN16HDQ2mr6XTnImSb2o441GX4CCqthNkDc6K6p8VCJKcvTIxCXGTBpfkeDM9B1D
7ZYFMO6XFaC0gp8oU3b4aQfKss0/7mhKrtorFVHt2k0iEfAAKoyCTYCxYD9gDc6B
jDLulct5sYXz8hPG6z2xasPy1UgV22l4FjWBIykrLScBWaUQ+xMYiiyk1GOJSGeB
+l6JXFFy8VS+bmlz0wLzWBfF2tz7gHNJDD/Dbm7ujJVVNKvYXVjCaZCelf3ONayU
w6tIrFJulhqvLtz2FpdQkGB0/kNCR3EOuu1n5UqW5ABR4Sgd3KF+pMu0fxHL1x4V
bFBW5+pZeaa/pehxobXDDvtQBjbUH/Liqvr1H3c63nk0sbFo8iIyRefW0l4jx2Vk
irtcnqzo5NJsAwaxS+rF7xuhoKV1xRW9jSFznhQJzpaEeQoz0KzoMj/oVkAOcDzy
dsgmMay92AqdqqAA1y+2UAydReShFVsVVix9MATcoGzKkwv/EN7fqMk8nCt2b4a5
iLfIWu2NtQp5pp/TmdNM3RzL6Ffn6xNwDnJCp6lDpU1uzho3nWNmfayEOWmXxSZz
W+v89L4wRsoi9EHGJlr6PIhblAQcoYGvOl3H+t7a0r0g4Y/CAAj5pAHHMn6nsDm7
036uJqGxF1S1I611/YLxartzTjn/tbc/qhbD+FElbEYhPvXYG70AdaVpSHguVaky
zyHZwCVmggiDzgxMK1F0ap9YRfThXApcy5hCo25sia+K9+6a+/stb/dOGly8aOPf
HUYX1tHRfVdQMKoMny6i+Tc3Sch2n1+IxTulrUnOHNKUt0NJQ0PQvKmtdodpVOKu
offBo8lA7fMMNOesrEQRvfn1r6TTm5/SpYyEYEyYwo30tvoLaNXNQkiHuQVSmBZ8
O4SySdqiAXVpjKIOUdjQeJ9r0JT70I7ra3bT5faOGbHjk+YQJZZBJeQJ4fo2Ui/w
/GIByvZylEeKHbg52G35hdDpLqZ0GapyTp/0oaa/BkXiryJQfBitBH7qKiaoDcSp
+TaoJZQ7FfukRY+xO8x4eK0uYUXrR2GvFBs54fujnU5q7mar+PkPpb6JynQrERL2
gY3uV+xPEAk51cTJTmEhlhCWylGYCpumqF/CWbrqbRtneg/z6CpeXPlij3E9tNYa
s+fIvS4vqk94LVGiqYaCn1w+NRVch9JjiFDBJR3b9FhFch0BQ1MvwgTXZNgS5dxS
1dfn+yMdA/wCg4kW1D/iaZNdoV9vX/E9cMV8LbPbdJsaoVVUWgU0JqK4Uios+fNq
nL8N4ZsKvFi+lTeTAJ26XQXSER7EX/XlkesEw7aM6QkgvKOgMm1CKef+iGYCOgAJ
yhB/cPYLYcDc86ODtxI6u56xM5tGe3tP1dDqKjwt1eL/cJ2TC8xSzGuhBMowewIi
2DQ46zL5CNP7WnNmvgLA5zR/sEmRCqTweykzUyzuftvA5Vxkv2WeB6JRyoCmwSzm
IurIztK/mYDbzfoKpwT0i0ApJAJSATYDl8IUf5MwDWMzNyI2pdnashSO0DKiQLMe
BCDxs1lFn2LpQkX6wYQVSaIu7yFfcD7wSPLN7sW9mDugj0UMkTymZgWrUKY4D8w5
M8EzOJZUExwOf8QnE+clgTgCph8LTWmDYBA4ocQDH/Qio3oLHkLv59xKCr7xA/70
F7eK+PkUfRK+RwxiSaX8OePJqQ1qrxx9DwRa0YASizuC01vDVEoW8OsE0iZXNtNT
eudyjcu3KwyNyP6do40AdfShPfoVLL230aV3/pkapCJ8d71ZdECMiPAlGmsInt5e
5KpHoPbYrHWAPhNZRcYGAIMsKEzMcPd9zdr+YDuQFG63hOZAFWGJ08fIZF0Vp1D+
fGc79Lbge0QG2xXxJHJEXnLr7RPnUbs4v2ZLh2FTv6hFxnZCVoAEe3sQwlWmkhLk
ixLGRWu9zJ1bk+Dts+Seo5/5JQ0bnNTjh6m3AX1PZXXnNWx/9qPvZvs+UNb0Nlzw
+59SAPmvYeoGKVpOedKtpmfaPI23QSYsF4mjiOdIUcbyEgN/oQRZZ5L/NoGGs1ME
T4rgyRUNlRz9y7Dwuv60XfJu/Xu61O7KHqahbRRB9MMFqnOrMe8kJeCsF+cNpi0b
Dm471AikJ86F+puh0DxG9jbSz8Qs/k5XW+eylsxyZs32BCazkg+a7vmxn8vlFK99
CX2U7oG5Kg8ZIotzpZUZqqxWjFUWkzQ0PNxa79tBt9VaaqLc3C/O/tVU4QxXD7ZQ
gapTFP0WNyvG/2i4OJ0TwQrmV5N6YZ8L50yP8kLDN0NsjBc8xS9RbGFgpkGkdQRV
2x7Ui7asSA9xP6YCluLpxTWUq1v0Hae5hcR34KnmHcLCN8L3ZOcTHan3JiQ8vLTh
zmmj5zAjmkR5JrP8upELI+DrkN10ipPAo7O60sPsixk9EyeHm9dqWtkuOm86H69D
NsxN6qxMXiMna++IsDD2zh4VtptbXldSTD3B50nS9eQ1O8cCmhLvCjqAJnbb21HK
BXHfTj/YoagZOTy7C7kCu6TSVqr+njRuHUXw13cIl06gIa4YAtJK68DuDkXeEDRb
G5za5QHOBlUGNe4UcdZy+PuGhKmGZzXqMypuyd3Z7QypsY29tQXXHoAh+Crs6gaM
TpSncByDi9wDl1tRLYMJ2OTv6+vkBBSwUXAW4Z3/dwgbE4dVgzZVE9wskZ+Cmprw
wFljbD2nsvePSu3MAyFyCJMzpaMhSWXyH1DEZtVgJDbTsZKoHK84sIXVK/sKqI4B
2RlM33ERjSaqbxvvX9fGOcmdpTEcx+D0GZ7Ff0Bp5fQUbuwODXAHyy/XUHLi+Tjp
3sSKcw0gtQLgR7tJSO+XLf+a3fnn/Bq1nk/g8/TBAKtDuOy8dDTr5HG4YhZo4mYB
tlj+LcOIUY7AfgE22jT3tv+7oMZ1P+4wj6ue5+82MAmsDYhLSWa+u8syYTCqvjx3
Nq48BPOCjlW4WHjfpgLelD9PjIeo2Gi2wVSH3lYNnVeimGPKzGvgNCsmdIoHdty5
zFcQOcWc65bcW80BTnyePbF6WPh5nmxEXbMUImXN1pmIzkmoSrw08XEGE87uGKBE
xoKFtknlAHLGJr5Jr452xCjAW3L4s3fc3XRZoV4M+J94poAPHz0CuEbhkQB5O6G0
ui45qjRnKYtDMFeu0v/PjKaocTzA6otLtJX6SRud7IOeJhRMNM4FsZYfVtNCxZRA
2MFZtdcIU/tetUCW0RD2HqcutxGoGdZCUoj1qyzXFJ47WHltMqXZa2moSpm1OZ2H
9CIeB2Il/WXUgD8sEO3ZDi2ildzFkR8o3O0aJr1RWu3jF4aDzyH6YtnuLoI9Qw/4
XEaBuZ+wd8aiVXUTS9RrrSDGCRWvH5Sd3uBe3G++yosyasijbH3c285WQXyzkPNe
J5ptyKvq8m0aQkS/mSdu4K2qO3/nGHxX+i/DvoSheNCCwi0Aq+L5/kMlrZf+gB/Z
Ny/60MiLQSzmb6TEYzYssr9DQ/ijytZBzEiKsW82b7wZ3E6PJENO9xZSEVySpMBy
8Qkil8XQ9H4WOYx+Bvbfs43Hbfm7T+oQOxwV/M9cHmRtpMgZCippL4/0OUTCKxDf
4JmgiHLi0duD+8ZN38EBBWapJSQ73FwKflppLfbCCucyoHMrUV2cB7JWSdus0xoa
4bTo90SoVoe0+RFYmDZzUWvC3tC3DJ9xYCKKxASdNlYnlt2PeA4Kcf+dgm7FGk8h
w2NWcSTZHMKRudAZx4+wLwkyWM+dp+9OZbKjp0KEsHTdiT9QxZjLJ7Ve3l/WV0Pm
sKj+IM1t/Zxa2mnBLiuJSWfDDwZBxyihUWz1vUsWys/7JBJXMRMccJI+ifuZu3r9
+x1XpS3B6BqpoHJRjlJjWbvLS3EWKpJ3ahX8FLmdTDqrKnVrvvV2pQj1Mk/3xNa1
ZDuoT/TgZ/4XVOwrYtpsZXKV5YikRPWrV2KwhmjvRf5tA/vQBw1dxKPya6SeWa3g
s1b4gJaGpK0tuUtTY4Z7lRKQFZ2x/BvKE7CuM6EQ0wEWAX7o7YVNSqKw8l56kmzt
fwo/kVyoW9eoAui8SQP4FCEOmOl5m66OaThEgnVHmPllxfEizebsUllwQbjIPzTl
qZpJnjJRTf0U2hccogZWl/AknUp68MkdJVe22hAPmKGKed6r9OFIyVGsA/dTdlQX
I9e54YFy0TgVDGeJb1rxwvGkrRWqqHdM75ltsLA03r6DAMi9U+upE9ea4aTV2Qtj
Ii2BfRJpO3zqLWGs3eHE396wTTTYNM8fzXotzBkkeY6bOLpG2sZIqJWXIKrvaeQ5
UXl1dAW9STm7TcIeVnh/YZLe7e2thbAoIwIBK2Q92P2xNzQYUXBwsIlSmP5QAXfj
xPoRZ9fplBuk7dTl/5MN1DW748Kks0PjlzP4GEkRqWbzSBHYmRdb3OPdP4tAqoqn
dwRmurw+L/7SMM9g3vclXBzxJb0SQL4tWsbGs5sWEiXJbCs97KU5IBfGOK0lPXr5
A6LRfuhBErv0ihRo7GOanmZIgkz4YeV/DLw4nFvNWvPXwA4z9Tq7dR/jJZIXH5eQ
3IcYKEprjO2bJENIPY08WfWZnBXXaoQLszMzD1K/QBOv5XdVzMjpptWZfRO/+k8O
WCSUlzAiFUmmkYWlnKcVa9eS2GR7J9Ky3bBBeIMjYDq3l0YXrZoJC2nqX7PLrZOL
eiKbb+TjsZ83Hx89An86ybbiquInKZmeY120VI7ePG3ImqLuhxxy1iS0bhfzdDyg
EJxzMjJ+lv5IbqyijnaBG7HGkAoAmBa46eZlvzwDDXGugIMxKp9lNAHseyD15uBL
9PnHaXDs/2YbZedr+6oHBKuxYXhAqnJOrdF/fmwjXfk9YeAk0WlI+2cGCPsH0WQ2
QBilXGI97ezkgqN14RTNfnY7gOXsJ53lLan2YHCeCJec6DzE2vvlNWIbJI5CS9jq
N713tZZPX9AO+wQGaZTgtJnqm0qHng8aBCxSkyQPLIJe+DQT9utoNJNEzPQEaI5u
C9RIkfFb+H7AC/c8PzwiqNg1t0FafbikjkFFsykXGXQyBwFjJV0A+ZJ6/PZC4tiR
L2nz260rWY3FNkbTiRF6N6YrsV4GCIsg4OV27TFh5xRmlKKqDTkPG6rL4dinxmP+
Wwu2bpodIMxIsqe3xXTA+ZuD0g74uDhD90geTGjeuKa5/adyh1oC+SVTL6p6a5Uj
CSKCfAguwqUFmNLTFkjY+6s4JBruvVSA5P2HxvIRSGf39GNhm4gqSfOjNvFFwoNe
yzXqU4FNZjRZhv3fmfIyvTqa5KHITDhCA79IhQfy4LXqJiMQv+4KFBpIvvK08cQp
eQhriCmftXJDy+BeffsW8EvV99T9F/Hbd4rLvAZcqhLvUizpKoBVCwiGg49IZS53
hi257Xa19JPPELmSN/MAhDY/lhk0iWy/FSUGbIUEJ63y61O1iig+mMdvuG0V9bLD
AADRhO3Z8nsMHCwOXrdRTPyd9XjWQ5CP2d1KlJwYZMShD2IpIjijwpkco8YQYVjT
KI6BSlTyFytF1K2M69lTU6POnyS6nSg4DUxI6dUuEaPhxxX3GxYwiQOlVZ/bzl5q
EsPzruZ2AO8Y0csqOO0VP29WzyiNW2DIA6XY5qRMBp9PrjfX9DHRIbiTo75n1QSo
CFj+RqUt+E6kIfLh4I+HFi+hgvrsAAMDIMAaRAVn2yJoEj2Ijn5hdr8OyG5uXME4
4hrm2tjj458yRcWKuN0/PpM1olBq3GPg0te2ugdUFrLHfzCuAOjoAJvDgfx2N/lq
Du2Z0acxm9PckU7sTwJJioiia0VWzbWV41Qobh/fUWGCT3to6qvkTb+MT7Y9ANDS
qgEhWZo+G8shodNrAMlkYFL9knqHn80zX9gsLX5nsXi/HYrQyot+8ZjMSHTQzYiE
DCRbxASYX9CAHRphMje3iPT+mxADbqVsO5EFW28hpUziXHnGBFSpRQ9ql9l+fz03
VvL1b5CBmXlEnQG05i+GV7hk2tHywvLyE1bl62W26aMtgdm4e7qUqVMO6B/4GTnU
MQsjmtlfKpzzEN4DfeXf8OvGEgkJ6KrbF8u7+JmC9C218xqzN3/739ToCH4/XHuf
jYqpzdQnD5QCqJeE7kVdIyG0b+oqejoYLNCRTylHuS6F0xLR8Rloq8mpyhIRiOTY
qWh9Dk/ENC8heKNRbwxoSy9j8F8ImjA+bC08vZWmBRPkCIOoQBxQyZkR5hrsB2TM
Fone0M/PsN/Z5jz4ByhNz2ymZeVCO3gr4Vo6W4H5U8NEcruyRT/qQyFvfWZBKrPR
n8sXrjbCTmR5/pKb0CPKipJamrx2GFbkgn71Lm10fnEG31qsoP6OQL4Xl7PCIm4O
sb4SFLXnD4hdXhOJW8AU633YZ+QwloOiNtr0KdrceqCusa1+fYpNsZ2bPG0l+IQU
MtUiW/1dHC8u3RM05OP0Hneu0ZLaztAOvZ1V6v0FG8vYV9P9dmeKmw0g8i4fWIIv
vrB2/tm8BGblAW9U3Xo2ryc/jOB522KpqMLJcrWrqgkPYJjN0hUvQtt/n/CAcBf2
46RsCBYhsQWqoB2JynGQgqKD/t44otJtWuIBF/HroM+csWGs6DiG+SPg5UAAk73e
NFnbXZRvqg5ZALvjS6jU26Od4DKoJ5iY5h5ggDOc2zFFJznEiVPiPbG1bprY1xvl
4sKqQYXjDMseaY2THiFEjKBtspG5QqSkiiNoHCV6QOUxA+qAACobjCbKGQFVM67D
ot45DiLUzxUl57ILfwbRV4YueMuKLmaSQRDx7M0BLZ/qvr9DYT1XkBCHq5w1p+aY
b7YrCEXRMBhEICmNUxpzqR5V1U2JHG8RrHAqPp5uv3KkFXtNcOMuuNOj1Ka0sc1L
3cbPeV2mdfwh7InaHmh9YU+zUXKsPM6+ELicc6XQoouYlKdy+n7OjeCBvjmS0TDb
eVG25Cj1MPIx90sqj413sKsltBSgtvOhvoFnVCrPEF8vzExBFfFTWBqG+lQxtnnG
8B7nDMha8fc5MpUZNzWITNgaguA/mDv3+vmWpe2+WOqqVeN1YN/A2AKEcm3hVK81
upci0IdKmGRa7jOylIUL67yrcRbrWPq5/dJGLlij3fyxgnOBP30zrnvEOhAO/lEY
PKMVHpVL7gVYKxLAty8+QACp8s3t3hlkB2y6tNWPDBW2nF7DGgJCtIIwx2IkPRrD
wXXJaEizW3hmXG1rBRyiwgDg/WoIN9hqJD2R8gIRKdmssMNIcY9e7VM1GyJncR6t
LaFPQjwpvdLgWl9aWMvAZign7r5ToGHg8Oe7BlpggEhyvlh+tS9xOUDeXNtySHmU
jyxocz8nm6qI4ttCJjFEBjJed9/1mVT9mEXytYj9B7RMM/iS0E5Tb/xh4U2MnicF
0iv/s61Q8tD7Pk6bi9iVGBhm6Yo3y+BhGniITezyXwElhZYcEGFe0W+mEOnBHNK6
b/vAcCqYp4y2lFLdmJdv0NJOZRyRMSg05S7ApVaGQDSLyebvfWQp+o8f5bfu3Fmm
Jtq14qJdg85cI5XqRarlYKet+TBGnl65qjbXhyuLD4Y5f2bW8rH4KD8sgPZ8CKGo
Q02kppTQxRQXf2gHbvhMlyFMIbexu+1ERwjqUDDg73p7SEUEMDLPHDFuOZSg+eWR
TxMtDf6EMdycmKz+doYyg60+g+/A/GrMZPn7B8OAcL2CcHMOn9J4NedLodJVj1W8
AHfSEw/7FVLs+QGLzTer34bZDul4jcsY+NJmsjZGzJn+bAHqLFwZgw2p54X+oVzq
KxJYwcWBq+iVHtg0V4UuqsMNoAa/z4CP2ptEWKdIzYqIScf6XkQe5ChHwhwefBw9
iWxvV3Td3+etjam3cQnhcdjBi8KxDDu5FRxRM53itX/hMAHxB+mNYlw8J0wF0bMO
xE4ITBjB0f8sNzcxjMu42nbUz7mV8O1uaGUOl8f4FHqFuIXulolJ6zhzjFNAIrNp
ZDAewK9X8jnGd8iw0h3vGY8QQoUlvUJN7xziUsYkuPqRAEVMhpuuYnkMTjgQzdUW
KvU3JfxYLGgKjtflfcI+ubw+tDoan081xxheePHRU8NIUw1dUfQyXyxPAnVwBruZ
oNsMSz//LclcAhUkxeDfHmX0CO01g3vyn5Ixwz5ZezvufwLb8/bZbqcqX0LEECL8
QRdeDu0UIM1g4cePsyc4vczaq3fm7wMZZcSID7IQhDkQVn9vhetWnCiq/MHJ1XbS
4u4K76Tcu2zQRmlsECsCrt984UVAwnXKuiL55JzrdhMjIEo3cESOGbdwdmZUkyWZ
drE3n+Dmy2ex4hA9T1ifpjo9rfjZJkfxaWrqETmh8cKLPUDpmOmPykaw73WuEyXF
ZIDqB3d7B9K9t4jmF7CwT/pmEJNT9CpXrdu/L+WQidlg8uM1d3lABQ3tURXMNSAA
8GDI1+S/+Qzrek5toUyAvi6aanN+faEF6VPvex1Z01wLLhm0H5w8uZjDIvNK2+MF
LW7EzeyXymCCsMe+2T8BD2Ko884i0sE/1w89/jflRBdt2VONp/l9XCpuAeckgjwP
zR+30Xh0kfUZa4qtD9Dz8qCH/efS4RNl3Xq3Gm1okrE6Wp0/wZl54Bv0XsdQZHsB
qjV48Eq7cJfIHCj5G5rnsD3WG40/WL4VvumnIE+zXrZFFqbxgK7UhGSb6v0Yt4H2
69XfKSBFp+XwzBcvg5bKMy7kpL2isiihk6wvJCojoRQnPpsi7iqFOTzBy6EN+sYz
9omThWgzJTyFRuVq8VofSc1E1o5Rxv7vWj0U6sy1BUN0BxhLwzwu34l8/heJCYNg
JKGQdFgwEiFAe9oyupov0mHPgZztQYlWEUHATH8zMxPHxJRD1j325Rz5letZGvHN
2B8bB05c0ypBCY1fQjTK8Wdb3i0NmNCLo14KDmRgxvCmz7xOJKPysp9IIf5XRsBz
2XqY+3MwRS2ODujDiChxy+IcsynzrFQB5dUvUYCUgyVN2x91Yi2viu4wmKPWpgId
OkzAC6YrywjQB2fh0ZK7wY6mGD8qHXYSRJJlnkEZZu0oObhwXsXu66Xr/uPy6L9+
pZ0CxNIhSd92iVIB/nlTB7EtYSXNj91P0B+/kYCONz/OZ2J7AzpcFfwvPglmiP9v
w73mbX9rpMv5+uEZZLdM39nWK/OURtYt2qOXTYzcWVM/rUQDwc0P2FakiB6SFwIp
N2JTZCLcdxJUfrrPPD09zbweAbq2nWix8er6XqFo5sDUHtAZF5WgpsDZgcDLts4v
cLHIHHxGZNz5UCgJ2hU0VXLEavY2ayyaBWYHFzuDaMXniObtEtwdqocRX7yjbvRX
TJ6SuFhtfP8Ba8vgzvy8wMhWD5ank44We3t+fT1VFDeWj8++US/B0pqltYS/XHT5
tldrHhnHA6uAILbuSJgcoQF1xxbGE95tUzB2P59qcU4miJsJyuWOmMZtCgswLsd7
3PNEjQAdi7TntYf9sMgWQ7qvexOw1tfl5F2qIFKQzm4Qny4C8zAJCwha3oBi5j9L
LcdAUHLSRrzdtN9KTlbpbMcGFRUtLL8spH+VokB+FcgqEArX7Y7j1cgOWgDNmW+p
gSBMI3cIm2c72NxWv63lRHKkDh/ZzzQcZgF5O2+Xz3NHPfeVvNrWsddTn14KCSV9
aGe46l8mYDvm6kf5H7PhFxXKQNtCXutV7yWupA+BcuKLV6vQSA3JL6uniwOLcn9H
hPQ2OUdQsQGDX9P2dLTLpyFqwmKJMGH3FNnnmId/GvxHatdz7IMjb3ddlgnN9orD
1uIFhl/DvYN4F+d58VFLh8tqvOnySbdsPWt3gDyWp8ydojnytdoJvhpEKoqZgFoV
LFWvo9XizMagsO+R226yZ4MunqpFDPNluAQxrja6xP53nmf70tX45bbdZDc0Iqr8
5s2jbNV9iP2HVuyEkW6rfWc2P4gmsoOXuXbbxMTVEnRHvTvmAxi513AnR2Z4RGSu
sI96VMq60eqkeDtFxUqwh17Fq/pFmDqK7sYUytp79CPZZ+g9Miw7BhSpUsgUmsuj
6yRJzYL/BS7X3svfS2JVnDrinV3SninOkcskfzzQqIlw7vlTh0Fdx8+W49K6mWsO
ktQzm3uLk7ybQWg+uhl6//WBuJr54XaUh7M0f9L27nX4KXaR/HIPSckZhe8vT7GB
QcKGqmaU8ZiD4ubEu3WDQMSKsuYoEplg1uU6wcAhQdADy05/BHMnr4EJi9ygfxUZ
HcRbLJYHSC8Imzw6YBi7jGutmuu2pwZlDPAEYRuJOFF7xUWJaV78CbXcc9IwWrYW
cYzryLgJ1kFCdg/+1tgLL1RtwEbKGI0jbSgeJiJBBr8B5tkWKC3IFYKIrXs77JSf
tp2yLIdjGkrT3goHmakuV7GuKpWP1yD/0QnL9rinXCb8hfclqCg7EsWOs4zzXY+t
THazoH9Xr0SoSosOdOdcLo60bntunl4Ma+OBRPwRJi6+jh9y5gWZOm7/D+QSzstl
g30mPm/ovi2U7H4gFB2NMhmE3IYR8NyhpFYObQxQsrdPJVG1Ow7HL7Lu0QXTMw06
zmnTq0hupWpx64BiD4qIv7UDwPD/9bEnwKbi7WuBbiLk64uwuynH+jk0EyKXvngX
wICdYh0MXRG65tHEvMUUnvvSmoHP4S6vNnpZlw1b+cGN1v4JZlJlh/zlKQ8eQDIh
YjPJqpaUZ/px2lIbp936X7ZqwYkf3zCS7kxJgpGa8tofVe3gm9XdEGIAiBQfwUax
Djr6lINQdRabVgpN1nO98G8GRkI3Q/yuf32WZv/g4MNPX6eRj8yy4CBfO/XYwTiQ
cYA9ONsvGH256Dgu4qcUPatQ7iYQJJtzEA+rOvnZd9Be6tw9bm3lKHUGrwlj4WjS
54wSF17ArKpmwWTiT9EQMdoCIZKZWEhg4IqYbwu8i2GnVdEZeGpZM9aNHcs9K0RJ
dhfiDgWL/mJjQdC6Wyuayn8brnfFsguxZccPclxdhco/maBM+YTu3KnL+5kYcwTu
dLk3YOz0iVOsE+HJghUZOURx0i0sO6Oh5FnhIrSgJamV6Omk6UtNRpAPNAKZwP8w
0nHOMAr+rAIW7A/I7guklzQTt81EgmWsI1fF8PF9hwkkpR8HLUUbMHOEodgKhk0i
cGoV4nysyqSTC0t+BN+nFAPV0nbHUqjJWQL1A/VRMaG3Zr1VRE7skwjANgcrsywa
iqDuVjbnReyUBaU4Fe+DT9EX8aEjAJQpQB+yDnwK3jMVj/RIXUiDQ8vosf9MINDJ
ZT1HOdmHnq4j9AC+Y7aGHB10UjMrJbfuaNG2V7wf1GA4gqYXTmlEZl2IR5h3SIeg
s2Wen7D1XNv3xokNrjTqUCVd6CjO9g999nkmEogkKbdOb/zS54/eDK9cJzmZpZjb
3c2mkhAeIAbgJLxKnF+b38lXpCLdVVzrcGHUmziKBOcwzBOdhBowPSf5DIn5St3x
5J9A90JKePp+Jay4cAVRwyxECQ5z6osBTtPhWCRM5DB5iRpFjkDNksYm82L2Yp6o
Surq/AfGmbqUok/s++zGKtenE4DsldsiGUllLhcjP1aivF8k7k2jWQCq/9oSo1FD
aNeB+7V7PVytFJ3znxbCkPELfO8gDVuKF605ugm2ZxGwNbY6V/60d2SXuG1B7V1Q
kulmYpvaEnWp8NmESXuM5dlWI4C8ova5MHZCz8/9CTxCnfiZDBPwAmO3sjrkG8C6
zKHxLQxOeSFolmpI7+bvqenw8uSdDLvPDDygA1tJIZF9QS3trF7Wk6zbBvC/mPWC
4rUcUdNWSqBnY99yJlUbBMEyuFJSNSpUbC0fjjzUSo4splx6Xmh+EEK0CIudvQLM
i1M4QvVhY7tvIDNflIXhUbeP6LVhHP0wncsVLZIuyrToRn+Lc0+Dg06mEyHXlhOQ
neMNxR6CzVRtNbtStqBq+kIHYpa+sfYZVbN3st4eSC3CldOFxbrIF/VgCpdF3l1K
sEnxKxG8/Uo31nE7Io95WKVO5lF9XBK6LezqnCszIyREdtX48EyglpbTo4nLjeTl
ZiH2O/xJB7sx2mg96+bfVurZzRCpOzuI4jJ55+upZttcKlE7fuRmRbxQUtyct03+
ugSPB+isbwB+4u3cYXMGDodUVFvwvDnyrmPHJ6dg6d4oP3gRUzSWofiI/Zsy8Lgf
/T4/KEdSmKFRghsZKRTXliW98ufj5J4sqW+JwjRP0CCJUZzJ8QYVXgQcX+oRTyht
TsTNtwfNIBaNYjfuWEZFQD7VE64sGlP6WKz2am8hCZsgT9eKQr4+EyVyYRbeGfR9
aQKu0yvIjV7U+4wU7N9cZZPKQZLID8VdBd1gDXOAQSoYntT9LNcWH2bTHs8yc7YU
sKi6rWfK/U711PhOZpsFf8Ko3CHIR99zhbH24/xe/wNnMUTfKi7a+QH2ExSkaB6C
lENqN0Jjo6cY/83K1jhlRmf/eejSPPQ/mR1AZzjIH3lp3B6FvE5w7CfcDMaU2Ts+
CQdy692J3vUBH0qMtyBZAGSFgPUDLaFcea6BfMCbT6mf9St4y3fjMWt7zZPuAsK+
WsXQbuOba5GbmICAx2lh7R3QFJO2jiudqiHNHb9TbP9aiIdn+aqCYpuUpaFEd8O3
wNSpbiL/WXEufw6Kl0QazCSi96x6sD/L1lJNiWEybD7Nnx6WmDwsD0yQ7woViGzR
eNSsF/5bp1z9SrwavEwVGz1n2WTSaCW4b834REzPvI+5IiU0AeJoURdYqZzABmsA
WwkZOj+mV9OIzj5kPKCvn5sHL4L8Um/WqSKCVKtpdamLOsM4rfeyr2Jr7C76oHhr
E1ZcRjvBAdK5IODDISmm8B0YUQJ7lO8kSTHM7MGLkqwWG3/zFjIRg67U3wL0am9E
JtIXcDkYJ8kP5Ai8rTGgSIhyXDHUrefhg9VX5SGQQs+rUGBovVa6jEtdqu/CdxT6
KTCcPe/ZEKOzf7ekhseQrMWhbh5A+HSytSD2jpTv0L98j2iAp1MfMa+3BnIuq8KC
hLm755iTVMA+GchX6e0+LT4x6nC6To7ZLal/8Bgob/rnL/RXOebH0H66xvnjiiu0
1MyZhmjLfLW5OJX+yT6RDEUzFH+gEil96ybr1Pe2GID41tWUQa16Do6R3I0/91OS
5Hd6Dc/CMAtAXIyeubpoL4IFlhNebPfxJNSc/1XgAbdi6dBAh3dsknCJ0tdoIysc
LZyxxC8vqwK87prgS+UfHZP1G58UXKs/gTD8yaNDyARmhsa9Y3xYGDfEmQSv5jcO
RazKbZbBmHWoGRjMRLtqZyPJ7bANyI/QglbJZKTAFNMskJmh2bZrQ+sAik1lyXFT
hfYGVS1xauPhz6npIQsgPb3kTWKI8gAj4PomhptbS+uQAnlR4TWBnN8KHIzKyvyN
bhk22KjsPbX1mcWM9E036Tk2/fDlAfJK6x9ptJ10swSN1hMAZxWcGoiFwiRxpMHf
gRP2ue5sFjiDEoz4tQG/7wYC8/4245cRVHBP3fsRH4PkJsCcowluYtKkOkBncDfL
Tqrqn1Y+h5RY0FHKHB+UNtyUOC98PSiItASnZwZe0C3d3Wapsz6bB0WuiWlGHMQy
Yta+j4NOF6jOSi3nU1iNebFId2uv7NvScak0XETD/quxPNEidvldGnTPWzKuTiJJ
Cq6xEicnM5aQkErxEt18u4BmtpbRLKQT7hWCDlpBy3a4gHDhkx96e9f1yoE1lg4I
Xw+SLPNdeWeFRIMcNUbppqBPz7tSn+WwKpDmuZJfa4czsuf9GMl2CY6AE/Dr8rdR
Do8BKrSo5TujRiwlYaHQDSVCTfp7dtR8o1YoO57npWMxHakVOpyy6hLqilQtvcTo
Kb6xmkF2p/s+v1jrDTi1bg3q73gDpkLYhMT6TquQZ4z0E/sZPtOPCk2/YRLRdZBg
kdTfektlWluF4Fv9CfBsqTnYidIBjUJ0GfK6R6yXstVuhLO9VFk/amNJTtgF4onC
tXA3IzJ7W00I+HSEyY6TAdyBrDM72IylBR2/hVfhnEaAjUeK942Re850pnVWNwtj
jS5PqIkWzXByoRHMSz2f4DW0on51Uv51UQOhEP33Gf7b2d6rOlEnfoQ8eI/j69QP
D8Qo71PWoguWNoto/xRy00z/S9Uh7uV/HPDRsfrwZzagsY/rso2MkMkzg9OAnLhj
29UQZK8GcgR5ClDtT688UajMjKTlkqnsbOlc+uMGWJxl9jQq0OS19Du2DGdd4hkh
u+Fab37CCgf2qT/im/3RiA0PohfXX+DvPJt2BI2t8zv8gZMMUBAHW6bqUqb0KHCr
8i3mTo/N0qKmzsch8qzKj50YQN6Vj+AZQbi1+5zfzWddkTfhPKM+iRqEfOoDzfR9
yEZE7SvnjD1MhNbMDviVoSIYcl+8z75lBgyJDY9w8R/OQQhv27lEZz5Tc9Y4sUNc
dY9c7KoWUwUSv1rX2hwI5Oa4WuZT2DMTdjH8Y13TMQNmuwz11eyHLY7IhR2o5ucO
8aYW5sS0dCnL/qTMF2aaUhi/OxHB6Z3UYKtWYkUuLfIKBZTEfEcRS2B2NLIQyyee
ZFPPatvqBw1Zv9rChgEPhh4FdlXBlpaMpqmMk57A/9dtjnkV0AdINYRfPNFjbSSn
yv/g3mS9MpDBsBqyBWAZnfJXrAcoIoOiTtSPclX+6IFHcmRVxArhruZ0m7q+VcgI
Dw1E5s9xuzx4FUH4geE9zLWq8rnVnc7ZTMRIzCOjI5aEZ4dN2O20FsRDLyML9Q/H
6w4t3FT4d3Rdvlwc8ZDwkVPn5dhNz/S/HvrL7J470W0C+eyGIuhl91eVl2+XpMgT
/dymfp7HopFLoUYE+NVKW1gOanLX3dTETnIjIls9pXLLBgCENcoFL56YDxgN3lUx
ny9Y3Dia/e0pqoEd7BHWwGXrHVhM6vAKD0JrAkmt/oguhHP6/I/FQeTS2Azu3ige
as4i02qoCOLXJeCRs5ubqYyYo1sJwI1xYo2AsBoU+8HAAzNG6EJbmyj+QeeCKGPl
Q27A1JvDmBb2Iyc8lx7Q0RkS/2XOqHK1vI8upMYQ9yueF8SiVZPYylcoNhTSWNbe
U8mAAg+KiJTkloKInYfc+SDUJbbBvIz+Gs160tIKuObYSYJxiLQjy+4VYga0kBvY
2oHTh/y+dIVT+CkwXI/bhT++qGU8lP8Mb85KMjbz3/ufiOjJ3vQDEbIFPS4igo0q
qyCID5+LLWxYxc7cy+RYO8SNxxbi44ICkhiPQFbk2Q3j1oSBiMofgqf3L/O8u819
4yo5HU/0ExtHnyoYqVWN0Q5Z5rUEPrMHLrTBYHblxaPOg1CTgpkoXCUYsPtTTZ2L
zX+bGjsGey4wPPEwB7Qd9P91yCv1E++TVaupphG6TduVCio2/c6dAvktBPeyxbow
Dh9WG+hwVz08PkrT8B+OPHI8EsF7fiNdq2+q6CABDgSoVQPB7lowJvU51jE0/YWw
86P1lApbLREdC11AZ4XNKiB4yPAk6fv1sP9YNbmUKBwgqDG0LZyTHdBQ/OmFO1QJ
nlMiY2tw+A0peC+eu5U1MdRXFT93igLuwWPxEUdIS/6EVUSPELsd0p0zX0w0uZu+
4+GV7iyXq5+oeP6HfAH/ePGpTS0fllmWS79jvM6KhZTr32uJl2aoqUsYRP6WVnx/
kuurGZnWpaaZ8AT2yr9st+plHVvQuV+75vSXfa0YNZJm5v/pKgs4Dsw+qH4DBcyL
sRrbbldsXANgp2HH2OBGB+e1gzo7WDrgqViItIZFbByUEgDHqlaXTLTt83xQgMDN
uu6IkgtrkjlCxudlY1YG+WM77ne5Ks+ZyztYBORXgOJg1ZXscTrDIwrmIdclNuON
xtOOk3B0u30sSwSy9gP4XTH0oJv8/ykRhT4uMRxR867/O4ZpRVzwcyRPR6KIBRxX
9Npeqj8efvLzCoWYUKvfMwgRX+eHzuSGl0LdgDgZueCQ2g8AdZzUClZFKcGGI9nZ
/ENHJHDtbcuEF0U9OuVLk6f1QIetfQ11i65+H420cz7T5yLt6U5GJQrEbKknLrjD
yWEjVfTvBrQd9IaHlATTGU7nkSq/SkBSGQIprlv3awEmP+Digaitq9yT6v9zvkL9
Q0bs9cSNTWdfBODiuF4DcNmbb31IrxMlpx3ZBafzb7zfsXc5GfXIGQmvnXNQMeoy
Oj0Wm72tV7TalKzd4S9njH+JVajDtZoECR+1dSEfS+m+OU9Ke7YnvZ5z6cvFkEUE
1LEKlfmdlk+65r2ia8qvqdEPnMulf0mxfRq5vLodpDUZEr7GAlzct1KPh9pOJOsA
DVjq7OVUPBXPjGtts3EH96PhKNCIpYlhU71FH9USW/PnPn2H0514vIm28aWtIp7G
d1tkJwPR90oOBngXnCL3AxEwLYNh4yRrBMh8/VdqP9dhLvcosCpUxjbbSM1BUiBo
zfIY9pYffMD2v6hDqvBh0BIGOD3gknwJDpLPTDLtIntBjirfWudQ8lDcxm4Qu54o
WB3U3I8htZcKbhGswSxU9lUHKyGWqkco67ARMFlOyejoHwRX1uUCRtpNSI1/kPK2
2bCj01wxAStkX1V1bpimPmhgPWkXDQkn7Vb6rh+QsZ0I5QeMi8WXu625hOeQ3fCp
JlhDLfAc1atYGFBKr7SyivLIkRyK5I7Qe+jYDNYDgVJl8Lm3Zbh+6f4r9T8YmIjb
8dCPqkQCVj2w5MhPi/fk5TuurpzCWoxl/rHTZvl86kwLAZsiLwHzb07oKwrwJhM3
Tz0SxsqAPPYEaTtAEjxe9KjJaLWua6XwnNQUKzuPM1UvUd6LQOmNLxCZW9daQdiV
rTc/Asr4gcmVuXxt74Mco+OCiZpdeR/J3dxKeCc3MIn3g+luvnWRlOwdjjqngJT4
olqrw8E2H3XZd5cOPHjLMBCbjN2VPz0CfXq0x267ISUg/ZVakRmeRH2vVeeka/gB
astD42cjYpwRlhZHBKCjny8XNhtoM582wpKdASvh5vwgPg+SZ8LBy/SlKP9Nftim
LIcjP1Je5dRKnT+He1auFyNFwNPCH/dXRTJ3VzdhwpxtFZ3bfhv+RUzx7YdTkg+9
mx3dkbDCTmhF/nu7bUgySahihC8h8kZol1Nu+vG24n72rjkWau3EqbmhqCJSCu9m
vv/Yy6FaEnup8W8SJLplyyPpvlYK1hS+X7JACLNcTkcrROkhPQ+IIzhBHLvaB4lD
LisigmP/OzCHMhefWRwSSIpnGv1cW7Zha3TtKHQjbh+NpbAQPY5aEdppDLhrkfog
CtfkPVoAiMy2t5xsBzq0X4zXr03A8jaF1Mxjmuk+4uOqMjHvKbtSxfOdt9mLPE+6
/fbBeThv2xkKwLE020HxCFWSPqETgCaGpACFwCATZedbxOHCq/EFhN9v5aCcuEd+
sfxO4wIlYB2kebH/AC+C82D6n92nah61ZE4Yk7ZNZMolDXSimC+G8ZlXXn3nuClG
+KQTbVYJk7JLazTR2VOC6ljn0/0dlFRFyu6H3B1lw8EiJ7sOxgbCWSt1e5UWhvNc
mVcH/UJUpLDJZKlx01vQa/VsO6HYqDPqytG2BmyRo1QgC+McfvTEDBURfjgytc9G
olpMGBwUH1bdBtRe0LcU3k8XJiBvgSgWklNFDtClSwXr3GJOrO5hnMlEIDoqZ833
2Lqo+1Ik6uCo0ywRFVf1bxFSUWUpfWsZJCF4TdlrJK+/mkFyZG4XFe/3J4TFeqWn
8RSvXRl4H7Rvt5lg44ODEjAca5M0GqUjPmqntksqIPDxkxaDJxJhwIbeW4niOvM5
cNVE5siC19DfODA2zaK6UDHSRc440rYlt/wjeDrs93Il3FHY35V9HZz5ZjmhR143
K4vuQBH4ADMqWzdL+GWYySVEMXoxXd227eVMeQ4yeJKma3IJlOkOp89mxi6agSU5
BSODHG3IE6PATimW0WKGFk4AIOjzCWGaxP8ouuQZlV7H5E/chGQN3tsmF+iwjCFS
pVmviKh5ArlxSyyqF8VtBL0/kWQ2v1Brz6RzDbsxTujbk55C6U/ggjNKIguvDda9
Eq29xMpgyuzq/QDUThjn6Zc9ZayVqNgYdtwRflih0MQo7JQKc6m9Ao8BJc1vp0m9
EnhsRdqoGP7B9vLP+RMYaf8hffCJJUfD/VLcLBddIYIam0k2G35BjPvClf4huTW8
4+d8s028uYpgJCbMBVZiMRyEPROZb5K+67uOMmpb5qdixYRiXmuCHcYQvwyAPgoX
mismRtfKjnJgH5iTWqthz0+lQnsJ6ZhHpYGScskhiaqW7dYPDd1QurdNVbUBTQR5
qOeNcGF87QBUnsg89G+qwrm62Acp3tVbRBJLiCuzL8OVE2BRSDqjhlE5gKulGdjp
iyWRb3cfIyN7Awi2MsxUvKZHxpN8T6Y2AdH/lv9hrDB7pbEacPQmscq0/wG7FjGk
15kH/KsVsPRPs4Zpvyb4LJBXc1Jb1lvX9cR0+R8b1ynKMuWAgDWqXKXrlpj/Ww2W
QLNsin6SlgXiRE6KGQBAyfpi9/oK0iMNxjRcp/z2HLXKL6s59XnNj3c7kzh3JiNs
hNx9kJK69E+0Ze1Fe9/nm2yUR2KFgyxqTd8htdECbYnodb24sDDpnd1x/E/8X9oS
GpeNvihKSAqmPIG/2Zlh5p7pxEHSX7Cc1YdGOqidCPUX0OgsjJX9Q4/QK0WH+U4C
dLcyESK62HDD4c7UIY5zPOASFQF3IlmH1o5n66m2fR0LOS9uuFbMvwypR20MXXYK
4SsdCWFVzxBDmS+yVdtDj3BBCA8v8ESkGtCWHl2inrqOOXJ+clPll1nQYSt/Y9gV
YYb//l/UA/RSEW8xu0O85F4Jcs9PTsEoiMwww7NDbrnIid2KlOwkiedlo802ZCLV
Hc5U69Da3wEeLU3VrPA4/YFDhbD9nnfuyb1ArnaUVkLUVRaj/Obd5/ixmoM3CamA
hrxwjqtL6kJh2LdVRNefPm1sbsGxcmVJ11e+nUw3TMrpiguoQnjD7yoiPHygM7Ri
n52+9i64QREoiCppU50Z+K9mk9fjqxKo1/zYEOOloMFiC4Xu15TzUXfks0lzOpTm
kXslQHCpqMyuT8IxadeI2G2hTJW+RLcE/N37g4DLCWmgGZmhqDPir+nTEhGNqRSg
5MJ7U2YheNTGUX5bUSFpuedSg3Xa9aFyTVEsemwrCerQEApkXxJDffZEJJ2XKC4/
xdGpMhd/JgHQ7EEoHDqGZMDBz/dQLDsBg2GqsZgwCQAdvDlvVYiPhMKQjJeyAqfc
ZyzbUCn9ZiIVVcrWtoMhd0jrhWJR4nb3X1JvA3Xjmur3NMs71lblM2Pt/ldWyttu
POjFi6eyN1lHGWWKnsx7jRs0m1J9hp9Lk0k1rOaxEIvX05tEn2N26wkmK5QHG8rU
4u0+ejgL9Rqql2kDcGbUfRKBhe0LdOLScx9AWUMfu0E+ScekACa/vHKZbPSHtq0W
b6DZjKKCA+6H+Vqx/X4llsvZWQnZeRQe642NsnIUsVGc6t/90aaRimlt8WEjqGLz
IhDTX9cxbvuvHXWt+wr+0NABAnEmQXwjo5qGw258AO0wGOv97f4O4rt8Qm1sLMME
AhUASkOFZy2qpZv+WGHcisUe/zUmC3ZLDlmdJplBTk16BXgJLumiNhfT0OMwW+Mh
PwWpa7lX14nr9sTe1r4B2+ZAWjbf9c1Cc5JTNwqtrZCUemrjMMDTzPL41tjbYdoT
DfrJGO4llDDdxYDOf7y7echJJWUGrRZT435oXTrxqudfg4eDVOEeZKnKV0YGu2e3
jNuEwOAF65LXkdK08TnRTEj//1ZKMcDkS8HAKl17MhFHP7AEbsj71PO5j/xaWZnU
WAzxOr4hIa5KXQ+9WDbSpZc8EfepLqHmCFK+lR9jolqInbWd2TdRyb7jIG+3GBQ+
SOwqvAGPv0KkKypJlQXYDGpaTWoXoZwRGYRUOz9E9s1N2G3swcHc0VC/+5MzW6X4
GXHD2H7Pe2NdlcDZvl27wtVTrN6Zh3B5KW7YQJQhITkJPCiEJGarL2zL4wE32UOu
Slm8WiRO2UGjwmQOAlc0dSih/xwO39kMF+B37gp86ugzznzi3BZYOg0518dRn1k4
rHRFFHloaE6sDy778HQTjdDmq6Wv1d259rCvD/Kqu8oE9CgUGbQWomXSBsSptyGB
qL4k+v6bCdOl+/hjh5Ou8B1l/K/SQSPenIN2NIGCugdejo6UmaThsnm+ON3vo2C1
a26qZMgLaVP+6jE1rFWUCiRELk0hoWwcz1nFYIFOVatC9fnEgSRD9zzRozFUxHrh
Pl4wn9f3n0y5sUIhurRZqua84G9BVhcVw8Lr+9sUcCs6l30MCPw/8Km5wxstDxiF
W4VaFNIYiNEYW5bWnBiJBoNkeP9LRoY07UJWPV6dcXQ1YLKDidZb9AEth1J2fvU/
AfVr6uwuz726rGP2EafTqOo9+Q1sb6T1mD9p4qd8ckpPTJqlQekSR9ATHEqVnSVo
wxVCWI6znOCH4aKAKPQGVf3ak0eZMpAlZeWk91LFm1n1Uk/X8KKo3tRucFT9VCSD
j+NocFlNQKdJhIIEsz+AWbl7613GRW2e17DqK2mKInJjwBKpj5VJTPmLjzSEpGoh
2EbYQLBgt7EKzBYeXFu43xlmIxoZGqWCaEst07mG+duhrERdENOyvSWidfETlt6L
yiKr2Su1fySlQwwkLmf1gfioU22Ukwv8zpoVe7vmwiUpIHXsKISsDsFQdiD+6iEI
rYW4ZygweYqqSyt+51L26eql5iVvkgVXY0hR506oqWDI8rTKjjdFVZjRFqeDL2pK
pBijh5e3preomXfBtR8PhgOhaDL+wieImWJornz2207nVIqn9YGvN6jSjaivut78
DkXX/qsDWeAFNq2b7uWLR9oJgiEWH2csEwfVuYY4wiZlxgYn+CsFQ6CwZQNmU+M8
F51iSOtdfqmVM0S5q5mYibtMcc2mMj9zXUkn2a2p76z01VPREOwJCyPa4TvP3Uml
A54zDWIzz0/lznRJBNOtQ5CiLnFM/lpIhif2ZdxOw5dNqdLdxjLhWprgkmEVoYWS
nX+Q8dVbuNu8/XSnmaIeLe7Kw6sMvgN7yv/2Xpzld6FFgHQU/ZwcZ4odScIWAu8o
V7CY30DSbnoBbAJ/yzuVhy5/ErF/OO2LmKLRexkMb3x8wBn4NzaSUtCaZpW1ijg+
k2HRkIbGaxnLH5EwWhrh68VI182ZcELP+eVZpDnarEoLrvpZMOkL/c4p930gSt+X
6J/0Cg5YpEGjw4+5MzVtmYnYIArWGVBvIVtyEj8+2maXskQ8iHUfKhi3Wjv6+if0
JZGaXroUN6XcfUjM7vBKDO9ZqQP5F63R5+XZzIntCtl/ny16Nww868TLNuQuXUVh
Kk3i5DUZZ+DXVcbaN6oVC+5jCj31oeTl1982YWzDTE+W5xy7i90X3hkz7BbxjLvz
XgiltWx0vttOgtOy9VgHDFVUDLAUa5wDizGqpBzFb1IzEDEXofrRKdlxZZZlIJKq
QhbQX+S9shWfSVslpfQPS849/z/qj7IANuHokMOswriFWl42eTvjWfjrop/LD48Z
vEX3zNZgDatW72CLgBavV8h8OlcPOrlILIonHLLiAvyAfu0Z4Iry00AfW4pNVlUB
LtAoDVreNg+/OUepOWJPR3GxyQfkPljEA1svKMSiW4iXBuWCqCBd7XGuki7xZXgl
9C9cQ3HFj5QX5uUhOtSBbfmj9OGfMXPa88sQg2Mw8kW14vAzzX4ZkX6WxWvXg5bt
UXlKpwAYzrE6CsR8eaMCnkk1xNVPJRuPfzGV1Fv90/NjwBqnypFRV0q5d50IAl77
6DR2eSC6p6/a0+wIYziZNs93qMS2c2ex5qygd/JXNjwbL0fgPZx3EBopVLkUvrFy
wPv5+1YH5MYcyG8T9TsKlEiylDa+iDNcVQrCJ5O3Svh4NC/XGPfVvaySri2gs9OS
IcPkgz7ud3A9624vWz8garSN1aulHVtiHWSiG0+38ycyvIE+u9c4oNYywQdfLz0s
kE+eZ+1+aHuOeb5X+G8WVfPeWKGPKDiF1sW1//+MyB1u7UKOig48cV373RB7g895
UaZ0vcOafVgk1Xtvi2teXCLdY4MqVEZFfXj/VyK5+er7SjL5B1pmh7ccocVsZt2h
2KrL4NNkD5l/C3FkgfMxmLC9ZTWuhWRlmyQ+oXnCS8xFz5Q7EGZISeYxtdnce7Xu
GPp5M2l25hzWhncjXUPOIu/yJrf0WaJB4XsqPyLjZR5I6Tyf6rKDB7eZ6OfKNpHK
nNjo9MdPZOcRpxOiJ6fSxfmzNxgwjtm6T2BbeTAfhoxss05tduzvPN+oW8Th8OF9
mp5rhELXZPf0UAz4MjUsYX2u2n1KgclllHQSehG0vX2xJ2U6TG0Van+aIQb/elJc
ovEdUQSNws+kq1Y6l/EEdBXqkGoh8NO6KH/P66YyIROpWT2fWX5FjGPWec60O/2B
2oN7qk0WuG3VpRj1rapPnscf/qRaq8dxfeViZ9ze28CJG59VAAY5w51jdIGdoK+B
U1lRqMx5PsiV273Kwrcq02hNiRwLWLyeF8/EXUkYaaHKHfx7BbRM4l4pK2BvlXOq
BCVm5qDaVVTKVjLRDLSQTsq8dANWU6TPjeSlQAjF7NRJ7GZbqGbPdme18UNW0ZMZ
0gLXEVR+dPFpfwW0Z5dTcznyIzCwxlNxcJZwdi/bYrmDJxxpdY3kP+e4zjymrd18
3Q26Z9gZUb6MPxrDwRBFAfc/5IXnLgZz2LcS+lQZxlj07Jd1LeK2OZ9L3r0QyMru
uLpKJD1dFBm+EF7n7cXUZyamiqq7Adt9LCd0Ug+4HG8tAW7Y6RdBjCqTpq1BEmpu
G+huAHiRDNLeB9VIJ87oA4SeYudOAvGy64aQGD15fPMO1fLt0COTzwGnXDIR72um
uzLkm+dcR1uBblOnBrXpdMgWiM+vE1hrf5Aw46MakGY6CJGUcw47f2wgOLvvDlcS
iAS7txkGcNrOy5QVLGVors2NqBiZ1tI/vgGnpptIgNYsv8opXp0Xmv02jbVZMGMh
qa5P2usLx9xgdqwm1lEJLizYw4YvoK62q3t1GvcRBPDmqTMyvwckh0P1Ud/RspdW
EnZB0gHBWcOIOgsXse3ia01tVGj9HLOLKTK1TJP8nYBMDTpZAVr5Dnk9oVwyV6bQ
/dt/v3yYUYOyI740XK/RjACCa22Vf7aJS5Q9iGI0ifLZ3OP01UO2I+26VfTWF+YH
LMRJcVH635J7XJwbjysF5b+Z47i8XuwF5A8Kc2y6pxHW+7w06+RNBiy90nKHefg3
LNI0iTBhA891pi0M/gd3XCKo+MgzqyhFLWuWgUZZHcygiogzOi/oUv2j/XiFoD8o
Dw+huDuMuLKwoBKzlkPyShOeVlyIKQJsbMEhrjieMOx37PP0uJuyytbxWKX3c/5G
Yd04vg5I2USyqJ+FyUCn1N/o7dbV6oprJT0O76GLFsXWVP6u/BIdahZ9GHJvcaA3
TMK6o7tLMW0hzhGv/RVxwHKX39/iz+9/5+9Fi43wNQA1k7xzcPB5FpcmujsURv5v
cgSZ05ilY4+eHi6sqiEY9ft6TMLOGbb0+jFlb2pddxF+BO9Uz55vW/tHFez2c+CS
DMfnU49y3zPT9teBhbTmy3tlxPUXLfjVA0yzq+fusZKcs008VdObe8ahXgrr2uNC
WWlkXZvhroQ+sXWYtYAQkTGquDkGEP3+KullIrmo1QG2T1SAouSY7SjdIT71VO8A
2kcga1fttRmPoadJ/cBrjCrNIWoCgEaXSuaNmhrf8AD5gB6nd8KxHBSObdLaluty
IL/5cFhkm8lPPhXcH2Z9T2dzc/7ddn6xTNyuu/V4yRg3eHHm5uciIGUa4VrgizZC
+h9tW0AnK+GzdkkmWdVOnu2Zk1llMUecYVn1xEOhelt00Ta182rZqjloItoaXwHk
ErZpTq+Y7w4mMzQlqPTdTu/0cKPC9Jjrwy/SM0HtqC8DhxHGFqpRSSfclL3V3PBb
hD5ocmAdEb73uWPzgVpqyex8lcGVRdi0X8IIQTf6mmIEdyQ1zruP9CqcRVoPVWi1
ZN6cqK2g8gMiIGQ+vEXsC0NeoHe2C40UW8pEAyGr2Py04tpuhK6mUvGRkzXZFxuF
buBrXJirFh5J42wI9UYSeDWCqfR2cLwRZI7/e50bWYsbch4IzTXf0OUeKu5iprAs
SQbwpZ5u+rgOVPodUY5l3+PbgOjqXgB97Uvwn8J0gOAJVdpLNJI0VawhPJbXgPFK
KO+2cXTLS9ROUAe8rzLXQ9ZgX6OM8TFToHoZENR5SblKoM6QZ6biSj7ivoW5XyAt
0Jnqih36cBia7LyopbDBKE3DKNgK/v2XL3GlkEmsRFSox48ie3WVSbl08ugKKsjF
gJ4/rW7OuL2UhDPQcVwDWdFqmhWwcz8qibnKdNDq2OBcARkJUq1uHc7soE6dTC35
5ypcnQ+yzjyh7wmcv74RIB1h2CMhT8ihEtGJK8oDUI2BRM0e3r1UoWojzDgeIkSg
NZFKBc6EQx/6vg+2r3D72GcTjlW0fO366/WY0KqWIwaalLQOAScem4XyLVvEOFN7
0AX6Y/Qr2XYsfZs/k0iES6CI6+f7AkoHecTxGnCXZnA73geuO/u7Lh9fk0Gf8Ydm
dsPDG/ymAVpAn0es+iUbOZLqcxKbLDWudXY47663fOmvopYCWuXUw+El5vWvrvL5
zK/PN+beeu4y1uOuqDfoxBdk2x88H3oxYaTz9fLkr2dxb9lURCLSgWnhiUEDRfQ9
meoaKXPlI+hJuKys+N3RTO7HyAGOuF3RRL3dtRLPGqetueL6wN6jWuouuURi1C4K
UQ47mmU7KPTnuOb8cknFuVzFq2QhmDluSwz9Ksp9y6nCvrRq5xSWfuWv3KWJlsTl
edT9z0MCn/HW2S8bJ0XwhBXr+q8AAsAPb6kzeNth3Vhj8pcwaMLMWZu7ZPNvk0uK
xnql4qhvRypAyN8sWn5Er7smnvJJvOrleIsGTnjTbfZxJ2Pm3ya1E6ASATxLaVZx
hDDlRsSXQoys+0/E969/fvHM33Au9T+uCga1jWjOLbA1TykBl3c29Qbip26sqhgR
dkL3PZsqzrrLFAk3XR5JRoei/FkIdSMAxBbhJLbLJPyXB3RPP+PDpXY5gjvckQCO
Ifn7XWtV63bwZTVYP8VOByJ0LigKU5LKef9ILK7ByCKyssynT3j+eaxCVXOWZZDK
ahlW2xvCQU9PU0ArxNjcXSU+l/3kd+LtCbxg1BDGhDda6kn+cOU05vjYG4J1XC94
eg/ZBXe3GRvFGtT9zAo/HSG3G+BYRQDBgEfj5v3G32TGtsGTkfCyaXD/ckdQz5zX
7r8SI9Objht3hWxPThhowMZ3amF/q/xrZSdDyX0SA/qJH7Hru4pUhRTKEFx+kXcf
oAq9RTKltO30myrOSeGbpg9P3H0e5sGlstkklHU+cwzJ4gOdQHc75j6ydKmkPt8k
WeKBHP+M5AaGywKpvMz8cgpv2VBdA67C6BO6muQE4UatPqcklMejOQzTJsksr8wV
T8ozj+8ksGeOVmNn35QdlN6wT68Srf0MJ+wyAYYg8v0yDlmRHPy2ltRz23yWE/74
XIh60nQj0LwNd+J1alWLLzyGzhwt2r3JRR475c2w8OXbH2qBrhfx2NDLlhsdaeuo
ErLfkuv+IHqb07gDbyeoDnnsB7G9ymB8uaNZxFvgK5Q/VkWUMeUtFhbPwPTTrTah
Rha9sXPQ3Euqxuh4F/MQccmBYGfZ5G4d6Y3uAAJNa1IvEzoap0SkvnLA5LTe+2Nr
XpwrKC7we4DS0XGSYp3gnen1UkG8YZK5rMSNWtVp06crNhPoIrS095Uzru1HQkaI
FaB6UEPkbNBu8+DNjSsPT6jrU2eyrft6M/X/7FJ2dPM/IKgjTmoKZ6hcWX5O7CII
//Xhhur88fpGcEagMJMV+6eWVZU0JSYDkkw6KIFXPdW5vGJFpA/B7e+gvsNAnXE7
I6jDZT+yAeUg1MAV34uXs6kfd0OrqNcwWW8sWt9VAM+CFDgKVfJ/q27dgk/XSGtU
01qdOdza16vUQIVHz6NnGYSabwQvgis+plLOS+iUZAspjyjIdGUBvIgSB1wawh/Z
DJi1ukuZimXJh6uucYphCB1p15JD7tl+/Y2/3tiXOgm1zeV5xPcztXXsk7kyrOWT
rA8SkaTaL0+qpflxKuRDvEFY/ZTXjmGF6VH5RRRZSSQDD6UpGm9zJIU9n1JfpJyq
ubDrCfTxUAGR4ASSmR1cCTUIyg5s69YZiHchRXR/mAtAgphrwkBP0rOdD/j+aGSl
hKI77w/Ya5PsWsCSk0WEA0kKN7CBtLBdlZG8xfUU6f/qvXyr4rZtWx82QQbzHq24
/p1lMGMcymdrEr9Inr1TCHiuqf+/ZEx6N9a5LaA/9nYFmn+phSSVkyHvPEVEYFLy
uDREhp/NQLIM7L51FLJl06OO2mrwsuIdpuHjHuOiPv/xtFKP7Mk6ymWlv3bEdLYe
TSRfmtc9OKGj8YZajr0+VQyac41v4AGwzpHU2MYXY5L+ueO9C6m7MAz5DLcabt6g
5PPDy5QqhHFrJoRfpOj9cfkBPvABHep7e7tucFCH2nPoFyobn8Z83zyQ9LMlYZgr
NcqFimOPzPumTV4LiH8CHdOpMgfaUN1PzetTTgtsb9lKgazegrOXRI+myk1cMW7l
OXg/XTROtBGqe85yl2V8PkBxQfMRiq2mbtHk2XMvfM9t//yBZHL7HtORIdBmxyNg
qLyXJTcT761AaaDFfzX22UUPGel/yTTJFkOV/zeEmuJdTkmTZxGiuSwgmv4HeDMt
pJBTj3Mq7fQY95/n6eDHKGJ1NSxAcKzK7YP1s+mTfUL57JwuuQjWIt34ICq36W9a
h1x34SCObjqvgy0Vjcn8yuEcp9Xy6pL4RfQCnRSF0uy8dfc4/2XAfEpqeBXPWJrx
jlWyMrVSb0qNcoZ1+5LeNU6v5Ky5IJ7oNL9CHz1xTeuGsstzKxUjwfVdf8aoPI8i
NI48Pb7WcDeRfSDXMJXSwAFEzJB4s6EZrrCRSv2R8URyWOmwbk1gYkWBDnsrLSxB
nmKWDoI7Ncf4u2MO3Y6caC+DFKUo0sIoJcMRdrNcyG3N03/g0cdx49lME6Z3Vkyp
nfC62DHB29nW3G1e97FoPyZKzJoAVw3NTyvW4I0enlsHOdUIbGZBToDryFXzIe7T
KQ/af5E1wOheqASs55vn9y128P29qGUo7mp6GhBanVPR3amSGW9FeiGbiaGmz511
/rgYFfeAeRvxVSOZDt0zOsOEHBw1T9WLVvtA0UoBuHDSxYPZ/Gz29oKOk1MWYeEI
UVxrUxB709GDNUfBZ/4foENpo6w++5/up68S7M43mAD9yALr4WnRcXgMhzAogOQD
MpIy2lVG0Dn8vBkHBP2VLdQg60HbmckMjGE0noZ/Y4YdISwF+tu8ILI/nf/kqe1D
5RhhUSHMPZmhg94KLIcqRGTSF+ycHrcYd7nhmilqW2WIrhQkA2OCQU+V3U2XsbD2
+mzAr6e4aF7BVNvxCF8SshuPUKxtrzDTOY/5cdTThiZ1rRA5INSF6mx/RWXjOUVU
ibqg7n8yalxAWXdQkywZAbYSbTz7aAi2qL0T3eXnGUpYEP4xYWUif9yIhsM46wAg
2bOD2D4QpIj2ndkOQgaYDUUKqOpHloVeDsS07yh9op8sNi5QxNSQEnfj0UT8Rx4M
RMmZdbHT3EiPOn6BUGgqgepqlH09rjiuM4LhWVdwGLiMlJey8I8xBAi7U12uFwTF
ow+969qgdl84Fw/pRAxz+8GCakYr8la+l3aAQ+5ObeWEFGSx1aOMFZOL7BIAMydh
ulP4eAlaLadFWvPJxW6YzBFYB5B+gnUh5jdNOvoP1Ojggx3gHA3/6Vb3vxbPMe9v
nbHQF9pe+zVfx1IxrJIIwb+fxmrkS496lpa+OB+ocUzo//Rf6UldniT49oftMUZm
8hgGR/9qiMNv1SSf1eD8AKH+pJxPDpch7DjRfa+awBqfZ08LbG/acoicqSklyUXu
XozqfbT8EicmntR31lzly17roJKnBRU9LwR0l/zQc4JftqVYR4rbYz6k4JVEV8J5
Z/Dl/u2ptsDvsrYY5SZY4nvJRQwo6pwvEzWRW/6kzsTS2kZwWluKluXUX1bix5w9
E4zdK/se2vKMEn5bGPhclY2OYIgaX/+AUNWie19fSnROcT0m0hOwy9TTXQt62hhR
wNJin/1iE9/YtTeQrtnua4YbF8v/UouVoNIoWyCcPQAKgQDPOlxVwt+KkwQ4ZI/7
dMtQiLSBi7waAt5iMFNn3zLG36qQz5towDeLMQbPuhSZ8wiTh0oByUlk+wfougIr
r0528mN951ESvG/9+KI2lO7ZZK/Me5NjAWQYyLtTf6Boak2Usvn9D3OlRihgqGwv
2We/xDkoDjy8TC+1sddzG5BmJDbWPVmfT4U/Gm5rVPSKKNEvbX2il0oP5lgus+Mp
LXTLDjoXLYVnYTYFEoXossLmPTsx5c4BqESCe6vCUPSwVX1JnRLWBo7ZbXxU49uh
HmFkdgTBkFzcP0gUttkETw7I2sqIr3DkQztxXdD+ZmLpUq0ueORokDvTW2Yr7FjD
jbxWPFjN7OpJVHSH21bEdKUhv5jiCZynm+cVL/RW7O8j685lUBs7iUBDjdihznbb
6TYHRh5WyazBNjpOw96DlFV+qgCH3jNxPf+FFvCmtZtyrF20Een1yDgFv/1CG1Cm
7JbLC4ikdRrQi6aGEorzl3rrQiSx02dinUbf1Meq0sY92MMzAPfIET46ZcR3Iitv
YgcWTSQH1UndRdNULjisGWTur3m1arLzjNTjUw3D5T60WWr9RgsoWEnugVR+5MZf
21gWhhpRe+iv3+h5m6XRQPDE7lOugdmKcPjxgqr5JAvyA9x7vasrBT8oMQ3zWVfq
wPlJm5bXRLjNdplGXqzArlp7Fk8xE2tyz/PxG5Ort3RGIuz2eBzpcdnjjqYBACBj
UL4XWuF2ULCh/IbcQ1o6o6zuqcHAvy17snkvX+6ghGYmFEBRXQsNsKCMcmNwXdR1
YgKogE/tLuRUcIeO8jLsgg486sN2Zl5FtdwL7/B1EwJm/apaKTb9Q7zzyHMN3Li/
QbXQ/7VSMBEqDqhLb6W4KDNcrP/wniqk2/7Nmp1Fx2pa9uQM8Wp4HHOrx7T5WqaI
vqXNjNAL55xmPqKgFPQeNc3yvP2G+14ULYhPvozLCOMOEeyXmmSv14rTO5hl1bFv
UdQuDpxCBkP48CNtHBicyq0q13ZMPite1vx/8b86tJ6ghKP5PAPrhtNCfmBxnREN
O5vuEq40IKNHnzsL+S025+x8YsVR5I76LlQ26LhhF5lAJ15mqD+At9i3mxNTERL0
rI75ycbxAIOWDLXvZmogg3n+dDj6BKB8GYX9LJEN3HyYbVYQxKpyjUKizltgADw3
0vPcBD5nTeOYtqf+4O+2/Mvcn3wnfwBmzH0rcFu2Wr58AF133n7vUKHVl41/Yjz8
qpXmLCZuAoL2PkkLv6CBiCoJFE4q9ogb5p4FiUpS0pP+9VM/150nSYnysp3xagNf
deUr/ExBrU97gWUp6qA3lQ327o0cuhy/531z9HrCXDHVekXuc7OqjKbN7dFlQi+C
RMWTflSoCEdjULdiHRNMuHEvUNtlCXQA5mIOSXe5OQ9XvqlDOT7T4W+20vf+PPsV
E408rTTby2ePmAhMC5lc0YDegXR0RQBSHF5gLZ/Qrq1PGip6niZAyI6obUhyGlv4
VBaUikpkE8qnAhXBBOXSYVEGOTiJ4aXDWY1CztY37pNK2vB/j0ACOxq22IAjHO3X
uEi12eGz5ucgxk1xB/juzJJJV9j0ufQBIMSSzdIx0IAaCWT1FzYRoCT0+AyH2krU
ur7Z333TRRgIneK0RCd2LUMniPYPLOdjkSLDMKa1ickFuBttuS/SZKEBBxI+1Hcj
uyEuUJGG7aENUhUfL1nZVZIqAyUbwUpNOqOIkzgWRC8ZSLwWG/sf90U5wWun/RZh
F6HZ96ls8fc7PArvmpDxgxxrqMDqkkfthnNBPeQaz4GSt+OIAbPFlFvWgzGYNfaa
dbhGKZlOqEBdF7A0mqcb9ITkQYBxHuCL6kaigWVEozC3AnkA9HMhJMtpJZJI4dOQ
wxtJdcp8ranOORQH7+rw17D33uUObjfdoad5g0uTE0RJVFMy8o8onzdy7T75ZwOv
tTubx5XSdSMMUMNqs3o3qa3Y+S2oXy7a2uxBnQO1tyc3pNaGhX31lKlAzWQe/IjA
GePGal6UlI9sacc556frZTm6TIifJ/Tg4Bf+NMjFelOGdnRHmBzpFYRxdmXAlV7w
TaeaDrw6zVb+c8EkDfKSeRCQiTrm83QKdQ+JVVvqW2w6MZOId+MbPu7yBpTH4XLO
ZrNZQkRW8yCQ/KE9ga7DegaD7nCEcgGphFZGXeH1QIcbhHjSWWJjAlt7OPScE68J
nMjLiIH9wpYBBGBNPWmcJ3k/ahRo+4pNRB9z70+Qr0/I54UPkAm6ASl8dhF+hrRq
n1NrqZYvYPbt2cwvcKQBrDf97de9obB7TPi8CHCe2YhywDcJctVQN8dJoRCUAznj
nPFoYKUiWoidKbIU54Fa6A0nWXfNY89IJF+sua1Sv+K4W29IJS1e7HQ9F0gwlKp6
21Rj0/ksvRbp6qnx15TnrPF/iWCBw6iRE9UFJcK3tKii2kDkbFehtxdZ2R782/Zy
xZwNNEAPm+Yl6ax7sGRlxWGxYH/GZM0ABkVj1DZ27XfQ0U/Mripz1xIHhYQ26k1I
2DV5XPlHQ2dVr2kK2/GbW8eSBK46md4aoNkLv7YB0gfXXFeCcuhJDKBdFzBp3g5A
MW0yXKhKHOfxzVE8TjBCh6N4h69oRJQAAMZqUHJn34ne17zz8rSozJ7HFJma2H0I
hKORpaB598wv5uz9dI8hGMRhF/Inc6VCQviA7fUqDqwQb4WR13NKaZUGb120kkq7
xjX4KOA8mUMvyQnRsy7f6/0c8zrozHM5jj9ln8TDU6aeqEkblTnyxUxNUkvsOKks
67k6KBwWRG6k17imHqu8To7an5FOnSO8pajRR6Ta3BJM9pyUbzVdsyip4YmHqsJ+
HEWgNDhu/Xd/WD5wb9vp/eiU95eALX13hrQ5LI3PsvOu1KLsDxfUzbgaWgBXbI20
XD1n/vTV0+sNEewLnWPOsUZzWPMjCTU6BudLIpJMZ8ubGDgLL3A3bEOHc5Z/x6Ol
rgOZaBIyXptwgAmGJJXEhvrUdjKfYp0F8KniwKXC+CChQp2plDgN6QpOR/B7o0fn
iL4DsopAlPkLc0r/FN/MzGxs3F1G+szi38I14lbI9M+eHPywRo3QzAcklgVzdMtx
2Tb5LwcKENf84xDEqeDt/cl7+i++sjrAj95J+kftELiLFz3pjkVebr06EH6lzKaF
UQ9gvpUMFwxNYZ9XrhJgA6yD3OJfQJSY/k8gtefsU45hiJo+2ZGM4GF3FWSYvKPA
mey9Lrmw+WmK/h1Uo47ifrsngiS5jtStSqO7VwlPvnqSYoJfpeN8PPP4iL8QzvBh
PaVFlNkE3uFVuEnAVtC8ELxg1aobcJin7ZirUWnsCtM/ILkUM+dZ1sWyFIgY35Fo
xitW60z/nfEFrCs/R/uq6YeZFfUi77jAv15p2sdfHwRbcT/xF1WhkPhL0MQleWXM
uXZf+YW/j/fSZpFijt/O2DVBI8K4jfYjYh+KU2WrZ2OiV0nHCAcxg/n//bvLQcPp
ZEYkPlmE/IHcUs9K6yhbhiOF9TPUE6/gDZrj9N2VY2hhzHIj9x7AYlPOhVcjgvhB
KDINZ5I1eaLc46mfQSfOpQR36qQgLtsNAUmi6SNKA7C//VYWoSGcHSgZ+NGGgRBr
x3wpG9vfPWyIplYvrL02uqAV5erftIKxVv1S4BkSd0FZGqnJOECQXWTZQ2uWookY
TXiw8zCsQ2yCatNedXz0JIJpX/j8B3zXbKZQ9ErozNzA6NmUH2v9KIxb4ZxGyArc
l9IZkUODMcwB8nUJR16218aE094WxPcGAN4KdjXHL+UVL+0Ds3BBLXEyaOYgxHV0
xXrYHDtMfa6ToXg7SWU1M4rB4jcV8VJeoPZdEoqwMc5y5XwxF7YuXjq+jmyEL39j
bxzPdXUdHCodlM+wFkpu0WQxLezvCA42C+LY27hoMlXO6jlgeXj/lzCMhV11MFb+
uyEQTPWDnjwwxCkTqddjxoKwTQ396T9WxFct+q9jWjyjIGfvSIw4ruEzRXapIaf3
c9TdG+U6H2CorCrL/DiQpUy6Xue+mw7PTAV9shWdmER4vSKRKd4p5WNP6DMGrjTn
SZzljtKkJ5EO/g9HtNJxh44EYXNlnuFM6yOuwoJLQW+VzbuIYFm2ovOpdPSv9gHG
OIFiLc1Y2DT+asb530KSEv+d3jIab6Pj7DrJUldLLNJbExj7baAvG0YewfVF8NHD
NVEK0T7QsgY8bAD+a3Fk95GHdbwUvwfh5SxgbvvP8p5RkKW2lIruFRZ7llhBeUv3
kwfDGdteD9sY3/+Zl4WLSls3yILGKvaNCCjuQM9amx9cp+tQu20u2oRNyBxccSZp
k37/1hf1hU4cwIpjJulY2tv0Mo5ElnuZhKQmecYqxpxU+xq2srC19YTx5EAVX5vt
FzFqNYYnlqLM/fIWOZX5hXZFiH4NZWS6hU6a1Iu/bjtHzVsHttycxs4F08/LUGHf
eSAnq2g9XHtyUeLzYZeZi/SCRfNRiYfYtMrJrnYZwc1weg3oOqhYXvpCuZxV62HO
L1vo2AS9kbgHVJbyvwKZFxMD3hZJyzlNlC2jJg842+ACXDCYovm9GtzOATrBAGjW
sHSBkHsYZR2quuwS9lSoQw0NZAQb9dq2T8lfp8BDSVpfYrUfEl2NehBRfioX/ByF
datjzC9cTgI7b5fvkjm6hoJhru5TZ503F1vKdA/ueLmcA1qCj4RkOMreBrDxIjTN
mo0ItYkl23tOAKWVx4SJQ9Wc3JFnurXYcq2mAZhNKRJo3yb7Xxr1BRIjqDefkau+
67v1JCF7I/eRI/8gASUhA4JVNY5Cb55at5nmNdfZGUkeOtO/FOOXOtMUbh4GOotC
iUb8ABhpGm2qXxm5hqZpAuS2S/jC03L5FGbniAP/IL8CzuX2SgpV4ENVlkgpkuj9
RJczDEk04BK/nzNXIQ8gqUDIgA9Qy1OPFxa6m80e1bncGPqNOYmuM1F4dxVMktNs
IzV9zBzKudtUNCwKp2sMBq814L9mVYLg6I1naCSfBgRoiQIpB71gb8WxP+iqvO3S
n7voPwrLZxjo6k/2Fso+ZLTZvyxoQj4yzuRq3AEmaG8lTSxFqATif4JnzNjZ/xoF
FSH/kcp7KVD2tV+L/DxzeBB/NhzLYmzuZf6fc2ln/3saY4C354GNIIW4yz0l/19g
+YMv95FI/pEzqJvB+zw3k0pIuTf7TJUpKXdnNNItfQ5ujUY8/S8dboI8hlcW7csi
qW6nqng3T2rlMaGCnJNetevJHGokqOTXVOklWVHOhjy1kVJix1DDpLmh77ipElXy
wB4A/bIXO7Cje12Cuoj2jsF6kgtkU2s8lEEDE5OnRq7pS9n0v2HKbjY1OiT1VmH6
iT8MdPYnkBWZpimmvBKwV0EqtOjtK7lR/pyvH9CtqSyAa09ga8YD/cNgr4vLE3li
o7iCtXdBI5lqyfR9+loM03H5sAigbve1rpsX7gmAgh32/et9J/zVv+8HrFcdADRc
3H8Xa2zdHJpIOGY+xQg27arg2nTY3XbFeRjH9T3QtQM11mOZlmIBdTikdraDfcGq
nXH5fC/0arWUqc3ExdCiJXH3TseCbiHR2YHq5MI72AIonoGiGBxuHLy6yA2e2jn5
Qfdg2KaIfVJgzoSkLqaYy0aUaERKxopz0tTX0sHRrVDri1FgqGuRzt0se0l3aAhP
ugJeu89eDRfWVK09pMf1khEaiyRRuycvBVxLV8wOnMxjC0fN8UBAtVwNdioEI0rD
+GdoKJ87ttswL1hiM3MzQsoeLDrQdQQEvH4B24wp1G8wSAHFp9txFIx73kCkH+7g
r65MmttlJbwkVHnI2dksjetjnM7zSKvPzY4BazRZqUMCHO/Dgv3BZ0RQj8+T3k/5
utX1ROTL/Vxae9oPIiEBst9fd5vQGnGmNB5m/HALk+vRWaHIN6eRz+GHIPCNSaMS
mmrd2SUqSZeETvBdk8LZCyi9o8pmBYGZIgTjNDKtjo9IGGrgWCCx+NvCpdum3I7s
qWqO1S6dnugvsiWomRhpCokplmZ7cmTGyKPhaobjHsH8AcghtVVjXoyCcJfJjlck
X1PYFaHJXhEBBCVugH9M0r1CFU1FLWQlv8oBfs9J36KEXuyBa6mS5yRCaedNkjNR
tXrdpteid0GVl6donGLb+qIrGempN7+6p10GVd18m4moBBXWaZwcNlEB9iSR5TUR
hyh5OcjGIB9DJI4z/EKvyifWgphN3r2eG8iiiV4elHTzrzEsKKp9J7G3GdBSJxWi
E4in+zWKRSuTPJKmk32lkHGVxG8bIfIdkXyGOx6HIsTTI5lLuFAOkWg+NlVM6esu
051/s+MGUY7+ra+TDHLDLV3IwdKRlF4QTrypdHsE8+Xss8Kt8y+hFgPAxZDIhhFD
77AIEQK+Nb6xpIPNrczoaQ4PHbF79pjRzPuW683v5hyXMBJ1g9/shrPIU11vkvdr
8df+I//fFDT7MbL+8mwXDkbGELck1FH6LD0kovCMEkM7YNaaTy4EuuVXeu+FVMbm
kA1H90Uj7+LzaHe+iA8cR4ExlAgpsJwxkhGux4UZeZElQ7yn7iWjMV7AzGbneu8J
9I/8Y/9NlW7HCQRudSGR9QV9O+TLoxJ12sydr9kAS/Npm60t/Y3ume2V/z5FTcIY
aW6EJPhSEqjOWCRSNh/70qdrTcjjyHD5BSWusAOQdwJXI4ano2QX23hTRJKinSSE
GoBLS5a9uGD80yJYylCRmLnJv29eFYjjtbAuZUED78t8+CkZZ1uYdTnsjquhmApt
wa8+Fj1s2cksHZdJTjZLQ9+CDo+16rDGkW3o6FyGqCNFtyWL7gw+E9HUB/QRRTI6
iVNMnWJHVlYI/ZgT/wwnnx9uuLVLanMOirj1qOe4cXKB++TiZH647i+z5nEuOebm
whef/+xm5Z+Vmee6O1vUH4xjb5dmovcmJDZB7v/yWmGG99OMnn/jKAgz5e0MLZE3
nUcO4DHnsm3y33pVwgw3tXWNLTTclAu14RnalhKQvmBfdQdqZgWVYFHiEMQyTcif
YISRL4r9MK3QezbQ6T//D6GV0Q7H++4ocbAmwDtSlNAF18WC1NXMNeRR2CqPLw37
8LX9lzWRUm5Yf2CZAPlWV7EJUZf4cpORoq/Rwd4m3o9bdXUUON3aA1pESEL9b5bt
cW5Sw/nzvuCbV49/Dsq6HPu3IyOaPf3n/eWZz9VeSi3o/3vPX5GUYMzd2zBTz1gC
XAbWQOc1TAUiAtlW4ioXYxc5lzm6y4svSBdaoElL7m0Mcnqfmeu0aqO10mRrJnwH
dkzRmBcm6sXJsokQONIsF8/4ctS2EdNekVN5YFz6RPOUnLmUPvY0gFkVU0IUNX+I
N8mMuCxLPyq4CZUVti7GTJiNjkvY9c0eEMV5vn6fDnvaTkIXCnuqyXZCN38v6pYU
T9dbsbuEgY8fBF0LB6Vzc1y2ciIAMM6CwY3AILj2DwkAUGJKn2EJSYQ9e5ra9XgP
n5xevMxa5v0sP21P73UjzAkX9oc80OPMS4WcHu6bJoBxujgMN1EmtIFQ2F+PbnfA
FRhIFEG2p5HauMa20poWISd+Jcv/25q5TPeXM1hLKyTptTi1T7z79CmFRZz4eoiN
L0ykIXxDPCwIHnjlybs+xHiHKPQuVe8d9wEVF1mIvCpmDiaD+JHyKLdgL1CvM7oT
wgYm/R4IxqVvJVhUwoEkgvz6CTFap5pAjB+WoqVIikKmTX9yOTEUeFWlSw5DCaXP
65dET0DEnqOVaIpgfaJ2BXRHnanTfk+vRBfXoS7CYD4g7C6sUHN+XJjcuU1NpFFP
jW2lLUgICI4hnwduPLLPDsJ+wULWecME5ypEEstGyvVeDuBHm0Mv4rm1wtbp2Rxy
siy+oDrIDaP0UBGkdq6h0uy4aQfRbvCLWHwj8nuKyeB//+wjxv3EYQaNzZlsO24C
7z9ka9uAwj1mOevU1IbJOTsKcDiOXMYwBkS/fweNyfv1yADfdDUFD265/IXkaN7f
fsI6n/HniWn4p707xtU+yGMVrKXgQ/NHk5qTVgKJ0Z+dvz84HKa27K1xGEW/zG4V
xF4Abpjj7OFrGh+Va5eOCMQlACE3RK91jB8rGDNu+npKSmnJvEvI4Foyzgn1xAav
gQnqUFqHMnBvbR7M1W+keq6BSBPq9PsauExg7znboRZyZ0pPAhwe23Ak9ACl4KXH
kkOtaVD8z+pA2ekdT4+ac98+VIwyXJtmXiF1Y+3a7HgmoOHtXUM1ITpU5DajjpCK
IE1kmnxUx4U6rGRwDRu3R3BgVZvSEitQK+fsKPgDUKM878y7qa4mwHAix9n/QnZB
Lx2Ihc3dSLrjAqeo6qbbzj04Gdp1KClSSXEhsdV5tNfQPiB+gFazJoqisf49fMZ7
ldiv6sEFuOnlWJHzwO9BibEyKZRTEQ0E/Mvajd1CCrx4snDo3ANiMgROYCxYMGvr
A6M+LDC+lpMW6jegw6LpWI7VBs57bkw0uS6lPljl4+uUeyVlJ7efdjoQE3cQoXgk
fTVRMODPVCjiAMUhCiWB29PZSCZzlYSSZnyo2Dp1WeUCX10tbelv+3Bcs1OLHXqE
dx4PHIDJlQfVMeDVa8s4mMUXxVne1GC85o1j7cMuvr1aBW5vOvRHnxwXBUFgpJPu
R6LnFm81d3DpCGdRdyb6tqIR1MxjelQVQ3qwmUQl/dtOLYM7tjKmuzFfjC1jT0F7
6lzPtL65xM33NJdLs4zVgyqfbZBaQo9WIUVVyGtm0L0J6Mf3KzzdvNNIi2DyIbNF
rXl14IqyLkDILsf9k8NmfwX7t8A49bloJoEQ97Jr9bxTqPm/KYRcbZ8egRyIWY2M
MXwM/r9loAd4nxlaoQvs8Y9kyl5vnJTGm0nlIoutvkFXsjOrc4G2tXp3L5OLLPfT
IRMj7kNGJr5dnE4O+ZllYH2qZZH+5Ow3HtqjHfI/B7CMGeRzez6yh8LRpxYEc9m0
mwlbcKhOikwAPUkEX94PyAunjaYeyuArznsWfqYmVtmOQvIv4v5exWLDRNXwp4xo
PbpQ970P0zDSn0fY1hUf/mZ1PXKvlMotJKigiyJGzjPSh+VGXHDfKziwlEFrAGOc
M8YN4J9IWYhqsOBTcLm5qflSJ/EHeedtGPfWirVn3d/UWWuErC7Y8kT2eqR6W4Ug
fI0VhOA9oU8VdAMgqhexxDCU6VZqwUGwB6Q9i/eW4PJgJPICq2eXaxAHv4/6Tpkw
kK3rtd4Dn273RPGnRM989C+tgelFekY6Y9ooglkjgrEJNsxkW+tf+5xyDfFPjETB
qjzd4zZwsI2IE+u817CrhKXZtp/+/+fqa1/Vl6eYXORP6V+g0COFdsJbKKNEXY6A
aWdwqVQdNz3DTpH85IP7UdTizjgUQbLizPcHhr/Pqc4yG43Y8Z+e6QGI798k5VNU
AoIiKur4CEWeT1ZCR5/7ec+bnJpYWngpYYp6N19SAI1AcUnrUmIBmTEHG+Ge0KYn
WiQG9vnRfVMV+ZnQfgsYKi6I3gKomLR/zq84vJnVhKBXGFI/y2Q7fxEe9zkoLdEf
M9u55kiNMPMIzpCW9x9oJa3nd9lRJb2+6Vi5gVHFUJyJzEaXtnkwZTFyi6SpA8/D
RyFeTXtJRgi1roMaWdk5c9rR2Ix7wM0o6gF+wUkmmK+R+Yfz1LWnyQS8Jy9Ilp9j
6q8zSrGkBTkB+Vn7XJ0CTtA/0xJDB4H5GDEvLKp16Oq0GPuHzXxY++8NrPVWm1y8
BNN7V3OPBOjYf+XQgW3jNwC/mB7q9KUi7SyOvbsZC0p9TuvZlWS8SjI5Kudu9vR1
UeOLeRDHhMG6Lrbb9wnV8lgaXSXnUdxk+6IIQ57SBMVZPiCAFNFMO5xDaELwT6dP
DktUvqIzO46fP7HMk33k3IuvInftUdLXWB/YHNGIJJJTSAmeHAZx/1KgJddmcNF4
u2Q/pQ3PsItZX6JFfkI9OMqjMEsmbssNlvIhurt9oyQCl99hNz50YXu7HphalKOR
owjx6xyQ/1EW2CMtgEy07m06BcxAJFQ44dDLRDVnmvmozARV6qFesIuOM7ctYNVg
aljwoBVF5wFyUxb+KzIwrKMRi4BGuIiXIogzDueUHe9WGUoksYYPe89yhZzq5qWt
j6o44GEb9ZjvuPhWzqR4QYrjS7lLDaE31pW0D1njNfVxrz5OARRMOU038WN5EzDF
hj0SCNFmefGIEm06JPz0YoD1QXhZGcl4tTfUmSnFDODGZN3flPJlaHluLQShlRB2
h/b1+I5kE5u+sbJZeyfUHJEfeBfvRi1UFzhAlmDuFOsQq8jFTFN0majXdwGRtoh0
x/sAkgxXeAx0l0RTSJd9KaDkojoFDpSh2sM5PZd7IfUrstOp5xSXVQzY2Zq/NS7D
IUENJQAfLObB1IE2N2d9Jq23i1dCH4EhMRTCRahwKI9xNt3TcFJrkaoy7ju87ah6
+J+IbiM11UtPoLVbV1G4s0TT8/TW4c6Pt7sWc3k2tO0AJ8y9N1pw9sUjNXYoAODF
pGtg79QV3KSIBflprEiPxJHweBUZCnbd/AXuxvm1+KCJIDyQlasEuqSZG0+NERJH
EP349AlawJqiggNV8lCHFtNT2dOeAtZ8g7xi5wXkhhKF52C7UeIn+9HBL9+pgZxl
1eLcqYROEpkMIs+mlbM3X6ixauF1H5xl0/kGe5Yhwh68JXmcFR9d4r6SsX0zWSg4
YDBiUagsgrZwGsDZnuvLnMP+XLUlMTGZCTl18l9p007oM3xLL/3DTSXQ3MyipEJ4
3T7K7+fBUELzZM9AnHvsxwHlzQeBvKqE/HYXaW4GJ2OhgFlgYtSvDproNl2ejgQy
DvQDa4hnSa2RcXPME7ARmPk9VcM/LOj2o86H0L/pdXpzGBiGIRUcWxz5L7gM8REG
rAi3TFW0pAA1BTy/eZs+gpeSB96+19VYjfp+FtJh4jmMyDUqYsYfgR5FL2hnRSko
WGA5aNp3uKm4BMn/Fau+qVh01Zc6Gobh5DYrPuQYAEZqYlxdBrQbEm5fcCe9nHZr
R2Y1aClAmgwAyAaWrKr3GZt25XbN7/O5XqUsNBwObjf23jtl46uL3fIMP4Ec6Ixy
OlmAwi8hU1IlADOAwsDwkPMQTFFrswnabnSdipSU+5PXPC1CkZs/bK6KwmvVbXCI
f+9JxQ+cbSw+pMmtDcNtk9n3ICpsHeoCPbm31bXPGugy0DjlR7BkYkVm3KRMl+A3
71SjJ6WBLi+6Ojrx4HSvNpI+293oOjWDOLpYtPvu1YEb9RKZVyfG85yG1aLZ9XxB
U48CzMe+yc2Hjdr6IrSqqiNB645NXLsy0jA5ElJR1gGRjWdygwB/5WAg4U8ZXVBI
Md5FeAvXTuhB0Dynqen0keiTrZHWdwfTpt6Cek9LgV0NhxXmt323QCsu4MhH9ycv
7POPGypAXh5nOq9DwbRmfk1JQ4N11UCGDXVACa2zWSTepNrXoVrzxp+37uc+axUO
yHIZP2/HQ0g/GhSlJhvETpVT2ZPGN1O4AIsrCmNm9LjL4x0RD6cW+3gcFirvkIKy
scy37V3c+sxQFyd/e8VS4eZ653hRv6gapxkxA0bruhVAFsOK2Q6/tQUWs7Rr8mz/
lwZMDt5RM5o5bCm+23uWKms6W/5fpBhBGQcByJKwp3gyXFLQX32ulqNWiraTMVAn
RyXYtKn+2TbUH/F5dy0V80gOsztaY/sY5V3+/ZGlv86OuFh99CCqGcSuf2uDkMX8
rhOBw0u4qYA/X3oC96W7fnAX0KX0s6Snx2hL+N8OgQ6q0vd28Xlpf8VxXxx5TKNa
PdN+mDPxC4ZFoARka6AIYZW9Eby83jCzsmFh/JwqRvzbkg/g+2DwniEcWUwsJxeT
wp94irjjweteDabT+kj3V4xhhs1K93Obfsms04RbEGNBBkMa+wZ8lbndCUOJNqcP
s8TTCz08SMFXWP7EMK1aw+ww047YGm2NQ+T7V635f7awuLhC93MDK34K2u1L5bgO
TfLnyAbkejRp9F04t1HF+cKvYA1SQNSBAEvaBe6CLCmWJxhHaq+z7Z5ItqpvqIpG
r2VSgCRJLrJTdZLvYhVOXxQKsziGHogkXMcYYTMfrqL2H2Hn56Elvs19EsIPFdeS
y7uR38b0dgqfroOeGseZuxzdCQPj845hWi8RVYpm5BFquaegFNWc8blYgBC1oco8
T4YPK8ry9ObPN0ecNSqqWEuDOkzzrl8ayExdhrDfsFgSjfDxwH1MdZKxsdSYobqY
R7jawrEEbEiKlEmAOFO7gcHuopFIgVIWgx4jp1qDkI9F+aAiuv7f+ZQjZPqGJSR/
WI61GGoxdrUrgXQjhyXCks++foXAsjJPBjahNHb7pTmW7k/mYF8B7DrL/XyuvbE7
ockpeW+ziKnJ53fXu1r6TJiQt+cuRccZYKWIzh9QwPN7z90Gofv17iLCb5oS/Aph
Eg/VwxYZHye8hePk90QzFafqZNWEY1Rrs9apcMwBK8Keq9h8GcxcHDHGMynGJGd/
kpFD6stGABZTOcOp6ha4Gpi+3PiqDqN4WgmUYGMFLGHUUMXCtmHWTYKAoAc/1rYV
XrQFfCJT6S8Js7CahFUAvN2W6DCyjzRXloYw3nARTktQKLMUxrax/10UPIOgbPzE
cg6Au3FxLUNKcHWtPwGedTFywlf8FLYlqapEtu4sSr4/oNRvUQ2ZNQEvONCjceZI
mksW83oh1/ohN+oBZdZSrk5oP4jiIwNTqU1HecydgECcaVMIXTrjaT+WJtKvSRKl
Ap3ZzEvvtV57JE769gNU/8swixaJd17Ub3kcmFQhGlfkGy+/vEmJBjJdPW0BYE6c
lUTVHlEdIrULeERYMMZYjC3zImeYrJYg0L+M4GOdwc9TEi2ecAROcJDPlBOQHXfz
v25taraEDAMhdSw+1S5FINPu9D74i7GTHm/dqKOQJWyUYfl0FoGg1IUuTriaDAPg
IVGPmIQBDn7FRZylLaClraCPyeHWB6Qb/dS/v24T54oY5+Yu4wNEBvMNUu1SaRhj
7rEd2BY2q6ObmWg9rHKkb5tbO4G4GjebHViB2op9Xw8ZV4MBelFJHVpFe5g9/5RN
JSFXd/MrHYt0F+cISRWQcYOaqdg9VJdJBmswa2FdVOhZJzgc2T9hXyctKsY1Mj3c
S5qLMTgMZpFVyMvK6/8oB8/rufw+yMVRwWymKfF4St8hkbQvh+8teVOmTVVMBLDQ
3NznGVJGdb4Di++oVUFGmXWU6xAksp3sfDFiDSLOiJuMCpALo50g8n1YUxNqRuVj
Lu7OsJTa0ToxsPNpKbjaCtglEFkoywXT54vi9TIpvAcgrulVDRNIhgzaotvvwle+
ccRQsX2Z8m6ObaBuq26x/6huiQTmIXF8LuU2bzM91hHxCnc5ev9x1pczSrwYWRh8
niwiXf8vQPGARsv4I3PPUZQJIG0dqZdvkY0nogkNRMbP3Kcz8IVgX4KtWQHQFCiD
vpSvACU+r8wnooxeH4xowmQGdA1BKizymqGpk73q9lfizRl0Fe9nwE8CxItA6and
hgxyWoZ3dOFqOf8T4t30Q+QxPqt7yPcf2VNLNvfHM88McVZDIFJyguy8MjQY9Fug
XRyeXZZITdiiBf7uzdXU7ikBVQ/UPvuVN0iG+wzDzfMoeeQX36rr3uXLyCuKUEze
t1sxmH0JoDg74YN4tGXkFOHa6yvqiomaCyrrYtRDuPm0kzuZkGbjqBEnDpz73mqf
23GF1qYg+NWWWCwzMHZV6yVzyc0zW530JIxraiLCu741UOwN4s4WN+Q/3wgRuqlS
NNcOWgTT4jxZgmlNqAFOgguXKYJK+ulBa2dyPzDEg0CatRUWZFsCzZI4S44kQI11
Qm8zbkXXiN9l2+6y62WVlaSUOnkf0GnIbO+CdVF+HLMxPkJ4Ka0bL4xaFGMBi96i
EMTqxwJvAQHR/vurAiGbCMABuwd5n3S8mSEsOdtEqIaCmbzmqG5/iG2xHV4rcr82
Av7AZ3vaeDbO/mZCEEDdsb9ZssoZu8ALORAEQfQfjnKKmZxUqBZ0rbqshhIc9bF2
tG1wtD9DtZv5Yk1ZOu+y2OyWfVSWIWJXhakFoLflpKE9YIoQOSDUfrqR7/zS9FW+
hk+YFcLLvMXDV3bA6KT9fkWokKlyyaYrgpBVWsFWP2BM3ZvebZHU0YdXO5KqznP4
581Xf9sOW+IIVtuVFOmpCQVCxw5aBsq3e3B5YIDLAGefAKP2mapJwUcmOZTDkO59
xfXlnvloGfG4iX6k7/wglmDg4MnewsEV94KNA42TxLyDt7EGpKGJXWHGkpo1Mjvq
oi9Z3cekMVkj4K85dY3cmULHi7MAt/eEkkTv1ZvplOTFbvjm7cJGbSaYpxI5goPu
U4jpEEYFLE4nMl4MxomQJHj6evqYnAyZlBn3y1lzDJIT39IQEaCVWmQrWL2hN1Fy
aOp3bX2jX2VEux40Gb1qOX0e6fBi2Z5rUymBlR4jGa5S/Na202/2EEb/xES1xuvA
PRQHSRZ7wsKeiwOL7mWbeeT1SQM0ediEbFOpt4Vom3vJQjBsFmwoS6x010ZVNN04
grjgPKSZbxWNypaheUm2mY6Kpl9K90al/+/S5CN2z+zehjPP4jA1Kg/4nPP6Fk8k
KV/X6Tg5dHin3G6Om/LHrkN2KWcOTKW9KJw8dx4VqSfkxNlX4fnBab1z71MYTLbv
AknztsLoON5f/e9jYgY396EMp4xHnISCSAnqFjAF5RIQ3GJlLq7yHWPFsx4yzEW1
mMTELZcDIRhaQI9DyNDCdLJGdQJkQy86A8nhCFEopSFgANf6nWncO2Z4NmEOkOz+
A9q7CHiyRjXVVWjGMl37xKrN3d4rCz48kipgWw3wglzk/ceCh/E0gZCCp5okyM4/
z9KMKuEE+SBNw6rgjaRolvcfiQAjbk70TjNItGEnlF/2DXFL5s2oWHGVNA+StFC2
aT0fETV9zt7C2WCKXjg4ysgO2TbH7U/n5tpadoF1rxwTZvQzyD40Z+E3CN2/h19m
lVYoORbybaCZTAo7r9fvNPKrgoavPBOBdzel3IgXBj1tVviwy+tOssptBL43Xall
/3fqmBh/r3zp98fZuekkBplLxEm0imFZii13TDN/R19vob9M2o1CDfk2c0dg/8LI
fC+VZ1f7TJ0u+yasej9/kDt+lGLjnL46MbT46jxRlw+spulfZKZNxAGEF0/KF6V8
ZHdZSB+jq/viQJa0EjpZP5fVDaXEJc6Ufn8Db+N4SksIDL/Fw8+wHbRc0o2on6Ic
v0wc5yOvK6yIoKbAxMnRPmf+qKEhTJl3WyCHiFKVexlMgfnishGT2XqtV3cGXAzI
w5W9uOLqrDcXzC5w6ElDcIJbQ7ScKliey0c1ggBe4d7Gkoy8g7Z2+bb0S9TMZEXh
dynwHAUlZD0cAW0cTxdoxVcP2M1qRRzgS3NPZ5ehxpRZpY+kEx7CRtsYSycDOmxO
Z+Vc1Z5mcyqtOd+vCwsh7Xrb9tmmCpFXZj8w/ZA4ZqmWmg8Dfcwf+tB0gKZuHZnV
TZM5FuGJGFR0G/ypGFWJAk6vLUwgGqRohTXc2nrC/WKIyUt3xV8cSQPPGsC/lRCj
OlkeE4wTr2QFRNTby4jijoQYClXDi+uhh+t0xIbOp7iUwcpCkSfAxP20XC4tyslE
fNbjilrrc4d4/p5TrlvlbOcXyFceSrzdkAxpMWAY390hNEVMS8B3pol6ai/jEg/L
tFkenmTqCRpERTUPqteowBEJfCHzCyn6QxMDNCMCkiQOgzbdiJN2THYWJIlMayyX
wrA+Ch5iym6FGL2cUydX3Cn9L41i6DU93j6AWxvt+uzxx6WxvSESNixLoE2CV6iX
vfguL3KwSuPMKza+AsJTTTC0F2uEuVibCS5Tnh8D1Z8y4plzXV2MbVwPFXjrGiW2
OBAMR2/sXE04FvZIoH1XsHEmK1LL8c34DcYqIAl6JP3df9XBPOzcoS7YjaYKHzNW
E1BXGwAXMZYM/9rKFXPc5l3Q2F+nbx9XCNCz3u3bjph/jeMYtj1Lf4IIx17Y7tVE
aNY2lsbeamfHAvrKV7tMogKwkmiqHSw2sJKJY6FZfMW+118VOnevSgF4qfY4IsO6
v38THCw/71iHX7LgrvAmMWa5KOXQkx8HTV91vKgNZB3NBsd8FMM1L/r37E0J+1jt
icKCQd51y4a2mrX070XMKegVPdIGv3WcVwgPzmsAqMd9VxGUDQA9MN7MCGowtbnP
EQW/XTAMq8Anj1M287GxI+7svguBWld9BHvlWa+TJyKtm4DoxFUT9UUbLeb4YVN7
WrKAnULrKi+c+FobvAl3ICZYFeReZke1rP0BZMv4Es/MStUvZeMBbz8+T37UdIVH
/JUDL8wajmKjzFgIzdL1Fep2R3eTG5D3V0m2oiT68ZKJvj74/qVChEtj1UqpMW+P
dnYmpGHYr7OKX+KPqAwOp56eUUzSTOxkyYHh/L0yGB3/ha0Qy+hIOUAbxE/shi8H
ecjwB3OVmgCp67+Ua/g5J/CIVfp9Nk/HLoV7cuFQBoN+7v87f9koWqtGpjHTUm+Q
F4viwBVN7+E8fyrkdcNzvwtgW3wHIzxWmf9PsyyVAg4IVJdZi0HCARyf3ZY6XEdx
+RNKYJem4Ncfg2I1LrMqA8Mpw4y3VM4gP9lKH5ZY1tE6F3+X5iv7A/CVkzC2dtu7
SkJ8W9l8UWAB7khMWDCOrKcTyoonokjloeGhvZG+eEWkVTZ6k7CigexUoWt2+Lb1
Ex3TknH5cCJMvc9WScaYMMGr6ha1dTMh+ArxGig1RD8Uyhm6ml7X5GPTfSf81ofU
qLn5+G5pEC6eX9zuOwzm3VYd7nVmkq5VLWTlJSjKRRu/eNcvp4rfqtauf8MrJlGQ
3bbF9mnZSaL6Hz/ZAwV+GoVXjcSS3hTeCGfokk0SiyK5+L8MRu6twRWVgBV7FplQ
DQvgE83bei6ylXQfH7+FWMMb9zKIFf0hbQb0IFSQ8dmKskPBqeYoWUNCbJ6MgZNs
WtHDJPgElhZOapKJu49hoORfMip4ilJRQaLgrEvd9GRG6Ga7Zdmz7hyZCASMuv7c
V4Wn66uvGgaOu4sXjiQWfjH/kecUwlgT6JvRh49BnOSLh1deim5H1UNrJ3Oc4tZP
m49vvDM5iZWs0SulbGDtHKkn+IulH786gLqnp02Ow9NTWb8LsMt23gQ/mm60q5FC
QGi6NLKjpAvecHGPIAtYeoo4YUrA8gpj1YwHZoEaxfkyl9J8/RsCkT8XuanRL+WM
blObq4aOishh8rHSsUKLDOX6N21/iGMi9YwqC68g9mGq8n+0BENTaqGALPdw7Y6N
Msj0q07Qf0qzDOkbOH1d2Z0Eq65YXYuUcLb6jTX9ypxzoe0fLKuu5KbsLn9x5ULA
LXpXeHq7RSbKvZ96Cyhdgr15azJWjRZKGMsU62PKAR8vMIOG2XS/lLTawV1QyxVO
C5CYSCftxkx5ofvJo5GwbrTX9SF0vNXRggbZEDy4letjBZMtBRr65LOOqKKtGbbB
O6nZls2jz91Lde2c42SeQoKjgWQoBa/T+BipBgg2vIClJwdNJbA/34XrQ6eikQB0
1Q3u6HVwlDT1a9nf/8S75pRtTyuzWBlYOsqGrVzeR3JhSAjg8hf6S+1XoZk2rynj
50swrp6k+7KKYgBJX3/+/nckrJurJkuT6/kEydN9OqPSL1mSFeoAltViZn6jNPak
docRN0DuOb6zXnRq+o1x33BFbMF7w9bu6Nn4dchYi3QZWZbJpIW+PcXF9pEFNCm+
ndiAxfv8QL9tSm7FgdbJcTLM65qQklFQMW4V/2oPJ4Cj3VNu7s+gSs7wEfPSBBVC
eQNRcKDfut+6XblDf6BeW9IhDhm0pkDZU2qpNuJ5MLjPPP+nVKC5nVgii/Pn69+3
n6CPFwJrVHqd8hf879HoN2ewAuj/uXm7ALGZqWG53WRlu7cqq8ehY7T6uxzZQCli
cDpjD+zbq5Mt8PWIK4prHwjMnvvDuYK6GLXZgceBJRILG8lpdStnGJHYlOyf4LMb
1wMwWjh8t0vddKIqQ87TUBs6Kj5Ijqey2F0f6R+ut/fj7j0Pmrm55Jix/DdEPmxy
NWH674mx10XO6rVHeccs5RvXtIVwnXYlLZqu0zKpXpnHnimFQRGURGi5SElNyul7
RAHdBOgT7PiSe1fCnNuPs5ZG1T4NXNiQUB59RiszVN9xnCNrmIglfapHDZeO3Mk2
XEitZARdz1EuQ8F2xhJhHtikwMIMDsfxlLa+a92PeuqXSCFRFRmcIgzfoxT2cn5B
1+oe8CHUmnEaeKXwoRrFc/rCCSgT8ny7cpBqgm5Y6ZMptcWloFDHaDkDKb3abJ8I
+i5ImzhAfBsQhRBzkvsKQX3md/ZSgbLynD78Ilx2d4LNP2r28oODwn257VQ1qk53
D+J/zSQdDhqhpgHAJ5+ETowfklWMRYJoaOJGHnG/UTb+ja1mxgFaxera85Ue5eD4
1yrdaymc008rwSZC47quggD0Wqk13DLYFsUgNeJa/IYWvetj4bJiluMh3QI5qXzB
LHz+6UQQ0pCue/NTTtL1zeeHFSjYMhjNZHWjUXd+VAn71rpXIS+SenvPtl+28dUE
o0qo301WRddP32KFY3GgUwt+yGodHHUb6Ca4VcxPoItSnQSgV7Z5VSuZyX1WyHe0
xBRMtb2OoeLPlWRxcy01VpeDY8T3Ga4MHiX9BxP/Bm00WshaxaOzQXMpf4K1bMD1
N+vu+geleh01vZfRSouSsmTHOJkWgGs//NKYjhLY/QgRj8YzOhqQ+NNbpN5pP25q
75v2Cs6mSgM97oxn0wPM2+CSo/hUVxOBFn51LeQwxuiv0vPv/aB12cufbxjU+9HE
a3LlLGaIC+jbIfqYwHsNFFc5CaINC26+qEz3mP23119oVXpC47m2AURmGhHcOVzz
OchWIhL3+xmS6ghW7WiFrztPIV3BMQWmHHpk+CyNFVf1EcQ3UQ06izamsShvaU/I
dIj99izX6rqUurYwrCeHmAQe4jDla4xdbxfSPF6kpGEK2Kf0HfyO6hgl4TKqd+Cl
D6Ts2t9I+Qs7m/0vFxd7I6ZK/1oYXDvWVRLXQfU7dWMx/lE8Q5Tm0yCpJFF3JzJU
pVP6CBInYiIEnMmg7v1MUEWIqIpxsO6f8PGH/tFfOC7nHDDruErMkGt2iavY+WVl
YlIf8rg4ShGutlUHQrgMgGR2sjnNceJdEyG8enAoklqP/4eEdDmq3EH/yzZRTJvQ
2QB+uzZ04Gkvpe0M6oVSzmIxeNsJyQfGJNQN9NaxFCz75SlLzs3QbrCZiimN5NBp
G36kYlchj8bVAFVRSTdpvHmAeP191lkgzzo9uqwzEqAjzTYvuWe/nIzz5PLPphX8
LQtqp9LiOOdpYdTBu2EHTNwB3aaVVKHNvHmYMaOe417emJl6rdhkFSyWDt69VJjw
v7FiDUEmqzXP2DRsUfvUuX4NaAvfDbQnPz0Ig5vkf/3wFsDCLH6tAQ3p54PIUb7Z
T3vtyByo7SwJnnaeNVyxsZ5la6rSL07cRHQV3V9OB6tBD+yIH6vJh3aJwuG216Wx
iI/weDySj41RZR6tDOVAT177ISaTdt9wZnTlkoRERJnwIeLiPtEc4N+cWwtGkzb3
3l/tOeNb6opCUaIniFOXeUCTpoLISIgn8Q3rqNqs3/xUKn3zQ2kwj/7Dqr6aTiUe
k11+egGesEwE/9mWBXBCy+UIES42BQrj4loI+ZkJ6mK+w0IImGsAGzPgYRkljv5n
T1nHjyodb7R7OX7rOwtUNZAjeycuTZztPznEJEcxmAcFByWas4TYMO6AfjDSVGiT
SJiy3ec4DOx/FPwULU+9VYkV71kZSoVPiqmocUziChrsZC6m1DnWR94bCD+mebi5
9p4spm9r4pgNh92ILzkI4kC5OWaOEKF+jDLIZOP9Sz3KWAAxiHpkdh7Aowhe7lmZ
Bhbeyjj0bjzO6TwFp/iP4P3pTMXqbw1pRJRF3YVVSHX/MZSwr5NBAmaZ5kw/eivF
GDSOluMfJm9zB4qvPS3dgauV/MBy9zaO6uOkV2faDArWMelmOdC7XZTtn7Hrv0dt
jVHe0z8eC6cHwdj816qXkXHiDyNAs32+z76SusKPvS2VaJk0hRJfp/C2qdFjVwEg
NOU4mNAuVvDjcBSXAAMWqzhYkU9isa3pnxRxHbqa2j9YO+WWGvfH7JnnQ7m2ulEc
jbpNTSHlGaYYwTa0St/G5TEm+t3KPZ0gyZrfqYw+u1yhMLYcpcCIHZobgXN4ICiC
rTwfvI50cLoqpLpMrIUXFHJ7j76f25a5Q1+btdfRnPxYykDigTnOwNnQVeEqOurX
lsR1Up7Wrd9coF/vj57tph6LBZHnhMfGuA+GzJMJlWGo9994xchgLtGhptFHyp9u
/FkMxXKqLWWldC08yw7i/bVYKb6mRjCWboMPWJoPDFQLY9TQQG0XU3atlOC2uEAY
D7GswCC5bbmhm7mI8HADFllg/jvIQh0NKQ8OMIwAkRkOCDctrwdyzKvuKi5antxS
L9hieKCwAC8dVvOrv5SG4XTeRyNMviJ6feoELMnU7Vvdb0HOnRD7BW+rHDdDh7yV
aVFXk0whLiYEqg6B0RlLWUXBaQRhXLK4erGRJFjpk3NG7uf3+DDKd08I0PfsRhJB
FExpmyjEqjhWX/nSH9yAln0e5wjRkUGm45eUSyIlzUpNieSlrOWTsPmOzyDWx1+7
9oRQFYNRLxl78JLQyIkkqOFzKmQrikxB9uPjE3eQ6UCD+Fx5BEd2mJOVtHKOUaHx
pAGAuvDqZx0j/yUFwOTjEUwf+4w4q+xpm9d1guR9KbYSxzikK14iHWf2WjhgALeC
kR0IdAy0kOH4Jkr4k0SvjvrXbQ0R+YfGab/q56zDJN2YCtsg1M4kl9Ov/GkX6a4N
9MUm839dNfs+TOFdCcWXShAYjtF1vbM8fl9gUDZCCfgPFKCSjc3k9LzkPSOuugBF
uPkG+t6j7brkciN+vnY0APXiG15bNI9JhrNG8aw8vUbmIe7r6zj95EHByQovP4zx
DUkrSMc1EysmSLeDNPgRxfhGIHGlASuHeBLDWtS9E1v36CRZ4rzUu/aD0/kbl2ij
6dTYg112i0SuGQQ4nti0qRLirQE7RzaUbGHBpAoCK93Q8PYEOEiRwa3s4MM/U/s8
2pPGFJaitWDcoFnwxyor6rGUydNoFME1xGRRCVaf1+SuSQabqcoPL9ePLScMUJa4
PT0cVtCza2MuvWwI4LoVVwJridv7cPqOcFXDUSlUOGHNRCt7d+SBn9CBHg0/QUWu
zOVcQRnFjOvOGF3rIKnD/HYd8sD4y4W6zBiIZwCrbSvXT5CxRRktXopw5NMX4WTu
TtEeMR18b+93iWaENWVEq7buZmFYRYdymaL3jo5Q1sNu2W4i5vvdosOcWMUocl9J
FN94El6hOkCzegtLDm0fzvLpr6kuj/Ule9WjYI+t+0YEnBiTNM9hYjFuK+oTKF+5
6dLw2srog3XhZ/G5U+VZC1Ph6Ff7nXNTN+odpMZETymfFhxy7anu2ZlFz/gDEcUt
8abA8xqGLEe1BCrtOSjdoLZMkGP1ZCYlR7EQsHbhQZtZ9sMBd8Y944UoJp4T8AZu
kBeAVVt3TL7R8AB04A5xXUfFtC0XgtBOZdICNH11CPEdzt2L0v2r0gCUyvp37XJT
RcA9ghHOzADNgCEq6K/6dUnv4heboDhXUA7gDOeCet7/VFzrEl0LoP60Z13s/Iiw
0uqlk45UVo8JK/3muSXn+8CZmS9YVRfUsHnypHU2XmuUF3ZOjUNGWWceIEDbVzJs
hKKiuypv1t7Is5OF9Rs8P+ErHmR+/azJNuOI18zlwnvRFd+pGcNqiJbtUI3jiGuF
95DJq++bGLvwU/YDRrRRreIZ9+QbstQJ2kKA/9zMaJvA0Rh6khWGYJfMoDHC77e3
+hYT29Xr7ouEEJewxYMiON7ccTlxs4D9bJqZ8swaflgqyHnc10XBxJorv1jXsQm7
csoEK5zxRyvPWsc1h4aJl7HWwOnCzI4NB0g7+fX39mmsykfZcHiLbW6yvSY+RLvp
8tEARJGH6kHTwVpuI2+VvN182DfcinIUGikpdQ6L315N/h8mM8rW1XD2DnMtZe/L
KSwoze8X0/SVJXgXhO8nK8POwKmxw2OG2oE0k0bmgosmUh7YW3rUIWPiwpX5iEqB
FTU+NguuMqk/dKVHbRHXwgirwcNVHJmAHYXf6mKAUtfMXF+Yp1aSAv09dAh9DLpe
p3gms5JWrfHFbNuOobn5bas3HKhTnFB3QK1AYmmiM1+9NyLeYjvibQBSb3TM3OPo
3tNR3IjMzCw+g9NHksSb+29cOb28Nbbvh03jlICtrxtCgSrDnZQaDvZsPAEy3xRb
fowHt/eNKzTbEJRH7uNZn2WEqMB6AIrr7VgG+BZyQYzrJ0IV+hsMT1G95fVm6k3P
dLP7uQni1bcOEhQB7LiSwMaUS13EqTbXgcnueGJQCYAeVNHljO/9tVx++FQmNkN3
67hkIB83twqeTzk10h3ymGCcpJbSAAuXC2l+hh4wAG9XglzVJnkUiunmYvzG1m3u
yC+whPj+JRuGeCO7JwYjTMUWMcq2at09nqnjliBbsMKMlyP3o5lK3oF5hh6oIT+C
+takGbP+qV4vzx7+SfEfh4iZ8sByPaGouIuXjdmK2bDzxaja3FS8wRdq6R0gOn/B
BAWtl1bGiN49mdg3fEokzHjxQe/s0hHIa4qU7GhHALNHFLk6gAXdCjVtf0MKGm7E
qlLjzGpuydBE3TcV3PGTO0Dz24seFMKaT07Xmg8vpCD8uAAQmlFPl00FUOIupfi1
BRdvcf0tWgex7vbEgkoUIN3x+hMzrSs4PY5t0vf4CeUaC0EeGWTGbmLQeCRxrYWP
4AKRpFOui7OnmAk70OBL9YREqXrR8XNEXpW+XdfTolQyR1V+yifwS7oo2Nv84rmm
kwNg8LzoRVIZITxpsaufJpgQwfGK42PimO5lKbN9aJ24qr7mjbEgAjQtZA4qNO8P
s6Tw5xTjJ/ADyGH+tW3eWjcMeU+z+C4Sl9WYVcM6gSc5wiOitxxB7qruyGRVQ/+G
LDvqEDlZ/ti/7swHJJf/tTRMKCT4aJuYbqyRyc3g8U8pvkUWAgJAIEWkRzsSN9KI
x5Uv0fsrU8QDgG+Io1zqm0E4rUxOKLqyhKqxeTbAlH4n4A20fY3MsKUMLewpUxWR
1+JVLUZ977S6mFoZdI9X9nGtKkgCrsOFD9qrbfxVy3ssiozQ9J8B5V9TfBPI0jf9
7wze85sK4Y05Cs+fR40KmCOwtZFVeMds37I347rEXSH7TlkUgo+3s7dJxeKNXqCl
EnDCJZ9CNTCpB9F9/hDwU58p001+lz2vfuUA/ldJC/158EpSDRfd03hLKcnyKzW2
5YvYBBnXt1h5wsNuOWQGExsoazS/monf89w0coIxx6mb0qDy/INtZww876+znVik
7vAEHJC/ZGQI1Hw6TGmZGHwvCcBfkGTHBZLlBEiqu8vN+YWBOv56nSPtA5it575M
3sCI8VXUAtAg/JH8ff2dgO/KfmLEadWEhXFhLA75lHRleCc1Ec2ZiO0XMKk+Anmk
ktpbqukvz1CZFLIAHXt1PnzKIx9vz/jjHGtpc4lY+whtGfva7lz+LtvmS/kaZkZM
U9MC5dFHOo6af9ULF7qzn+Qlxn6BNs/Ouf0eCOo3SvrHkJVG/xzjTkKDHLwQg59d
tTaBXKdBfQVCJER7F7mp1dtG/7JGk09wnWV34NWzjwfuOhj/pSJMvLLQBuHAsJP+
8Fx2g3aD6dMDZe/a9JbeOcNYHOyrFNX3JsWpJKjS3KK9+Ga8V+65zsCktUsr8zjI
qoA8Y9bzL+fFVgqldZnzHWeLSyE74rMdivDWALTQSbjGS0ItOh08l4QMhs2EKdPZ
waV5biQSwgv6KiadQQgMTNGNsmc0iyOdyjkwRRI8JWyjy7FzBZT9+b+SnpefZd6p
TRtagD6PNg+xvJF6qwZgIvVJ+75gVp3hZZky73IFHozmNkcHTVfdnGYK3oxNNnkZ
VNSfqySIgInFcUK+dduVLApb3tBtxjfhGyPqN0JPDLeCgOxE1fpFXbyABI9ad2IH
OedlKFQWxwg/Zq5D9+FdX1bQkvVvGoNOnYjX3SwyGvHf0BtoW95nslGUlgWDTmm3
5v4hbp1N0UxoFl78vmkNMRXFA5P+SISAazn05My19+gEGrsLb7bKji8OaLFhGL1G
VIEa7YFntXrybaznv2qRELJuRITG9MyotMf1Afz5IV8O3zU+MTvkm9Y0MA8bTJr9
0Dw1tSL1KGG2OT8LungHF3ND1GAUesLL6REBV0zl698xutnIL6+CsCydAPuD+WIG
RUMsMF5Vq6dBByoD2Ya0ky8HAfJtf6GYPmiOV6/MPZoq8BfvQ6+D+2DCZrsuvSN0
V8L9axux8i1xkj4PAc1MHkvxmLSR9T46xQVkyc4vKt/t7ACrzezXAMkdwnq5WQxk
AMu8s8h+iBcG8UPnU9tmNmV5VaW4JsII+SHphh8Vby1VdnPG1vMXLLMBQXqme5l/
NYUu4yC+g/pr8Ud0pBut1NzHbueBXLzK7P9vwSiGIueWrG67cDUJGPDWT30cjXa0
bZ41ulpk0dJqzaHLpzfne9vZj0Izyf7HgjlXM+btdI17N7UoYBDVDhuBce9k8jrP
Mq5vYnj35eQqMOk9e7JYBusyKy6ml2j4EsryI4jeXmlymyiU5BH3eJupk0utkwfi
kr9jzzgG3nKc0pJpK3/xVeliO6uHh/4KDStw5xTmIw4AFNyctT7+zPaiP9htKFmO
/wuo415vFQotlJd4HGOZytFR9pRW8a+L33h9PvE/EZTOaR5BKhT6AuskIGnoWme/
e5Mui6aBElB0rF/yXIMgfxyaD00dlZT5m34iDzKb5yamF9Sjb8Bwf61mk6ZBblEb
PNWC50O47K7iPUO2QFYqIJKHyejBcZBXvC4QoYPcYjqcqFik8USEzkOtj+8ngupQ
x0kZjYHQ0Y5IkSavBFnLrhtUFjNPIvpYAgppfBUrzKkfqfk6PEJPiuZ1aAhSFK1h
YKKTKR+HyZGYEiUM7BjOL9K5ssFh7xevprubNMq4MIj+1h/eZoUE6GXcj9wzL20/
4kDvQHNg9Ot4Ld1k746sTmDFripE6MhRhO1RjYzKZ4wz9MgdgwbF/leg/RsXr3eg
eGwvgpj0Gd7PYZmo0jSKYAk2kxPT0k2S/MKi0sY0bqtJTNMdbIa3NopxIinxhVKO
0+kaX/mNXLgTe0YIAx9WVE+xsMb92uFNjSvbUmWoqCjaByeosMrtCDpaQXZoAZ4M
MtOs6hwf9ntcJKrpo6ISb0tGK5cIGpR5/+u0R/VM8nXC8VBIN0Ag+/7AL90Ign3U
/bUR1NKIfRMKA79/yg9FX9C1FUdwnUV6HPgpYbbAG5d1eyYk/jxD+2WTlWlgu+Xg
Q/TBz9A0WwavUoFMSXIojSTvTtdH0pOpJl1On/agcXDKPOlarevZEoxTQb0E3LEa
Um/GNFTVejwk+5IszlULUw2ThcOylxt7oeldSlhZDPH9fC//Ww5G75YZSwWUBwgl
ek+4mdmMZTpPFJJhLC8J2VjyGE6Ntym/Q8Df02zBViL/Kv4x+bycLMkh0/Rgz249
898kqWmc6WWq5Frn5kh+PFMAMUBeA9zJ0pTXrma6yI1fjVWiCGp8QpZcuOxjmtHh
dnWOgwtAqS0PbfFhh753jMIzZkAtvVazR6n22nV4LHlkhcS1jSeDIq7w/EgbZs5k
ElZkduLSRm36iH4gpmnh2Ps2VgHHqf1zhTJIy1q3I9jG7US9zL1tJp48vUsoazwp
LyUnEsHJDpoT4lnLS4KOtKBB6eUnYBiOyg6g7pGhtHg8eQWsSH8vI21JeLpXM7S9
Gxl4AGzb5XWxt5srwwipxjpAuf5l9pF/zyEGclDy8i7a435mkfWY0U6YcB2jCQQB
8QsVXA5QP+KyLZjyvVfhdjBfz3OQD/1jzDqfkD8lC0DyXE5UgvSTIRu2ROmLKyoX
HjzuRodNcSbgSVCNlEcUfmHaxFlMhM5AVGoAxDXeETwvKFc99BqSPvul6DNsk2J5
Vyom1yzuP8AeIFP9EAxKMxa7xyf31a/CtVakCtWylBIRpCrtmLXV4TLAqmhIzbCb
u5712m7ijleH1511cP8VVXF3AX/k25jnct8Gx4kXA6RRZS6bcZVWi+wzAt/RW63j
/STT3rwQKA+uq1DDlfRRjm2fuCzGM0sB2yw5N4uuodF4509Wmm+pxFx6l+sK3WNP
eJ5PFQ89xCAwLaR3qjlmLktEqJ2scsfdKkWdohR0LtcmjnpN9MLXDh6zWI7FgDcG
srC2qpPQ8IZihHeZZBLIH6nySdLqeC8x4Rd1bWGqO135vVc4KBg9IdLfkKpttjKu
CHJYErAkp/m4t5iDkVcX39OLQi+ea1DqVelWuc+9mlaESQhsVpa0J0EmhGjcKCR2
J7PMce7fBgo181t8Hoak/qYhObIgpOB+3RGiI4z5OvrYf415v+iovPRXLV11SnaO
ovFGx8uSMEu6noMqbhIgFVZOjfPrYsrVPsF7pVfwynqpsVLcm9slCIkTys/fzi0S
NXxb2VDLtUMPnQKc5YfrQhLsvJKcfmFB33Px602pEACnF3BnSa7sW6bpNi/l0IOS
bwIHXsCXWeHFyZICCYXQDoJ8AqOtITH+rFbYB0+syRzSeVYF4BOm7HtITY8nIqXk
lqv7GU6pS6RujhB+9VYy6gi5drdO95S1DUCn2E3u8AwYMOVM572OuuBgTcVgrkD2
BbO5L96L7c4gEihuLn3u/9bqaJvO8YSC5uLYKUaMXTu5vrOEVMDhPiiBcQZboLKG
+ZMXL5D8HI15NNAfVx6Z/5IZTrIvgZRzLMEfpz2b5EmeIyA6naBMSALY2HAkzx1u
fJj7pb1fqJVycKDdvGzVUytmaq5B63puapXqEJJuXZI9jCHJ7VBHe+OmvUqJqy2/
5N5tdobI9V783QnwAHMyUU0a53MspUGkX0XVSAtM6eMoR0cRsYE5Le2c6Sbef8x3
llWJHbych9l3+/ulOHKmFakY3oChqYl4KMWfQob/dow2VLa9ecyyZ5kyvpFvnRO9
XuNv6ImSh1hBjOEJ4LStGO0EuUsN6Q1VYA09++NMMkRHfSTJyApg07yhij9+tguH
plnc2tTeEmLSKPfEFuLRH4E9hFQyKqz1K60znz8LsaRx9pCu990cz8z15QSXVQYi
YRhlVkX6AFw04y7B1dMVnBrnWZ8UOxz71lCJfeAJc/xoH7rNuskf1Xhvp/9uWwkD
Ul9HT3S69VSSFy/uaz6x/8/mVdzxZEKTbTBWIP/fwRpAt7vGTYfJFlyz4MhDrqvX
1KG6Hp96rsY22ulJcb6FpIZoCnUIInYUqM5qVHVnW6rwop1GNDCcjXe0Xu5TBThZ
xjBM3mZ3zD3k7tR4R3h27DAizyQDKRbtLflXCFfPTITxYa8vmvFZ3wII+gdJOceL
kmLOifc66bb+Ef/LNWftLx2z0lRWUnnxcF++3nPFPi4Rpgfhfd+hD2V+wRbzKX0D
ab+o9vFp+juVidqWMrflph9hkJVLuxmwNuXx4UzxvctdiNMi4QupYXtAJ2jWPNPa
FOpUFSEDl6Xb2MVSzwdcBsCCLyMtRP4zI21z9Up0N8Fhq/a43RAvOmKRrLNa7CKq
ws03M00eLeb2IQBBeUEv645VPeopCzVQc5g2G6TzZcHkxY4M10C26eueAlzowW2c
XCuWB3iWUwKA7UZUrnYcfjeCDZy5kjmmLX5hqi88YQL6hqUtIGVHiTYLibC9fMg6
oAaGvJRuNVbeP69Z7R01lJ0HoVLQaVTXg7ZO4Kz0O0I6Zn+2eueT89k414tIjAS8
CLJ7si25cmV2UzEiYuecqfAkGVaD1e7mJp0slwv2UnsbMpNJFWCERJw1+bkLeWaX
jvFKp+f+PshzWsJ1bV7l2b+yQ+fdyIRLLbM+/YY8skJUisP54ICjoq7dUkcqDCOL
Rdkm6OT/wxHOC1BSfcy6YPigCAnxZ9Ju308DDOn1cHC+zw68vyziwlEVwo0vjEdl
Z7oMZmIZpMWV0P52tt90Kd8qcNZNUkG2sTC3Y6aGTtWDpq3fKS9MB+XCatw1natb
RZD55CTiZsoyq/Yvuv1RI89uY/vzZ0ruEO9HLyiZlDpJWGBJxR48Fqv8QEjuwD+u
tATxNVs+dorFOy8erLPu+145aRUZBPcNBHSJeqyPr5x30sXVxhgOaH6kBLqYFFka
VwkQJyIDa6i5gcg3FqDbaoRXN9NIIk4RVG8AGRd2frr547Ll5/KMn8R+CY1Oat9n
HK73qhrmQWheMs+40cgGU3TGKr52lxPvQ466pvBX9tSCGzXFj63Rf5tQG9qJXXjN
NEUYo4dN31lfJNjClWYZE88vn43PZrZYJYroH0JBsSf7jjDxRojxnOEivcZt7Al7
+esGDDUgJUFT0gIixr8dTU9LwR3PNhlqUFBn9J7karFzRHiQrsrvPSYFhzc5SjvY
2OZuWgkxlqUBeSlTZlUXIpUcE4GF3PoOlR4GfJ5VjjGWjnS5HXWXKgx5a5N+L7ci
3/H32LFiaHXVZqw2WX0ehv2l7ui3nY2BBTFX39aMzpPwKraWhpkw8E0DhCU8zpRI
ROckQ/dIJerqpyTORABoBc/iBGITs2CGi/tnhmREQQ7Bxq+uEY3L3p4nPzM8Aytv
9iCqBRhefn/9iFW84/MSALcHhseB1xxV/0jjNEanNAXTo9fhGQVNvqRBjp9KfU6x
ik9phEFe++iBr1rUZ7GtNF/1d1DOA6p6EiTnuEjZhg7leukLV1yGi0hDv/zLH61M
3yD+/a104g/1sqDFQghOo5cqN5ncOYrAbi9P8mKh6JGwcN/jNuGRm1fxMpIG59IO
9fneaUie7pY3FM44EJ94SjB8gnaDVTdZSsBUfIi5w5521st+igBCOhoVZPClMoq9
uO5PaPfFc8S+S3n+1GQ8dGJmXT0ONJilz14EsXWLLZbDa/um18AgAQYqPO06bk42
u2mXXi0MXtae579czFuZa0GCClww0wxnnsz0rUg/SHka4XFax5Pv86zPgP3vgDPD
srp071l4bc2deau7/CsVNSTm5hhqZ/YZCWOV993YQvrw8MVerLxPc4TG2NWji3sF
Vpx/FzDfLsbS9SWC4kCLnAB6D6LfINszZfGNN0PnxJaaqMWpP88OWvkkrnFidTMT
go3UM8W0Rn3ilitGO4IUeu754JA3X2rZTupLLm5Jz6UNhVKmLN+Y390EXCJIhR5Y
n24p+y4Wa9b8F6KTq27hSUCpIHLynoDFR/zJebOKCA49th66yuOcKMJ2gXjWGC9x
3jDC6IydmLYMjzy0n2UKY4jS/UJJYJRnpGWl3PAPOQ5Cfb4bu1VrWX2ONyGpO3pc
UDft8oQMnpRAqSr27Wl2QuzXylZ75JQRI3CfvyAXUh3pgiRZHiBrr++RWgigqtnM
//FwsWFRggqK99yIbSFDc5+842+AXh8pf1HNRW5zlBBjnsO/MA3Q1vBtj+dAOH48
wwxhBzflIfORxdZcRGyha+W8A6DscFhXi5s4qjGTSJcF1+y5VqO6b09iV+P7Oyuc
aZM/OmrT1HkWhVZISHc4XGGMB8o1f6mQHD+97UbTuPHYzbzy1QhzgA5zCL8Gcp60
MiXFq+NrDCX33DG8TN1mapkZTLboTQs9fpYej8JOXhuB1GGOXBh23P1gN/0vIJ2O
0W6OkPstz6t9I30CwGKHQbeLrY2awD2nx4bxXRaJ1dbzgeaT3JL3vHH0b58qwSmQ
flpDhIaOQeM3h87+yQIrd9RQXdRk44tXT7m0s5KsOyMmJOg2LbwJkyre0sk8li6E
L4EIWGe9wNUriQpjBvdupZ2xgV1wLCkeVCNmaj3FIdyLtYaKO0jYwZBEIhnQVFAW
CDbpRTpWKwC79wbjj7gACyuG8zzsXQ+Q1ywxttc21+pDAbEVxFrXRsswNcw6AS0y
2g/MRknSfoBoYLCKSbFGc6ETidPGMOa80+19GHyw4+WBmukDHNyJ6p7AaU9Z3NxW
suCIffkQx2pH/mSSbgIFcMGQG0DLwy9UQ6MzFM8VUicdlg7yBzUAcqMGln1yrqNX
WvDXNWWALIJQ3b/1XD3PBfXlQQi3030rCnap2FtmO5+Losq4JPmXlIDxRa0qGyh2
D33fcvxffoljpXW8PD7hI2F9T9RBC432V4Z0s8hD58LgXRCpboo0clUg1knwQGyH
VO/hLTNUdKZs+m1NBescjUTNGWAqtLkHGI1ggs+m3mfEgO3dJqfFw2AaQK/4kgca
zDFotynNGduOcUiaCk079oX/U5FO2+dG9Px5HCwEAGdaitMRqGFtB4Ph6bVv0O3u
wYXyNgFi5Q6Y3z4MyVpThhrYTQse4Ow4O66cuTfiLdSW7iuV/e4A+Kwe6L0E1DC6
C7NeiB2iXKaPxUw5d2c/pVaMYhPYe0/52n/ghVYj4u0K4l7uTAvcG3sClfKNBXkK
0/cbXq3KGcjGm92quIPWi3OhF4ynAmnVUqJLjdGSSunEl+Zmd8KcXkwZLTDPehIG
FStQjt3FLWobv40tvsuNvzzUphsZdudTbK+11xKPf2u02STtPP3RkuhQhtAAeRa1
kPTloynqFtCcapUdxOnzr7ctn4eJoYNKB+naBBaGwmxRrJ8LgyRusPjaMDcuqdIm
ApI3qgMdVsgoa5LTvnXNloYiR7F67aaISij4eDLMn0heBivl0JasFX5ssLSnurHQ
LEnGuFkBM9WpM57ssyYuiEGwKG/Y44Uo53aib3RyyzyhHBv7zYnwp+h4IgiWvky0
pTNNx3QahfQLNFBneZ4UUkdxWheU+Mj5hBpef5ItLWcfXSBWQVr4HUsyMepcGZIz
2nWHI7dNvS5O1Cb5CeHS7MEUdbn5KWmjp9z9U+g/LzYAzZ3k4h+gy4AvG97ynUgo
EbiPWh6lLoPj5in7PRx7+JLB19qzykBsd0W7at5K3+GCaBz3atQGfjvUIjXMipdv
XdN5FNEMYAUPrjkarhqDr+kf5ksDvQEj+VfXxNduQWvGTp1ai4n93JElO0OI1hgS
GTghxh1Mir3y5rvDC0JhtmmOfGS25P+/gw6RjsN2BkJLQd0BR8O8dLSRY026QHxJ
yVO35Tra6mqAQe+37BLfQkvwPgjU1SXzQhfOwYxI3IwC6ELXHWVIuT3cV3utFvXj
oiQz31GwgHNRYipR+pxILbBLGiH+TPvn+SkJ8RofP2Qdz5JCl6RuUAcCsumOqsJD
Eid0MGeRD8y3NCREjSmpqhIKGC701S8l228Do6yCm1xMqGn3tkNJDSm/dYwCV22B
1+slWJP1Ca/Et88u3V037OCg4yIaT7m/QQrpNkoEDKpxvnxxSZIwM2uDkL2k/rhl
1skF2LYdJu2M5qktOppk5oeCavP2JebNSDwrlTJBwjNcR2+h6LjMUkDtwCOGBNRo
pVsIsZLS1gZOszj3EKGbgHG18j1N4ssg7O+mvGv0E7FloxfQo8+8pOTyitl3Vvkm
xr7+RTbf4Mt3QZkCBxSJIewQUk3kEZcPUS20sLv+K8jzA7h48i2EQvopNtydTs2T
elqyqdGoWRc5euCosgmz/wHy2XeFKJSsqdm+nlKyGnyJXZaghh8PFGli7+/NDdyS
CpWFzBKg+M8eBOZhFXXcKuY6t/IwqhGiIlYHdsbIgUm6urCeV6Wa68uRq4s2DSpR
CzFv4fXpl3aCrh1jWyGincV45tjInrZrW8cLkmCSpgdjlfeJwLIAQgB6qidkSWk+
eQafsp0BRIrZx/DLrfrt2zGnkzQnyOaeaQrk9XVCn+sgOrseiRFhmPBPQWPyiSk7
3wjg2hSlKUsoNOeCJXikhmhUtsp2uiFuIMAUCoRvkhOmtSdDB5lcVPfRPvuk3Tqo
HmdKgefnBXFCfgtDNRnAdqFQivKoBCYms2O/eOJJbWlBt9u/yYx0iaF8R4WYCcpP
AqGBMoBN652XNC6+2fh15LWzHWZpkGh/qhhw6waSikFuH8vTRXuVErNJ+jnxpRX7
JdqAEAYDH/cPcFnHOPMSqgPh6/NLeekgHOVlMBn6WjxHlOv/HvZktehAdBnrYB/k
gIbpxBiI3jq1lMk7HrAgwFkmOfFTN+f/fOAflFoy4PvFE5CMs1hr9YhhSbN7PZRK
dIa8MIQGKe1+2FUOqru4mcG85D20jIltD8qGXWP+l2fapHmrKNNM4Hwy4lK+bK32
haIeK3dhUI7+NTqU7a7W6p0wd4xGOtQsbtGmHgEqUVhFf/o9VBS6fSW2i0/HzfTo
UIuFsZqM/tDuuAbuVt8AVfaS/sF16sPAtYgqCH77bZC5bpM+7pN22bwa+ku406gC
GbcZffosgwFC7A0dARlWkFCjqqlnB+XxF/Hx5KQ8ar7MVbNE8pTH0Sdhe43bzHVY
xe9shftBnQoli609xMCYd2zFqQZBkwlhUS+f9wVXcWpC/esrpHjcujGrpoMMVNN2
Bq0cYAmfv8XOfH0LJBZcHwwuLXn2SS6+bxgwZvn5q5kjqWWlDAojlgZdW5aE0zAb
ftDED7lsJYKGCNBOSMRQ3J4A5YJHQE7lJGx2L8KVnGlbvNgKJO/ZgVwDSPAWKjvW
Jyo+r5NVr3+mwoQaL3c/OhO0dPVf6bOXKRhiNEnrkOQK/78V7qPoGwafmuhtlBhQ
6A2BigXYOO8Cr0LMfD95IH4N2+NEsJoErD6Ud5xIEuKR0mlgD5M3CiEDh3AEz3zk
OH2GHHbldZ09BjoEIYMtSHR7V1o9n7rPbzefzSjykPxZv9CtYQQFMvFB4o+a5eT/
khqJfIBJG36eqX/QuN1lHxuCP/v0jzsbp7yaCsrscnWcREEkE3252faqbzUVTrBz
v+TdVPyxfepooB7rfroK9qDmRUL0msFsIDa49aHv6Utrzz0fl4daftxcFYCD1dXv
gZbP8nx71xEKJl6XQA3SBY7SjE5WHXWRtVYAOBKpxuMpdZaJMUzdWOY2vBptW3ca
qufg8K2O6DwXJldUHvTsHoNvjE9EHIpetl15hgHpmJRWIDYxS6UEO4rkIGEWoBzk
vd/2orCPULJb9i/r8tu5WH2BN2xgrFuZSZMG1DK1w3TkPV1y427vPhDHxPX+CLsJ
t7W/5rLwP7HBlvKPdAhp54vwqe5qp5RjMAbjUUqSAx5WQqtbxJ5kPQrdJddbyhv6
8WSNvAS6uK6BU8GrniHQyIJFrhKgE5XttAumZMqSo57uIw9TuNSBbHC1lASTVT6m
zA5tdNDN2AwCF8gXM0ouMA/y/edMQ2GzyCxl0bIK0IqSahAPdvA+M7sDVOL5WhwQ
4cEnUAcXsxwp2fW+g+s4AWP+lopIlimZ/QnVqNvTzKThMZA3bx8G1DqfJCDHs1RN
ruVZTHrZURPgWozSig+VpO8ISNLyYeJns2rDH8AqsqoV2UglOQ9WBlGzWJDI7VKh
BaycKEwoQv5UA1UwpmqqSm0zmQ4fmVCygQCTocchM6DwAKRv3Z40GFKuuF/tJBFW
aDju7NRtWbovlOei6sUESVnBxw4UbHzKYxQMqIDHpu+0lWv6GQD5auxbZLvt7eoG
j9uxQoR99YXDebQN/3EzpndxJcGu2LsdycOab9JiEF+lmScer6KRZUt3L30IPbg/
97sTw8/sRKoYeJZwNVTq+A+axX7ixNYMCl8U38I6pNF4a7zcdL4qCTS4IoutQYL9
vun/E+wa8gqt7Q8LvzOMjxX2AVGZXjCNQE+AtTNnxnBZ4mJtXFBPsAHsjPO8J7sT
QmeuNcmWcCaabeIgrjoTXQwtbxlfeSC/4D1yC9qlOTi+5zy6ivKSOLiflLa/SrbZ
RWftpidBgwieFgJ+hL1fIEK2zFubxKtrBTxE2V5UL//lCZ/6QtWh2mk6i2t6tW59
y3MwP2sIT1KNIXRgQ6TdnB9gUZgMFgCvenGTCcQOnJNZiekvpwev6ZyrUa253cYs
7uV7hhhn6/hAD5AQbJ2v0itAkMgyMWEAoOXt9jpyEoQWbKvrf8Yo/BuwlJ7OyUsE
v56HhUZxIr6NKEoySRvv0d0yA2JL6xfc1KBWezM5M9WxdUdaIHHP5Aiw64I5MiLx
jpHvoLZyUOzJOA7UbdZWuFR7lrg6Bjc3cxF4Gg1QFDGpXEZJ5ofFVsBw9CzGj4av
M7PvJsLYiWTyPWd+et0YH5J5CDn/d1ugc6S67VtJ3kfmUyc4wVB4fns08PeHw2ry
4MmA3zwUxGmpcFw0kDfasyTIZmgdtfMhdvC2zYT/XK9+00JtnY0XY8ouB7GqF/l1
w4GzIhPnUhk0kqhqSuo+3bZyO95iCrq5t2cKBf0ZgV+jQXizOLLJbt2frHUj/7wT
1YTIA7pAzPvd0LCsjfS/VjvPbQu+2VOxh1De5DkjItzucaNrOI3Q7glrrJBd/7LG
8bgTJXqZVBN+54QM2W+SQr3NkkFyIbV8IramlZkaIwQRl5pTHF6BbwGualgUnzRw
+Le7nj3yplEnEJ0usDrWmp9YRu2vYd9K790Ljwti3UOR0XRbS2Ppi3N0O2/Y7Jv3
9hrNk+IJRSELqkaiFCq3V683rH17RvOm8+C1w6nhYi02RvzEgWXE92PnmstWWfVx
TaNephk1typ5FuGBNiOu7QoIKjq1zzf2feWTKFXv/yHWm3CbDP45ZtXXk5l/HgKe
mbuIHyz35F9c0rb/XprlSXnmPmYYvVQ8B5ziFLFrxjnt/f1Xy8b/ISKvyArmgSiR
ccEqQQ0aQ6QInz4gXk6ezACjpmBYrP5/4DtXv2tT+adtbn/hW0UiEwkBqNub1ezB
P/M+P+RJ4ltIhc+PZTrHSyv6lq685EN5hNIazIC6L4K9Fzfg3zI4uzjqi7Mm3NMx
Z3Pf0cmFCrRMLFIneV3aQ1RYbXqnw3aQqxCTK91Rroe4EV+mBn1ZVuUO1IvTxMyp
EFPBbDnfBV9RUM+LEodHH8q+NNWA5cyoUCU4pca6aX4pRMm0GqdiUUGSEDRUcYPx
GJsx42/8IfgyJ6xfh6CIBc0kE3GOjZ/3SIhCySYw849m9zlubvs7E0eBUxHkBHg9
ExK9kTrHLo59yOQLGSz3sVEf5e1CJovGfauXldGA1fCaCCJFcuM/Hc+1dztbnaUK
Gx0VeKpmsI/tgNfAIFhSZpubqGdCCNzbFlWGM9t2bkE7eRGBm2Uhdh9L37SP9Pfs
h8JHo6cOmtOp9udbfnbAJDGWRNe9+bs/spkoeokOUreObOnWAjOswmRMCQjisfu6
BeMlBwqcv30ddMEZidMsYeelyHwiW/dm1f8lzYJ7R7XX5Kr2HNpRtoFCjCmaNwtM
C8rg+fMQfqKSupaaEZE22nVpoo0y4njOvCQY2D8BILa9iutoLfFl2Db9pF0MXnPu
hVM933ECN47So3jsgCRWH2iJVuv4bEmvetTg/9mKrs5fPVl48dxPO6/jHCimlkAJ
EFaoV3qusr4UIJMfVen0FEm5eEF0cOKAtVQN21aMu0HT74VBd1q8Bww3ONsqHzM6
BrYrTKMk2j00T/fhrNlG+/qHLYDzHYnPZlvG0Ee9YoQkCMVJNFBAqVU8uxJX4hwv
GhHwWeju5StUqoFnyKLMp35g6hTn7G3dwugdrxXRnbKl3kmYDPc2/kx08M3bNAqK
CfM9gKNou7davLvPmDUlsXj72BG+22+YxZfeTAK8y2kVR6da6To8m0WUIkWo1VGD
Vb1g5INOCPe9lUnjRM2e8KEDXAoab/1uGXvkbca1XAdJlsJNvafuA2kDO7ivOuD4
+lB42IQIg79kLtwgFMH4yFFcxZrcT1eVPj/iBj7K7AyaGk+PBr6jfKuSPQ5HE8Ys
StEYgr1CaDfgzxkhg9x7b0ObRH/7NrUkjbsowYOYSXs4rc7cM3wJ227fn0sKZ8RL
yPdPWGGeuJSlNwLpZfOjCJplucHy4MSZJ+7tTLgmhGSGO3uPtDWkwoTp+sku7Zyc
yWyNF3SUfR2MspD2QTIzFQMKOQE1ynXXTpIGdBDM6Zr9mG5qq3EiIvfpvQZ/46uK
UHjWTFkTp+QX+i0YV5CkuPmyhT+iV6cgHXnf4qnKvF5zwUXn2VPWflx4PVuJ9zf8
2ZE6LQZXmFX9BsgTAFJzLP7n++cXcBU1AGiPsiguSEO+V3MeZy/62iSWyNsJuFST
5b20K9frmJPft9gwWaVW9tCSD6kFULHyPIkJanbsbBgzbrG6gOUslagPW6uHuz1n
c08T7MwJb9G+QRo99noedl1+A04KamSjddOk4oOrrQy91t3a2cfPUdFluKgxluLu
S7lHugh6NEiIl9KdVVmbzJ5PPD0ftbtEv5ascH6PGDKtLXU6RyNtT5e2zVqwJGkY
TiGhaxhiaFe/9hqV3Qjf/rYglqMD3k4wzff6oIrkssQeH6wcfks47pvckj6QmAzI
SBMghTkB+r+aiUC0+JGXh4YkPQN/NmLpB2v9qx0s0ViS71tUC0MK0d11hzUc9lkh
gS1UE+TCaSr84C+kCiQ5PVmM3g38+ljaE0o/lCT1M9R2nHwY9xTrFPDm5SCqBDBB
zJDuewiGBDs4n2d7hk6MVNhcZXxyIP+il1kQqy8i01Ax9v6zxoHJQGIRK0ocgoGn
XdUNHdQVLHn1vXAnZzEROea7jZ93pV5wlJlvr6QWnClq2OB13ZOLr2HZ0sIDPzLY
kiLXHJS5hE5lg82SaBdx4JFanGPWMe7stlExqShZKPP93ybfM2KthORo+ImqgXHJ
bJl2iDIZi42Ng6p1ihRlk1C7bIInjfHb7fl8x6IUoUp6ul1uc2dvpVgeL4FcY4EJ
by1+JlP+NTexmKfuPC62RoMrtRmSoiGE8eNvDimEbXmOvP/hUJOEG2Gc9yFFn+tM
SxJ7gfZty3FL2B84dCb+OTyai9AdHn6uC5wWYNM9f9KrQuls4fd8IpkuMCOB9zcj
LCY8PZvN+pUXpHLM1xvw01ngfsyE+y877z30aRppNPDkdymo2L/WOLvZNZsMYhGz
GrtdPxUZDG3kgUM+Hxo0mtzd1x98fziEXqVmkvzW+7aStOyJMRg1X02aCfEu1W+i
Xghv42xtOr+37AK2Rjb1ZS8xeW9xhXjYTovIbB98LmER8HBxC35NJmTjY5FA4tpe
4s6x9K1HwGYrmioVywa7+8zcVEtn3Szz4EqIQL6OOLtOlULdqorM3FsITKYhkWl5
+xcYmBVP22mqWhzLj6UGh1/W7vunJcxtX5dMq+8DoO+NH3DDcQaB6Rk25z8JIYAP
x/cwAqMoqcTmK/hbQpx6gSNpBrg1M0kB3Fz+ihs9zX76U1Ly598ZsKdZ4wrbvRSM
U+43xvgOH8UDkGNLFwTsXMFoylqsQC8SdgnQI3f0XOtBKrHGCW/GrFlwmCJ2mi8f
6wnNBn9hJsReeIUUN7LfBs8mL1v+k9DsOJ9i/hE0hn1WeFBBnVQZTpq4JkzEzIEt
nYYLMPhi9PShBI9s78PAfboyvp2Elfw9J6rfdx/LXDoVqIDJLjBv+D2Au6g+O3ht
wTBX5Pg/QPyYXOBdQ/8GsylwFjIL4/cC+WAMZf5ZfTzLR2oTz1oByj5OeLwYHf1J
YPoutK4f2BnhXIGyCIX/odNr1SNZFjwNqVCctyqWP1qFnfgGrp3rbQLg1M3+Ab1i
OL2l36M02ApgGm2bTPQOQ6uaAA3yZQCBPw6wU3WxpfzPZml9qXS4fxsXzuv7+gAS
0XPxCJO8SOwBlO7A6p1ntFAl5E7aKuUTeZuJn4fnATU8mEbzUCK47+nSdyitL6Gm
8PDnLqGUZKJUWtggIy4Tb57ilm3CoSLhjWec5fY+bpshN6V7Pg5bVViMcRhMTS0d
+NDO4BhU9RC/DRCKVku2Zg484Xpuzj+Ro56TelpEpu69Egj7Qd1O4/sWkfhCgW+V
bpMkP5Sg4nRTMT2blOcQ4pn+CYV/u5hIytK0YnprgWPCddVpT4QcVxK6v60HMSew
iSAsZFLsYNkYSWareFBWaQpB+D2xdbPXTwVoi2p9WtB6N7DYWFKHA8H6C7Fj8Qr3
urifdZ0nYQ2MDYpUlwdb5nH/GRKqXYmwRAKO6YLuJ6+nJO1UAf2kfhyU20XP0ubn
BOh0z+sRTbqqR78FQPrYvc0L5sLZZ8Tspbto8PXmH/8ID7JDlGj7yRevt3a8R3fL
/w32rfiP/oQlIh6hn7YaBoo6H2vLxMBvQxL4Uqum++fDDurxCpUR65O/YOUizhq0
Lfsbj53sE7ZlHLv1FwGjDGUjPELMW3r2rxAegVCwQ7IUofPz2opVBdwuzsgxUl5k
M+XhIKY3zycNVF38xt+TrnLiJWTx1aiqcvg0Gow4hpBl5BsJmUz8HYIUEXsuQKtR
HDtJNejEwQd7S3pzA/jv75AF2KWPsvoiEoB0EuDsXKJR73Cb4LYs41gxA40+p2tT
8N+QPk0wdqF2fkDUBZxzappbHlgm4zBmAJQNRyt+DQ7LEABC2jo0nzdsj/g9Dz78
OfDyFpgZCMwuuQ88RAAJA6DPyL1Qxf9QIAnKSksEwYdwBwjzrsG1G5Ph046A05hv
Ap+sn3rct613wsWK4x1p1E6IJdo9QCOCDU0535pkZsrSWYdp+kz8srib6cAQjHaH
OmHYsemhdhakSXGkfiZrpRnbV7EPpg9h1WAhytbngYlaKdZ15JsFbyvKUUotYJnF
BywqQ547q9tRmUBFPKqAmHAJYuI1/2JrnDP4YEJwxbK9ce5Ygxuos9rc9EIZnPyd
QKaINIXMs66AOcUtumZf7xqkyPHgqCnzX3utjNxgztBywSTpesuTLbIBC9tJS2oA
xDdEQPAxNwLHFRObRWjqUkOu6FZZDJ5r9Ug2L4Pfb5ys1Ka8kW0oycNF3yuQLHRR
qaXJzRr0yP9LInT5gYmZJrM9eHGtqtpJnNoeCDZ+eODnALT2eHN5H6nqL3eCyAEP
7g6QSQ5SNhoNhTRECLD+F5ZM+IbRyjn12PywmV9K555vOSZjFy8gg/oHq0T+P8P9
cYCErmslsAByl+XsRLEOVDoUORl735HF0PRPt2hzFKXLmz7cRAz1cZF/Wq87dA92
+Wp2z/WArpRKz6OVCQI3jUeRzp1P8mkjpoQde9G0Sb2NWYdIDacI9TbguLcmnQ4s
qHkW83PE6L547xJgp6AjsI+qOYMSOh2SoiPH620l4bCNAFt/gGpD3rfDK3RGNEjb
wpBIKSGmwNRdTLucCkOwS1CcWSP4pKYlFt1A2KV4Q+2iGGBOi/6jybuqUGINeY+r
1/7tage5PtJkPa9hyFV0obn4+m4GuroqgfpHWR+ylDJsDw5FdxKsbA4kJ1VPqtCN
9a2Oqv12BFAFllR6nqF3qVNhCyJDT+O2JaCZYGA2imOk8SUS8thVCqELIntIgALc
cIoJerlibVXaKJ+C+eeypyTNRiROmVhkDw5Q/fKJUMmLIjkbFnAv0DmjS0r7vBOZ
KTaq8yVhlc4VV+huJ0eOo9w06/bwLi0VwD1EU+QOlMIOmAtAqIOAcCZJ1jPZilYN
e9BXJ7ORJkq3kQSnULPuqjYytObOzlxYbXjjmSFNjcOLiqAR7iwTRRggOwE9ArMJ
jxLSylrtX/VwcG7Qa4OW7IFYmremZgEDS1pu7tN24xo7MJluMWTsc3cRNh/W8BZy
HEFTjA60NmAeykf1K3VjCi1/eAEE2KvStbfe/zsm9N9bWxfWzQxeR8uLdNK53WpP
vORCuyI99u06Skus7Wc4Hzi9bjR+bJ1qRQ30jaqdw5iciRri6StV9diqyOr3o+Ok
5QORDl6cQhOivwHJRbk5L3mEPozJpiRPDo7lmTngcWjzgmgcm5WDOEC7xSGCl7Yo
JEPx0y9XfCzz/pv2Ka6g8WeHtX+hh4hGtT+29WF7U3fozy95Xm0JOAxOKybUGHUe
31YaGMHUbmYdYGkTQ+ao831V3wjVpOItpm2MQTStt6BSIdw1sLzzdXPQiurycVZB
/RKHkp8uLRRddjBAjQwjU83mseYQq9dZT0oMDlnjvCq6TLaMz7TTW07nB6CGT/+p
hMb1MGS7RdoMtAguLlZLCP/qA9EwjNma/8Z+a2jCgei/Qp6rq4ujzLqkqJQGSZqv
K1jyYSZxD7YjCZ65MRsrsFGv3py9z2JoCIV7joriCr6LD52oYNPVKsCMNKNA2DSJ
Ik2uqgydCEEAHGsyWFuJtPRv1KBQzRgVeUCbZemyPwThhMda/2zemxHRMtKBnnTO
E2YCfBYoD9aULh3E2if0OTFPPrQ5O1+tDJMSHOsTXq4rQxCza2YbCHAOjbfm+tfx
5b1ntfE2nC/2PIoamaOgZ1gsj0PR85SLcFWomNRD9ZIZEYcNuaCPFuD68O0HgM2M
DKeTgUdtowo33eEAJixq3V9QBaSwK/079/L08Df3Q+XAnod/nsNMIfBV5o8/Yrqa
D8FVwC5an7BBG8drqfRDbqX11oryrWQLx/jvdda+2fsfpaRtBYqgcceOlGqFid8s
qpO87OntM450wFB9h4v9YW8aDs+zAKOZ5tmhervXtEhLEXwh1jHt/FOZLlF6T452
5vfTHNeTTxWsKdsPmdP4dR1il4/5cbYM0v61MZgv8AEuxwUJK2kj6h2aTPv2mIV7
BVwWjcnY6ZbwcWGIPamirhkFOTrPDTmkIFj66TJSPIU8AnDlXu5eG2PJ+to0Zp7W
8ujPiYB8j1U16iDMMvb8LGfxsP8cWy/yZ7+6Y2+uJ2Y32C2CsmZsHtm3ziBeCCEO
9kDnZ/1Lm+oLFTAnVyBvbyIerF8pXGhRu64x1jMCjNaWFPfWIsGtru4j/9P0QB3z
1HtKOyBK8Id4pI1dsZcxh1Uv3JUaSNcnMRT5CLS01FuLBJDbr7DY07I1owGtm1K+
UeZkXDmGuxfo1U518nFiU++y4WowftnUdAIknMZ1nz/EPnINsZfU10niYl5hUx64
OlXZAkO/MQNjO2iqYqX60IWf6eq8tiV8Jpr/CP2mC/GsriLTG3h0iPd1YnO3pi1f
c0KywDTNFYfaOneiQazdJP5sTPiAIHYbe9mE9yDLllFdXEWTJbe6mBAIKYCUljZk
kJ5HsPgSsYywARqF5VqrNdKImcSK08m7QbVoK+hpTrV6JvdnoZF+tVnPL0C2H3G4
/tIxlVFDhTVOIKAbjHhmAXffY8U5sIx3nAY1taawKXBM8p+e4HXF2hqOhuQlIIU+
BDXYxgpxNW5J1r9Xvs8+NxhHPwhMsiyeiTd3wtBSTJKQrnhQ3ebNTQmsWjcF0V1+
b/Ez+84qyCe9qaVUf/6ky8G33RiwoRN+i4fX/Aqr12Clb8pHaBsuEThd0Ld6nzvc
F0/nd34YYZyo5qWb63oINaOgfEAzRaJjVRCVq+6Vr5pqzMLy7Vmk/PdGlDtygYsy
C8mCpxlMZLRcfAL7DR5nwv9WN64T3BupZs6RvM6gMEB4bhcTuIj223t4od2Zf0bj
ut2tT4ouv6gPopFptH++6tjq1E7AMtVQbmCx8ZxVZCEjfqUBn2QDMPrMDJEk4aWc
WfjqSIlXJxJEjTuoYagDxlSBN/d2M/IPk55Lis3chEk8kq+dlCmNX9AdS2rUl3j2
9aPF7ZDTBLDCkpmSCpPV2UP2JBteKX0Gg4Ss7D4MFZUgX+r4zAGfQeQxFRVoT475
Fm8tiveSW/rzOXMDrmNIKF0AQy2OSdTpRLH5SSsXHj3sx9SDBlTryQ+MmnOKNXjj
j8ua1R1MEUkvlD0/XC1kM2cnfIoksqwNA1Ur8zwygoPna0Jm48eL58KHQ4lGnZ4G
8vMGeAunY1it+aiul9j+uoal66Jr2fV/UfbQJ/cMx68h0xiigVbJ57hbVliYTQ/o
EWwVCX7Ae+d21CGUbFGG+vVZrWQG8iu29DVVGdyEw/xG1DyJzeFKWOmyeFcWIYTd
fqYSsdbU/G5RuU1sC73Bo/cpLUsALM+VTrD95kqCWE9aQduefwiE//nyXfj+GSFC
VCXPqKTUk8BPLH6u90dmCbfrR8kt/ygG8ZA20hmQZHx6d3ziDz3QQGnd8XycWxcJ
gKp0f4tipTiE8Fs2Xb2uVaIpcIVszTJszCAY2RIedOHRea07a/mhzvS0zGrF/I6c
3+0Ee1Wo0d8q7gA+9ozqr8p/6u6FoHSl6WG5fzm7mCCK/veiqzrawlxXRENh9G+q
783ipU2WJPoEDqGzCUAAGIWYtojWsvoIo/Lt+6ICO9yQRDrSPkZDZiNQKFgI4vFJ
E/+mEbpPse0htuD4D8DBU9YLuLdwel7oBzPaYAd32AdbE2w22p7okbpDhIRuW72N
DIikstz9WFkuOzcHjB0W1NZommG1mY9+r8JQVqJAbsGoAxVUlJO3pJMgS+auiEPw
AgulVlU19OKMvIboHK9FZrziCaFIZa+pjriIzEyRcgy1m5jgExwqYzEWjK8frylM
imzRUsptmNouBssDoo7YIvgY9dgczrsg5+10tXLb/w41tBg2PuMk7SEqgDqoFOXc
AH++Wy92bJd9wwok2i2sFOcH5zs2nhip47vQyPbi1dhPDCPIIPWTxkPZ2WYHkOaw
jyDhmCtcglkP4Espbn4DgKLge7qDHFyo07R5vvj4JNSXLg5z2LQNgTHNjbmguuoJ
nLz6DywY295Vn3F1oFZP3ISN9sKgGwjmr7VbstIGlRLVhtcYgrFeVr0YoBQ8qCad
VMM0Vq6rRUvLhRmSVuHuocIfoZc39i9UI+OAT4wjb69k6D85/FaHWqyaZ8mQdLBz
cqdMFOFeehNYni2nueJURswqbZYjBJzS4WfDCh39VXJryfHnNS9IjhQLwfOBqx7Y
/mLFhGVuRIW61KEdj5GbvfULSE3qwV3FBtMKaOCf/3xqbY4K3Fj5gJodq9QqFtu8
STxp0wvVAkTrTaQx+NHxKGn9xUa67bf918ppW2Ntq5qIZM6z77KtNDCNTMhY2BmH
0k8bzfY4gv7fxqJshazThUdAAo+O6630pcLCknmL6mbwz8d7xgiR9XFxwR61Yg42
1QPuee1sdVmmTPoiVzcQLoceoVIO2gk+XzmAxBMP4Swl3tvtakSfcQknLalq+58Y
HTBeB4JtMp8m44sSCh4EO4ubNiB/Xbpy4MpOkQxgW4YaYnBbKZuRHxs/Mg/jw55l
nelZD9657jHfSF9Gm80iMEi3RRR+Lf5gsu1MOKEYzGjh4AM6p92mtowLD+iwFLAV
30A+nF8nc7008a0H4cnwfQ5Nlw5HJn/fE+mBvGGJ4+HNg00ysVut8ph+3VTQeyu1
T4rgvL0mwNaczKYLlKIdFXkmT2MUbIIBEMLwqcCvmIsELeV3yQuiEr0oHKvpxFkz
v5K5z1XYKAEtYAbXWOZToav+CYNrblVFQjjAyvmrBzEFXs+LHpBDVqXd6ROPvmAT
dgnr/dd9WTSQAmh0YC9vXqesn9DKWWcEV3wEQi5qWudbsgzoNuSEFCuIwemseTY+
hObMGX1mrfmsb/OEQdXiZhxzBML5YVU6Q306wo/Rlc9uQA5Q4n0gvYtWUhaTsp4X
nFza1jk3As8xqg/UiZ3f1rHBFsbTOCH5drfsvelIr09rjvpazwy70nH6seQaU2/Q
rno2ko2vwm0mPXtGLmpgROVcmeqaERK/oKD1IigVsl8MpJjiLPrNI6wuw9HgUT30
0ou2UlKLjmaiyMIeffsDStAXDMFS9MqK+KmoajsKiUo6adPldLQRXe/OziPIc4QN
uNQlMVA8+yNUuTElMScx3L9VtjBgWO07il8WAbYJaRbC00SpSG5CpmgOE5XbN15d
O9k6C0Fc7RNgYUSsJFVnPEVOh/tTVtUrO5bUKw/rvboPre6aXW8Vc2K8XXd/vQrz
AgS/DeeRpiY9i/KNtr1bVQJZH0qN2gTb/jHUovbfZGzzUHbmPch1YmKXTTlVQTZc
2Ef1PU18iXCXnSwJnduBUI0O0hueab3/Iy7RSqMqdMeVzWk+F+xZsgNE8Dz2/nx0
Zoms6xsZCZK2uFIbRQC4BpyJoT3LJPMuqePQHiTP+RB5jfpE3Te/ZvfMuADPcunW
S3OE8y1XhWwimx0Eldx8XLnDCFHdufc/GxzlrV8vG2KN2+RBguBqQKNmMRjr884f
SqwTbYg0WXVkItVdoNZVLZfyebvl59r6iJMTQCB86q3VRyjjfoLQ3PoViTnKCstd
YtBL6UU9yScfSqJ+j5h35jYrbz0pvi5Q3D4czpX7qXNUQaggGB5d+JOROUFhuOZz
Yjq3josgPr0E3Pd00GTeo3urVN4w2iDLKDgrwXqJJGsLcKHog7fNg9jbvwygPFMI
rXabt/cFAntlwv2mRmXxiztkBBQM78aT+85UixDt2un0n+RgOvM2LLdaXKcNFN1/
98+HnEEMxcNwjJx3cVowbn+wAJE+AVo7XwXFuPn2REwuBkvzmSXuhgVEzaOxwV/u
asKVD7R3FV4NzGLEKUsoGzgqiA03jVPnqyhwDUIWzs3KDCq7z859SP5XSS5Q0qmY
APqitUDNJ0Kdq26xTdYg/k77P7mPc6dR2BP+PHQEI34mXz72SE7cKsaWjJoozKUr
7iwYRatx6IaOG+WWMU3lMpV62FFTKIEpdtt+T4Wn1W4dSAcEvfrMz1oxmNJ/36VK
4HJo31Pr3eipe4dxrG4lX9rQ46dtip+9iXCIgnSueJ/61Pn8A3FCZmOEE0JYncLa
1aJdSd1jByceVaAKSrR1N88QpQ5tD+ODl9sRAJMKaHcxkXY/d/AD0y6/+jOpSTCS
fx8Zw3FAKF2IMAsWPPDYMHv+8fYUd+STBdSV2stiFPcsaN+RmWIejt8qLu8xI1LE
DY2/fVOIAm5lHSXt2YZwM1OkkmzhkaNUvbksXWVtiSmSy1rmKinapCBBGZUUcxoK
NK5QFIl/M0FBKxF6YIuGDJRRJ7fo/vXRXY8cQUOtZeAFaJujM4XGyBcF4lAVCKJy
InFJSzCcpuCe8AAoieRnYgqeVrdPTiaMmhaBqet/HkJT2NfQZgyW+5ydyDP+hy6U
i2WJlUFgj5PLrE6dovw59l365yIaG5R4E0V+EuD2PeTnBupIghSBbfXcGxCVfgMj
qyKjkKSzcWrvS59SEHmbWyFPv5etneHyjgOxtFtn9D9sx10IhKHHqSSM1B5o+wZa
kK13IE+ELQ1NxRxxp7k5MFvtKxzzL6ZwFCr2npVfUNAtDBvQrOKEOfGjZphUo7dz
t+hk3A3ML0ZVtA+kyjGbhAiGXLKRfxQxdyMFxK9OMLguQxlTyJIiKe8Fwb3BI9ob
VbpGgvKb5/2dWJyvT8zDB/aGVhAITlbyxPo3Uuuzp25Hzh9WdW7j0eCy/sQoZrxM
ND/d9B3paZceod2hwhqtTveGH1Zvex/xMYzSrLkvSy6K+pvvEY8W1qcTl0dGpQAB
OilFCqatVd+VxJL5IZhppUrbnOe4jfsdOTidXQ5SDHEFcwqi5ZW5JMpkrwNvbXLL
/6j3vF83zZvnebQCti2axgLNe7Y8tmjstW04B+U42+2RnLgbXP0umIt0fk/BWlSB
921a8s/hGqh40yGwfOmPWh59a8mbWNqTL0zVfqgZPdTGE4X5WeR4ulD2YAzNko0i
gr3YuIVAazYDsuVTGj9tgYObcgJ8HySAz/65wBL1glSrKFTqYmpdA7IPiA82eVkb
536XHtPGjl+vRQDwu3boTg6lGDxoxNNAK1Vl23SynesegzhHuI3+k5DBaKJ52iR9
NSr4ZoTR1zibfIUac91sSdXfF3HDJ2m5hvJdwMnPIa6yN+89G2c04cit8zo/20dG
Z58x12PuflsDew5wii8M61CrXMHsf4tr5v8Lm5qjrDEWI0abFCn35PlCXJ0AeQPN
90qxqcCBBBNvSYWemaYHVaU/xXzbyAXQMuFFDfwp0gAIyLzj68STy9qc80i3k73w
2MKfBgP63Z6XQw9kH4O+o6EoNqkuIu7wFVdjYae9EQ6a2qRB6gMqOpY53sza7nV3
+n96qljVLpgu4idsbwVGxGtUs/66sntXw15rzWr/Dysjow+RivaQo0oLxtZDC/yZ
BvO09Ks24z4r79VD9HQq8s4Ng3QQ+Xp46RnsI1cuCCBusBMe8Ci37C9wcPhqblP9
zk04TQs6Mw93cWOFGbiThOKvRK7qsmP74JNa5d/3+9yRBvNf9aZPzbMwj77ydvc6
pgW1FiNsawdM502TkUIY0ubVC4yLEPHnYsKtIhCudg5e1YUVgmqDu1uDB7+wN5we
3U24eF1vq/d5X6d4E+OvoNHFvnaYA0OBTIbvNo+8QIHQdcv6KMvIlj3Il/wZLO6C
7u1t2EnYMAbqD05JU6BgcXXfBtnhFnKzZpv33H+lShZ70s55U+ZjD1JSbQqrQIRV
ykpSeV+sEFd6CRitwuC0LO4i2bbTYMnyANl9N3UANyx+MUc1TKYtvL2TEpw/LIWa
lc5q6/ZmsVTVwqtalcRMCU1eoqyWPdlsNDzxaQlzenLhEs63Zj4exsvmJRLOSw/T
deNgmmlwZW++JZLxId02W7Rx2JRdxNbBP51CAbfII4W142lgUP3BrVs+dmYNV20k
yY/6u/KAcS0jLwIHdXl/x9mWSF060FvgoypNqhCLM7lN/vX/cBrfVU9H1PatuA3+
ZQyz74G6FUrJy3AJkHpg+WTa4ZpSevqDvegqRG6GxQEfsIg7InPTtepjPrvpwQ84
CpgdbiRAlAAQGbciCex3s3Hrx37FxLm5vPGpmckDgSobQVjyfrIezeJmEx2yhJrV
Rtmid+feCTiuXuWsM7/Ti0Jb0m3cuj5ZgUmqL4dBUh2E2QJHNEA2pzr6Jl/NE1lR
W/JJ6IfjdKIVkRCZB8aApfXAkREdvbwHnEvwsoabBvk1pKvbFy70xCPrtr6E9VMo
sKx3F97nMNosamy9/LaxCpzeRZaCClcwPP2UqkGHVpgAfussy+kfvk9MZL2FH9jQ
NQVMtTD0hHEp0ewbh9RhpQLjcvZpR+qG16mdXVJAfxeYkGb7atQ8tODikF2Ra4F5
Emh1BIMp5EmL30hGAJWwgfILe9TSQUPdW4j/3djsQWyOPHeY1YKStMDKpjaBdzpu
U55BsbTgYBH1p3tVp36j65bSPegd8pRlcesWEsVBPaaC8nor78b/n5x3Qal6pAR7
ZPDzepARLPN49bwSIDPdFeJx1SFZy3MGI8Vyh3vzHqi1VXYGyCuIVeGLb55v0kkj
os+Ch3JArF/ZR989pdAv1gq3xrcZuIC3iL547bl8Va9MZ1j4LFyobj8Id6K/wl2b
Bx9moj4ry2bjzBeBP+52iUm5G2+Gf1ETnZhPxRt0U4VI2xa8VVfd89LmEshK1zI/
1voKBIZXzOjDW3hxmc4TIldrQedDyijHx9lAaVHCh9YueCdTxWWEFXSCQL+mNflo
sH8q2B99/+84Bq+jU1LioGf467flQPZb1tb4qkp9s4n8zr649lAcmfECu7lIJi+K
9O3Jl0iutkEaERJUoTne35GTLiesA39eu+nawTE51ebf7P5bY+UjWOgP6X86US4e
gMDOFaEHXbzx61OBNxKqbR3SuHAQfjXIdAZXkdtG2DUT5cac7g9jMFE6KUPWUpVb
vjv0QXQyV3TlSw8SvoIs/bk8CUgvVtizZi0O0PnNWxLKV7mmSBxRfp/2BTjTsNdE
Pys6XzERy4wMT4bPu+LKKP9EejhzBoc+NPdXHJF4CxUI1chyyLD+6PtzToIFmknh
AUPUywJGvbKqH2Fe1jTXlWZUWnvYRrRbDn1zpal8/z71SXIKMtsNhvHtsCWYkIwW
GkUrqSUuX+QThaTLFnginQGYad+BsAJ3UIv4wV8P2KV9LNF/vD3UNQsrJRwg7KTD
oTRepSRMTLDke0P+C74rAyFrKpoda40ttk2jkhqrNrZEFiUCFZNvnNU5sahfqwzW
PjtvpxBD8osUzTgIr0k8O+B5iRI+6FUgIck3ojP1nomqLtHqd9PW0MBolrJogZWV
aKsPtH2Pdb2aMgPG3T93m164M55GlSZxsm9aWHoJcwZzkh4xMkAosDg77QLd1bkw
x3nv1Xlx2Vh0nVQ77Khg4X8bmdrEauOjV/6gWG2FY8rfdIELYUukbHXlRpppLjNW
gqXxBMLRa0KJallukSF+ank9uqBwf9P4P+b4JNpOOYJ9mOF8dUjLyMwB1R7FgG/P
iBXsAZOVFMho+xoqfMb2NeegEnrr9U9leIraBo2X9kU9sRun0TOVmWDC0MIFbRHf
3U4vNJVax8EicwCtSwnk2k+LNTtsDO43bNnlMwF/58Km1cw/jjMTvXUaykikyYtE
nrxPq+QTlTlOZjluXm8a5DnjiQJGKyZuIYUSigwsQWLICcFgnRF96ejaL4lXxWH1
i3ip2pIymy80TnpTdSrJ211elMW+zMSIL5JxfsgfTn0HIFqowkDoCICEwdVZOT4I
13lGxsuBnVpzgiAyfhEQn1SEjCnjdTqN1a31oGl5RNLa6IBRMKTz1LwxbsHNHe/J
ow2Yv3ZUf7+HKRrqIOKLYV1GPOvqIRtFd/SX1q5HO3zuTJ/NQCwKhKgISkImVmfG
2NPdc2wj1K+yzwTUZPC7Y2F8dwcFkTiDUrgGmGfVYeX0g6uPzh0EzLfHQfAok9a3
BcRO6e+veu2bjGkC29V6hSNctgnpWCQ8CL17wwDmpq+ics+KqoT2F335hsAD+hEj
c10kuYZACvutOTU9ejvpF2OzGcw4vVyRUiA4VDPqlMemzWBRnrhuufwlDZSbA2jS
9W3rlJscQYnmH6hUgAfNBnNJDjgUpiYhSajociKUQmbh9EYmYs5nszq64JzopLse
eldlcOm2vSaMpqazgMstLLdhKnE0odu4/oH/QdN/Jm8KgrOcfW8rbXt2Tt+t7VWy
3cYFptsyhNeno8re7E9foNXz6uJCPCD/WUCf4w5NnDZ/T9lCKzIrm3EdhlFUpe/x
co/c5eoWruij4f3cgc4ZJAbiXYLu3TO4zVty4LRkQWd0efj4z7+9FTk9mR0h4YfH
AAKkRv38mX/JRb0N/UnjmDbhijzSpyWh2hoLXrb+xJhYoqg+/5mG6Pp4o0Obmt9K
kU9knL9kVTWRnKQ4dGAN7dObDgKMRei54eXFdVrKwWnvCAvt+s7qol625/a9D/zM
2K9A344bwVzdEg2AZNd2CnrdyEQI7nqn6N++m3TZV5nl1ii9onlq8b5fcL/1/zVQ
2OYtuL0Q7Br5n+ue2uzqZYaIo4g01E93y1Mit1eLfn7218dEjmEJPVksDvhFynyJ
eYa4Z1vW7UWNAg+bRpLb+zZdvVwfxSyKyQ83rmDGqfLVBBrVqvc+zfXvxs4j5XpO
4vTQFvSP9i/uuZ6397OK/B8SlH5B8KzXd8/EntKXa7JW+9KGsLNCeUDs5JUaL0SP
ePd8fEf2ARanX/uLfBVvbjFELrrD1XgrN3wgX4MLKhdVIXkhdaRYvfE2LGjO6bTf
/pw2JkZsD6lqV31lzTqyW4YhssWqu6+VSFmZoT3nqp3R7Xzj2Wi1g1lWITNSWEXi
BdcrsoePQU/7uIaa00cXJza+w5+WPuAyQo+qftL8YbKcwkpF4B/fx7KXku/VScsV
/9dIPD1l4QUgnXRrEeMhvFGnRER7Jd4gXbFJsPd9yjC6IIvy1fBbkOUIE12I8Rxa
UjsWyR+HH/T5v7QJGLRHHdFsSeQN4gvajuMIk7PEDvFoxmPUhyZJlxg08sa9NS6T
OqzmCqQS4Z2Tfwl8e7o9g3M51Mt6gnoe/i8Zpf6OXFDVCqIRpgAw19iiLRzzLVWn
JA4ZyNKEIGNUAHElJKDkvnHxI78evS3EJkh+aYOOiSWuvP8H1mU01oTCfeGYBwBR
20rxvUlmfuc+VcPNWdijSJakfCi9W6tzX3dKvWXwUOpwe9zRz4fEBJkAcAnrYRn8
RTnw0VtYFvN/TtfVxnAng+gnGyd9Gr0DZDShxLqZ8/6dlFUMSoRwh9E/ajkAlhsy
RoRwam6pKDWK0fRFDoKHo/Ce2ATVm/T8au6HRQBKCpExj0fxMElHYxoz4V2vg/Fh
1fsUKhcGH1FpZZrJ+LMVXKcyuKIyhyAmoxB+blF3TZzOgqulNT82VjKOI79n9CO8
vae+EamXQAHg/MFT+lMLC9SyImeGYSAfmS0/suwsQt+XoDAdUBqM5+wQoA+nAqkz
Xurpmk90c2UZcckNOob4qeZ24DPiFSqBCzExDAVt1MTU2W7G56hT8ReDqgvkYJSA
GyqcPHPo7gRZXZ9ThfEqkVWxGHE451PwC7/uf08faULSncl1pHMPKd8RlL3uoYUP
i8BfocHcPLlnA/HNpiTJzLUGqdu37dGsE2ZaPO/eXuyUpu6j0jqHdhv86deuxoxE
p2aKT1H+mTrZBxmxJlFrUxzSMQj9viZ/xf4IUdgTcMtZa04CAy6NR1rAteC2Hz9R
Jmf9oQRVStmg05+onrvqA7831FPDWqf9n3Xto/aQTe7Y3FBuX9y/NQb51gnD22N/
X5pdLX7jYQGi5iEHMfX3vsuk6F8jXzYRbZ5Sbc1hwGsLUj5+aaP6JTWjh76V0lSz
+uO++qvbqF/5SmjWJetlqzde4YZr5SQGhO4UZouM2CxuWsYZGmM8PuS4Nk9KpEUQ
KvHrvn4imAOG4uuuRwI2W8B187dljAvVWP2bj2qBDupmwJwABlDE4jaTIBaAOem0
BhkeZyCHXet4BvN1XsUaybNvVI5wCPmRbUsuDO0iWbcy+/0RRrRlWU3+HCCQzD1B
zl0VeoU2dxL4jmi76vS4ihNXLhakU2790ELv3NwDFHBtxflooc8hw4Qyj5WETfxB
hc2TM/H3Qc4R3yms6fASx2Hq+Eqq6NOE9bVcvM/Uqirhax8DjPi+fLkLqN6p7nmF
4VwPhTdvHPJmttCz0EmMi9bc7xENaFhOIjgvYnGcNQNZDVtIOqF3P6bQ/4jROkj4
HWOUamZ3159C7wBGEnX285otn1qyqfcGA2i89Nq8Jyr8bKeEXojTr/zupGxs20Xs
iCgmAQE6HoVENhK7ybaGC3u41Sge6QzDnTb3CbcMKSqcqRqNBRvpfNAXxcR+BORk
mh0kdKQo8zA8etz47bmo5DDS9YGVS1lQik6frUH/NB9pc0jasAERAR+6v2jLuh+x
8EUx7w07v3YdBwYC57LmnbhHUNB/IdXrJs1MIltgecZjd0ns5W/rO6zDEZ+KwRtN
vZfv52tLwiMfUnFGvTMiXpcMCpju2VkD3oE1r8cSb2loRLGBi55ChP5bV/uY7MeR
lc+UU4ULx5wM0BlOTjd0DYla0luiAuIJtNm/lS3zlnrACP5xpX6amaifQM66uBAd
tH02UlcaYXEwNsR3FazIsizC/0U//qptYX1QuAKJvZbZpLZTQKjZIX/upz1JdTAG
feGj3gDDU5PihMJJDHigXS0tUaRBB3p+44g9v5y6AEYcEXqMLW4oNpqSRTS3kYL0
RD43cr5cP+W5bkR2k5sZGkvAYHDeueekEW9UVH/f93NVew42RZz3tGw89TacfCMm
KNP/rriU3AV6SvU3ODiLxlNHYwicpEsB5sirzjbZMDOtwe9zkJNUA5ezb/ECMC+g
laO47A3Bi1cFwsT3p/9OzQ8BuTyBtAtztZpaipouT3HSs6duDP2AtfonRZkzPEDj
4W72JLIE3myWzjB0FI+3FwrX7ABRuM7HpzPBmCl3Ll94OV3dQ3cYFOh9aT8sa4mP
QeYDT9PaBGZFJFWzgV7qEKgP9wy2B1Fy/01UyzOz5MiYnv+2Ho46UygyM8kLKotS
5PAi9KPebBIvFiQQ/x4DiN5LSrdWTOaKiKkPeIj5JekrqKOPQl5wHwJclxqGGn5u
AMj+AIaA34RlDRyJIHjGuUl/2qguzkIiZGx+7TykD1OmqNzCA0pEgapcRMDBN4An
WRIRBG+4m0YSEq9oPD6Vt2RVkLFRcGQy/UePNyQL6nllg/pPqCGfWrOE9reNPql/
WU3MRHvm2VzM86hxbZU+dVKgmRljKOAjLevZC8+eEPym53+O8kCgg33czoHukd3O
YxDWHtc2YfwiaiQY+ApR4w3iRLnMGcSG9Cqvcl6XVULY1O5t5PYfcVUzBClw2mud
u1iS1csR6D2s30ObEOPf8Jkqfuaga4LONo4RngJRMRbM7hFqXIC1/IJwD9bJLlHs
misY/Uyexw/zZGDphkVmxLs8EVYU6rQK3XQdCJCS8uzRX2W3v4qoD6KEBqwqch3T
EB2KJsRwESLubIGywwZQXDSyGal4xXXHoJ8KPmMzBpbBPNdfBNPGVHxN5KJRU8q+
/CjaNm8g/GiVD90TZD+X7ql82R+WJRBcpFC0Kk40EPnxHdosFU8oXSAELFFF1nFr
iJEEQsjhQI+7AN6AKmTnIOwHN+pZN7e3CwBSAsMiyZWqPEM1Wot3YbQcIu5lINvk
KVkR/U3hAUIx8lsEicMs8pc32GsOB/kprrAxxuCgf+lwBURMaBLFP2jMDg99ctDa
/PodZT1EslggT+joYgpTpeWoSfsvt5hHMa9fBAo70sfokKfJnAJzy9JLeheFTJ12
9EHilP4M8JJxKhLXdORjl90Nq9yR38RcdCoknLXgtBxVisN+T6YW5Q8DQx5lwkSd
QxEhRSLmySMrlqBvHCDGUI0uFiBpkpcE+jATRGYY93g7G/Fb/HL9gi7P1DBq88ra
KG1XPoPwhyFqBBEY8MDKAHmbkAtlqrh3jHV3GexGGcdyoVCSFY8PCtNk3o2JMYq0
/Gzhxsnrk1uFfmVb+2oO7jcAxW88dI7GexCDzG2jXg0NWTRBxwc9BBeqy09aBqCE
cI6rFsLxRY6l8E55H5nWxcg9uTHjPzzv1iA0RvnGejrxVEYs2FrUrm7n3iRKSwgt
GvBKFVYze5d4AxNr/rsjw3b+0s36KIoAPKSbSQyXapJrFcbICCuZCLgOGitid67W
QD8FydWnsYFxT9gPyU7vudDo0TNXHlbh2ZaKZ7mXygQcyie6fY9H3taT5lXtMi9u
m2qujMbIjjQv9DFHsu4F4Xd4fCL6QffeiAUkE+J7d25kHTJW3ohfHQRPieEREP7f
QD7+gG4Z0OVWG3C37KllZtrL81iVE9M5lp3sXSxmeA+WwZC6TXa2GstFte2sCEiU
EjD9KDaB+yJpPHEGZGH65Qd3IIr9sgDlliXMfNwnpnfqBGjKdaY9TmdRi0HlGILR
ed6uzNH0F3XeRLnuKtkpHc1DDyDiGGiT46TOCjydHJvqzPybSs9fopvTkJgR6XZy
kBTdXqRSqdYJbvbKdI5babEuQ6+Z9SRkaKeg2JL0xUMdGGuCDjvrmvXuc1wV9y/t
99AiUqdN8GNqvn0eg7qXJww+rLSteCZR6wkdwjbd0x0FmCkiAWzvXmJ0thdvwhEY
cxNXQAKT6jmx2B3VfkgEWmzoPoEnMUALwFRsHYOEDca4Eea5m+KJt/kbSORdOgUl
2L2eRlDkuPvAooYrU2CY2PmmSUi3MKXtzWSwqfIxAm9G/ZfAxnf32w+qGyD75WHw
eel1heXLLSomHkDviPUkC5rGRoY5Uhmt60TUMoY39MR0mRWkJC9MT6C7L/iw4K9p
UAvZjEUmu9RaixjQ/hEWJslgRNZqycWtj80SGWIhKGMcQohMrGdIjE2iZ+oPohkq
3vrjZmQMcnPwyc33zWPsX0+jrGkwTtuKFWAnQE2crNZK0uXG3WD00IHEyUMNWk6i
o/l+zYjLU5PCD5KDGfYaDMYZU9SFRrGALFE3bVkgSt2ggQT9jSY3T1su1cuuwWo0
lg4zuVpa2uJYLMlGuAM7pouYQxTXWM3O8VLDmn6mcJUVbsQhD+NBlFtzDpksh5OO
t6r9KTW61Nx08GBpMsEv5QMa0aZXhtEz1xEjzgx3FfV0SZL5epcKQDLrDAGSTPC8
mcbmnM+I7kfZM6s7RYvCCqPSiCJ4eTcsPD/93VRfetVSmrepEwJvJU+3q+MTK/TC
pGXdf8jdxSuS9whuM0N0M8o0dgJEpA8GnalQSkgASm/TmdSaXMmX+ZCIgvxxR4HM
aeYO5mXMQY3HP+rY4NGK9He5bmE3gm0f3P+gdYKf7kJkHHdbXV9ujPKPLknDYLkp
V8oPs62awA795w9HkN1+G/SSbjJcAFGaNIqbp6ABM2nbxvW9TGpmbzI7A3TyViUP
Dq1h/AIqA7PxiK1iZqY27cZRVluj7dugyPDRlXBMq3m3Cb1q2Xk1pPOcpqsxeMo+
wNLvCmlNLezp39pN3RUaDQdKv5jPa+LJTqo+LCsChIqmq68P6QkSWkjoGiGgL9h4
KboSIo8Q7wP62raMoYTAdL8MwAix0/CZQ1ROJqWApsDTdH5VYDMaRPDUVI8OgJGE
YrvdhIhOytj5Yut80vCvOpPI3RdNe/hJTPzFpR1Af90GvoZFhnm8VBPQfYApzJpx
ia3Yi3uD3oJacnlwFEjjvloeCGRJYQFsI69aTiCKu5YsmT0hJgmxnqWVIzwB0bRw
geMgjyWTF4sSCyIHMDJYzyIgP+WI5u57SZ5Qba1AI0lw59b2yyfrvaxybiwwyXz8
hc9whiEA+VmNVbIODMqvI9TfVYeSQG0XwYRiNGlNjyumpjpUV+cIVYfLieDNXqge
GcM8FKN6Js3aJYSY1O2CdJIxGci/wvqg9S4ABxfWtLVxDob3y6Epm8TVWsVnVtHT
7e2xf3DTSasLrtjVe9ogadzl09SukhAJjlFCsJVgYwhzCgw9xuqmw9UbgU77X6vd
nVRY/ggnQNQStg7Zlyr+cyPxkzs8bk+gt3w0SmQmTG3MPmiHx17shdDH2RbxMRWI
9ToKpeLEj603V7YIHVdVhQ2hAzr2MRQHl+ygsTndEdeoJ3M33KsF1RTSgFEdqKfq
D4hDdwrxhCQ++fEtlHNd6vyvNMKbgqxrKhhKy1DiyMSFVPIC3M/9Q8DrweIjYzP3
ciu+Q1YPiL3xE5WsLGBpbVQpDORzCSkPNNLhDplCpIr9ulrZLFKwO8UFiBlUJmgo
afX2gAkuxsAJ4Y9pSXLJZC+LS/U29uNQPS/VqLxiqOrdYjg+EMJ8DPsAiH0kvKrZ
Zr6009ct2ddKUqj1WQcLX9S8aLnNwP5bJI9H1pI1ChRSaCtlsKLsBD1CKZ5tewmB
GS+chZ8cmEd6AAcpvcQD3Lv8gmlVdElYey4wDS1QNKimmeDOegKLR58q9DGp116u
j1lAear6yv/ncllz4zjHLW/v7EUmaUhUqPwQ9EuOUekDptClGvvnGOBIlOEP9GbU
sHEQ2soJBRrawf48nlUqdZsTpRB7vDv3Cxyt9ifiBVSh8/TgacdE0tCQHCWQtrpv
Ml4KId1HvZOxd6MKrYbeL9MF0kieoGpIfZYqhlbNDl7QkehNTePT/4RPQic9NaCg
A6IKXD82OkA0GNa5Uk7YHyPnBWfR5eZGi5ckryVrWFp8YWlMKPE6XqyJWsvu2U3k
3Nbu5tPcHJjWPIEXgvhqMaoqw7HDQgNcHbZHI7tVAdIHAP5i4pQ4U6584QMkpc30
DWvUsIqfpufnx+qYmmJZs2l0A3/rGfeyiXy8qUnFomgNM1iCyPa2KZWGQoI1gIOC
VIhc5tXRYgwt5JgufxX0xRrjOl4rgzWNU5XXtCaAotLuU812ITVkbNFYy7U+b1+x
Q6pDg/d30O14X6jW21a7CW3AfEuUeAZVj85sz2cwQLBoGOV2JbGeVyaDkJG/l8Rz
AKY8MUEBM8mpUSL33YMlcaIkVt5mgPkCRAc+RxITuPevuTtj5Wqn8NZttc2rVkCc
W56Kk7Nv9eC2rEyGCaFmlBs0HTQmx7qZl4XTdPTimHBqYy94aitYjVr0k2dEHB32
A0qQ4I7le0JBBEpzBVj0/2FrhRf3hbonD/3CqP05UX3mN/5e4yohLyJwmFhXRr7j
cWtHB4aRQP4aARStWXlnJKzZOzp+1gr7aNv7NvuOl4g6Axc3FPbr99SVrfJf/3Fx
mAEOfAT0a1DJNNg/iobVZW0P2mS/mrjM2lG9lnHp5NCqtui+iCEIzSTnf7/9oflg
zA9CZo773jUPFLhkQ39rGcT1PSDTJ3A8SsTXesroV2GM5J4+TjCDYyH5pPsqjY2Z
fWidRlOQD1iDUlC5lIUNAbp74K/RWPRoqsuAsRYNhyxKnW8h6qZh2+S/tGeYQ1qu
vhE79GQZ9lOscMSLgH6HOobhc2e7fVMeSR5gegeM0ykBja++YwH5T2TbEIDQc6fb
3uHWe6kouRrTX5C0TxB/WJFc6W+ScWApONmdE5X9HvplhGgyLfTJHh0xdbdu19wH
SOb+PurYi08yDEJMfpZqHyo9eHBznM+RxdiP3TmvEefhMfvrEO73h5j9JGwuVNLC
ao9Jk7WtKkSfrstLLtVZcOhEPpc2I96citHzZJDDQMLJHOl/xOryngiCFX1e/+PM
1Ig2OjFVExuvNIEtLgEt1i+sTpl/ILbwmDSVV3VQsGoPzb6r2VpsAxAxKNjo/dY8
x/qEhIVtDKwhAmlP56uZVESDdnrz5Gtf3MPRWK9h0tzXx7vaRrnGJYvPS90mKS2g
fxvduIpVB/mravNFwkbozj6e4+31a+a5oDaiArWsXbImvwR2nuov8Aj6CaPuMLyF
Zg7Ln7StR2dsVH36zVgwUAnHlB4BZybYWhNDsFZdyBmRSkiqdW+s9E4ZGVx139kA
oDQA0ScgWxnfvPbXzLMAcjiLGwhBio+MsyjiSvs0CgleFD/RJpzpZEmVNg0tzIFv
tFrra1bqICqyfiALHvd9D66FbuzGQh8RPFBUz/I58x7ap9dd3HCh41tAL2XaLRar
li0raock4EUMggaeYf8xWouSJlBlEdYlPggmvzMUuYInpTQ9nSGyfBnWs44RZet4
Jp1bzO4OdtU25XJhnfktLP1N74KN6ATqFDsOjE23/UOBZNggFR1Bqy26gGYaQY2l
fux5DL9O0CLaZCuD03Do8D4THuKAvrf12Sp3xARVx59G3fZ83J4gPofiPW9Z4oeq
DTfdf/Azt4zohXeMWOSoc4hbro7tLAHi/TJASFrHcJZiAuQcwaHGBo40gv4ptUNI
x9FlN6V6p3swzETIC9nOgPP3Xy360l6k7WrNnZK3EDzaSIokDNSmmnEnJvHuipSi
uYmpMjF5ww136aZZUizPWHuGFXiSoSDL0SDV7408nFM8tronLAZ4h50FAlfHGxnQ
VxamxpvN1hnsiaw6mxWUG2ui4gfOpt5Cxl6mSCO3iCG7xr2k9ngWUicrdlSvNEmN
ogi5zLuz2oIgZy4Ocu2QEN1BwgpIJ7QVwo3yiXjBc1Oyr+KVomvBxsRVEC6Cw53g
6kyaMy2M/euBBUFcuabG1eYt7ENhAaaPNw2rZLQwkfXObmKBREY1NOZTSHE3ipD9
utmns/ZAjzwBDdREAfwWovAdvxYPdPR2s6WUmDOEgowszsXOG1hzHpCv0NlFZ+IG
mUCjvKBnFI/Cq83xilGAy6pnLSFDxOwPE6b/gaCQ/g3580ge6ssqMNPor1Is6MMt
IUSxpBGkwq7FY+gKVktN16VDUDyamw1FfJDEinE/wOuZPokdcPBIlx5A/wC3flBj
q+RJ33tWvaSTGXEXW2JN1Jy/KyH4YauoNny5HYDWsFXiolQCq2ALt2Csah08gXam
WIh/rml3yBtj0vN7nBQxIgj/d2fzMfjxKZjJc/eEiswCW/kaIQ1NUPTyCBwkLuG1
KHUG8WwuC+/zfJMLQiXiV/MZmkX3UAi2Mo146TDu5Uhb0EGMXjuedkSGES3TuJ4o
Lr7mfLWW85njxHqJ0Sv1uyB8ptPP9raZG8yxbk0YudSgJjz2C7f75M1n8xLqnZZW
LZvbZS0T8Tw6E+ESThMhpE6oUF8A9QXs/VlYA8DaBR5VP48v4lz1zHmwsYj4IV/W
EvOeTcXTBb/pnvcgs9Bivx4d7nZuxBM9DKomJcNKLtHavP58zQzJkzyQJjX9540F
UwFq/YpNoCL5izfV5zFdJBSmucbczfnnLnvs4rPpq2g+15e/DnLk+DGLo55+W8b2
YVaz4XIGVkjuXYyvfQXVpmt+IVkjj5TgTnKMOB7Xj6eyr16s7/H4GK31Uwx1v2Y7
1/z5an0Vqi8OgbuIWNnZqA5oVymniui3vRblkxBvrBX224j5K8XJk+Aemq4OEKU0
sri6QGoRgbc9KZcfyrhWMlk0PG1pWZIJPr85FyWIhMrbuUPqlU5dLqEym5gg0Oo0
7Y8pCX7Op9GSCFIjnm3zF2ikB8hiyxFA1Haw88uOMI1TXEThqxRyj/67GNppTYGx
4Zcw5rpRHN3CSr2qW9Yn6X4AE1sv0RcXCzvScwhWKSBJ2yUkgmIim4fNmJf0xYGe
FHfcjuM3JByKMmGNeVQG9nvR2+3KXBkNXx7IEq4GvJ1Dwx8OAtMPPQyP7UAwijWm
xPvB27VTRxQyW8lhXqpXD5bzTTgsrUOEb950QpLYDhjgLnLFFKBL36LfcI2y/LtS
Si/SJ1seKzFtiVhAxmCGBEsi4m1MbdXwBD5dcSHeRikzaq7P5Lf+00RxZqt5nWXp
L86p0OqA7nWvXoRduOBXSCfxkB9JIIfDHUtKXRPioGCgkA9I1g9eUjK6x7Fst7h9
9HQbZuFdH7mfEIRuaTIO5dvZTdfISXab8S9Q9lMvRO5hbK36zFkEGeEQcGa+BcGQ
2FOl0TMRmRZRiG5vNEYT5pnHxgZyuiBuTIm3UjJ0sq0uesSuOGIjcUOA/TuC2kLD
YeIeqHpgKf1M4jl2lMvKGSTFIJ4j2JIF6ySIqSZcPcty1Xy1xTAFRk4IDm7r46/u
PE+1xsiZeIH5KqPY8IgendJiEJ5E+ebnIGBuX2pXJ/LllDoV4Wt6e3iHdWakpGPX
SdMCwlL136PBg5iHWCRj/thucdgPEu/BYQ/w6rliG7s0NXrlInNuCodIY8a9PV3H
AzSvH6/OS/WLgu7uvZV5lyTWFR1HNZ6YIFctHfpLXqE040PBNSoVPtcKMNar3GtN
US6+HhN16xu1Zaczt/N1eh16MTiratYLyZbyApthYgsNxS3HF6etpvuO809/putm
8zi2NH4gErSQ0rpqOkM3JS78dUqO/bDJ6XDByVofubv/wM9On9CW4GY6Cg+EAXBP
vGtubUDNxNzYso9fKEWlr3olYANVIEw3TZzPsh22hZPhXNmKsd3odX2Qsx7H+xVH
V+GpJ/IkJlStv2W6XqqXhdJKn1Bwqek974lrUVy/wDxNeiUs563uAZZ4dm1ZR5yL
UD8irbuWHs3vAECJ+5Bs4LWkhV2NCpNVsZtrbPHt/IepYZ8RJxgHm8lFv4cLDwUp
N7HwXnpUbRhbtqdIB88eLo3u3mRRGGu/md6W5lBZTXrIbFUSwoxxvAOBXLlbK95d
wqrPu4LG7HIvl5WBcrdfR9Wgt7NVN+jVkCZuI6OZUhVa4xeX8gUjloQUeerJnpE5
dJLoS0NrOa0K8Nqx/rajmZV371FZe+WaavpAEIyD5i+kNnE/dGk1AVwYjQ1quL+5
LBY7cSORfu927bpSiA40ufxlegixw76fdVsxLX4fbAjpp2sLUoXIaoXhDspSy9DX
w8+AtFJmyjjXx9z17t889+52MBvkoBP2CbyHQzVrHgGQP58zvFMijpZlmX0nYpYD
7+n3uNOrRiPgJVNpWbOPxxZQMgHexe759JtsGnRPuq2/NfJhFckN6+xYN+nwc4My
t2dFX/uxq23hiMKAnu1eHTMn+bUPhHw1O1nDSRCA1ZSfUx/m0Z4jxWB1rVlrQsE9
3m6+35hwStaElIhOpx15V5dSOiVQ5JD1qhp6nK/q5cRtDEb3rE1F5hktX1m75ZPm
HTAtvhzRzxxOtyFOQdNx8yxfNBILZt6cNnm/t2BWGbi3yyL83kjWZjU70mweebEe
X+6Jf21SrCENduAtx0mN3H2G3hzZVfpz5Ol4bjF59Ph9udSn3l+a+hN13lzkrU6j
rclV3fvIIC09wRl+EvAsYZA+QcB3mS++QcRz3bk0b7ZCcenGIYLDTcnBLmfqriFZ
+nYaRQlCsPuSOXSfKm3JYEaZHjvv4QBSjw+rXZE5SdELpuGTKq2EZ4mUkJaN5QjI
jaZ6R6rkJE9MJSwh1UfWn20dDJw3nrkeEkCThzUWtSf3lb6p8nr5WNOl4vgnsB/U
LPqoxpgZEblXPF9zDEtPtR/49yzA7qh7zRTHDZRT6/LyYqgSdfJbpUeJptxhm0TV
71tS4Y1xbFCqI6ApLRvUy1c62X1LyW+Y5UzITPywL5qGJOftwniWHzhIogR/nDBn
PyOSf/o69Ye/Z+iErQQ0Cs/dsv2qFnQDfaXYhzGRK9yvtsdrxitSK0cCNh2ja8dX
f/47Qun8CgyWJQua09Drs210QeMxJcVQXB3uPl6MdIdQKDrBlhMmEAl3w+5X3b7u
n9u7sNNZlP6fm68beKYlAAmYlBuLqpap8rCC8Ebm6yRJdT++FPDw9xKTh/wCFLST
il1Ufe8AJJ252eQ1G0WlN2wE0e6ja8EmSAxsaeAGr87OZY6u3BppipNgjrkn5wRZ
rlmqokuwPzeUZfnpME/ZnN0G9iIpP3ac2+ysCnAGb5Hw5DKRLoaqq8VnkZ25JX62
HfqGWgDahrKkJS2pSSQZmKVrK7i+9Ur/WZHARDH5qgQLbRcHvXauHV1syJk/8JRS
s71Zw3BVvne6gD/IvnKOWzy7olWkrJW2zVIyDyMJwAJgh6f2lu0OK7tBSstQvzyQ
aBrSyV85EPoPdUg0DgwYYKzBgLIe8eQQXNJ4Q3/lD9/szXSXLMJtAS3NGwD5sc2W
jhR4Vv0ECACc6wCzg92ZJb5Ea+VwX4/TmLx52isYezD4i8xwDFSUE/phOraacGRw
8zk3k1kKiGphzLQmU6ie3RSCnIY2s2itUNSMU/IDOIy2h0AxOMxShqBXnfQ16eJ6
4KnrChU2eYXkHoRpYrm4HUucZ+voNp8zy+m/8brRsCECv1sNV+joHo7n9a5mj6KU
c9VBePbHVKWLjEnkwIMLy+higcKTmVLx/uAO2E0nHvp3lem8thCRRy+PlF95S+0U
36HOERLyBX3XOmGcMm9megPytMfb5hU2CKM+3PjD2sDO2RtgMt0Uf7/hi2kSo+0W
wr9/nU9FRuFIW+qlmbQjI61yik0fpWNW5JzBEFqjx6EIHSmfqdKlNC2isYqYSvvR
gz69t+uAFpsF+YTJqZOgEYdUugBwScMIUJg5J4HmVSiAJvlgN07j3JM0ZZ39e4Re
AvFOMniLZStRnuOJVL+BAQw02U5929VcQLJy8jReHYh2+X5Gmji6bP7+Amkwy8uW
EzoetAW19ZrTHD1joxo7Z0t/ZC95T5HKFoU4N+B1uVHyOXxu49Jibwp8bMNq2G36
wCZ+P4+oxLzbMuJ1PqVVe5SR035fg9tPNFtKuAX9K+jT87LE9dZ40Egm0r8VN6jc
Tk+H+v+oFlvY2lsWOyhGUksYowHFROM6BIFH0CwfA70JlVG37yl5kiFoeMpHeBRA
4jFr4cK6ePxsPyI0TY4IyAbUdo8oj3m+1WO+djn2yECbKBwMdS+dij9zXMgo8sO4
mhvZJcSqgMEmg6y5A58lnSNkss0n6iMLjI3GWqOlgU5MJP1j1+nxYPZuXceSX666
Gbac9mAr2aWldOcR5CkcKP79OJn1s5GZhX/qvrLvhntYMYGIvJik+3L7gkjIKnbI
nbuls6nBED0V4GeuVzJRmA2DJA5XbG77B58d41INObN3oKwqw/7SIma0QKITfnGA
Hghbv3yG2T/sJX4jaInOhxOEovSTpUbjj0pjhoBhUQmaMeLTyq2v0brAWqFf3Wb2
BdmAKGrK6jMgVRazPo3Yk3IOPVeEcAoBPNOd9ILZB0lHQq0h+WVYrq38QPXtGpD9
LgE9ZQW7oKJG3ic9dOa4+iYy6UsD+ZeAZCiqNdR9XOJvEtzKrojXzScyniU2TeSp
tUkEfmvjB76c9zPX3q8wWYN54nVp/Z1SsawYz1a9BbgmdRjNQJBoNKiZhhRUnySr
5DGDaggkMO8kh3c29UWpi31D10N+FEC07Rr+LUTPPoYSFN5iVfpSp8sRwxfqHnX/
7KS1VKZKrTs4bfTNuNffaotX6VOSL2URqRLzVtSGQAY2ETTmQlBT456vQzCXNv/l
c0TpkkSlVy91C42dsDVWsRYfPZXK+tTnR4EClpcIQ6u4p8RTsDb9J3z8nKVp2y8O
UVQ62WKaYHJvoLU+1YM2Zxd0rJFAc+baESAskF7nMHW/GpcV5ZW6f1LQp/1/nRvA
Jc6+2GPxp/nNYxovpItNoMVGEKZ4Zmj1u/3gSJM4FYadlj/nWJ4viCy3fgfwPN5z
NajqY2NM3l7euXwx6m8aHfWnpR4eFDCqGFcQlwxWjByI+Ohgm3IJSKDzM+Qk0gIM
dB9v2zw0nX/JA5hopEj9nrk4vUgyZLpozOeCPpbA1LwnxgKHXmBR5Q6QTWi4HpDc
EODRl8adPRjledmgtx6sVCZVVbk3v9oc/dNXIek08fDuYNxB03P1rmspmoz4iEu+
UhF45xP1Qv/W3wOGRiD/9KjqYVnG59StNzJcAVO6jAmlwEsH0QmruUL3cLqaiwJO
i/p8ND2nPkfcQl9afIECKUmONFZuuCbt05J2cf3rjZjF8qOGWde+O1JQ/LfY4u3e
gzPT/cVzF+6dYf9fvz/8tKLXzj0/3xPmQOWiquiEIpp7VzBxqieLzpKfJxJcVpNY
vUKNadpDbESYq6i7a0gOJA8HkcOxn6xDmQUE/BzSMVgpimwNwPGm4x+b6dvv+L/3
+RcyQj8gTFd22P+i59h1AKFP2YKeapJmHtu0MkLCopRbvBhotwH51V384q3zNkfJ
Xa1oUBcM1sqUrex1OAdwwubqwUboBHXyi/CX5APpEvVs/ghF3zDKUi6eSZtPyTkR
h1QXolq5AMQngPP+9k53r8skYvyWgmR7Q/37Y84OTxh+9Dmir2eNfxi6YH/71ZlW
BSzCkADWJkD/rEcwyeb+d0trU3Ngu2hAnZcOA4+5CUb8Pg/09MkOAH43o1BJ5ywz
wdzUJfBk/K/M5oJX6xGW3k2uslJPExP7gXYdQ37xlt7dY8mVojkzJwMdiGhrtZ/D
9QnlyJXdPx5FLTMKH5h3GzXzyozHPE5Fo1l5xQcqixrXOqQ5mzIFzdisKLhuXASU
T/BpYCMTigA3TDbRO/Kb+nbNtME5WVp9R2paDOwsJ8vfj+dMpXnLKlrxoNaocc/b
8YFjMN4yocymSEgYum6AL0RQ81uZyKL6if9Zb9JXcjm4TAfUbmX23G5txcNpmdlh
MwzaFawrquWhTGln54GVX66aF4EM3hX77BuvKYiAZR51rHKuacL6CSQA4qwINti+
ZajRbQJTa/71emifQ31HYzL9S9NE5XAE3/QzHg4x3lcXfJHN1B8PVB8QI4YN8tSe
Yz7BjirsIhOUaQl2J8goo/slhVK1x5dKLTWCM9rWM2DJfeEcuHxnB/ip6+j2ZYqP
/Biwxfl4mcEMwm+v/LDHkGiWurVJmAgl34PYEVeyDethsqojG6mWGM9SxAw7EdK4
eQlpHquVQJwM8pgq+BDvsvd8xmOT/ZJN1+skhH163+ELwH9iiwBUjw7ey3/fzQBX
OZfwVaelhvOyc1a0PjFHdn/SrlOOvP3opBiXS2wM17UKKiZzJnjUtr2tLtZqGpzV
gAOQuXwwDe8JQXmSlgOfRrVgOq9ixpigLT4ohRFdjQalMtfk7h98Y5xljzt+fsLc
yetZVw1GlAfuJY1JX/KEkEqCdToGONg3x3f27mZc5sLqbkUpNj/5bIfvsJzHCkSg
pVMpCj4FBjgy/ZK33GhUn82VQ/6fDw5eXhEDy0l2ml9e1KBV1SSa9fmxAvZWMlIr
QxGRlTM7DJftOjOnPglqzg/Rpr14GG8AHBR2YIwdGnGiz+xKxlGc+jXJDRN1Kjvb
qhcxY0r87UjBVA1vloLIkS3rt5k915Xt7OYQvvVDUNkXYpDR52GgG3UHd8OTWIPR
iwCUtXzw0Jbf+d0f+jKyma2148hv4h107Maa5W0j3A8k+RaHvVfmgH1yhxk8IzVW
pr0OUFGVevIqeZEEkMUj7XjkbFfAiC1GvKiMVSalwuKoqyyKiNuPlVWnA5TG9KCf
SnSz7Kt1rm9y655gJvAxxA+zLU9dHcWgD+XBqFoJWmQZX+vxu2ul6LHJktdnXr0l
Nr98wZuBOOGPWdS2kdU7UGrG+413aRVhnXhYG2erVO5viBH+awPYLklogaiooc9R
SR/wCrQwcvXtwDZFP4MKUEPINfh2h55Ozv60e6C3Ge1ypFg23CAo0WFbhh2e9dBo
3eeEVVrluaDjswJZKUD/v8R8m7oX+MNMQTgr0jCV1Dov0hnU0thTSaPx4LnORHzn
5dBRp8jxG+UFOLiMoaqojMwVRChwD1AQc0p8f7KsJwls5HTRoTwsXdkxJUEKYflM
pA7MdAda3MpntSurNgzljTUTW549emX8IqVNhthgoMR/AE1F2sLHqP5q61IRPxim
JWSpK8gpZ3SBkhPZ6clnThv3QoILrxONV4uEN3hXvygukZrkG/pRFQIKTFemfCYD
fsWeSdod+HWTBg1EkgJUmRPiLjC9dfsKmTxrl+DPQrV4rFHFYZJ8PLGTfU8FgVkw
djcnoaZzGbW83wuLd1Z+Yu+4OIiAbkvx48fmamPtNFY9qjFq/0HQXJLvKF98ZHpP
soH9HC0u9Q0pBI1eE+69g7C1Eo1ceSkwqBnh+e3Di4j3PKaddYIdjqVKWUP3uPu+
hE5mut5elgTdzvVBOUwrhT1+qWJiM2uyz8Vd2jRgEd0dL7h5UbR+ZqMnkn34T8Yj
XAq0d3ilOMRMkXm80MngcsP1IM8aEDJXKobMa/7kPjnltGsCxA1CWk3W+JT62LnL
pn3wXAxwDTD+PluGhl4SqY7BnEhTyt+XwS72waTuVf07oV/Q+FuwfcHd+L6GidLU
0YYn4i8Jg7BdGxM1ccDQqdWBlJJONNqMuyIFyjLO1qWmKhCO39EfQ5gOvJ54/ho+
DMDNKbRon0yN8vBzZMkOhWWEACzdVetid7bfSjZtgaywGeFQ4gDIhtnn1tSHo9WZ
Z0v0gDFL5Kcg8FYSt4ZqdzHbRuULmFgJZ4jHjF9sXXEZonRbY6J10ob/DICyJ13N
Pt4T7RRSrDCXU6NF/CUYtCNuEG1kCVyCWM0hQ1azv0CAh1+4nTpLHkJaXy0wdhWr
2n5/e1a0O0cHmgH0ZIeie12YdahG/ig558ANO/a2Zt/M2DlSqDWdz5lrr23ONaGN
J5qLs5mRXZVqPXzsWu4KIa1MR8m6IRhH+wu9HpNgA9bebm5XwdZpVWKfdHgGCEHc
9T6o+RY37jRwqBc+s8wdNxBRIIhXKCse60FkSoSngpTSCDgisQB8Q7W3xT4vvcXm
KIInj6+Q9gJpXFgFKrP3ENmCrSsydZViymTVkN3e/KGo7QwzHvhOSwiB7bIn3Yuf
/PSxSIGfq36fLk0F7FJhHqtunUBE4ZzLZkJh8eX6ttedeG7oG3+FarxpwUIxVBZ+
M/rvf3sJ0Ot1TJp8jfDis+WzmB8U0MNFYlWfIpfQ900h3fDFvhAo3aRXbNY0HMoF
C1xtN859ii+uCknBebkHom+vO3k+rhF/hKePn9H4DupgTFyOaQjLVYA7DeO1bXvF
3h4xaArsqojHs576L9lWM0R+Uu6LlbFezxy6oHF4S+2mPLZjo1iQBO3IbGGOFPWt
vOgcTeBmEbxWi4TogQ7pZi44YzjXkcJYchiikFyosoKrBMYCP+2vSbJ6MN95/kLI
6x0V6IB2oTyAoTLWyWsv7+ZeLK3vYY4uYXw9PGpTIbFLSO8HglGxueUHD1Q5MBkw
alM6Y65/BpUsGnA7A8kOeUTBBOw1rgmKpkGPgibmJGcCMmHkXDlr4DEaGhauOi7p
xTvDvQhIrWnm0CWHKFilvjtkeVnCUnmYYugxQy6SI//gK9IeaV67jMjVIaC32XDi
8Jq3xLURnX7klafcQngA4m7cA009Kz9+Xv5QaiSueQVJbKjew9fPinSvjqRDRR39
KBOwmf4Y6NPvn4cPZtT3NLDl5int0NYOcSqqkALZ5WBbzswYlv5aB3eO8Qp33XaV
1CBiHl+hO2BHQgV0Wt8g6K8QqTnzUzx8NHmq8CE6bqDq8zW73oXwA5YFL/pZAIjw
hTUt+3kPfg3uPsq7g+MyhouCyhx9hJj7faR2lNltDZVKd/fTlLKYevcJnqdSuCcl
dpP3erbljt9FLoEas23dtDnVH87dJm8iw9Dk6EtL1i18TRO33YJBwZu4pFs64DDd
c94TzkYEEp3NoN8YBlEyvQ0Ku+KrmjujQaLOhx5vLGyvQ7BeDC+Iqrj96WQMrZNW
XdisDLjQwAA1gMU/0qbbybsas8VRwVpYSTRW3En3nYi0gRgrpBRqJhNd1xaXTeCU
68NJ5XYWXnwdFPtxVzndy+zAL5d8CwyLlwWGIhB2tdqWJ6LlboIXgoYepcI0VA/9
xmzsmBzRo9u+MRme/B8Q4ZKisA1mWlx7ePU8rfiJociyrqlmqf2fAoxbQcKv0jXh
EK4xXW6Ve7J4h8dM0RdwjVkGFYRrK0j17U+v5ByVBsKGj60SxU7ZwToNxosdu6+U
9ce4XUzFafNMXdab4j9yXdQQagoxkABLFd6ic2Y8/vH3T7k8FaNEIEueBgeU1Vve
4psg5nNFeBFoZSFqmaAfvQMU3qakx6d+/iYwphg3xURBxb+Pnwb9GZIm52N+9/91
So97dECi0wSP4VLHpnLfV7zQzNgvPhrnK8W2HRtP4EEqxR8hLwVGVMFhTY9By1w0
yuIzIbyWybjurhEiN5/GkP0y7Uex5wyxwsemRy0e9oS0KezvB0LWKhq2927IfVu6
rllo3hlxKmdh4uNnPMdBu0OGMGK2U9q8MBkerHpvDfDxtxkyEX5ifW0d37Bw5pLM
d6ETpLAQOI32CiwQmBuEffVDuchJmtYEBJP5NxarBxATqx3wAdcxdo8vfDq/AbHp
34OVmxEt6heX2sSytCzIX2nJhq5Mn/s/sNI6geMzxYb4sPR5N+pLfYwFiEwpmOnb
UHaUsJOJu7N8fKHLlPx3kvQfrF4Nck5fZ1UnusM7czBWRlGqowb0t0LsdasVkpyb
y4P9E7QBjc9WOdcQEVWbxw7bMCulBKWWhWOHQ8B8O+xXUcZLsPLtNZmDxRqlgU4X
m3igo5Ei/IU9rF5kuXQpNUGBEM1c/T5qsHDJHSD6ta9Yk7tXv446M4k/6JKRNAuZ
BPndD+BD2z/ZxcD7jgF64d/oIx0TUsXU7bcBQsR1nbCfP23/KAslem9RTm+70dWL
ZLsmXJKkNuxi2B0Z1udBvCv+FR1inj9Plog5UG1nsG6L+Y5fYowKo3KahEElLkxk
dZJTY3xBOM5HwwuWrgLwrmlKyuwlVZam1q34kUkpUGV5ZDTkeLeNRkDTVfkarnRf
Nx6wXTJb065Jsx29Mlc30RqvrmKe9+MyKQ9L8YzICZdkNluNkvyOng/IfMDAYxVX
c/tRePnCC59mJfLA4zKOLgoeQgEBAtgYeyAV/MLhh/ZdJKkhB7pXVXj3v26ff65l
94up7Dk26QMt+reh18+zP+4MoT3XZ4AX2yERdql1+Vz5NjN3OFVi093xRm+1LkPb
8Z0BYp+Nfd38i6BswJa9+ZsE25mkYGox4e1cj6AdIObmglmVB25U8ZMPGgZm16kR
kMTsDRv0w5no5geGYd7BKRYLI6zBMt7tzLXNGxbpY4dog7cc0gnUqDzb4ug1tuyJ
Rs1RsyFm9YYFsKfhdbPsVD3mx8JxfnH7YpXtpwQuH+eUq9YN7tfIDuecIkRmokQv
0bbTwMRNE2hmfLRsrWPiKtf7FSOmpJiT5GUrjkGUy1nLvJ3NeeueFhc1nDU4TcVy
2t23dfQaK92v+B7A1xf/0yeVTHoK4hTk0SkEz7zRzgJILQPzPBTsDrIVon5rinV8
zGYqf3n1bYL8RTDdb7+lxIT2wPrkM5NDbcV3/hgf3TfeRXPljshlV1sFWgY7oywg
PXFozubU8HW1LgoQjPiv2mUWD5SA/AU5OBTU73r8t4tUKm3SJylEIXBGd8IwhTHt
vzqLT5dOBGoCt2NkTFUPjkHPF121l/hvd9bgP97cN7riaj9kyJSOUu0mVNpF3PRT
BANbGg3hTbda+AkzuT6A9rYsqb+aZaUxI/Q5bawXuJZsFks2cpypPN5975oxkTIP
bE47I+BmmjWdHpnPNp9TZhK/J/c0k+5v3y4yKATVxFolbJipoczjDy6lSw3f/WT/
84SVljZeixk7taH8h3Er7vkD7hPBGI6IkIY6IIPo6kXryB3I/06AppEP4HtOKj1d
ULyTspmJdjQhmM68tfTnbleLLSKfYm8D8nWaj9RgCMXW2ZXFUkSRuI+/OVOfdHQJ
drd4C2HZvQbjtjHngqVGsFi2WQNDiHOKOHYWjrbF9W/idB7h/ZKRn20+QAje2bq8
5AuY8EvvhQxeUZzAjc8Erw4V4ksgB+m94FM0bN239yCn+nd2DDJgW2+YJS8tnRUK
tCRcH/YNoE+KXYf41Vf3y79OR5weIxZJ5AuixvbgdKdvbczjY4YLL92NPtB35QGa
jnNXebqOnfANtKg7+Nsztkt4nkeouvCEihOqEdjq+XsVAABm+VT8NVfuDcdXgc/X
3lLMV4GIWYk3hf4KuqV5qyuRSWEpYfiPTiDHe8L+fXAilQSjbI3otn+sSOIOOSZv
RczQS3Y7mQKMF1Qt3BA4aqEdBiudvjm34XTnpwaaxjq8VOAfBZB8LdynsNsDrf5u
3+t6282jkivZM7tCsmTLm7s0ov/RiLlJFUt4QtnScnF09x4uJh5rvEIQsCvnCpl0
pwQ5wW8sHnVd/aZa8WlY6xKXZ7aWgGGHBQeD4+wG0f/GJ+m9nSStjnE4z7LVeCM4
X4oavStn6tZ0TkfFAzV1aG+lkP0N8CUGf0Ly7YHiznf6RL0PlJoJ4lAaRPrldPiZ
bs0mYwgvAAdmT55pUuusm8p/uFQt4KrOeXriUTy6CpjptLRcgQgYuirNIcPxzdJf
4y3jo7419ETqMNvy1PGyqV7wDK/qVjKzq2ZIP6LpZZYkegcBttOA6/SStxGfqCYF
PKVhrJI+1NItrBhkfePGNFvNA7QlSYnIow5/P0JyWbNB8tLPKhXimnsdpOo60MBk
22q8sCqZ5B8C2qWJ6XIEZxknVH4DySTKObqndl96TsYQwXln6JXmpH3b+igGgFuY
eaE36Be0DZYlNp1qivwK1SzvDrvF/Ks3B0m60lxwRuIW6p/jSCkw83C/oaNTMQTX
TPs7AE62FvHZx7kcZdJqoLWgpLcdWE4Lq4pWwzP4hFwowydALdGeKgp2ctJrdEOV
LvqGT0NSHB/3NAREKW9GzHjv+yeV7oS+K60gw7ZuMzBN4NQ6wbH37uNeJfFPZphE
zwr0gABVW3UhFiMYGy5gDtER+hkg91p3lWwhuvHbEunnWjoM5ls4dboOUwpNeV1v
nbjW6Mbf19+9kmBWcbD8OrFfu8KA0iwj/OeT8dyvXVYp6z+DasqONFID0W8z7uUC
50xO0rpETeBr+rLbz6K9mWs0XqznVEOgbNeIRzQyjoZULv+HfOgzJX3UMMKQ6zie
7vzuKfnhYj0N8ujbMf2YXAFH6HZAFD2mweKMztMPru67yHWNMIjzsN/sln2bvs3I
mqCEwQouqr4WObGxKnWpemQH1hFn/CvEPaLnChocx9Hzd/gjvZKUCscOcrSplVxZ
HIyafz1M9mHGgAfA9GzZk24OUyiiuQUFcJaiHkJmN+ROyc2voh7N30cP1CqCp2kq
0YY81h4XTvVmF07G21h0vzrQs7uPhGCLD7tVZ5dte13XO8UXNzWWwFTccBclGNxz
MSs3hslpCLFDgf69veVYs28nn7kW5b7nbK0vrLakbck8EMj62+WfUVt5GSfrqJCE
PhSNVJ5WmD+TaU9G1rRw7UKJBhJGVHCBN4kbDlrle3vDjiEwsV9zFiZe3146/rMu
LuJiNKI+h5Q+Die+vIE6hK3FBkFzP+TZ/NRSFs+iFcH0Jt5eabK4CH85mXdLVInf
nOjMBv31iHJ8TDoZylIqE4K2a6kcuHSfmXEizXS/6XiTWCqX1SROaq84SsfAM9nX
D+G1HMY51F9vdLH171xkHkNzuD4tutoov63pVK6sryKP7BlB5oMb1yOXB7HEQ7Jl
b+tX/OZnWTQRGWvRECMiWDQDvKktye14bd1teE7aLSaG4F6j4Uv2ezPkC5ASYSeU
dKfqveCgKlv3gPB95/K7g2SueAH/hduFLLBowOMgsP9R28H9PJyaw5kFlX2dvhOH
hhRVrsVHsRYkrfWumF2WKD+DKAhguPqMg5NIjR4W8gubyGoEtW/y1Q5Q5kJxYnoF
lO5aenqg+ab4g5lbYIf0E06RX4oGB7rSfuaE9QAQ5vxRRmjKSyEB7rHg5MFtCRuz
Jx5wC8SPwM9+tuOXgt6SEuRQ2B+vE1R526DFwFKHo+PwuZy0pkp+AguXgEXFVO7c
U5czpKrGv+gRx2fsmYPnzDJGVG/bPSESFS+thmDYBIF2A58d6pRuUZ8NO5FO/4OM
qzXABh+gJvRQIQLX4qZu8jYTSjzVn7YN19TqwDEJzIcaXTpwcziB/dTiuxjSjLxp
lUcpj8Ww+/h4c9aHhl/P0DSa8+PHciej4XQHfmX22bjig2w+N3qzoWbOxmldTQ+0
1xm2J9AdqECvMA3rcEnhVglU+1B/C1gj/gj4bD92C+pdZSQerMp5+uXCv07zX8XQ
je13WBMmIussZrZXgsGl7sqx8avOxhMwu6wbVmyzt6uZw4QlcnMCZFdk9XZSCVas
Gn9YTtpTEOQcWveRaKxF1+XHxccGsQkqvZWAtZJby0RW2a2JQkRniCni2Fi8KcjR
iAJaerTFjY3ZMpzVpVwIgDAO3PCQomPo984lx/+fx9VYEKPdB6HDg5RO1pyzN8Al
0TwaxuR9AUMdjRY8staSZcJTzb/j4EKqrWjOoLGfqhNfHSJD77p2DttL0iAcANHo
W1sDx2rMyOajT5LFlXNoI4y5zyINEuuMeO2gvl25efwwg1fogBJnOS7r5N0fv+6r
xr3OtDCV+u+R7fyH5EEQVfuY3BZnZl3oZVfq1QO5tVU9b4zrPR7qJ+IIVscdC9s0
Cca2kaq0ApkANJAyQ8ve2rv7n8v8DgiVU91fKa7hjRGSQRT2uUZAz1HQtQ5nvl6j
dcdWxspQe9H7oFydpwbIbFIqkfrYVyBEgRJs7j8GCcHI5WdiFWRj2hcnNxRlXhwl
x0j3QyexhvAdxumkB0ldQOPjNi3TgRKRYZRXP4rCp1VfekpNXR3HYhv/aOBNfbKe
VZO9bSIrE7zTc32nZu5qinSizz9qwJMDdcrCyrPOlSCrYWW9baXTKXLdQw4ZE+K2
kiM5I24rDLrlnf0rn/1mOlthuhRTmNyoxyBvAk4zqHtGcdScX5RMk16in79milmY
Q8YRHL97ljyGbCjTawgaapD88O6LcGIVymBBli1o8mIylvjEBXyeW43Bo/o5gYHR
fwDWofFjeN7CGJrEaVrzOapSSMXhXOLdKVxsIPBOXSWeTejH19MV31/T6G0EdFL+
0sucJRAhEKLAgOhyqVCUealcvLWheGy0Ts1BToVDZ2SWMWvykeBrdhj00RABGLie
8v1FN5xvKpPZPwl3Gw+E9xbXONIKdeqpLOoJQaeudzAwAW8mxW0RJ1QzyrcETr2x
PuPRr42vZ/x3E3yR9apl6Y+BWeDFppmIkDrzqr9SpoEM5nPlVEWc63pyPaMHuo//
bqsxNZ9eLE1yC1OLT6G1HY3Th02nVqI41XmIlJhO+6sRegnWHczoi1KqtL8w9FLN
QKI5L/xHiU287lThksbPvAj+qr/DQiI/ZCtLNOW3nx18eg8JkfgsK7UNBq20gOhj
e/+7AxAzrrIpm96bR/8mt+i15GMPa1FFrrAIIoe0ZkQDsGQHqdcV6U/5+e1Vtcbf
cmz5aHH6HgzYrbQ4iBv4lOFUvQtROOQO1HIqCP8Q5eaZyFz3xlAdfdOOx8Zy/dTk
L+oIpsEFjL0lReu3gmzccNaBtdTSKIq9S7Q4FvCijo/g/cK/qelUZ18X6kuDehBc
gD2BIHGNk8jKXixvVyoGFZP8sth3iB3X7TM0M4vwBxvbwE1fcLxhqBicRhteGW/O
schZdIa+RNEhY42s3GXzalg3kvJzraemPrQRJR7Hxzu/YiS7zWFKI2Hr11Q7KTxi
70ZQYpNt2fQrX/dMn/HJAdbCp2DSRq36EpUB7Tz8w8/kzHUTD9JuUW3vIh7kWYiq
7RpYGMgitVJVGWKVvGV1W/MTQayy6q039PcMFNL9ZCoeUIQm8LtdXCOQuH4Oh5lT
vWKJMXahwG2ou3ukLj1zippS8/Y6PT9cidmUDk38GE7hH1zm4rQlUGYpAyRJoMIS
0NnOtl9nno4GxiH0XDf+YME+FZj5Yt97len4cmCfUyfqiEJWnb/vGzXibS4CPCH5
azKTZh6Rl0UmQe/W/cVgGMST0aKUCT1/wjOmDlamRLNwyIn9enDfdf8ZTGsU0EcD
NubVUk3KadV/eXkgGNB8mSaKu0+sWG41kUxi9sF/R/iMmOD0OnZ5gNeh2U2xUux1
4oMYt4BBufcKyjvCSMIL5tzfs77y+UnT8qUz/gWW8bzKQ1K6QpmKpWUlAZSnM5KX
VIGMnjSaxBkrM381sPxueYlHx8O99MbLVgobqNq5FvZIgZ7dgZd7Wmmwc5X58JhV
7G8LK86YfDN/Bk3djOcZ8n80J9TkYGkjCykr04n/v8D0bIFtxLW6Yp3uduM4CSJ1
igpn0Q/8eW7nyUbQFsCmwVl3J1AfGWjEFjroQGbr3398zM+YYtyNZZajCxfI2bdG
POFcsf+GQMCy52c6lvPNLckJmq5gm0MpR8H3bJ4Tv4VcFlzaGlCwqUyWAvF2n+l7
wo6BjYQhyNArTL62TQOSYy666L3L8WefKqO68p8mQXQdI2X84R/BUCfyB6NOj3sE
ROKYkRTC3wA3j7JDUAGne0JLPcyvTcEBqWzfqXb91HXULkX2fbwd0ra0d1bt+u31
K2PDRyUDniFDX7EcKtLZ5SkbB15NotGKUcoQjyKtaZzFa/SOPQg0Wgn2hGMsi3oX
t9yNFWlJ0X8x9+y7c8tJo33ahRmaJADjTlxyyhWwG/kacQYMzc3FiFPsNBKvAj3E
z0RjCWL7eAKd6G5vmvQv+pABZl+tA1N4yPSDmPzLV/ZHZ5603AXw53bwgo43XDmy
hlCKGLfE7EZ6khpkgk7jamWf9RT/JvIhPWx1MNLUEDFvFp5wF23jNGWEjH5Xa+9Q
73fniBaqz3oZJNpqd7EKna/MvmTGP5zx9EDVCwWbuneuKar+kl0Tovp1jhgDEr0R
qegyPJopkuE0p0n9c0UNrMeiyabX6v/90soDqm4IJFmZdIfOtsR0brVIvU7OLQXp
PWfevgveIqsR0CJ00FxPED/IOguF5Iqed9MtPlpAtIuvaWJk2fGXV2/je0aNnXuu
6n2rIB3lbQGrlb8MRmdkQBxBNG/ofpFSfPFsUB0L09FkBHc7CV/BcAzbuHiT8EYe
qtNzqqm/iXTo6dkIiPUY1xsodcWMZpIMUJn1zAgNHejD8Q+GSnKtvhQkgc8nkZrQ
ILNqi4EpepYiQoFWH1FEIUwqYSvTkyYVo0ERnuVF8Jx+jGS4nO33vnsXRENov0qC
MZ6lqWcfsakup10G24cLfCHa89P3b/yIJVT8/FqgFtRnHTiuV+ZWHtAeyqnE3R2Q
QBUObLLfI4NkmZsCJxlEkWrsaEdTCKRSNoaeVcBLRkDY6l6N9CWjxn+yVo1f5xIK
3tA3Ckq8PhTpvCFjq1HG3q1/4QBiFUIcCfml5nVf/kSQ7QrUc7IOcb7t6jk80+Aa
aLiGU9LzmZYKI7FIHPQQnfqJNCPSTH/mvA2zygqiLl6W7AjYtMxHYmtxMT5IiGGH
YyVlSAxvc/vHjlKu0YbiuFnArFbI+UtWoxjiU8ErkF056ztoqy8JSCRLsw8dHfY3
4IbN3crbfiutBaycIKUJ42H+ISnqBXq1CnpGNZaUyKCfpBQ1ol76NLvBbU/fLmws
ooSOR36AEz/i3O4P6J2vBs+ronrwXR0oYHUK/S8EiRW/sx2a9/u+6KiNmgLAwcRC
lETc4EMc6NQb09iktSHBYgEzu+dKK7dEJ+9dGJmwbWB1JeX7Vub16McZOsof+VTC
szd802rWA/wnRPipZMVuHJjCCQ2g0KGx2u9VZ4kDRv+h/bWOkQOtOLIztIKWO9NN
JpdMRQ9xSmld43C5phswGEcJuB3zmg4waVFOFYyAQDtXmKTSRSjFWPDEaVkkRg9I
2Xw6rsoYR6noPB02O2s3+mxQkVSjVGYa/DG5wD8qoQ4/c70RG4+lPXIA+ujbaD8w
cGgkQfzbVI+rqlV8lbYa8uZtXnBHnptLSl/A14/pSqnllIYcIl6vFyZUYYas7/yk
LF/SNsZzC24/cDV5/PLIQThCa5zKOE3LPvamckaDiSgv6UVHQUeL09ep7R/JxGMO
CAH9oQoQzdgB7VcGRtPKFbwHusMdcGxOcz6qAofe/lHPH0l4pctod+HlXu3UPj2v
tbe1L/7kz7waJI883KCg4V+gJ3Ox9Py7J5hWTcc7XWF3Q9EFfV4T72vRnO/Dkc+X
k29nPJcJzmyvZa/kLrZHuuefcItdBowK3yHXpcjP6QAV0/K15Dn+Kd9pBBXr7Apz
/7bxjVEVRZYImIEvcKnag9bYFp+rUjflxYQ5ZlV93gJkVmyTgff0FV3vPJFbsLUa
KJo6BJWvG/8CTBRsSOzqv+h7Oc9cNsLnMs0wU+d8BuBgxGgHH5AeDDlt6xcFeMGB
Fop6quFZoGKqQP0YPHnpftAYrzGeWG+zxKYWu/NYLJ44oufvD30BXgNfj6VA9r/g
PiE76geoTNwFRAoEkQjlJpafi+XJPOegQocaRZorfqPnJFrX93+JMibbPNC9zovz
0LxkDggVb/pXsi3pKwEnHj2cLsUGc+w64PC4IBmgW3UojjfK8wa4EbU8EBBk+QCU
1EkwmM6KS7+PFiRhHMuMPC6Rj8EgMOEmn9lVCTaIgQLWXCoNsPMJ1JF1RT+2WwjY
vhMW3j4dFDDnYk+oQ4bhAb/06B+cccRwjpjj41KgD22PL0dYH9adGe5zvj9FpwDx
Gz+An24KLHKL/E9YfjMNbpxfFrqR+r5TO0aAUQARzQiLo7ls42s3ku8iPYcugnm3
U74wBxODsMO5aPgld2yL9MnsRkCiclv3DTUl8V5nMMKcYJweVCVen/+WB0RMQlUR
LAnmt4R+jzBbZxjTFKmaiqf2oB6alyQFhiQ7W0IuStZFL1BvXZpnneP0SCJEapSZ
dOO5XSi6K1lOgMgPlhXOj1pZ7U8sADemvp5e2kk+vUEt2YDntjUMehi694znclwX
xqH5v5vzW7zBgwbrgO+BZUHtX6v6UQlRG1cseNOae64KsnycMo8jCsru3dcPCDzi
uk/Kg5EPuYYrinK5pCAr3iNQjnbDLQbgqPhYGl/ZTWMhHYBQj3WHBPGaBoELJbSc
0OgjUVLxW0ZqEVuhdmiYKvce7658uxA7Dm9utmynchcDkgZSrPRs2uFJ8dRKfYeP
p2FKCIn949gM8JD8AlIBMlhXGI1rGxVZ16fnNK9tNrg93O+lnBk362gEc95OgwgZ
+Nbp/ELDoZ4/4RUGwCHYAFtwssO71exIfUwSoJWl3xmqbkquT6EP/rY2QkuFJ3Ed
lNI00EfYHam0AP4N4Ww7/VqN6oSudO0p6RvJ/PYPeBuxxUjvoSiX2LrPD3sy9qOF
n7TIrOx/KzPKyfIzhxFBTpZNXrplpdC8orVdC7YMkI9llI9MDPAOdpjkFv319vWy
NpUTfIJEp5dbKKLNoMrx+IVCPoc5bgdyqip8kuYu0BQLXd1jy37iPgfK3tDUvrR1
XxCvNtV6U6cGDxfajXBe6sML8Tku9erz4b1XOmValVRTztEvtYB8SWsRBwB6FU4Y
APeLnRRSztMJHIZsvhE5T29L6UVAB/MoW7mnEPHAW63Ggy/ZiQvTGcU1iVOdv913
0VfgSgX2R048EItTkYK79+ChwOXQlpcpShNsEuUZUs9ZrynUEQZDVBI8Vv2GWegc
50/nOFB+2ZsZJxszFtJThGZbVVYvagpGHzntu7baRrn7bpNMYvtDUdmO86KNfor4
DxlZO213UJRzSjwlZynogZzyvZSF8RnXian0hVJfJfPSb+8e6DVVVs34yOSSGhap
vBNh2u8iB+2m/JgDfZ48HopN3b5Mdu8yyd64J7ycBM2nPosBtE90Ebr5bNeAFX4n
IaIev9IOzsItA4lCWDVMNZuJTjB/cOWHGTeiFz2pPkGqRlzcS3DpRR9HaZXaslL0
tvH5BXXMFJr0VCxSPgRd5poWf5fNSAR3wpgiZOl3INnCjXBmqiCWqsLSAleuxhIg
seqwPHzAm6V+po6owUqFCFmu4/QaJFVi60j4JJmbTqZPlati7mWboOyOf/urFZfN
Wmpkstxd7O9YuINYvZHiYZkYfXGivUcSLQMSjZC/IKf0y88o37hPxNOf4me9uKQd
Xm87UouBTD12TQr6GABGAlUUrbFbHRMv6rpXS8yzIKjwi0I7y+0kL9Bh2NIl2CPq
dosAWivN8QS+whNE4EZpiGPF3vQAe/xiwr2uZxEbWFvjCGBIApvlq4FAIrjGps1M
1tBeDw9Oio1EZHpGXr+wkA+I+Yb5UewvVEOCzWP4We5CunzFndpAYNZbDn+OShvA
VPw96F39orZnq2A28leq+s+YTgpeQflY+/3ooJjr/4qrWDseLIPEjY2LjblrT0ia
1tYYG9PUvuXJyE5W+Bo0M9pdjM9y+q+CjUBvOh5ik2v+C0B4z1PtDnM//rpDdI66
gdhyd+30wG3jfAatKDJXXezaqUtqZAMY0jsmnieuCNi1n8QtMetLOy5Ovyv5wrLp
YLNPS9GoGRIU8COwsLYfcANRjs1wKsZzBOdPy1/C4Kuzpv556cSr3OBXWGShRXMR
srCzXEluZA2uzL28NcVnEKf+MeFq394j9e+MsJgAWIwGiL5dgWg5YtezMfQEkW5E
KZMl8paJC5b7bj+qlGrTFatSyPjLbGguujBBvP57/kFWKJkv/8dHHwUjla8Qqodq
ZFVQAFJEz4lNHartuz8UzE/Z9aPAMCGtJZGOHQDvNJYDptFtG+nNudwkvPrwyVgG
hSSL68gxGiLc0xgXXM7v+8jZF28j1CeRF4aKPd3r2FfbjzUst33Nq5Cm5JOA/Y9T
B2qK0SqIL1NeKMsAJkg/8T3B/E4S8UAciyK2UJ3G2lott5FM5dXE632a7udtLIq9
xhnOJSb5jN0HX3jT8QNEawp9u9iuv1PoFBJUNYoEjJI/IoQufGj3gddc2tTz2wv6
taDDphL0/xbSKX5IrWVjmfULnokQ+ZWhPFJ0KbTZwsPF9Pvw7Q7mK1t3RDCkexOi
On8atdfMVgiHjZKs9q1FdUiGsUrFfVSOZLvA8Du+PVHP2k4ukPea88Dvr08hnJgf
LwziPjQVvruoCqQgsG0cC/RN5hmnSreQloMAmM9POLTK34rXN3cgMCZI62VCOPHM
tb7hPdUPIDryTZoaKFgyHXldv1fvnqmJQvc8bbGu5cs4jRp0DuGJXlzdZMe9UkQn
/HoTGP1aye9077HiLIG1WaiU8FuKd4IB9QlLpb/0lYEcyO540Zc+TKduDTy//5DO
m4sT8It4NSFS9cY/wbM+g9cdLm0mJjcJR9trENo+iBptexULSvaUj9n1zU1MC8gy
B9sd6JTILOaE/sm7skFQssJImLRb8MDfrhPWyZsCWJ2W74eYrUwcQF1jKxXwdBT/
63jrVQCbLhfL76/rvseCToxA6KiP3y4hfYPkx15NQRfS6pLor4Qq+D4wdWeIm+4I
eX6QoEDAcCpAipg25oQg7RDKTJStx4tQTel5Lcxk2lC8SZd/o6qJFSmTyy9uwc+9
0EUCx/2cLkG2fDR2CwGrc7QgQxRBQcae56TdSJuby6GRmpDNECC6cM1uaHSoVhj+
GWnrWV9PStbjFogcJ0Cc0032rQUeAgApr4eW6qZskK8fp6zAGWVOymoQDAA3GyOT
8AkJGgRsACYnLDatOUgBUAaDwKFWaHWundoLUjR5RNgOV1Aq7xu3vm6W3o+CjGsI
YSxp6TQxGXbJiCYTuoLwoe71B6Vx3EgM9v6v96VTm01nGngIMBK4jhh+c0F/PMBD
s6h0letQYvGnFL7PBLIVQfnGqzTfbgqHrfc38wAH9EOuN6g+1iLzy0FdISYqWRoS
srPAWmg4stcUzny8tg/RssaztIbcq8Vy2Pikn5tnVfhD/gBeTyQ2i6jR2K1cA/zT
YuIdiC6MHmY6fOPmNO+q1lXq9aCwe+Fk+hKVFk+JG7kOXhS2AZbwmMpOrN4IjIRb
AYnnJ569Ict/0A0ubEaXYfgKdCp31Z4UYAhbcf2kexxIvcdbU1p8dixPgp5BKSq/
DqNrpiy21uiWcIQlISaGpqukUhX4nGjx/aga+boZwnJI4zDq6vZPXKfgaoZPZ/Re
zB2UnPsFRMAvGlP+LxFYluEqhqYJ0u1T9CQjE8cLt6QdigLqDL3szUgY3RE1D5n2
MsJysm/BQ8Q2nmHUo5SNN9p939/CE0dcnmoLEmV8yJxw+2hcOSSDC+BLVyqV5xLf
trsHB0/xlAoq7yazMVUwm7GoLLYJrPJKRAEnHhMN23lEf6l07SGwVFXjRaxb9RMO
liImP+ZINtVetn+bywMI5dgLbl5GlWedavTjkJQtnNZ1gpVeBQfcROpXhjQsHiTr
2FVYeUwmhOColsaTz/Sc3z2EhuBD/3Tq9N0Ncc9Vp0O0GFInKBKl+82Jes6aQTUW
cO/6Ct5cA9Pl4V5f/2WbKZsKVQaQGK+jToDnSL2jBom6Mkj6P8C8vD6ANKvRSDFS
dJOHxu8XC+dngDUg1RQiXNbyVHOST08vArftjGQ4uJ/DZd7XXgAHrQIXNkdijk9j
WjzsvA8UJV3+8S5Q/nLRUQXUzNM2rGB3M5nO2hzz63huOWl5pEgQ1F/oVDPZbnOH
SBaxiIXzRl+JMnCgpMFf5PAcBsLmFzTEcwwbjB9+3R5uhT0Ropz7niWMoLRsiT5E
Toj9cVv/1zAx4ZXjY0PnmgZ4JcQ5ByTrIugQQV4jJEvTok+Uwvzt4OFBQ4GO7UM8
zDgK2B1mQoo62hDv+K0wRpzUZdh0TXIk3dOfUn6nQuyxVINAhRjYYhLtaxIaP284
i/RGrN7XHm0jRtfpuXLKPBJv0u8inHo5gh8HW2Bw6LAi2cFVyYP0HZPB+h+WdfrJ
deBO2yCiJnFxnWWGXC2YXrlqw9pXL3KRAG2VKiWBs12N+uK0KyUbjVhDDewvmysK
KmOLdI2aw/pUZAramR7/T6BTBEHi0acl6NBD27MkGRweld0bkMRVISeEb8HinOsD
anmJVsqBfxPxS8wv7kYCTRLLuMwo19LvlfD+NC5ioG7CqOd42akxq9GGD23tQSfJ
W1+PebAr+CUHzaQ4JoR/WER76pymEHa33qwAi4opGqfXQDVkrMRZuYWk1x9t7Rh1
CWcejOOWb2is58PERD22fJTBE0SbIKgp2Cf6bq6IcCoEtYMxdt+PTeXQpWWRHuVO
I3gef5kpAQ6rExTLVlRcrfw3QqMiaBnjqYfcy4U2wmfn5zDwjqiHfVIgR8habcX0
CBbwzgQhQ5AYS6jUpnHfCIpGcMdxVSAW3xse/h3ol97gkOHn6NVQSnv5K7eV7MHK
AiZA40mYqVMUWEF8MEiRdj/9SM/Su1IpSv0++LfmN/TXt4lQWCACvxJkgvgOlRXj
1wXvive3AT+e6SZ9YEA/jHYFkjUeC1yFmKu5vBAmDKbF1HxdvEEOR9vXao9najcR
rsRe3BH52PAtlhc8d5Y09sFmg05pyAREgw/7CzX4t0Lebh+vCrX/Ox3p3wxo8iDO
CKPOyhRYf18xrCTNNFzWGjfIgzwmpLIL9cWzIG7gN4wjRNdooRcIHCuaLQKX9NOr
aiGUMjnzYvWB4RBpFv3a3dMvMmbM2qCsJzVp1E/HbrmLtGxo2CwhesLDGsREfxrn
1QoaCad54MF35pzAzI+hPtqOsb7ZreJgafmOQX1hrj7dj83Wtr1TSXYhn8TxcolO
EQkicpYPXUihqBAtYb2V1Y36Fms0DfLLb05Li3lk4qkvGkmJTWt9Ajl6IUBQoAeZ
Xkw7hiYfpGumGilRG9oet+q3nBH3/aP8oI1oeB3gwW94wpcj/OSvenwsUluMDbog
8gSoy6LQi49qftVowgEZqZGIZqNehJU4q3ZJdQ/44+I/Qt8dOfZb6a+HX8mD6OQ1
Mbe3KMcWvl54GP5Czv0UNF2mP/FLlolD1nlY+VnA/rLLF4S1JDSNKAkMj34Kobdl
ugSnjGlj0YfgGl8cY/1WlCoX7mzYUkvyTCn+WCKs3w/JRTYRN8Y4skz/IrMjzR6p
3FnCPCdUqZxEd0tKJG/BoXk/mV3QbonslL2T2pvazGLApMx68i3zbgWPizuE70MR
HcZ8OEMpDixsmLmPU+gN/irzpXz43W6a3B4sFC9Sw73ElFFAFAHDHdJGhIlrMU9D
1KW3iUPlzjX6E8U3N3skoI8A9m9LCpsglDSkfyD89bOAKNR/lM0d6M+jYFIs+pho
15aeoPfC9z+VG0cI0S28dNmT9jUEPOl5GrcGQajD1jsG2k4RgLWoYc+acJiTrWeZ
jlmfgraakRj8UoC/tA/034Oa5d9mkuc0X1UbAoSDHiZfRgY+TryZcym+L7Cd0WgM
s2Vfhk34I/vltDFxNTcNhNHEEw1S4EkNoIrD6xnJp3xHDgjPo0lxqZbgWuTOD6yX
uSDwNsZf55Zkrw5QrbPb1OHQUCeDmeX6GZF6QWLJ16iwrna7egFiOVmqVN4+iD0M
xAggEVfIqCy/CXaNp4zt32nkBqtG7nHXGXdRfzZ0mEe4C+2ORTBu01iN84+PCJjP
HidyDbFbkDgZ+V92YewILaXq364cPCRp8LSGR20BbxK09WWQCfSQkVPoEHeG7awS
ohgDEOq4ciIJZYjdk89+0ebnCdUCfA+Bf9M7BWPfQ8jqBW1DOhEppctHrYKW8vzR
yBPCBYdC1rK3vWcci6CZxIoQpHYJtGZkJvvMpUs5DFhf9xKpWYFaM7/3Po+qu94G
saG9mIae6jZ0s4gQTTKuqMfxuVk4pvZGwtzOLVsTc0uSx46lkv+C0b65IdtXGJXm
7BUdXggYKuXanBy5jn6EtoautnTjnwNEmUq6XoQO149INkJEOJZ7QDe2s2IoFR2p
NyCjAnXrTeVZWQ5r16nJMamYgWHdYS0kHAtd9yqhNDZrCltgXPnEDCvt5DxQ9TrJ
8AkDkXME4aLLykm6B4tdqeyWcsv0YVfCReqwJi7ajJEafY1F7sr3DxiP0qDA5LPr
WwfGyZOjA2n7dextN9qGAGga1/36/I6wdrlI00mruDmsGy5j54nYaFkzxLlShDyp
2opmVUPvrVGPd12V9MEGM4Co92gyp7lX+iWXX9JzsRzz8yZv1PFG1zPBWIAHXy09
JIHNV2mOFpvCpq6kz40LpYofZuAGfk5fTqONRby45vjZ/6l3yKEElLirnq9m/K7M
5d2TCWhSrMqbA3GwpjNRoMcQiRtymExxriaO6Y1hjyZQG7R6zNYigiUIp71wzWzC
GWDUxgR9FvEjSZ2G/1SquZByQ94i+PKG7O2FjuZ1Gy/u8YG1YtCw/ZmJ1uwIjpYB
jXG6fcDdcrRFwiXFYWCepqNxEavZsLy+wolQArZpf9H1SlDqrL3qCVrpaSpQiqNt
QaDOIFTs1DHELRUgLp3AHxZXQ4jN6yyiYBxznu86XhNM/G/qOqStHtdePV+9380p
VxHbj08At+V/t8wq8QHj9kFO6RFJZovKqQ0nBmCBvoJlq5iD7vCxe9VN1i0WFye0
c5+50orONl4ZnX1FM9TseW7KC8SqCOTOTCeAQK3KPmz5I2x3DCLsOYm98xK4ouN0
T2TFfVxy4lQhSTBAbKLT1S38ldoD1RYrURSRG6s/FHwZtffszY9VW6HEMLPhNHBO
MsY+ik6OaA+hNRrpmqFNE9Ds27qgFdmxVrBqYRV1jr5SD78Z4gUDxCRjyaT77oQ2
FdCK702Wk4Az4i4jIrBLzei4rDYUQXkOsfeHGETqyvbCzIcPR9xxqEEPOtslPnt3
nGaYR5geC+5WhxyeAlDWwjf1e09aH1qswdYzuNv8s4IUuyn4NKLYlmAcfCf6t+Tc
72amCgz4uw4umxwxcw60joofbjCdKeOgQixZuW6+TYJg/PPgDsM4ojRJdAr+Audk
V1NE4ZuaYE5mt/A+4eH7bSfz7nbOaab/i4A2N5sWV2ybxp9C9gkuR6jaX88yE6Fi
iinzgtgEnxmlVIZ7QDE7+7usPSZ1GgO7UhfKgOUqKI7FwMMRi+j53mpZgCSuRqjB
xvrjKYFGLI1V+HDRPquEd3Gz4OI9Uq4aozzN7AuB0KTHD7F2rHFL5qXEZlmSwyaY
ZXyVvToX0pKcdG5hx+LnYAOHBqPoBIvU0BlL60SdB1yeB1m2FLohFAkAF6N8TvyB
o5Xq1IgMhnXT/kFN42LH936XY7aVwMYM6DLKtFMpUhLB38ULoGAVMwLJIP3BsmLY
rCb1zPB0UfOn9xihQdBEnR2JIWYqScal7klGhhkYDMjjqiJZVnKPa8cKLFGfoOld
g8pBQx6+wAl9H5C9JJJp/81muqsG6j3ppdV3qt8BiUIfaDYODoUskx2ywAVd4KPI
UE69XgSqWN/5Ee+IpI4eU/piAaju00iWNO8H13I5byODgxMQ89tcdaBXl75C6H2a
gnwcusbRrPkT/IWd3U8Dd0cfXvRSNVvR08JeR5M/gNAoYCNOK8D01yxHssnXteBb
KibhGuAk1IQppHiPIDpfEwthsyPFLgAFzahaJ8kUOQKR9zib4gDCqCBYzdKwOxCz
ou/KnDbGnHftAySC/DGdKgIsNRVOvRvN2n53stiO43RCwUVJwJBMMxqkUB9PpKhz
KTN2WqZlf+4RuPCyAXkYB6TWWyz8YpCaNqmpnPiKRpZRFjcpa/wQgIUniBK8kgwW
qUaYvVrXxqVgag+QlUSSbA5j9F2ib1h8SG1VQs0tWXgnn2Mhx/LyiU09/Zz8Ei5S
Dw6+s2XJZmmuf4em2+FVdodYbNtfPdhPM8bjfBKb2JDj+/iwAwIm3b8l6b7q9VrP
7GmPpWX4+WRPcm7bcAehwg7uZG0JUdx5WoH1uRWnSK9GEaF7zWA6Q1+kxUfuBeo6
kU+Z+t99vvPzs2QBwuXFnLbs9Kwq57rXworpD1bSFLa1IHFfTy7If1S7q5ZuKaCd
0pWvmwawxKYTxxyoAnbo+evk3WGC9cSZAFf5nCh0Gb638zsbgfjQ9AcSMmHGnD7z
0EXZO8sj5KOZymORcZVYBk6ad4eim31osE0DdqKz44pZXp39a0qbBfsblysH6lwB
w8FBxFl14G34d2aRvPKlTDI0pSoMUM5bfU9AYSyp+6hqqPkq4untyV8Gf1z2shxL
t94FVWXrw/83M6RtY9LzO6wqdxy+gjlVTdx3j5xRVjMj3VEozXSwH5xnDTh1nHRL
k5Jzmzx/ac7K27VkWW0SpTj2Ta9sLNFFgP7I3XF/LT1UaOWVfK4zhjDN3hWTwbW+
Me6KJ5RhDNyIjEbWBlOAo/RwuyTq3guLlieS9+zwkdBlLUKeOfU1qe5m736QAHCc
912If2JPZruAu/9F5VJBWtdrrdJojzz6q48/yzecDjlbaOFHMn5Z8tHLLbRLb0S5
XXJNeXPb5kYRotFuWshLnt+SktmzR/yHBsukd5K5e87RvnssKmkphmY9rFUFTKk9
sJvj2g2Cds/IW4vYR1hLYnTdOKFUHnKYRWIAMrup+Ft/ZFNfDAiHc7g+jLnFor8j
PzDN5TCMxtJXkIk6hU3pxjoruGlMT9cZ/Y9KuMtjbwmdUmkkTHCcSd+i6giZ0DcE
pAYoojH+uVuv0lRyg5ny+tmUMAxFX2hyvX9mWHp5QJfLN6RO0ZwNRRxfKILtrTvv
/vlSlQP4DTKW/+3lZKuH3BX7zY2gz3hvI93KBSHUpc8nms3v3HblMS130Pn01460
M+XOThwoC+ekC65FucSQyaDe7ZLaB6638AfMszi/2KuOleI0mYWP9uAd/VCQ3T4Q
LqLZOzRB/2FbAE580gWtYn2udbfyhQTu6d9wBwH04lstpslbiP4Vft3GRJjTiQ4I
QuDLm2uILcWdQ3Xi+096azmm6x6iqMHGHKMlOn44W199pTbrQ8CfOD1FjzL2aldx
STSXS0E85vwV4i+r6b5Un1fyT6AEYxHViNII8W+Iaygl3KC+wscoGf8q+ia9pzgp
AJGjiFbn5A/+y6xg/z39/5p0oRN0k/7aWQ6uqfoJXb28gkydDReHTN1KarfFemc6
egYndc+YZZj6IQYdW309l/R0kqU4YLLOArC6uD6n5BN3VKMGz74txpFgfPOvjZmv
WzmwAM3tv5qkKDMxFidz/0QURcjsx0we7E4mCEsvLKXLFhBJZRqqFf0da0xxGbwM
xFFctuG2dAHJH2gjrXP3unbfSTnVQWrhfFFmzrb3XgoxVG/3wHTVZ6/5IbTXuzIK
o97zlNDJG4HPQqh49HNIJYLSbUH9IKaFXheswBBTVrbMgZS/XJuDa0Tmx4P1lATd
LRKaneT46B3CAi5UlGqWgTj7x4U1QnJdA2nEuc9O0h5vZop/MW9W0grjKqR3aMxQ
+0UdFCCbCwQRQW/0npX95Wh2d4Hu1fpNsEHc0a3aPRI2AKCuvV7JmKzfflAnC+AN
xQ3D/RZPrfZIVO8o9u94+iC6qjmiwoZ/GO4igDDteLhsPvFUgBE4od2DK1Zol4VG
qPn+xj1nI7qgGg8U2Di4qziAINxlon/w1rmVZDC3TPI8PL2uoXOSsX5NBEkf/mdC
fuENz4oYqXNeRrIrPXUgIyka99Uejmkz2cVsnPVMishOle/tISFG5dKZ7luP1vku
GhICsZu5MEWby2DNqiZTVIpX17ohkEzN9WAM4IKyRj/f+kBCCq2nuotuZ8oNoFA3
eXPsdqWiWhtzKIrtWXNimE0X3bkotnlEdB9H++2LfauuM7YW8Pc2Rq/WoFsj1Uxv
e7itpJtPcFgtb6IAZS93zNPwMaWu/LlTYO1AAbd989LhkibM1wgC7MOlMepiM1mP
ZNi7RYumz2JYGZDkgSzVrXreTk81bDQrsdfsGMjlNVBIvWY7L0YleiR15GvMDskS
rgpWx/klT37BBQBJR8WiqYcK26W7fC96RpWa23PvH4xnvpksbkw3QR/kN5y44ev9
5a8VpoC8ftxXFsEwwY7jJ4wpJHAnnpdUqTVzVdQdcXb4lEEC3hKTkuJiEJmkmJlZ
UF3KwywDac2kQRDEqUVQ2GYFBnaidJZYmFwcJJInGycivpD0+J8QLUgmj4qY3nzS
enCb11okkcwlKh31l77cG4VGSwXos+jW+0yZ9Q0y9yIp1oY96q+uk89lY8wYJBwE
qeYVo7k57zorEyyaTzeu0bsVRM392VF5ZSi8cH4LAhJMPBpA/y7d6Ss+yuABxUNU
DOEI7ZNUWFCoWoLQCElbOrPwed6V7wmCPpATLcxxrf/woRYqZIwl90Py1wVqk7FK
GkCOOn8ASoFpdrRdOQOdnAdJe8wCccnDcEpmafWuJA1WcoDo0SnJ+2uFOfKUhMwi
y7iOPWLKhYAr12K4sCCUASnQgSXGxmyZNzkXKF1bRD7B1eD6ZHpsGkvHdw1kIuoT
ZbIS5AXvxYtutmQdpuZvgrtSenbcOTrhv6cKMTwbuLvynMcgxppeNaELNB8NHBlo
Nt23t1Wz6sMOnF+VDWnSE7p7nrX90bPTPJDJAaQ4QG4KWWe138ibZ5YMa9p8km5D
7vk2KQxZovsX9BdW4zlh2NN+TstWcU9HeR79deLSXBjgUbjeqbEx6jCnnsca8Kh+
gGS10tGpJvFphlnu6S0s5TbX2CilytqhnH7ElcXuLG0rRbWCjzLZANanQEWT2OwT
f/2dIWOmkDhSVwgTQe2q6vlOnuyM12lgj4B96bz48+r/UFa8x0sDUVlUczKSknpi
LgXL9I6EnmQrENjgR4YYfBR6z7NCg7+Nk0uhfdkiFh8IEFpD03s/SSdCK0iPFVHA
x2J3Heh/HA2mCzqOTML5rFzwh8OVmNegiqX4BvH/uXoYMtKh6Uc1wkURNiojF0dX
10SHpnhZ64+TQVm2uJWOZRuI+pxrVr5ubhdGBmjno9xSqPHYH3iQytRqF8mLD4CR
0POZZjjVSEQPWEHPmCgM8ownmhSJjfyEP7Ww6uFUTbzE7ph2+6eq4dwcyJsFjHV1
FwmXiIVkg3Ciki+P4cv2Rwh+sXIFzFYoOEnIPflPykqZSEAtUob5yM26MS0bR2OP
ojugYlqxsmCdXbTBnuqMTwjjB0FgvDh9kiO/6lipsRQudhOtJMawZVGB9ExC7Z9j
0knTzUSIIgXMjjgzd/GSiD9g77S5Fis0hauNjw6lMK8YU6OyIv1QqdA6dsJNw2Cc
+ilFWOfEOwdxa6XX03tb06Vjc6QfgJIhvpXGew0Oi1KaGkwSiEqjrxkYGRLL8Mvc
S3jLBuW5EUtXBm8D5X949BdtR6UcrbAuzvaD5jEAqje9pmjavPIEfLnCcAVJWIf3
OkU+s4EnzjKXygyPPkdrepyNPaore1ms3KlkoTg53oc8kNqvj82MyC4Pk7JVyFQ1
xV/3EC5a67LYQz0hC2qse1uOrP50zQ0KWWoY4dRH/+m+V9YvMgbAGSQjiYhVjKvw
RvZ8gVDotInuH2085EG1cJRiyvyLCNhCfmOHRwQG7uPUykRGMcbmNVT/KOfH+Mve
GKDmLB2w4ae3w9eCTRUVoJp6qzXnJ6pIXkVB65bHQLO7g+JuRH54aXIbmzQJa6SI
ScvHBc2fcE4Ptmht/OMwSiA26cDc9Z3TR293cIipIOACyoUjwpcfQ3RGEOcduTAr
bMlj9qg0+oLXO6q9T9Ri1URPqN1lLZmTLzwrh/4QVAQ8+gi8SMoyGxOQKNyRhitT
54Mv6TI4n0R3P5g5+DBVbHxUjcpFv/uh5YGBmUW3ifrTnOvWyXiKlp7+a4DgVjuq
WuwauZBlfDBHmN7THdilRYAQtpRRxER1FMqajhNLmm6+L5HPDT7CVqTO3xvJ/b9x
QUqhC3AHxRBoJMFdaodLhgjpq9nXm0AZw0Z5CkhhGXJRUA82g+O9iDfuhBy4XIKV
A/ycdovvcSfFnSHlNJwvlRsu7kp8bAnU1SsarjTbUVPv59kLloWbGFHyuD20JjgG
R7Z+UPIusKu/oQ76/jsQ5ZNfS6XS3nDHV5ciHPUSt45CJZWDH5PMHJHDIVKqN6zm
aeW0UVM9I9+RjLI6uf2uC7MCZmHPYmKKORNIqWKyFJeFeX3ORFX6XDPPkO54f+dj
/LOsB2vLhfwOHebqR9gBjT44pCAkrJj6ep/JIRJ2/iajcWYOoLrP2TP9D/EUuZo1
R6JGwCdR4U4OKo1e00Aw0YXZgmt/dfhIaleL6rF4oFcM5phMWPN4Rqj/N5A5LDOj
xnGDXgg3jdI7tX3dvstxRMgO875fl5gUpeA1YTWYZohd2qdMjrhUDun3vpq1OKyy
6hrTEyH2cVCZT5lHF0RJOF8TdMBD+3BHgpiPgioB9NrLv6KFbizrvUlfFE4bkPkU
EGcYb4TkzV21wGigO8Enl/iHaJyZLh3rbJE/qbn6XiYWItEZRXo0KSnw0TKAIz9z
Ltaw/X8arQV7Hpm/5hwDnWQ/plilJnRRstyKMXQzCY+0cRdlBDPJPFZHk5hikHSL
eQVEZ5WfKB4pOVtKc5nNxrkgmrIPDmBT7dy1Rc0b48QZ2sypzXr8i1bKRV74z+h6
AvCpAcNA0UE7bs9dBIXWvJC6DEWdq9nYDLi/nmdpec/hZAdwS/xL+emfvj+P7eY+
dSHAnDVeLZ4b/nRAmDQ+evw/MHoJofzGTBsFfIcE+M+22ev4k4UtBhoKiZLbJpLL
LL3HjSQBzkGF1uZRfuNvRxmw8WJfPwbcyQGdpXTM8OEuUmtLvrpVXlNJr58xSfh3
K+61GWHeDNfSktz7+kSoVJ/3zHfc0ky7VHrf/7+EZ/ZpnQXqaEXsf9bbIniiUNIa
g/rwj5qGTPj2lV4RRu8s7u8gdCwrvbn0pvCn3h3QLDnqgUtgmzoUQgcdcMvvG1b9
2ZJjfYgRrqrT/6p+wU0zjpFhF+9k2fvEloTUoGFeCHVT/Iz3LECreGAOYKJQ3FIY
0vfCRBskBZpzTBC1H+cnqCTjXrqQLuCJ37dh0+ym0FRxppMDxwywJoVwDQu3vOIf
OzgEZbAanoaMaM2SbDnvjkUbu3nbHHqYPJAFZGKZNNDI/FOTN2ObSyIJULf4b2y8
MQ3BZqPxmprCP0JRnPO0Z2O0h50gRVo+hMWEJLEqg8a96d5pk7V6d9+kTwh6lPh+
N/F2R9vQAIXkOzr1ngFccnMPOOWEmx1ZYG37K1nmUTiR/Nol8myTjN5swRunC+JQ
dmP6Uo3V47WmnfnY/81l2+TqPcdvYejHWy3s+nUkZ3QH5Am3vSE2s6Wnyvnl6Pqr
LA5swGaMDxLuHrUjB1KKILEXdfzil8JYWnkdNH8CqSu82BbZDS6Xc+KDUYY6dI4m
IkINxcBTkB3DXFeYz2Dsc4L8Cj3LQVh0rDwrk6Q/gL6BGtRfaOREIS1gBOWSRGLz
pVz5aXyBGguCBroXpuR7fhlsyP3qdeD6h8lrEJ3B1APItYpogYXJDsT3Np5J+xPu
cK5NTfOE15UfaU2QcYd/hwPFSmrXI+oeeuV1co2O4Rj5wSxUTAwGmr5J6fBF3LFy
OUk/GnH0ZsWN+QUxKaOxMYxVp1j8GCbl8Oj8CfPKnW947dxO2lMaYc6Z0WxTQKAX
qg0s7gMG1nU+371Rxyo2aAn8mzlNKa+A97NC5qN3UNJhQXtYP0PCg8lzRc6Ol3yF
vSFIYIVVeQv9ykna8BroPhWP0lT07sHuvkFwMxD9fd+5EBNrVNasyaliNNWVWVCj
IdrnIr9KBFy4ViTQ9hw/blZni2kXr+gDbUP1ODUongyN1f7TLc4SzOV28JWf/n4f
obAGQAxus1KOtgKzrkeerDkqBv+GcgYgggZ9MuCIX2arno7Y3hVfY8ZQPM8/b8sK
9XTrUL2EU7o5SNQTzdCluMi98KRoW2LRLQtMK52mAWy9igaPqEeiJHW96TtDB1A/
KcouvamZy4GhVgrXhtaaHHcMqklWPsBlVwxTpO6P2nt1VkN4BvH39sA8s8+z3LMX
CMAkkexgpN2GwcJOOTsPp8o6g/Bk+85yjztquyh5wken97/sltiwLPZ1jvBZh9V4
Pz6lsufUf15QIBC0fP8WUP03nJPdD4kcMV0VGTjE6qLb1hkhHTlYWaxyJeWbqzI5
t4h+38tMYmRAl8Ci5enwvMeJWOK9hGzxEbz95qwRsJzcKwukt0VLBvyTQ/64mXFL
nIyK93eFYl5iP/fIBRVmg5WlKbSIlp37kt+QTppi4+66yG4ngPZ2+KDC0VqTsSv2
BIDDlOH+MEowB9xqKHu+P7i5J/rFOsvhc6q4DIjs8YczGTfmfUQBVsRAXTCZqJI0
baChtxutz8WQSrQOpqOKD4OYYdl/zceWO1ju/JEqeXOndmQty+p3in32ySJR7lWB
VV9J6bndBCPmgkQqXtqhlQXyEArN4dwuOdLO2wLQoEXO1D8PofBrLqOuKIG3z6T+
ViBU7O0L2wbo/NVYwzMT+IJBCJqMdz99dT/v9kM90sQTN3j8j4GDLcv8vTk/BlAn
6B6srqGOGHSXkEx8Anegnb5MhR/1WLoO1iR4tJ1Qax8g2JNjtsNGqSc4yfqBKty7
Xnm/ahEsLVtRQUN75WXQvVDA5VZ8sAJbeR6HzOYHtCMMG9GVHhZaSKPUJ5Wn3IBC
oRFRumUe2di0LduJkIKdMukvpCuVIXC49Woc3tUSdqXcgL4yHZo/pzboN2QYvlVj
rnKC8Ni4+TACxFlXW1VniI39K2FWJpzPJSeb6Iaz3XlY8EHPQDRCllpqKXWRjrAE
wvp+vcBqAQqRVvIKW+gjTubnwPO/WRRwUsOpxli/ErtWjX2gKgilsxfI2zvMyMpS
ub3Ooq/OmcSyNxSpkOzwq30WpDgOF2q3uo03MNIv+wpR9xqK0b+s44KfrfOnub0P
+C/HapWLAP2Tj4Fk8fA9AAotmvrz6rjdThiGGVr1zk0fQs7vdFJ1Xb62VxeujYYp
IFpJ62n5ySt2Nrxt5Jh6DCilId4DyI6bWzh2ouuIHcASDeMGNJ6hh2yqI7lcCzPt
XgnFBs3zMQ9Kap/PUU73KKx6zAlfW5GuIL5tjKS55fMrYZYCIK2Cl/+Ldr6KkvaE
msp3My1R1j8XpGJbm/0OVfCxyBDVuOqOMpjCm1Gw0A6uWXvR7BSXQ3igmpLB/DKg
bk7Sg2Odf2YqEyEquI9rD0hooErc8giT4ctzOBuDXtllpvwF6Jp3QIQKEmR7pwu7
trupJioQ0IZmF8BolTNbpWEOyw2032tK1R1huS4+wx9Tv0nLJfQlPlRKRAoPFL23
Vo9qL293vv3VIK/004lT3F7CxzoyOe3VijWysMjxLWSE6DFaZBReBySgT+cM0E2G
CoTfpQKEhHQujGJHGMKoipA7Y/ru0jpLmAEEghKid7Ok1UJmYAuQ+DWxI+Fz4UR3
ddEhv345kVL/t97FbvnWbJcUsZStf9TMB7PCWvHKf9hcZrHibvmDNS2j4r/C2QTS
P/5dOqL6O3a9CD5eowrR+2IJOfvnBgrKQZVEKZaOQbfsj5p4q1pMKl68u57qjdyz
W4d8DuO3X/26chhBo/YFJkzbmW3jY4SLzgNczEb3FDAkqxdpIzPEPusNJxqz0MQT
jMQ/Sr1NdsNc90nxw1L+3FfS/RDCRWbh1q5OIUc39vi56bPqQ8OOxaD7vmadeWFi
1yqiAuG40JFgWiw1n5M2nWH1Mj5u6gt6lPhKuj/Ust6rENw3DN/C36CXFugUbthM
g8eE614cKZ1uqo8kcJaIyj1dlzAANixkI4J1PbfywEdlQaCFIj6JuVFqhit37gM1
Ut4kU2vkr7NIgwJE6bHg2gp1cddIPDWxuU7PC7OgcSc3HksGoRAdjpkWAWlRapPh
bULi8f1Kwpm+F39w0kxhUsErQDRcpSaDoJO/ete4VjzaGy7M1b/gx1Fjj3u+2Oiz
2HCbNkyPBe+AshElYHRku0dAjswRaBh7ZRrYNb3bWHr8Z/zBsfxR/X0tSNUouaoe
72oxnDZt1dgLjKrkFlmgJvEMqER4TrvrjUBnjPnILb7wBZvxrfWwys1DLU5QnWgj
6NaUR7kSPGNxW7zD0a+Qy+0JGFgwPwSme99wdqqX1Aaxlgy5asUsd6ipnawMbq9t
rFRLy+VdyuBrmMvOMNxJHNEUQ2ddqx8+5jp+82kERJbUaUL8AruU937JpeHruj71
r6FsBAhXmqFiC/hsXMwtZRSx8cUo0Mk4/ri3rUbbFCjEBSUNJikv6hhFb1YiQ/Vl
SeCqmRKyDDxAor2oYEnvEunveTve/7j7V2067JjMW6do2DEE33ppiYo4BcDh8VpU
htWHlZPl1yTK+BDudDRgBtM6P4+y+806gIHfuUVfjml/mHURI+trulKfImontbzK
TsBFWb/qgNnuqTQ3ezIVhz51q1UqKCUBAeAvPS6sJHzgl9jQvDfP9cnS8825uIp0
Tt4j7CDhLMScZsaAeBVc6cbVbxVhPU/4sJbH2yV6KbU45rnCaAObog2VK/8oXZvH
b9MBGV5MkWtZLphuWIo7NIQdUYE7hi8YqfzR3jXET9sjhJAcxrypF9IfiPYt8+8L
a0wMSpu00baGpjw0srhEoZtGrtlY3zmlw8nnmwNgdtgwb3+QlzkQqzenJ46H83vD
O6YFsOlmW1Q7+NmW8OqohJwQAiHHc9z1YaqvD/No05ByX9nwVHo9HaQNT0FGt7kY
1nEoIXIe1Zvb5A3vcmx9DgipECFtwpOSt0nnoSCsxZ8zUbq+9L/rFCi8uf64qCr7
Zxgk+VoMozwUnaZiR802aUlVFE87jbVlyr039fMox7nuFcgTGPjxQW/eUmMxGMg/
1pvT8+hKXrPao56n2OV2NZkvaMOyvcM99SGrdJ0nT89gnqKOSm9tmyd9r2Bu4wiy
xU2Dw9WmEHlHELoYMHp4KvSTdzSvNCZHUz4Dt9yNkO2utMpRmmL0l0l3taykqyB2
3n0P5ekZ1XCJ9Ny5+qHbdZ8KsrowWfVkX8B9egaprx1WH0dV2Xd96l/EkpD9OXS5
cKGECrWvp7P6i00D+uou+2TkVlWZrV3tEwd5MHuty4sp9lfX+9NzEHt9aCGf8uA5
A6iFDgReKa5CDeCO2SpMTaEWVWrpUI2A7FTK0cy99+6xp3UWhXR68wTewx5lyARp
k+lQAN3DYkp0qe6OrZzvHy/OTlW4n7cM6kkK53FrDrJd6HUPSOy55iJG+J+l1Nab
azKyeecQuCpHCtrYhUQlTdKWU/FWqefsPYODzzjAg4x4JqZAVOCPPCHcUNrIbMlG
jFjUL5CuFMH9VbSgL6iBxsNPmumq9KB/qo799H6RBcuM/gHxK65C7qLgmqBzzmH+
KqrgT5//jMYmUE9tUty2lR5hV9nGsT9phqiSI5U2Qu2mq7zbv9Qu/B/oY9Oi/Wtj
DmfSFt2L4l7WoqgZOH7qesXscxRpMs8MKER0UiUNZyMVrptzdD2/gG+iyB75XLbB
toDtWWQpgVlEubTwSSr6lLspF8wCBPamJMbQ30g6MjeeJw/rUzk2OxJF7YPcvvOa
j77RsBE7tM3Z62gz7EsbjVshaTcbKuNWVsdCaevIeHIBbSglkQH7pHXJkfl2BVmC
gJ6YJScFUlgC8dsr+V4ND7KEunj4vzZjeyJ5HUPXn/GJ4WSJz92fSdE13lFmuVUV
nIM9UBpwh35E1+qlcvm6DJ23OvwEXKoOg2dpUIE+KTp+Cjy3i+OR1lc59i17Pif3
vJcc0Syuuflt/xdW7CZ20dKAbEGNtMWJplGJIP3vd2MHppcOsDIMMpNJYYIyCyzK
q+kWq+1HaL+D08OoiFxFhoWQm9/vWCQ6g9xLpGzynodCDQyCU7tStQnv+n5GHQIx
VlObwLKnblupKnz6/yWqwlf5eZ6aWx3XBo9dklnIrVAi1YNsbZpNAcH+sD9Wn6/2
jaJZgeh43nxw8eBdHYLUi1uQ5mFnMDGFvllT7pC4chkRmp9Eg9Aed1ZxH5lJxUNS
MLIuJ+3GSGcpOgTHGhsNxGdfO4WkIn5A+tyXMvtFhR6n2D+PPT0R625yKiFGR9ZQ
xBbQQHlHxVYyppT6c+k2pbZXrP9UdhqnFxVkkd7RFzcv4pSxFIeBF2sOSr0Pqdo5
M9PLNFVJGt3WZG7EmhGe9Igv+q7nfsYOpfUizqv1+yXZoeP+wft3FeVmEnPBEEfL
cnxurS9Aa12RVllg5vYUaJiqz8WgtHWiZAbnAZVP5uL0Dk/NJjcbcbPmU5pmUDbE
ZWGUCOG88I3n/AjTGMlbwEpygCDUoydv47I2mKXYCQEcCC4ap9DNlaGXMA0WT1Q5
E3zOHpPArM2EhO6fZnPDArU3SifzOnIh5U+RJ4jCaepNU7vcW8qdRLof2hIhKeob
9wrJ7IngMTsAxVXSkIPnPIGpaPqbWMh06wI/hXhQAIRNGS7WPq9py36OaW8MKCYL
vq56R3+iyvmZjwSa/Q5tYTftuHiE3XGNcMoDdvqFuMYutb75ELHygNZpbyoCgLJ8
pLrEasIW7kBcyCRJRwYLP1o0rXIsPR6WcHuG6AWlp2JbSRjcawJgxe75ALjMgcyR
wBex9oFXDccbB3zJzELHDNjBTzStZmWN739PLPBAnOIaChhtpyBWUBWDKxCzTt7q
H+Mm5a9vSxn4VRcLwm2WdTOKqUx6sJ1A2gTfBWeDPgar/W/7lbgcHB4czHmFTJ5T
cigdEtyud8r7LlLuOdOy8sbs+woMSAlsP2bySK+H5RKLoXIcwrhwEp/0WRWkgnhn
JRAflLVhyUAo3hYYOPmmKbR6+c3rXbA22AnLsfyhoMIP4iXzwDXjh6uHJ6XPY47Y
ptmAFNyVXTYgqKebam0qsf0H1//sltRrANQxaikU9ujC0+VtKD1+ZWokLHbAbSMG
eWKAOG3Uv2AM3D0L1lbw5WXY/UWI2vwnVb2GN3ba7AtbdJCl49A5UlQIeGGUJW9E
E1orenA5FHkaSIHk3Vs9fGVaF+vx+q8MhQHl6Pb8Db938diN6k0QS1GUK5enOjKB
JNkU+LBt2RI9bp5voySl0Hv9Gqapy1g7habjmJo/CDn7FKJvAwI6X+UOfzez5HGL
ZHrXB0KEUG5XLsSw6WaWp9D0iwW6VOkr7YOx58Kg6K8hk2OzK8uv39SSqzf7yiOR
q6PIa0OwRdrywviEuW4sMA3ZBFcLis6m3jVGKMgXKwxEojSeFaKQ4HgrAQRUY17/
GIPALoKM9f6Ei4Z4w1Av9wEh/goqaf5ojpDPQwyNiGbxLkSJshhzVKRLr5TkKevg
4vkc9Y9VtTvrcuchKUyCclR5ZaGKZyTqLq70Cv0JOYNk9b6zUThxMXVI3LUdghpT
JkLYn4HJ+VXrQfEnKS2TIY7ApWlJnKwbbrAfH9ixk+w2dDDOOIxpIX2lfkTTZXcd
V1Z/upBflUYeQhtc0ImOcH2/q15kJET7eTo72yU5sUfYXa/agDE1RAw0SS07c19o
1oe5GMjeKHzTd5lh5Pg/WaXmRE1u42zuncMgBvOC68/0BP6XPmydom+3Wqh0MwKf
5Id8y4KqUu/sv5vagP9L2izOziWNxXiSPCXTxB0tyaHai+OzZcqwHxC6noNa8cYQ
T6jbgQjZ64RNuNbcQAGKH6fEqkklNlEdT8DgT96Hr5oafewhIx9AInyzx/1DWxZI
eRmYkcuOLATnGLDCZdi1OM5DdClToeIQAOMsZS+PlbOExPGpICRHhvikFY797cLx
OCapNSo2T8F9jDi1gsrnMQLRQ2JV9IzRRM9QYe4ZGhk4PctNIYfC8zJLCZXPi1BY
T62k01CLjrT9sQd3bfVcN0qhpee34byVaBPmaBLXunt6y3U/KLB6wdEPqFC+aD0w
rs1JwI12KvAGj4uEjMnu9DYhKUT/YEdr4JbzJRJWB8ZrNDbZiU7gea/hAG+oP+CD
j3N4JOQDNlfOboLL9z3ajGdk3aBUmHbJGbALTm3AGzqsXkEnUrqLOKqOJ1wCnfjX
1jPOjHPR5cDNnLHhJgN5ZhXR4//mPgBWtF3ucU71+u1xoKYvZqlf//IYgA319mwI
mwerteZuPdI4DZObxoH+b+E07ORCpTwpzPwcaLVuHzLlc9yAcJK9dcH2dn140SWe
GP8lC274wJBTw5MF3Hkri/LqxwYUaR6+1lllF77JYYcw48FsNT6NxDg1UWgHWPrL
Ie8pFRILI+fzLvlc0djxZ9kdDj3Pu4EuL4UfjiBdEnkVNcmeHvbxgqEQSaDtkcLb
NVOHsVmZTVL+TgauSi9mZX+Dp2bFyJfLuW1PKPR92Foci4a5jZF2Q0H4wUzlBFqq
LvretuORSJ6dw5GEgjTx7Qn1VkBlAdO+3H26xLzwPFtFpIkKoyss2V/nga0tj5ih
4CrzWqek68K8tkUx8WOyio/crlAyS0Tk9Hv0ITOIlkPgPNfXiNwLyM1Qghqd6z7G
lt4oq+mjjF3MO8mG3VGHnkR0dwNOEKRO2j1CQTYP4jep/ADxGMc7Sg6jPN5NMdyB
vS+me0+BCra2tN4tWSMR6c48yWWAUfO4sqq1InBNNv3805DXO8RmpSm8kuaujuAI
vZSuDeG8dRJvCYkp5koEK8GKjE7BeATKcNG+D7DE6Ps79szPmFF2BKchXfkyCLz3
aqR1LCKcDywyJ/+n8dAm/6KHU8hZeqgWDD3Tjz0RuXFQHGVpQR6OP8IOSCqzgLaF
tj9wLQD/xx7rPKLGgEGtURYSPBVWRjbfrjDUbKTUD0gwd8kryRyPv7NISBx7dQVt
6C6UQnJjHK1adRntEdZY5X9onp0hdtOqo51qa5U5DDHYcnztSbmqM8VUlZ5ET1LZ
4Hsjn+l7tWjPjbl3GmVKE655V000nOaIqXBru5HfBnZWvzhowiAKWGhReSrhmjKf
J+0/Jgd1G9SIi8KF8xy+nfiqFTQxXChJHC7zOleUbb/S+QH7oZn03Bt1/WPcVTxj
ILrKUDI1XA6LRI6NqpWfBusWHdFw+i159q2B7uk29rk3Ip+rp7e0kgA+PXM+euDS
SFaI+E/OxTzfjJZEf6AgpYcufqYca4ICVKA8uz5hdFFIfdH27yAR+rPbm6DQVKg/
/s3E95TUHSH/bdzZ3vkpv+WHRkM1bP1KSY5ACv5KZjgT1NV9cJMX4C6O/ISRcv9V
DCr2GgVmlnNRQ7ZSUe0JyQwu4ptukd2m7Pmc62lzWDL7l38NvB/q+uqSwfVLG19N
OEVCv/ZDIkh9UXlVAmBaY0YP93PlBGBT68ESPrQwqol85sYfJgL11dggricjybAK
rxMzT6Kvp73DRPCDm1l8NeEHB6mGOzcq4inEjsItdY0Zu/ctQ46U3rIIV8BvLElx
DQgSfqOelydwpDIY4s1rFdjTy0bw+gZ0RHTiRRG1FADLocJ8krwmXDC9XqPbz7Cy
dTZZSO1SOSxoNSyvTZgCTEOs2GBvLwkKD0Hoc2+U/R4AFie8ymQzmsIZBi6J+LgH
E2PcyCplAi76mxXUMhEFnn53cv+xuwtbELUmu0VK/A7hGJq5sESntVnTh18Tnjia
TWW5FEg9RDhKaIo+BET6/jaztNFo2ilxzBfFMVfYWiW7UFzWYqwPKTP3N5X/7cs/
DLIWwTs/601tFP+X3TK7W0JTayBi56vhDRfxhJpO/T64t+bMOdtq1Wv8LErrvT+2
Y3hMLbUusCa/8KwxUor6Io8aGErEd6Afze72w3pBfRpzZYBcjONajRLA5o4vWaO0
BaK0JGK5zOpjD5cu714+zx/q3k3XjuVf2ScudOHykhndUx56zaVFWgMNzpqJKBjM
Is0i/qiLk/ahOKTynng60T4rES8Jt52Y/vHflIVyW7NRgjZgXZd7fHHtJidsqe/v
Oy8UPjO9lPk8EnrKgkqoeOI4+Ih0k5AwpyTXMJcr9iVOP/XH7Tf3de8dBvT1+WfU
JTN3Lc48pKK7g/iC1QG/+IEkOUH+2IgzwVvMgvCcXZ2IBjqQ+JGPmNGB/aAedD9h
ieK2fA/HAbchiQHzLtH2P74X63200G9zVkq2FvyIis21n4Z/oLUKw7DAfc/L5BD2
m+tGZ3hxM/+3M69TK2AAkXK5/q1Sq6bWTZEDF11h98feAUofCK7oCJhMqmWtFDuS
6kLq8HMSGEGAaDzi1KkLN2fMUZwYH2VrPiskcishbRSZp1G1fov8Dr2Ywqnb5wlo
fzo+YCdQd8KImQS3iFHVZnGFRvdhfd+VsMv2SvsSCm3OXLz03+LkO4CpYT2iby8Y
ilKwmM5jy3iysJa5o0S36iP9zEe48aEfTKqtgoe7QYDEPwkA/P93XbTdIZaAF+dw
I7z9B2x6vIzstH8poT3MHCUh1Q7Cvv25s/hiIOGc0DKgJ2aVDbY/zTghEakNHDD/
x/6KZZAcy2gbhbGVGE0Qda8bJp1aWhLLrOsjggNhqx/srvHBNSRHaVsKAG3Vvm/W
pTsjpFKbmflLRRpvWamtvFmzplHjj8eXsn8tNHndKVfsxb66WQliL39gYkvX93yB
zfcyZmB51MS88fRNGED0XKwKil1sIWLUIfyjIP2PUUIgyrGgGzQ20cLWr/ZMbn3/
tjchCNx5i6K4of7j6/+Gn9GBUJ/8QCUah/BET1wZv7i2xmNA8+ajRbcOn/wZ4Xxn
hc3CWyKOhswNbaTdpqhUv949/njQy396fm95MYGXotSLErksE98Dkg3nf3jL/WBR
oIN9jPLd5TgoToGrO2nTOgYjNl/5SGhoGDCFC2iHQ+XEvEYKXAhKnKVuG4japBPP
7JIaXkEFIWW+vZbNAumxG3i1+49rekyBuLbZAWjcat+KpSkVuzu/cYdRqWW+3/6w
86Tk3t57diYp/c9rcAmEixz2QvwQnWiPDnq3p2CthfCBekNAR1BLss+DMuboPU5H
vuGW2BZFN70vUXusoofFVbh7+A7Vw2915hH6mf+LGmDV/DFLVZSAr4nPlcEsjSqh
mv/X2R/9oRaksJcla6DWzagawrjJP7tvocmdkLjG3ZHw5fYQOzMMxqXd0zRyk47T
jd1s99/VQab30HcfVJl51XjyBhNUAPVj94r5B3xd1R0z/N6++894B8S9z6oLAQQZ
5kdugr58V8nRerUAYbJZQ5it/fhZVrN6xt9QeuxIJpoUbSjm0NlvytmLIIa9+Si0
Ry8ThnSfkRns746ZiMy5TNwQ3jCAx969iSqV9nm8kD9+W/9ngQ/CWNe+QnM7y/vv
TsfPvPpGXhHPcVJLyD8LBKoHW5yr2+HmK/rytWsrlciQQmTn7KU+SidfAPUOXmJg
cmyoFXzx9rCmQ5+tfJakzZ95Z0p8SrQFdFZkbUb4PZKjatUZqqscfmA6J06bbVki
gevU0RbSAhVLDvwwszBczHkUDPV9L4IiWgHZypPPlLfXnXTEmRDTPCdO6M6CHfqz
vzNAnQt517fdduMeryPbnW9/gJHn9VylNDFBv3HMrd5YbpmS/6haJX8AI+QDftb1
zjd43oHda7Ysm19RFy42mELnGh0p8XpPigN4b5154Uf4m0TsT51DQVKNXk9zAGdV
MncKYnLw5zlfodIn3lK3Hy4jLIXaii20BzaeFNnTHCuHAb3cfsHI/ORSWMt3BTRc
g3pp0xICFyvim26ekRUrR0L4j8axk/LGtUo/iBfNc5o4QVdg9Kym/vdWnfp7bIPU
OLLP8P5Pe+T5tlIehEeSSkzIIKW0rNN1yoOa6xDo95a4MHsSbx1L2TGNqrir+Z85
ZDykduUWj2DWFRl9PxTj1AWTdB9ihRvQfx3LHH5mUPTAdbTjhtwbzGUUUROLBKcw
D7JJO9zVc4RDldgjjBKzKWd5hXEdYOJQfSCP8++vFx0R/5BjvuJG7ci6Bu9p/wvo
X85g5UU1MAupEkPYwi7MO59U0rUy0pr+Z4yWAFNCTsIeVFfr9Ve5PYFJBQ1fgIuA
F5qAeBldA2j3wgoSSbDHzSrcQ1ceB0hcIoko5iErBrsQLLSbXGYWJLtmkexbSbre
7Lpfg8kkvJ/l4HT5yzc2E1Ph6sqNoisZPBMzpknxvltHDNBggYKsvKqUUDDIe+fZ
Q0g96/c7QdZDeCy5ZjtDYb74i51Z2CHctnlbKGyv3sfe6l0fEAJtGmjhpSnj7QW5
GU98zSrXGJrQqOhuDhYtgtPVjDalldeC1UY8GpKgCvW6MxdWDZ1el1Di++UTXOaP
QMZG69i2e+Qf3AcFrbOPwely5VxxGw1bxOWKXAL9BzadvkN9xu2gzVGo/TcvIgBX
7/KQ7MMx0c0bWodlY03bhYvXRJ+vNxOj/IoF8Wsd428sEIJ0910Br0MIX9RL03ds
/YunFBS4IyHRoV1AVq5pBk0GQvoxwj1D8WDaDlHNfHb+9IxXFlE9ZtE1ze21E8gJ
4ZvG69d5Ld2yn5bRuzIzCc4/TYx4wdkaRTx+CFDGI32gmChQaYT9ZLCqa9EtKICH
24kUrXOskFMyrozfBpRlyqDO/bzp1ROrQ+hlbtzFMJsUdwRyKR9LN4OMKwBGUIw3
Ue43X3dtoAMr5RJ05si5YfYQn8XlD0w4Bvlp8HIZXG6syx1nCboYP/29PzpCAIS3
gpTTWOLHNJMq9hj92s8IEXxQ3RtvQbpzkk9L7fJB4n7Iy+Qsw97qgq7iLvtho1Ua
NH4pjv4BuspAhJG3yShOr12rlTbtCWqqyeQKwoXTPKICQxVd/ukqVQKJEhY9R1OT
hRNmCQs4NhsdzqR/oCAamZGNeoN7yfONHkUx/uCJLTmW3WKZmsQFfL0iF+Tm7tMf
3/yF9WlcChezWZ6NBvfjcxl9heIFaukpi8T4aMSOR7g0O15tXkFncgQkat/jbGbM
5LJ7lHskrbK37fCOnHSlSBXc80N2poiBQa55qG9lX3jpA0KrNeABWa7G0v0JyHlJ
ws3KF5hQOkLg66KM9dnF10DqPXl3Oq6BFTnlQeWZH+e5PAYX9ApaShv030RIgyHg
6kSPmHHbEXTWJgBzEFwlwhWUYmOIEi3jNIEz9G0hBxC3c/prkcPXdzhfocSxTx16
cfiaQ0VIIzu2yT/AYwdGXjy5kBY1kGZb/3XqnGazfMUqCxsEjeesHhdujDOCYK4H
6ma1JAexFsOUrpybxypbu+HyosozLUqDEDoY/Ex8PcLOnivRbQHERb4VlOeEY4IY
jS0Clo6WcPL/bwI/eqq1nDQc+TsPb8n0e4LD34bsLcPkDsluGGmfkBHpD1mUdKbC
1jSb6eouSMuSrOpVi6rxrbXIfrCLgJK3fwnEXFj79uu1698bW2MvVDDvP8qhHIhq
nYKlp3zn1hnLZI1w7a7rlBvDj3cZ0h5lX6U7l1Ge5ScqCkQ6A2Mu6O4nB0850lQm
9KnwIh71+YTNphkoqsbytrWgWZmLQJSRfcPEyINe0iIo5pu4IbDfjxOU1CbcVQ3Q
ncjHIe+k3t+j+mgmbZy48JB6RXcZ3XqDX37rktUkT1isBeg9Lz0uSK9JgqJENEix
aM7IzrQ0aWwKDU/Y8I9ZFZu80hoWDl71diFPb7n9c+Xs8pKRo/Xyw1FDAO8uDyGG
cfb7gXkxHGLB4ML2PQHV75xzUbDuKRUJ5yNPZICU+OVjRl3laS2Wl/dFyZOgjCLg
FNwSJILZ9kB1+lqqkh7vU43xxqlvNdhy9B1WqZxJl2sqo+HhLmEAr3lbcvIzdb2p
AXJ7uAiokmf4S6l6ALtPa3rwTlRE0eMHNwl0fgq6xp/AZLSsv+mCOAn+tMsgXr/j
lwKFLqfjkFmxB0AGr2DmwV84vs2hfyOiZov+RKoZgAo5bmE8GbdFujuP7jN5ul1Y
+/gpsvUzWu9hW4YmN+QdNIP9P9VpLryFIF/XBh1bDpQEH+NqAhbMYtKPSDMppBn4
1r3EehydttbS5moAZhYZuTbFHN3x05rOzGaErp7zqDWHT7FsdWQ/x1ZWOFYrIv+3
ChL/A9Al/IE/lNMeqAt7C6+Jv+xiAzje2RiUNDoBClimLirGmWHsUNr1LsrSPzK9
bkkPJukE+jdvdyDcbz6qynU+iGSs6Dl0YmMuMXIiuZAlNfJUPyJkqyD0xfTY0jM8
RjzIIbQVjgflwB9hkTPZRcIPk/pAG0hzvwIiM/i8VlD3mngXZPEsp/XE8S+9VIja
hgkk5Vg72jkN4MNIPrNgMTQOOz8jDXAgiIfvg+FYDJhHiCS25IPU7rAF8Ovqpcg5
d27hj+KfUUXa7YYI5tT0uHQGyoMm/Mfkf9/SdYmwSJNHZaLldLHnZqUW7Ek105Go
7+kYkaASuWktzbHzWPEqj1J4dHqDDzdye0Nl2CmjXfI2T7QNooKcj/UVNRsD68sH
91D2YixhmH9h04JMAO7fDfqptYRLXtPwsQDQp/rcuqZ9Hxs8svnBALNyNlABIhos
1MTMaueejXhrVnSSOo68Wv0UQHzi4+Rk3a9bPfkyFr9ktlpYNAwXYt07rvbeNQek
94QfF0iQ4ohD6mvm0M1JmALVHj4UdaBrp8YHPk1awalM/oO+utaLmbCnfU++Z/uY
NAebpzaNS4zGGjkPJFl8vwml7Ly1LPijmzoIqIFgxK9IzLSXb19GjyRosSTHTdAY
5my9h0gCbtcORma/X4jjf17/dAuj4skIVvs2Asuwy47SIfaqowAUwSqWVImSwsV/
tyPbOFH/666d3X9VMUib8wNGRRYQ3WM6ruTpgEAngswPpu9Ve2VLxrOU1u7wkL6C
+U7M0Yf2AsD5OMf+SxmOxy90STCBYZasHoPgp8prc8X2vkKk16fyjkj3QdNDGE1K
aJULkTRelOR+iHcs/RqE9+cS5Xv1i/sLI1bP3Ni/Ipad7I9U9mThPl45MvxvHvBy
nsXSIkkAtMlh4nRvMKtaLqRAeXqsJZjif+jVkA7M34QV8wfmVBkPfYqbvgO6toFI
LR/M/7Tl+inF20mFm1WO3H1NbFFflxWaP6pAP1J4wRQzNVP4ai6qPn6xGI4nkMiu
QSb8wUs6//UULTTulyKEF/yTY1splyXxbWx2bI/JTnhtH1P4xZflqd1ubKitdwjj
LSCmRad34YHCbRte1ALxKPIEg0FnleGNLFTyaNfv2W7qDOpFzLgmM7qBav3D25PL
1RwrnG7A5qorzNnAEaRz8owiPVhgR4hgHlLTWE+PVVw2xZ1NkVUHONzgOhF0htVK
Gkfr8FNtNfgI4UY/G4ppqBKQNk6XS6l95OQM/ThGPPcN3Rk7JfhUKEduRd8amEs6
dhOWBj1JnzXihAgZlzQ7xoy3xrQeJmDLhD8p4RVumgEFCKh61aNgJRiE329EVn9U
fURk1OQ8gUdyDtlLnG6OvCh7PxUhjo3FpRWptMQWcmdBtTbBU8VAPlc3wGjN7SyT
qx9opZfd6qGqquuYBmL9jvYnumGifeRWQ6G/B5G17B6Qq90y/qx+lZ2QplazfUDY
h7KXiQ3+jbvo6Eh93+XcLlFNq1jkjtgzuoa7HBDS6gX6MZ3LJudODW+hk4cyJn+4
S7UK9C0k95u4jZrpzc4k8V6lwFpHEGW/IhsVmwZ8jXFnA8r5dlxagV/xVgxHw/j1
VtO6PP1TDQ0hNYfz4/lvE7xX+iSkUD60GDyoPLK6vl4rj9b17Tbdm0cl+ZzLttut
UXMLihvcXAPTBjuc4OxMu0zkKARMW8QBam/NURkhZEM6L2BcHGLUpuxDd/nHsMFF
JcpX6GngqLgM5vwSPfsZ0HVKu2yINrUphNp21nNm3g8joKh+zlF1Ja3BV3Z4Qwsq
/t7uReLKm22lhf3ILzzlA1F3QcpMk6yZ5nwcEmnLSO6Rca4y0t02spLspYlv22D5
SzcmBvb/x/dUMwtH62E0B4xGX0hZh9siQz1kfveZ6YUOiZ+6osX/vrRX05pupiDs
amtbUWWUCJC8SFvuwBC1D02Nxtx4oUH+2x1yQIfM4c4FnHzMBldL2lBpEf3pc0+Q
wA0vbda1Jt7gcTYXOhGGLYxP8QG6iVyefOFmN9l7TZfuEo/W3vDx0cEphotBxF2z
tq/y0AX2CLuKk0fFQREQoFgx081hyS/7d168HROOOdNtt6HH4FDKbxlxPVczVX8v
KWrhBWpa1NalvL3W9rxQ/9kP2tm26zwgqLoWmJZYivCMXQ91//DZ2S9lQW+w5HAR
GAQwE1NCX7g2/6LQQURXqgaDe0UNVVkpnSlHm7Yz5Yg+k+JLQmZB5t6lKYMa+6/a
4kNbuo9ziQ9roSXZn56+kEzbFMzlvmpRQzMHGGxUjRg80oQTrkazOsylLPDIqZU+
gBbZOzwlNWQthoi3JKCzRgv9WSV2LBKNM8vzcridIG3VWaXDrEdZxH7PLZoNucfx
+eJYWmS2XccylZMqutwjYcyueJxivX9yQ9oshLASiYd4QMLM5P7jGRM1UQwCrrvW
JLEkcPWq1O8TXlI+TyOjw3HClQf84k8eYqObogHTd2aCTvCKh0WiLww8xcG32FAW
aUmV7Nx3ltjiSWOhCJHExJlP53u8iCQRDWATjkrNPRQcikgy8uvYu2kdTe/p/Wh+
Oi5GfDy10nNwHPg/08ZTjrhZbzlUKYe2O/ELo72RNofECZwA4+uwLV2QT9cG15/J
W3Mc9oj+E3aaE7DWo5HDVukLuv+9ZDSb9HQcoN05MBYb+7AFZcK0zZj8t2JwqNsd
3V+prRZ0I+sBBC+ua8dWz7FN+koqMlemJhiYRP8wv29RxQl7OYyiJWb8WI9kjvKl
dgk8YLe3RF5y4ub1wyEoQU300RXfyb23w5AO3H95HdrjbM1NAoOAIYC30EDgM+d5
KcFR+CP+Ef4Ezbjq0tHeXDlO8DdLZ0Ekxir9RaJxcBauEhmPUhUbKMAkaU+f3GxK
FvP1H5P7AAo732HLorC/O3qwe/6bIX3pEoSPaXKqYyk1InZy1A8i3CNknyspMm5n
itfZgh8ZhbIo17Vyo9ue7/dlIkCqtOR8YMZGLQiXnZ9fUhotXYhYSfYCXoExuPKZ
86QjjRK7+PHrK0h7jJLVt8olnAiIIRz7jfF5t13T/lz85RXHukkbU7Z2hV+Zu9iZ
UQW0HsO1oOVfgyR1ep0lzMEE3HZpXSuDm5ynWGDN+SVjJTjWa4WcmdOkLB1IN014
EqDuj5R+G8z06RE4HnzPUS98DwtTES8nuwZj2hIM+WPBZd1fqijNczhdstbGy4Ed
Tp27wz5iLwxW7novN5m75nQUEtOGGKyxDRf4crlA6cNoVgg3l8G9t78sacwTpsqG
LcNjtoXLs0577dJmp6h5by2oA/vF324nyoUQZTP9JBbH6nSHDLKmLHO9C7R5R4j2
nSebTDhIFgethwjXgxFDbVpFDg+ijbrOLoCxy/UeTFWMVbJuZCtTZvX8glIuiI74
o7a3cdpDug6MJU3ibC5sV2M5AVDvkKK5WG0AFeJqpHkooi1gQVEuADR823Ztx05H
Pm7d6yMo3esObTvabQLK7HhGVrnUeUhJvGLIhTviHE25+9IPmy67cZ+9Nfb6tS99
Yfg4hpCKUTLapXYC5GPQAVUL66OysjbU3kY6HafTSAiaUwubUKT5eiGpr/VhICFz
3TAb3M4A6nTKBs3L7hoVFghr1jX1qJHQpv/PM94aPgssgWsJxizeoz4EYU183vpW
dcasUwXO2m3+UFnJjeiqcUe8NgJHkYi/LPVdhAULNhQjcsPI48tpEDXYNjOFBKFV
H3L9dA41oP2QRN/NyUb6elYbik9oVwSWjBmPsqDpHvhBz9D2iCt7MyoUEopRgYO6
Qs6WuC/RcYCzYxW7VXrSBX3nbfFyNHpdMzb+3CDOww8cyw7NG4I7XtNtcFS6tPnX
D6dEcpDgK+29blyxr8YJPfvzZtzaE1OYJp+z9UGT6ABxGfzBXVfDt+DuGIaRChsc
dfqwoquIQGbk9C9rCLq5hWM4mEDc3upXUs5gUjnVJfvAyJIpI8RzT2NIGUE6Jy1j
H/+/BCYA/CsAED1jFGsgL5fvGChCjxskXY0VtLJB7PPL392e6NTNfE3QgVAjEmxF
vC0f8+ywKjElY9qVymKARi5Ff5viAB3/qYJDPCkRvO7tc1roB8VAzshrXoRtf81E
k3jDRODLTB0052WK3xhhLFQapnPJ2AXK+wH1km1iKQX+WZP/csljGX49LTB+D0ZO
9UoETja/G+TYiDaQxk7p7nD7Pje+s18mGL91eP95dBTv7ZiRCo9AOm5fnFL06SYz
TfizQ9+MfIev+0WmOCtNMpvLuVcQ0lv3gDnP/1QH8unsJwmqlriW1i6xES7TGehA
BNIIqQ3sb3SqBw4+pp4Q8bMMUGggxTSqup4nOMrqCGAgRaWm/oD6NlwmeD6E2n2+
Aw7+lv5Yv1OTXRHHOBksOFsLQ7jgZuwkfRmn/H0QsA7vX/CgJWkDQv4iYT1WhA/g
MeUX5gzJ9piXFuMiWlih4IgQivf7NaoPTHXfJmSTUFhjSJsUOGT4VN0byAB2GoiW
xU4FGC/A3J6qOs9MbjRxydN5ZazeVnwwGWPcSyAe+SvzFDW6JkLzVoK812gP9AG9
9yZPCTje76+oMn0T6s2Thh8DFdRv+uqTXM+SU2N13uMST9DIoOhuZpDb6Uku2wRE
/uHlhC8msJ311RCxE/Pgi+Ls4F4L3WBw+26NeCzGRnPn0yQqAn4b3Mg2lAyn1IEx
S+++S27wtO2PCAgMM9qJpoTDKTguRAlJOW0JV0BpdCO06DLCtj0yZC+FmGdWDFhF
0AkqAal+8MnbMhvwZHlXAObaHHAvnkViRE4kPBlPhE6oLCwDSj6/GXsK8I9Bjqib
EPI0ueOE3StV2CXLfKahZORN0B34kFAik3Dw2YWpiMN80VFTZvK39v7cEdwpR/Mk
mtgu4gRmuwJ7LGlbQATm0ngDOG5LXF/dPbTaiV8rjG9GJjvs0p0p79Np/6Kgzwf+
EbDVOgUA9wFY97Y3Bk4DTr2JcjSKBuvJlspTehad6U65D7Su1o88sr+zrAxM9L0n
El7IJ6BaQh6EONPcs5y9N2w2WMS/aaTTrZfbU84gNVo2prADa1LLjG4Pl7AorauM
HirE0X+QShIdet5AVDezVSUlCTGU/yp3w00YKWHkGnuvAGlxrVKR0kq4w03zgc9S
amxLQVPqKSlGND4nICLS4sTaoQS+Cto2R23/SuJ966GCZbwLNemQUwVkKlBu+pza
dEye/KegWzABl81LQwGob1eRii2864nMC2UuDaaYIE7rtByU1gsUOnj0uso0v9Ts
7AewPpge1xGfKXe4BW9fdRXyOzUH2z8G6u2iM41TzOhh2A1Dq3Rt0WSAdnIOHB1T
wjRM7U5Zz2xWQ/b1unsLjbMhmBEpeGL4oSjmKpce/vpwPa6Yvu9FRb93iYVTCTw5
NTry2LUcuzcef0NQNoLLsYRG2jA+HfaH6rnqsA9R8GnCwlGjIVhoOBBoreS8SjjS
7zpAUs9w/3o6Hno3WJOh5D10Sy97+6pVt/9nCjtKzDV1AL7by9fILfH6duFqbtX3
tHlR+8nLmYJ5U7hNTNixjRY1p+uDAoPwjdHX6BxScCsnPd3KwG8bvd6Ok1GsQyWc
IWpyhQcusoL8PqRXR9Ww2KucsSBXgmCwBLk6wKJlzZ8kTbxrAbLpGDrpfGWg3mA5
vWAg5fGNMJGzJtnI6Yrg2/Gvi0TGpokEMXi1YaXORye6hVEsOZe7ESMz/pYrzO8l
ozTuC5407GZ04bMelM6hdynhhHYWpfFiFpO8nIlivjdn4US6jB8X46QZsBJEEr6I
N0EP8+KyA1xRSEFmYmWX/m9sQJGrH3kK199EYnwNexGHlpNa8zne/24Bw5GJ+QOt
Itr7kT2EmiSAPz0pWpoTTT8wDh1SVpl0oL0LReKs16UQsx2Vk25GGDorKUXJ+4UO
8Nra+rQjsaoLieDwvzoRvM9CMFMJZthAqlRLGQAoN4pg+7dvdhMFyWrQ2dea6lKX
qCEAVi+tj7/0IGrHonX/Sg3/KzzYdcbiNceGauf8zFBJ+eWmc6AcBlpfVPTfP3/D
rq4zTlbJniBWPM1//pkE4TbxpoHWEW6p5zKq6sqC+e03NbLo5UYL7Vu1PQYL0psG
4ijYBude20b2KcjOobHmdZ80iu+JeoZVOjwsHwZ6Ih6+UFF1EAemX9xpqZKhQ+1y
owBGtnzvmFB+uU/JPP7y68R7fXyYJ4KdsiyfaYmzOWsEbjr9lhZM0lynsAUF/Vkx
Kx7QHhxAWP7evSac4hggmg==
`pragma protect end_protected
