// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:37:06 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
qtjRKVQeWAOJDhmqS1XCN8UGRkVzDy5LZcHDEB+OxsL5fha3UYlM+NMgwzKk5xOP
triVrzKO1T3yd7jQb1XVjsQZI8ryCUl77EpiJ78KE4pXIGaYC1oIifcrQWf0rcVD
LcYf8JFIRx4mi4WORbu9nvRg/TLbO2CPOvGdYkz3RpE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 17360)
e3Gbj7XWw4ONEJrG/8T0NnVjrzANLR+Mc1ETC0zw0CJX+TIlQyih87etabxeSwbZ
kr4/MpS1rnUnCKsXR/NXy4DofMXBb/YqqsExxp5p9eBXMAGNe7mSuSzV6P8nlpAb
JTQ7R0ZcD0zRh9X8k1stLHik9BK2ykLTmxporHaJiDhEypVCHZ29G/BpDZY+Zlon
1/KAZL4Gm3s5ltEaEPqURGWuoOkST9RhVSA+MU0WemV1Fsb9zdZ7Kv6h33EO9gVT
DuDvEozdz+CxdfP8ss8jKKw7yZQYIjWcHmWFXXIpVFVwsMgMkMu85gksLmxY/irN
0s4Y6G1nXeK48W9etZOPmt0FSubhZtyT2Fyz2fc5+LiGnlAM2coxlX5bwt7DEMIf
QimWs5R0DxKsPcXu1jOsuN+HoggXWNLXjpV107qR0CP3sacAxENp/6zQUGWCyJgQ
yV+htKEd7G6QNIiyuObO5IVxjyeQFW3RDf0wAnACtJ8Qe7H5P6vIgslekk8DxhkE
I9afqS/SwtLTVlzrZFGXmelSeHSwDHPnpHPM8VrE9rvHHnoJ6zshMCqe0SttW8JJ
nkgJmSS8HQlaWOf4EBRnPXiMNzwEoiFnDwZMXDnbFJLi+U72PhXktbMog5Jkb6k0
Fv1cl6agtD/nzVe0qIm9peSiX2DWU7/M0kbExy6i7IRfWPg9ztgS1UcoG+TMXkl3
XRvvSeAYPyqVb41lxOGskmg01KVIqhdn8da0iNQDIpsy6TJTeY00ZBupa/nlLDKM
LcfTBnJvRXnuH5bw4Uk59PLmN1Tt58ga6YsidSoPXk8Fp0AUbZubGABRrXaf1YZ7
vCCWjUw9OsrREK2k2HsRK3mk34p6mYFMvsX6UlYg+v6/MJhCRiUrU29EHnpmZrFm
F0u1B2lp8Mapj+cVuqHy9OQ6+uR5bItJOvHS2Yumhb+fKET5vhL8p8RfRIZsU3aM
iulVuI7qvRTY5sVH/3CLYXRNwB7p4dFmfRnL7IIxxgoPXM6rtLeOC0IvtPARc/0T
0M54bpuEtyGyDtES4MTZC9+w/6HFrcwYhBA3Tug+nPtr1jvJPFMuswwkzjH4HmqB
c+nDYa+RiolSVh5trOdzW5pMFY9yr8VVuh9aVTE/y8eOY8Nh8zOWnZbHMjqnLtts
2AXoj1aeFp7YHMJ+fIWgmjlZ/eA7bjWkFSOLEAbFCeTTR9i7xu4AufA7bBhpaeiK
4GXe3OlHRy8T5cxBX2Ye/MU3o9A/LV20vGS3/WqqdwI2jBZB8toLcogswCHYX+Sa
5xeHDGIlKkM8bKXqvYsdy9R76Q/eaDPsFRW8ZAWrMvHc9QkVqcaKUucg7G8HV0Do
1HDZI8sCtthl82FbHMEtA8oK3c1PBLXOGL7d2iAZf0yuek7NjYgRRRNh8gvz5afI
HDpKzekhmK6fYMB2TEO9nm3jfGesD36w5QHHtxQYoPvnbAXrN+2A08sdjppQ65u4
ssXsczvNnIIol9AYSqylMrxjRfblUVQSjEElwFEdN7ZA4dwI/xt18Y+naTDU7Bw3
8d5TySmtsF8IDSdKUzrRvAyFKrc+d0WpqBL6TdBsV9K5MA/jdF+mrwpGQPumQJoR
rIHmfu2w4l673zf1PAUSqp6FWPtHIxrdG3IbqKjaTPddZHWxGzV9v4yjUkny7pmX
Byccdp7BtxdJE9jaU7knPTVS5atNzvmoQs9Kz11i++Y3sZM1uoT+SGCjqRhjMulU
ZlpbPWnU5vqwDA5tiwVm7ws5Krcj2UeRUMNPvH8AgV3Bi3+oRHuBGff+OrmmaxFr
K/h0YMggDwQRMfMgyAcSOFHvPsdrmgWQa6vYBvRxgmjzEpKmYrXJ6bhhxsriMuOv
bAOd+iGECmaLjSljC0ZHXjKUX2y5pD2fnKwTmneHm1Jxam2+RVk4bjDW2Op6bVfK
pc8c6TyqWC5FE90XQbDUSWkFWyREgGCX0wxxrspG1LhmDiE3jJX15/sAbKWHMV9u
ykCwcjLJUJ66dbWcVAC3vqUaMgexRerV1lAU9iASxTFN5Df5q0b1I58YkmxpYLbN
gNm14uVKCJGpvUnEiUDixcoGUv2j74jq0/fnwQiLnwDTo9QPUXLNUsP+Gj6U+jVB
xPQ6kU04ML5THa6Ewid9mBMm3V8jSHWCgqxgzrK9VUW4Pke/PxyIOIrdZ0TK81TQ
9iz9cDANngD+hVmeGHmM0RKClDIMV23XFg0zFqvvMDBJiSu9L+8K5DqKULztYSU1
02LW97AapwQcg7dJCZ2hfXdZQWIG2a/an3nMiEpmrNCfyu6fnnQzKMzGlj7P3IWa
Oeh3CsHwIM59JqDkxvz1KMRaKD4R/F3/+af4jUvx4MPGgcsqU4YuL6yhnhkPs5rt
FpYeyM8BY7Ldl70JeqwqDV8gFwKC0hCh9ycv/o27aJ9t9ulPfN2awQE7dQd/NFru
/NfKVvIpl2gZ6GnNslSZlXWLD4qwpf7FdY6Pfv+3Zc3qvvDq18TTmOAf3saG8aKP
PAOXfmlwl2kkyzIga+T3gReTXDvkS3t6LGuNuBMXvRRGVHdB99GHu8vPd5SaPhqf
dd6ya4SGUk9Sxoz+Ev7CG20ALnO4S4+UWA/hAN+iYoo7RWPhz7kNm4/vzi9AcL7L
fRe8uz8USClkQ0Cxb0muRZh8fc1YWtJe0/QtKTAYbd3GITUHmpzPd/1xiP/tWxgD
y4DpRCPQutkYuBGjYvWNylMn3yZjRtXa/NGTR6Aff6+L8AzIA0+DBLE6Jxw9wKlN
ifOrtiLYGdnM21zK5vW+hzmABZl+M8JbHWnWU5O34qRjTiCvqAcE6IEjwauJk362
pRjX/iQ6cRMtCPKduvAElKW1KYSaJVghTTOxqKy6TF3393MYaLpNqw9hWfx4td1k
aYjveEyO5KGI9Ln0v4QqbonKDh/C+1SKMiwaggudcJnF3Cuezjz0921P1zTPz3pk
O5d+2syjmZxf1qUWLNGN6S3bPhI7fx3YFXf7FO+W7CNOjBgQeQoEeCKNZRgW9UUB
XlR7zlshh3hjUoG1VMPVNgTiwIAEuk4sdPhzX3K2gzZV/BsTyJDZn3OUEfhngAf0
y2tYO4PbRach4m15kpUcs0nNJnG6ZM7YrUOdxgJaitBelsMcxJsitWPE3T0eLYKK
KfmfJ60fDxfIJW8bhz8fm6qlxz9MRhNIUuyAAbE5+ln+6xZCjqaVqZAJvVhKOCts
3TO8MEuXxZifQQCv2mrEyJEAIlvN2PYj9JRWPsW5mgQBvSXy4IB1ZBJJhWMdrZ5A
/6Gd7w9Zf0VCJ7INw9C/BvcaCtF4NZUTnHwUSJIgMXP+ATC6fcfW0oyiUa0r2Yji
VXnoxubiDdJrgkBt+04FSZhCi+ETz1kUp3bcU4a013idWjk0J6MlUsJSl0weemQJ
wyitkyPwayyG3Ypcu/hpxg9x48ErLfAe5vkxbu/Es8TnGuW8HFWaqEHbMsLjVbsD
nvvvkoQUk20kTJAARzczuuXDQOwzOxPOqasPYG8S+gK3VswltarFZjBH230JJLJO
pVyshSrxARaqudPseDtQRjmsqIKIRK/x45ddUWLQSumukyUoUyypE0OtihLxU9Ce
Pjxs+ntiyb+ZBbPkoSIYI1OraY6vb493n83w0QP+tCgjLoKaUtkWbK4VNfWHO6iW
BTa8za7H9x9HGlYPEy4mVuYJZyMcoVms8KHoaY+alNJNugfLvUZ+Kv2KDw1SMmcR
1d5y5WlbDnY6dWO96rlYmZ4vSJQslcXgXErkxhcai0F8D1sxI8PQAowX8BSfd6UJ
7S24g4VmdDoo3X+dblZBpN8QlHz03PcrlvZqp9t63tu+CV6Yh+kkk4Mlkp123o8z
edLYYtADWWz/kA1mtD4Mcrfv2ytn96ybsERZxTcOYKGNhbVghCUvnPJyzt6bz3rz
dapm04WnitVbHL4CnYzj19j9Qt5PO4uXjJQo4PZSsysrVrpQuwaj0Xh50eW+lUss
qSW63zFtySuSNrWzcjRXir4ndfFNA8CrhBgpUcAl28rztm4dtdk/hHETMweG8LEr
78An0Uz2vWLbwSaHQDq0WwoNR0X9/bBbOBrgCXroMqfCIaEjfpQhSmZc5FMe07Pz
PVpxLmTLUpPxBImGP53Ypkf/VJMvV0NImMaeybBvncOaBJzNpGVfuTUlhT/NbTho
QPZYIk7P6FPo9oUvXnh5ZOxCpx3+nRyJAxv7sIJjGyazvIET7k4Vn4sbX/FKgubJ
gl+9CeIIcK4KThKGwpUAS/mVyFEAjDk8y6jTUkc+3XRJSn4VZboVQrlG2iAv+Xzh
5oFUdlniHf9ovtGngIuPGIh46XyTWkN/Go1aXANWmeMCR3anGjpn1BofbHxQlYP+
BThQQ2MHT9JyPUN2MA0p8oZNyW+5UYJJSZoQdZtjnRdht8FCqpTAa96An6U3Nvp6
Kh8ZYcLQ+o8fBftQjvYLQMpZS6YVUeBLltuUXdy7gFjx9Z6lU77fDyRCrA31z78L
o8FXx0kN19MKqIVA75I08dykMC3UTG4LnlE8yAkx9L7Ukwpjk/3GhCqbrtbw1uHR
xVmaqHek+0HD928xChWCVbl00sFBVWwJ1bkQZ1kjF2IxYe0k2x3zIyyNgeE5hoqw
l4+gJfbiylE4d4DC6DJjEVCXfRFgjWim7HR1DcBwt3Y9pY5bIJhVGQp+nkGMlwdB
B/ld3qh6pe66rvIbrKKgfATKog2Dra+bL1vu2YOsNBtzJf2O/5+pX4s6fwUhdEs5
Y43/kJUIG4K2zo8wtYMK02dUfZIH7HRFvMUbPRpdHryYtB8OPbzTBSInuJ+p3xsX
orTQ9feJjfE6KdTD6xakU6YoPmemjuL8lcAm5gqqiMdS+F+JINMiAMiJsEdTu0Qa
DpqZl+akaMVB8PUZK9UflNWW8H+74Mto+mY+FgnFSs2HXspE7llN1heapMDv3G4b
yrj6/9RaOLmS58tM8sRcFuJYGI/jEdi+V+EbpeEQXSCI6mD3J1OrF9OkzGE8PnTb
So5ay0Sro+AguuVFtsqQ1cUmoHH0qilxOK8CcsUSXnLRcSbg++jBc628m/LprxGi
luddF0tMPB3r9qz2jmDAdgaovxtZAWmF+eu7sDESoKjaCVCwEZu9Xs1Rhec2LdRO
9ymdHiK0HrvrsSP5ivVLDH96Sjl1QKc8NsHMf5kVWELNGWzGSU7/LY11zjUNzNT6
SpQqhWn3ncJ//cDJ5JZMeGG6WlBdK6ZUa7s10D3fFDD2gMFbP8MAcADznk3XCvAW
QY7F/1K/jzscm1ig0FIj9olUs8ShkvDA7tIyVXOF+N4mrAKjH8t2trYtrhjlYMO9
wQoWewi23nF1bvOu2PJ0aMAlxPDoN+U4Ro9ZVRv6I4UVyGplleielKypwZJoi5Au
1WYtIZb806tsmo9Rh4Prd30rB0YF12+r+kVnFSk7Ll0ewYLhqViTbh8DIfvi7cEj
PIPxDKRGoh1Wmv8zC9JhHX9lkOcUhSk2rAtq6bOjUS1TUJnRI8Gh3DGZ4zqQfphK
2bNbO2ICMNESLZHqFv27EivUB2h6JhRV9972AQSKQHIaeDKatVBbMxjz0fnkUarg
YSSa5fSacIvp+IPZGpVJDizG/J8bWcC/TiwEDCt5LezgHfOYe6w9lD12PvFgJLvG
VxhAND6mVDzDUTE9hB9nDJCnuAkmrgM9sqzbGG6sttbS7e13RDFPJaAwzgJ2kaXc
RJoFI1GxVXUd2dZZEU3Q+paMSySqHgpHa6VhL5r09KXd0y54hpcBR5ETKspftoeI
bYHJtyQCZNVG068fFBuviZlq5r8y70BbiCbigmEpZ0sc6EgduT8gvkYfmdkTK0Ls
O4oADm9SIUCNIl0hUFbGXHdUd7mpFhi6ZdKaz82ZzcjwogFbhqbTaOaxvEDGH2FN
XgTjnOzyvLA8N3FDzzuFXIs6VolJXhDT+Woib2WTP8bB03B7gjPCH0FFSLQkz1Aj
I8n15DtVO3ntn6eZDVahE8G1pWKyMreYzf+6Bcs2ojxzHIusqFmL8gDOjeXPN7/1
9uPMLi01iAnky1XxrFH22mM+Lai+frH1TQLt7D3TsX/w3jAyrtbp8Kaw+6M2/2vQ
Vz4CajtbUPhIKmz30MVAj1R9++5vFCeZ7auyPcydSaV6zxWalaQ3a539GkKq/Eea
/nfi+HiKS/fV0SGpdWeoe1pIDNdWtgdCXfF3U0fb421qMa4ZyFHEM8sBdQwc/yTr
Abb6Xk7BC9lNSV8jkaWK8WA1BM+9MWdSEybObEGCK8+XM4UpcspHAZd58POqwS7W
xm8HhRBfU7levybX0R5m1T7d2qdiNWaJMELhxmwmJs3qYALZTtssCwpbhWCc23R4
kR1C44lrqiJds1p2cOQ4mClmLf49TdvStDnsD/6ZQuXhHtCfOcwH8hJ3LqCXZjtO
3y+HfsRIDF4rAAGvPn2liiR2diZvZOLJn3iCVt3Bv8wLlPnongYb35jneYs/Z93g
Pqb325BesaBaYiYkzMFZqnh5vEO0B1xBOy+KQJl5IZYP89TBgJlGa3Q597MiXWj2
grbTIetfsaDPoIhH6lYQJJs2zrfmDAiyZVoCQxzSm/lW6nKhbESR+3PzWQk5BfhN
1gZNdVQCAbcy6ZizbUmuvX52dWtpyz3WELL4FFJQRohvOLzVOkk1qtBjheqzHA/C
of7VBrPWXQngmD7cty6ZeGf9x1kg1rH+N7uMaXGdwigy/2W1wWxElOAmlTjsEJDP
FjWaqC0nT2qqookDr/4zhEQWxPdCbHae0TfMPulTtiuAdoZO9JWgr2pv9VXbMp1S
4aL2E6Kt8/entcS0kGsthAsgD/MculFywa+dXL/lBoKYw9STgTovSxjtHUuPF9x9
uiU4lCGWb+ZrYeD7J5y5+ZoldHPVsh5Q97GIQHOky3ZwNit7wRGHuU7NluntX3Q+
taZURb1ulN3Og+dOFL1rZ4dXu+6miVXHBYwKCKLhyFx4OnkPDqOpvMfMkXx4Zwhv
b/kvpzSbaY2OwLFYEGegNst9M3dvV3nI4BaMzwrS67frt831ZSFFRZWNM8V7PcCP
EzoUczCZp2v/JtfhlCUnGQHxrUMWdOfTHaRb80djCaLegEktucXhCwP9yo/URA0f
S4HWYT9KZPsV/fhINkM3BcPp3n/VjlaFAeGPApNZfBw+OEyG8+kpkuwQfUvfQsKm
bpEBdI5mKRd15LzkSfYh3qLGMY0Hy7UaKfHdC8aOZmcpzQj/YCvBsCvyX7Wy3fZK
k8fGC6XZNapsF7tGWFd+77HRyTs9DkR30PjBqg5QzrqZLr1P2btBK+KAoScHOw2a
OU0V9QFA37qQhlJDoUZynWP2IhBD+dF8iOZzkgec9toINTAJygl4/D2wiDjGm2jd
AJoTjhHUZ+xVO0pF4BTuG2O5f6PDLGiu1MCj0iUgDUpt/avC6N/HYj2oqrjdIoeq
zYP0BwVsAKS3XihKobMb9/MKuqjVDs0KiNsMpsXcuvdVWjGCWwUDLWI+U8/qJ5go
xfzU1w3AuVkQoDcLoMtjmL7n6RTx/CpHUBhSA2hMePX4C687dWQObmHrzOrKr+Xv
N4IvOP04XNrNxTfrHg+bwgnjH7KnL49KStiBbOAygOkCUiUUL5CxePJMPUCgPyjF
MiPdrR6dchng+McM9ts5U8W//32BTcWnV+yyhkdvEdv6/hkZgtNACTprZy6W/j7M
HVBq4YOE7d5K+ERWFxKhSRwD5eOv9AKn8MJgBIxxEWAF21E7d66qG48QmIG/2y4r
Z5brySKfRjsTRxjyB5DvXGW90Y8n/tuZM1o+qSXB24ukoPMHGYZoqBygTvABYgbc
Y8/CcvXeCUXOxQx1/XTjZMOqQx0SfTxi3Ij4o3jX9RSnuwYmeU2BcZaTvRx8l8Ep
1exmKgRjUWAnyD31HsiQeI8UqCpYRMXVB8GVBWRles8KXvqr2G5p4zRhd3x4eC3l
Vi+QMlfm83iRERSAST3gGoskLqYSHRDSclCP46MFbIXSmDpan56qH86pXhZGZ9ZE
XmBTEGSe9Np3yjyZuJwNyPihbXCt/bmYmavmdZiV/UmyG/WXbTrDtpEwWwn5YSWM
eesnprKDE8mqB/kUwo26q9KJNfDF0IkBtyKCzFOLBVyiktwd4xIM4qT8Ncx2/O2C
eHoXo2hjADoGwWk3wVi1heYBDzOLz5RT9SmLdTbvFHSKgkZr45Ge0EJUco3pIBu9
YuKhMGg5QYSDK1lRRD/qrRBWVr/AltrBu7nMmSwAet3vEJOXvqpINSRgwaPqnNKb
Kfq8zJntd36rVOT+934CVEHSoL/I2ppbuOuDYD9rid/plEXX3d3rOBOPby+eCdmx
YY08yoyx6K7Tj+wwpTdAY6AWUeBlW9N/dMevvP1VjdLxNyQ6GT+JrKBbAeRmZWtf
RFY1RV+rM9Tqd9Bib+euz/RtUPX6P1t7VdEH8ht2fXiT5yTXuKo7cROL3IMpyMOU
ByIF0eDOHCkqjMYNxoyoTBtt1n8jPFHgQyKrsNQsi2tZ+wt8YAEYz+55ZWresq4J
IDrG/EWolP+v9223Ezcqsa2Ui3dVJDhwMDhKTS8fIfbri/du6LlUN323sgsIdnXU
IOhhxSWtdhv4g4uhRZmHJo6++1v9Dqae4t2qRuGE9+6SYPUIUe2OePwVLMaRNAXh
Ps1qzg4E2RwJvOnwj2QItvosMIHIBlSad5+IxvAXiyt+7GW96D02R4Oq9ckBHhEj
fUxBrmLDpRoy4SQhKiNc1X2K5XtwqrRKjMgCMgG4CCRELSizH7kzJh4NSpPnX40B
yq3Xx/9fwm4PpupdH3ULL+uhJmMRjgwv0tu4oynpRgXEt2QWqcfUDK+eobOdx/tf
S7xJ8Q/vifBVxfSoCb19GcuiUPXgxEnE7g8CPA97YF+Y5SDLHfG2fmUSgf4iRWm5
/o6EsXiVv8ANVemJ+WG8dHFBxomgKPrwHQJuZStSkynlnahZVqiV3a4aeQpJpW3Z
QbLWlYoUeybp3p4bhXNhBEh+eQj9jl6/4qXfPHvIgpjdPwNoyUq4YOHtK8HvzpmC
b82QYIKiiwsvV27ZVlBJUJLtT8pI3KT+/gSBprYo99/bbrbaF766mqm0+7AgkewM
RchwTTbrb6k52BzLYPCMgnjx7H9Q+RXKhaNT6WpZXjChrM6a/nQCLNJ6AwglD/pA
0j4DTQPqwLVmcOjvQHUst4ehxUb9QmQPI2msaeZvd4gsDEV4ryS14GpMCYmHBuBH
LQ99LxiCyFbp520mezAc84IcMfz4G7WY8yFgl23bs5SClENqskv4PCNFgMl/u0Tv
VBcQoo7ESia38CULfwlce37ArWyPHyNPzzthq7ll7Rh4ggmRc+0nKqfu9R74/ipF
ZmpYh4EYUdgmRK0SVbfJ0+vMRanZLj+eviRAnNZxQKy53XMjVx9+GM1Vj4qXfGp3
Id6Y5ZzRR5TziKiwQtG5Z8fdwz2DUT+prE6nIEUr2bUBV+jBEULjamFk4HkUgBz3
FGtOiNYcRd4f0zew5NynfgaQw+nsiVmq7nLS9u1UU+UKGoXCt7JjjAchdRo4iHYC
N3mvCm9lJHXGjblwULYwpKlQ6Ab57u4GmMg5fYz8qIH0M+Mma7nZc5DZT/IqaUX7
k4RO7LVEcQjMGI1dWQDHT2/Tv865g8vhyz4+qvGON6EU1/GgBSA38MOo+/v4IZCa
TCtj6a8o87pb6Srmac4SDSHjKDm/udjY74XMtQ8+x+snhxO7T6lIZqGMm8C2XUma
2ochVIi3xd+gKiMyJ5kKUuNN2kgTYT6Fk047sTQgzcK9+RZiSfBxaicNsw9WJQA3
lq2EA6qfwX5zK805JGb3rzBpvuJP4xSpwf5hQbksJ5MF+b+QekcNxi0XV8GG/XVM
hGeKrZoq1GhFijCuV0XhvEKISMu+nXB3jLo3l4PgrQE1jTOTNwIMInB773K0mKep
bCLYOytqBnl8vJMxn2K8EQaxr5AcN80/CHIFukaOnU8n9phqB5r7lv1CC8GWzB8R
eUZLPM0JcsdGn9nZ6lamBuoVrwaCtmExPVbyIEcvYyKrelvOZ5tiYbcNw3RAbpP4
GqRlfwUWb4JPiuGnXmrERUsPwKxLEPfigwJapKXQCSSGPUfL5dorqyz3K2S255nJ
5XxWMTSxfVjV4a7vsEpKP1fbXII4RThsf0xwQ8/UCvT+hlz4A3s49EobB/mh6hfZ
z9RRqskLM07DTIxpKnqhg7IF/h9SIGO3/6hrOXpHLk1KcqM9T18p4OYHLPVNP0UZ
ul7mwTlU4WfbB8fhKcz3SMn4LOx6OfBKvgIxV4obozI0Kh6Ynyml6Gf0P2rLAwcS
IdSAI2eeFiD0/MIMS/6TQPJLZe08QbJDnaEsUMBenB5dr6U84UU75XczEodeXcws
AZcgzvgzDWzA+9sN02wFxJ9KfSZUmvhfgOCs/iCGJKyfmBZwK21Uq+ufZeGF60YF
E2bURtx85+5Ue807DhWRwLtPjF0fU9Rh2Z9G9IS6y6gUxQMVnyc3GqLTgghccKUR
32e7XEVxfMoI/HYDGgIO3J/bfhc7SGD/8l5n4z8NTbkZHR2HPO1WsV4N6VtPYxhy
KDp/LWdf/BDKEPmkI0HzCE7zEL/fs9vsoOOB/GSAl509Re3Z9jiZIKiPwMLMiyF+
vxLIEfP5I4KELsvaKFa1Urm5Lx2ydGpzJ7StuGklPIo/olehI4j2/PaE4fIhPP2C
3dbNiIWC0d8B0Ye9uKvt30R5hBsRYSJgDr2mXND8A5lZbsW6sDVMyeHNeklua6su
AIlzYE8JaAK1xvpqyePzS35qd8NCuPvDVNgYXDPl8lXZIVsaFlURUAvbksbZdRr7
8GvUSN8XYIg0v5mP15LrQNjuQVDlt4iT4nsGckMfzu/PyYW7Irxzu+g2vlKuMDeG
EX8TTK0ZmZVtDlwkcj+QdLm2SGaKXKS5gnwKAMja/LFO1DJdHEb+U5Ym6TDzUiRD
z3K5zYHEZ+xGE/bG2Poj7+dpbdBgAzJ3LoZM/Et3Xk+ulkdRLf975duze0oCF2AS
CBlTkp646VS8smUoOrKcShkkdIDGUl6yZBcAPDEc8W1fmrTOiYwXyFX7OYAatBKt
HyfwglkBnf7vzMqseZN4Enm3eHQotQdl5g2Zm/uO5wV8ssrPtclEQfrTt7o4UV3d
/M/njno0kXgyE/Mjh1CwXiQ4dST8SbYDhu2SmxY4TMJIUq4KvA7ZvolQvXewo0H3
a1oLhWEboYhdq63US82LHGECwPPRXpkhTygBVQO9CvjRKiS2UdIOazbgix/d+gwS
jXfe/sNnr1Vh09t6D/ojGg5kXh8FI5hEGD52lyRmyQtlFm7iJR1zQpZJiIpHcWKr
QxWgX//pT16LegAzW3HrnqEYlDccGYevIje5wu7lNua4IX/ku5aF4X4a45K7duqu
9SgZSN/ug7gO80HvKGYxNzfTUNMpMCBCvIWH2/zYuaFnXn7/wj3ps5Y6sed+gLpm
b02Rwgf+y8KoE8jHHbWYa6CEtTc/lRR7xpnjQ28kxiAb/tpw3l/lSUT1R0ogz1e4
F23nUkSCBwDksUh1kE/n8rHFKKdHN7DuGIO3t33H7d/3YQ4cjn4qWat8HBmfCqz6
qZ/0QcI0mChOH2vbH6sfjeIZI1QcO0QXsND5OWw0Mk3oO0gfRz5gs8cHAhbFt+pa
7m57bFpsftrSYCUrzmpBGQRcUPRFLK5Vb/iI5+MwXfa7o/vXSvkp639t/fOgvRHx
DGcqpYnditNQMCejksqlrhNrS2HjlhpHr8k60xXlALd7uviumFIV9XJUoNpeZINH
x8LQjmsFL/q1Ubry6aYdfVYiGPBBRE9TX0Glk/fPmey0POfvW+53l71q0+d7amlx
tbKuAG0O5wNd4PGqsG60R6FiLJSh4pJsUIVjGhTAq/G55p8Caa9G3LAo4cx4mtG2
C6hdBZkceg/uLHL+3IBCEdcjb5auSzIzV6Mm/+1rnz9ZwUEjlW33RKJVjnA+CRl2
omT4lVQ13g8HUHCoIWWruyD9dP+4rLN0uR2XmO6jdf6kanddSt/HMXWkeZT2Zch8
7boG0c2pxNpdi81CCWIrMHUy3QRaknCyh6zdF+8R23nLTFIYTbbpKFQgr6EyjApG
bolSQMkWelKSY66ce+hHGEJHqRr5DGnynRaSw9hHVfF5iQYhXjytQaEWfOGORA8h
0LGdy5tyhYqkfp4BvttMkeF+rs9UC0mlFnr7SrYYqBtn4W9MZhHR+YwYlVxf07wx
cHM8N+s7m5aJbWsqw/Kw0ltDw6lwtlW8wYES9UiQO/mJgnbGFaMkJEGX3NfPMOdV
ugeuZO28xcqeGnXfpAKu/1XY/A+QWzsG+RZkKi2vkZKZOcdO1A4Hd8tsjgM+usar
RezvTTZdY6/ajYviALTKSttrOOizJaywCVdbgq++CMMbUqjchP/JZJX6MHCvHqFN
moQ/xKmn9Izs+ZVJ0NRPUJboH1top2f2t8fVNlBwIkNhfIoGvOAWIw2OhTHnxP3I
MBy6m58PkWfoOEzxEyskNCCFIUqenfxBnUT7xk9NlaO+Qitoy1o5bKHSE/dQMWnM
T/BSj7ZcCpuvZTGi8LCiayNLLpWA65R+AwMdwQOnWKc984OmosJm7m76l2WcJE12
ijyuOCNXTESHfOU3pVwXZvL4Xx9wUuxcM700soAFmszQZL2m7VMkhgUM2VsXZBxZ
CXH5OqjDZmBhgcK4oPplRqrBYmtMqBy6RiIVGGrSKEx+ooUFss5DPC9IZjD2mrH1
kb1+txITTOMovx/APuqjRmzSc/emMx1j05Krz2n3m2HRWCQdg4tEiXL/JLDvbJrQ
LRiJSRdT3FOtQNSM5WkmlscAf5F6hAnrzMIKHFKvS0V9D+C9ckxZjycLa+AgsZNr
3jd5vhS8IvJBupajzGmg5+AmpFKjSbl8VTAqxHE/V/vRf064ynCsf3R4eff9hP0A
Ys5+gFY4pwVjfxzxnS1pTk1QS6mgd6h+kw1oiDGwnBtgqCX7TTZGssayu6fGjdOe
gAkrskTWI2AG4RpZop5Q1h2BbOBOgF2d2i4e2cnmZhR0U3UL9ih72W+Udxqdj/TH
Tq/lvP8vHF2pqsWUy748sD5PvlMmtpaZzmgAzZtwfJ72XA9kKW6R665O6pdLxMG1
xc6imEhaz71/bNZUlSTMkAW0OoLDLgjK9FHUbHX6y5vKITnCD9r32VsZFZ3Lc3rB
YQWU37s5HH4zXXOoDk8wN4Go1RozusgINiDT58zJzerN4sDaG7MmkObQs+w1k8hd
1sDE2ylkjvHIrFXl2lyRgo8k2CVevrCmPmwozExSB1lqmnQUG59t8E3v3sND0Am2
xmhRzbhCpfifTQDACp+MUZl9DPF79BY0eJ1IKyyPm1OlfFKbF0knWPzwzSzGfBd9
j7EHJ7fjIPH169Kse6eQbISjsNl+CsO0ZDlEN6bqXSz81FaiOKJmInSwf+k2NWeN
ac3jXp+avQSoFzoCcQ2V8dEydcKkSH9Drg/WNfJJlSTvhSVI4J049aPpsvhx1kF2
elFN6dN2NFb3gt9FuiW68JJKjsSTQ7S+WTBO37qYd2pKwQUajR3B5xXZQ+htu/fc
vb/+uDxi8otfDBbjor58oPGm+p6/f3JXzZLqcD8N9rRYf180rggqzY3iKZXLbr3H
O3NQZyG/FxnUlgrXf751yAnjtK4foRI8hMVmBtOwDAbe8RQ1DtUsLF1ZLzx1/Wpj
6NdHXycXDIGpMDaduycGmxKYfO75VarsKIrta0JyD6PHf8FQ4Q6K5GwmnSF7NaNr
G/AM7EK8aPmiUXxQI275XMLkSgzXZ0GsaqDWJZrHg/kPWOmuf/D8bqbYAXBRCmdl
lLxGVwPP4eeGaLMvgTDmj1x0AoBOcLvuRBPbDW+iVxQPjJU9Hu/JvVWfNzGWMYjo
vI3ca9en8gIYM9YnVhOhsG/SJbttYDMuZLo8awjWPaN9SaN1BgmUK5B12AkzVi4Z
Ystpv0P2uvib59O9t/Rtu21FjJ+ijAa0yKTZsakwyFl7R0j4qhEDdj4oNHcrfqbX
8Q3zPcEdhuq3s4Ut5nN7YUX5MlqrRKITQrnf2XURdvG9Hm+YGLw2uqg5lxP5GNI7
YwBMemVNvh8enBIm9Wc4tomjnSYW+g8/YXSP1nKbjREM4uTaRS28XpH3LTgz1TDp
5Pqu2QBk7ViDjQ8ulEaG1WH/v8oHUEfXlidjdrQzBO+1DiAUC2l+8e8yT+H16Tqf
InC4dBsUk6kdyygK5SnIU+LwnERjJA4FEVUEYWP0FThPJvetC+WQLuo2WjzOzN3r
TZ39n4QxxeMsjEznJntkLLvNx4sSZO7nrWVPmIHueJadVDOPMIV+IzlqUCRFHktl
yl/WcY9J9iJFZGm+3IjqvuLeuYTkK/QsVbxDY9RiOoBwDasmaiQg8ZBKOLqqqnd1
HO2seccWghTL/sVCCf7Ex4L4Gnew0eeul/8dvlAblk7wCL8ue+GXIHeiU01Vwl/9
Xa8VCdFU9WHbL4eR+W7cZtSI0Tk5Jp7OeSiqc6W29ezsCJ1emPlH9yJh6aKz0lZ3
GWUFNZKFygPy2PhXFLSn3E1MUtu4Q6AD2V9Wx3Gv3J3aeccQ/JbFsrMOOS7J8VOl
W7Ae9kirw+b85JbatGj2xf/+eN8P7G09foyL9VEgyTz1smr8t5QGkn1/a1nJUI7P
XzteaTruUHDqrWXdsOhtxot0DXjIJ0UR4OOZRYF7Qs+upc+L1eRuUu7+GJ84TvH0
S68kKPo5mYZ/HvR+8x7GJoXX3ab7K+imI/jfT6n8B8MTOV8f65LiHupqwQv+kpy1
WfVSSnE7ZkPjT+whdvO09CgKCYrvh0OSvRxOp8fL0v5x+DLpt+JprJ8ddot/bC5d
yIK9nMCir2I1QRxNxMfoalw8Y0g5Zwa2+xJM45shgFaj8SkL+TtimUAF7NHYZYEw
NCwAnKkaTp7EaZDFxNQYB6wfbH/ee/uiyoZS+grdSsQQLNzgjUXOgmr+/S+8Vd96
3ByBZxuHx8hQWERgeow7ipwX1fS/b4BH1jXGY/MCaeJWtIMPPoXOkN5qrwZIb87E
ILtkCQB9TMuODwiy811+VVOW4UfEIxk/M4/kgusz4eGWou7RPQEdUAQ6jjc8DLUt
VozfPmJozVOSnTxlWDCJsJEXNW7GIzdS2BCu3bMAdC6dqaINH6IhS0ZHSUvtmFiA
g5pmRP93BgDarBbgYmPifm+44y0LjFDCwhuDPzoxJOix0jhIRRtrP1Y6MPxp71lz
M7Zi8AorMRgyZPq/oEjn9KA7DQtVYokTOXSN/nt06tGQAFZm0l1C64jK9D7/z2mW
8knr8jYT1S5aSwoANp2yUdYkXfDEE4Ix13LSR/ghkvwD1wESChs9a8Ei5bqKyoWW
mwEJsTL+f61mcFRussqVEWQxq4/lFdFnKNa1KeMpcxLmbZ/IgdLUR3letOHZROPW
P5cO0WuX2KDJlyAS1nDG2nlTbQAruntMuiRTKkUZTbzXdFuMwRUOavq6OHz2fhVq
bNfAR6t4hjLZ3GCDXfd19+k/Dr6IXZCt44MvG2RDCEYMDGyzYpr2EmUqkBAegvJm
x5U+djQp/4U371iaGEf02H8O4zQt0nVMHa+bPmTo89GRkeu2ziuvYZNPqrrxGVUz
uzzpeXJDkMRz5gBTNhpBUrggjx2AqKd1HeOfDCnVpfeeAtBXAAV2OAlpH86axtUg
aIbO6sJec7a9OG/85lxLIcYfkq43zY+a9nnzsU4UMLr8qgHaDoXEN88cUUqQfvG3
Dhi1bwYLI29209NfVDCnIxYIw0qZEcwIYeWO4KMxOo9JmDiau5Mh6xADmCzqVJUX
Yb6xZVhwn9aTwL7nHyCMWVihoYuCSESDRE7jIwTpQgVx+Y1pyIG47y4k/HgWX8GK
q7lq9IT0nLkAy5NTD1jYLg0VcXKF1kahzHDhBqnT5tLNbKil1CLNKIt0cB5ImREO
2BbhYP+UTdFtWFfTWrS1APf/HbAElBRVsGosMH5x+h+o0GZVDejP7qzQqpoBdgT7
ewojj+W1vGSKJAU9wjL8yoYNb/P/f21VJk31un2cf0rTIZPI6GOZvXk/7oj2e4od
27T6UhKJ4RWB6U2RagoV0knD5kYx3cOT8NcmhgaLyGrKPwZ9W8M9djZ/Yf1xTc8w
jhXcvyyqRbabb/PvkLzDquA2VCE/vAC+olYp2taznOMERNGv6E94yJeVCbqh0ogd
rhD0iv4W72SohEhsVK3omhRTkQM8m2PSTfsHgC6drUanKwM8AsQJtxJH/0eJcKjU
Zt5lT+HHMz3OgbJpyw/Tjhni8b/k2cy30+7i0vTXMK2az5J7m2OKm0JwGLE9qccJ
798s5F1dRGGX8tPyEp7Tr7F91aQHHu+ZoQc0zC0GCNSR/N+6yMVTx7/BxaBuBfCE
iMVE2Jn1vGwf8cSJzCPcrSyPEyG5aa9wDPXm1ntyWRb0CPKG4+oXmOBIkmBYsh3l
dZs+WOYMFMW0Oz6VsJ28xk19eJDtgyxtJ1W59Yc+oXaxx9Jb4KY5gcKJ3pUtCQvz
UrLJWo3ZShCKucq1vgrSSd6SZl8UrdG8Y26PqnKDTqWtmp1fkGa2rQxLzI6W61Ar
Y6kG/eFC5nyy0aKjRrHIcb+gXJ1hypeJcxlasIB34ksioJBDRDaSGhPZ8tRBtsvP
oCSTwCOPvDHIf1XGih8nAzFklYm7R5O+et3CkRF0hE3Q588tHdVc/fT/XOhLiEiT
PkHdQcMaQetOR0mDp7M0r9N9UrJTLXdPkMdxltdomK7+HWtsLOLFDETUUoe35nCk
Ec+ZqhN8iOntm/C51KQ6J7b0Jf/eMEsw3UyMrBoBCTVjgwJXBFtxts6J3jQIn19g
CXf3lKtq44aOp+gFaax1L4hqameJLpNtYE2B1Bere3DDcYhysZln0lSifSCmC2vr
X/j3scbg6v235ZyROAbLy2ySnIacPmFNBJ4QltAmOa/iuh/HFOlXSvQqCCRxWess
6zFLQRAcXeFPjc3rNl7PYBGh2yCbHGU21HncEQ4ad0ED3hc6O0pb1yPDQ5xcGqf8
SZ0UM9Y9ZbfugIdp7qiOy611VDJPBOgUX4yDceqCDa8u5o9a6e/+BfqiIluupQ95
CI1qk0kpdRRlmsYiXvU+7m7kcmcNsdhCqrbPGyhLvT+Z+GyVW8pBqc9CaqPk3pdY
BpIPk2dhpJ/rXY++7Dq8qyL1h4guof46+cMJG8esDmplJ4llMGcbr/lcQoUwl4EW
oWD2XgQAn6h9ht25SQDfxGK2omnTEDfFYW2VfGu1r0O/wrI5ghHgrsC50JbrDryo
qDjpcIV/iBzzaBh0jatBJUOgrmfqZ8XWydYAu2E2iZn9bNyqsz8fjewoTE7dgAma
77j4AsdYZPgGsB4w3qLdqD9Cwbi6+NXMjmjRP1looNiySC3DV9CRY233gwZtyjPp
EGXw74ROgGgDW5dqo774mw3p+9sFDW8RqKYNN+5a/fiNCQXrm9X9YvmlWQzi0rXe
kP6K2pOxnSOCF68EPRE6S2X1n1yiktA+WeSfEcRn7imav7IRHG5ZO30ipy+oSelJ
HrgHMATgXQlto6bZIV2lOGebiJWEynLx3IT3U/P3xPei3Hgi2GuHVqIxTuEquHFv
cFbVhrrsKbta8/TyLYIGfH4Ob7KUcKF9TY6ufJY6dbxEgt7VVzsGhtWOqJvS0aV8
Xl2WR34PuGzFidSn9iuG412tTDBTQka1GeSFPYK/qHTv7FqKS1vNpVMl3fvkVOX+
ziHi3Tbvq7Ag3AHJfkBVN9Bmkhx6mY4Y6th4v9Ez5J1KedivomdOBKVSGRaRb6mf
gG3VW+FIzvVPd6c7sRXtAknnOFCqn4Wdur5m1gYtC0v1qQ7mVEKPSBFZZ0kesBQG
HTahuPw8dUweYAY+aHQyhupWKzzjEM8TPWEqtG9sYw4uOwaAK6mD2l1E+SsgF3aM
7I9ZIHkBRloIee9bIi5RvIZpvjA9GPOIhjYEe6WSpBzRdOsBud2UvrNRqoWJqn0r
h3MtEhf1buuRQKIHnwCmcvzsq5G9I2VUI/rLwZHF6YGXkIDWhlgk6+tIUCZuFyqK
5FTsZneVwuJzAj5put2QdiXvClxNFuvK4IZaWHDZdcOkneux4srjG6DHctcMgFll
UWyFJ/oYMwlugoHp5tAoZkW9A06gLg505WJYS3PYWe3N/8pkkvDleEYRU5cbhmsE
ClC9Eglnpx7wa+zhDWFAmgkrvrHI7p0A8/dUKrGbmj3ADDU2NLQfQNR18SsoBpkq
sbNvk9Xs1fB/sZFwndISSQE9N3XTQO0Fo6/pHmMUXPl7QRFWTnVf8LLpXrolpNWt
FDv9/W7UjHuFnbu6M0Nlr9+erbbkdySXzKCUc2qVOTKovNHg4r1xX2kFjkSqgW2j
v3p8kT53afmsrybmBnVM8rZvZxa8xcgeI5Sgj6+q6t6SBt+7QW8WaWB38pYkRyow
er4/qtSL9Eis8RlCf1B3gIoTQmxMyIaZLSc/GVuARC0ASyNGu6LCc71enxLd78ZD
OclOAQ1gDP6A+YQPMCoe/6m7f5AlZp7bO9EQ3545oUjSIkJv2Fw1c18f6R5LnC70
Iqsv4ip4FBSTOkDuQK6DboXeBiQCQROEXfq56fbvv9tlmN7X04AargjlFinPK9s4
vnZ2jzB8bqMm+pAtdW+tPomYm9B2WbZDeTFzhs2vyBTRWRLKaGwVccgodzeuPz+0
YmJn1frpF5O6JEsN8Rq97L4GMYo+/9+9qkg/eXDkHf7JL2kfkn6oGvcHytLSPPtW
JSDIspMTab12nA9JEesjCJPAsZTQpGyuPDFq1yEcpu0mPBYzhENDYBi9KQCA/DxG
VYHusaodWvZV2cvarp95+1eRTcoMBqaavsSpFaF65SSuIGXYzKak/mstXg5zdjWs
t1Hu8wFF1Roor3N0F1Oye4yBgCxBJJExwnJO+p37S5qBxkpc+jIlNF71htyg47Fc
FDQbdNb54l+ycmBskO7OWrdKtNxTG5fSLAoNcsNCyXRWEiTSfWELZK2iZPisAS9N
KCnJHwp/bk6cKmITacr5F+z1avbOryq2+z/1U58EactzF9r5d+te617LdeCEse3K
CMQTilp4ZJUBA44M7WuSMjgnqUfyKy+G2FWbg5xSC00ZxEMhQFM5lqIrM4Z9zLtY
eQ98ET74dIFW6aVk89O6C05Uu6qUsis6AJn54vnUn8d4fVFeoGmr6GtKSmG5CxIa
THzyl2qt4rgSow8PhciG6bqmQ2+nEEahhBDyuxcxsO8WSAqfc99Af7nNti9zTPcC
w7avbEtFzJkzKBCXs94w1H/k7WHMI7C3S2TSeecBHTrBocqMhAy+J+Vqvb13bL96
5RELTF9V3GRoI1VQYkTL4nehsgH+pso9CBnsQPX9f3cUiqEOI68eFtYRGppLm0Nn
J6PzzCMbsyLM85eVdr3lOIfep63yaM8UUA80qodlQsLukhPRvHxXL0Afmd0CAFvh
bMPcu5T0f+k4/OGrwqrvPPTbwgdftF+RJc2xbqPYrevHyFjynKWL2HjxVsA4bf+D
lc7DAEoHdt31L8vLvBBy14ZHSj0lGrQfOQ4wUgfNjZ88+o9VM3knKlYpdCYD7HVs
5aYd5BFrjfI/drSfZiOxVFDiilvUHcBFJqHgADWDCLHxxbSkGu8qJf4sGjItwlPo
KNHoWLoQwDQF0aWETgeIZlExbEyg7zP89wlA2U4ibSpSA2pt50nVTzVbNSD8yoPi
Zf9s9Tl78d+ZLP1YqqqrjPBHF/VxlqyqybCphpPgNeTmwQtjP2VJEhE3vYgFqptT
LegBxHz0nfN/r/wzOqv8VEIMCPFbdtiUBc9GEhtVigZufZ3Mu5Sf4LPdmg740izc
KmlRfnqbEXYCE9sDqnM5+sbHTCiMIinuNgtPLDc7t8+Ni+KStUyCYd0dJSxzzRgk
lwu5uOyWyDNMIsS9qOTeTeMwmzam3fjmkpRvCUAdbO3bPf5USzEuJHLLCjD1qrvh
uh0DUottZI4Qi+2+Q9Vuc6B/5OwpBFI9KmECzGd+Uv8oSE7VBnUliVwrETVaM0I5
Jlt3ZdyrzVyaB7qyI89ZYwAd09g1R64l0/i1VAuJA7VGNhrpG8+U41tndg1ayP96
bR1md10rEYDXjW9L6i5BUE+L7fGZLFre0OUooagkg6IumjqNHyVyBhLBECmPWnMT
TFzL4VdnD/5u3qIAbDG5J9Kq79+Q6bKVKQVh34g188WzX49R4YrfIOscVYzmvS97
D2O4fUYF5mVDRIesapdjpQPZDXNWqEUwu6RQkFSS1rvUrsAq6LKsTnmH7GSXueO5
P/jIUv7PUGZmOHntEa5FTr9so1QM1ieYtJHYrYcYv02VKxQBvz+/QexfcFJNFkvL
vHACZJ3SMrnaACaQ86d8Qerb2VXThLWOpIn3a5eqRLKg1mLrmRt/in8Nf6kvuOMd
FK3hvquk//UDLVZqhQD/24rPR3ZV/VSZ9V9LxjS0CA4Z/ie0Gevv7ZjrG5fZLDTs
unpLJ3H1Xfurwi6feEs7+eeq1NqCPg51Y4c+cAsL6jobJdGVNz0k6n3efcuoXUUs
lgqcINT85RMYLXO5oTfFnQOyVai8Jmp9C5nGadUFeiKcaxDUr73ojgxV6CNm/elP
DCOxG+nkIGenB7Ra5RMghnB7XbHOchp562AsXRqqIO8Y814PyQ5lvqY0tp63zbfP
BAEhQhyT/VwCaXzZLYV+jT9sggD5nLW0BCzRCK2XuST2kzJBlzLLH9kQcCTtC1VL
g/XhdTt6wREzhgGeMrR7qCLyGI/Wk407AfbaCHkM8FoENMJ8gAZ35cwnk5/Qr80+
bgb3jJMTElCryrxeMYsOE8ad6kX6NQnaEO6AvlGfg/8JPg21wGQgnlgfXSt5ZBx1
ANr25RKw5lHQVnQowfimEQQuC+WDwwAlo2uvnUOlGmydVsiiFtmTyJn91Q0tEWIu
eJQo/suzm75WX+A5KW7HP1c3ZjkbGPor5vh8yy8jiA1s2Fkgmq0JuDn1zTW0UbrT
Bi8GBVBk9B7bsWMjpLlMEZrQmVdAVPC1RzeaVmOVRdrbP8hDJ1D+wZb1ZYEzbFC/
EVWJlZz0YQ79Na7Cc+L0jRHKdWgUMrHRalNpSS5xsKCvkTqATIydTw+ULF4UspMu
3f7QUoBgFJ7OJIP23E5EOLp+vtOhz+N18nJL3rRmsefD4VjIhiDLKI+QWhzWypJu
PGPiyVp+ZBg1sjpGod8NTsqiqlU09AO0CrRBY3CGRMLZzbWTbBhv11ZGaUT2ue5C
5hSE4nqnR19xPGv61IAFT9F4WzShwNfneRa/esVPfxn6UWd2TsJlZUEC6LOUzQHB
T/I4THgAk7+LL4GH4+d7BrQs+AQHdh/OsH3ZKr7GqIaU5RqxWaJ+Lya+IR0f245E
NgLhIUkWOU4jdZwa8cFsjBd04yFpU4HFvhBOx+eHiimI+/52ymyK7DkZmvcwhglg
fmhknxOZLHAbGYbwv6hgVxo4+u6MaoBhqvu0srNyd9Bde7cJ6OMufTeS8DGxUqrF
jlKb2/tO4VKQP5Mit5hKxJh1EYDsW73gz55uvitQCMIrZ6l5aK31RJfBaNGiUQ4W
TxlCr+Ka9963xt3AW7k1e1QbluOE9Q8Pkm2DStFUBT0jtC8nkPE6ydhWMuBwyzNt
MXIYesdAJPZPf6xHrBXJQbQc8z72725t5jaIto1uaqPp0UvWgB2Z3DlLpqw1UEdJ
2FaW0VFKZimcIv090XonkC4E+p8P+j08rLxX83N5GfAvRJC70v7s/RensxFrwIzE
DmMgnoprEDCRztQoiMUcg03hJB0V+dflrczWbsdPx5BuMtPV/KOKcVjIKpxH5nAl
FNL45UQUpRDyFAV904kjlBAQkMvOpzlAiEk57CYsUOXSvFyFjvRt6sW8qRHMpyr+
4JC9rcflUF3fhtqPRJxJE9Lgrwc/suHgP9RwF5d2DXTHivJOXoAzNhcG6YSUIvs4
Rh38CG7605F2gAaB8vLHOtenaC+cbBWuPAjuAzvaA+zmWogt5AKsORko4r7G4k4a
anLzDxF+0zO9DTDZWrCL1GdrJ6wLoGclh8Oywa8wytYdLnFOq2tGtC9gOrYXSbLb
Dhv47fX4xu2avjiLCoJRqWtkRU6sBpgL+0FjUUz0RJQvFUc44JE8eZz2jf9NPuQK
SXUkSW7VSb9QGKLB8uG0+WVEx5CeG7DEqKFo52R6FssvLJARgyAndt+3Mz8exIIf
m685YrofzhFlpKEc9YhNhnbGBIaZyjjXAHU9oexzJUDamxUAfc9L1PP7NjYAuJcd
BcPXxdKbUBODxi0IsqwZdsTpMSfXI/vzIgpnYevF6DuUITq+l+LHg5hyhk/nNMdd
omcxiUXcZrrQphOMQ1xJVxzEm4QOkNepn+HbjZLdh8O3RTkTaGNLbgZH8toSpuiz
TU1cbr7DBklGY+6+sNi1gn9ZT9gBDJMzoIGQMQcz/ssLlYFNaDXxoNy1ciUJIOOx
aE20v0H4o6PRycaVEvS3VOOOvTzf8/fTcPCHpJA3MWYLxKHuH++lW4/ZvWlPQcVO
M16HNTjILr1S3LsXO9JaAEOCfKoH9QLRH+P4UIKYhc7r1tls0IoX6Ox77rKEWtGy
LI+BTT+4lKmbeAIWUPfX3hcL2oiKDw7RkwtAQ2uUMWdMPCv/DzXlOPCDPoAKkRKj
nWQejAE9kR61xbseDcyfcYn5UZQMKANMdf3wm0vsDnQpAJuJBOHJleve6TXz/j7X
w5mVnn4spuLp1VV+9BtUSV0HnZ8Dx/kAfTltBDvx2fdJfUYbC7K80bCnfIE8Pa6u
mYN8XCjh8y1jPbVn9ak4SaLP2Evt8MlM58KyMXEHzJXjONsnL3IkauOScConIx7n
3yNzYqS/twVeb9V33VO8/NfK0Hs+sVXpv/4jEFMLv6B0hkq3NyCYgcSlWl/Tu+l5
thcUaOb8CQQ+0eJpILYbypATOCwJC1e8KLIjk9EL84iQFLQhqGa3Nv/oZ8P3G7Lo
2bJHcXb6Z6wodMYNMJtzSzVqKUmFdlxnJdn+NqaGGDFsdnbZ6v2pNTTealIdCiPY
dYBeROzKuUcj1kwzuTBFGFc0dIKbBC20JLC62XskTZ8I5HTMg3KPgmOW7H7BH6b8
YtS7QIo/ARhafLKl8ymV8lDEKpmC5C7IAEWZqt/rTTw=
`pragma protect end_protected
