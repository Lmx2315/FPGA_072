// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:36:59 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
NalSVN2stJvMDNavH62s21chNNgGYc4rYPAJ+CfRpqeQv3ZNHAC1S8zwrHdh6rwX
AwMoJ56H5flnc6NUMKhNqaVLBSc916uTqhTexouYjh+AfV9zNttjyMzpTcQMhMcV
oqSecOWOCP8l6m/Jw3xZtF/E274AFcxeYO01rhqbZ44=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 32784)
UGD0EQsTZ14hTb6vjHuL0O6zxYPCl3gNMzstzmPdcTJcgxJmsFx3LHUl4VzyE8k1
o/mOfhFZrzmSj2n5gkU3Uoj4rFsoQ9eL6uI1leansEw3+i6uu4wHcweg07xSEp3n
UKgJ3EzPjd8+4gI7Q+AYk2VorKU8FEAIxuQyrsetluiZc+C5FK0mM+ATrjxrF8Od
zPscTPhrv43tstLsaCrpcJbMnO4oIvJPUFvKjnsj85LHGC91RINVgakqqoVV3Uvl
RhNK2YeNYJVf8IXbD3eJ8v19NSP8mcOpsJDQxWcxwC0SzCv3sC53n6nwbS5/q8yO
cHeO/+y8WQXoYHK3aglO/zZJEUdkFHf6J9Wd2mw5GoUaPCiHbgdfwy+kniRY4Ctc
g0RjmkbiLjQJuobU2Ig62Kv6gkgBcsJqvsxPHzh1dw0JGtRgb0Spr65hhS9bgkX/
GWXnD+1b791nci0Sg1346+sAubdCyeN0Mtl3D2pohRbPVlQympANF5+0mfu56Cso
uEEmsRdOZ1OAmxw2nthSQSPcAbyBYcsKxjGQQd//vGPzL5wJWIWoZVVnm1kTIlY+
lTwXfknSpg/xyWiNPlsX3ECi9Y+wASgojrOnFgGeNozbM/GGRNKqRv2tPsDJjN6k
DSOYWK2GYqk7USSw0fO0Wwdi+Y4riptZr/pZID3eckaXCZeyN0devEd8yfG/LV6H
AfL+h97bnHbFlEMKfVFP4AmFFh/TxpxB3DiavctSn4JtQw6Z3v8/TDL5gok+C/nU
TNS3SNn7WOeDvtOlE57E5139ypepU/l0FGKRZrZ99xOAbsY/HivlgaNrikrrYb0J
P2DJ+WKH0pUFI2ez8H4+SNZ2iNKPRfXLqBbk25KDhcI9NeoehBRNww2PBiK9eGcU
hLAItciXJeKoqX0mySXP4q4gbiOYBthOlgvTLiVjjx+FbFzM7lIvuVtCeP5nF67O
nU/Qq3+yXvqEMQ0aH6x9ElXsvEg12ael2CByjoeb4QA1exd+igS6LEcl3cXvWSHt
dgiiCyPwApK2mM61HyC1XrJSwWk84qBY9oQtywfPyGa0nr2wqhLdn5mJPczD8alG
H6DFEUITPoonu5dwYZ5rcuQgXSbtB370nN9XcDbQ2zV4WZn+Cg9KqMoB6wf1Zzf4
mA/z+B7VWi5a2udBs+gKvnCw3RTKhWisAvO5gXmEZD9wt72mAII8s3lB4G+TiyiL
KnxcUq/WZt+VGEIqxfuASshsHzDovss8C3fXg1NL2mQjSays1aX2VXNwuPXeXxR0
r7feGSdJi34dG88sD8AjlKunPgTtvEy/qOuKEwDqF0Pz2Ilu2xxG4N+VtUiJ3keQ
3RV6DzDaQTUvsCUyca6eqOrsAZJYIQ6mgcmI5TwhlhB4IcqnNjb87BIS5YSnHfaf
Kk4LM+rtSsAto8Wy409VO7qm5rUu/c2CVism+didEYfSTu48Uun1TwQZrnMvFLzS
NVrGWXBJ3qjunkGJUzGv7SRXvXmOW/eI1iQBqYLV1dx60AjV+etuHRt63RMEbL0a
hysqmNJNMX/mbZqnfi79/gbZKwadu0pneQjFUcXVepq4ktTiQXhgpsKTERilQ9nA
RyM07faKxzcw4V8EF30swBXf0+Qa/XI+GeDlIXebBObmdKHkfNrtqCL8HsdsTGyH
3UR0+o3T5UdH0iZ4r+zElrHDqBxmC69vPaL+JkFR5PuGGAzD+tJKXBDAiUX5SDyc
+FbWmTwItDc+xmjndOUPOXvdNFuuw8lImKPURtZLXf4C7kdHxqIGw4TAboo6LOUO
l50GTkyk09ZUhDBVD/YIZPDnGJuIPL5jDTOisSglOeUhIqzAJjBxCa1ioUJTH/QL
ZYJsrM+SG6e8pGl1U3iysp714og4iqO+/IQP4su86OjULtPEC5VmQCq6ACLifRRI
92N0XUTA/h8lKyE9HhAsFSrlOjxjJm6Y1pUtEBfbzxLpl+Dzp46yP49Q8aSboi5g
3dfoh8XQfnuSwXCNvxK9CeUCg541D3a4lP+1rHUbGT2UJdWb5O4Ghmciuz8SRgFd
xharLHphPxH0Ol3VmbLcuMZ8UuM3yj6zHD0LAOUXYzgjknPdcOpOuI3yg4G+dtjL
Jqc0NVvMQOjQaIatoNx0NxzaJeNfF395sVXmiQDVr4qiiL1yWtzzWkTgq4fCHa+L
gRuOT3LKUS2c7BCkNgp/aEomz6ewWBoN4/eDRKoFngH3Lr7kqQC4G4plfc2unud2
GV8mjf/9MI2IaeaavpRodAm/uz5LZIEZ8WudtA24njXqbbZFfC+mOwohfLJtZXa4
AvisFlir8hQjaTG6t+CFTPVCPOcucTM3GkHbKuuE9ahaVoODOVTqnpyAX4snGhSc
d+ZvN4v0Y2jynN1Sg15NMcAG1/T4iGk43H8e5YnF1ZfVxb98p5eLtFqZ3BBd4TPu
XVod7gE6kdZBAAOoPpJ6xh0I7LQ5ry1qRYk6PGP2FWYu3K+9DLz2oaVyATBwLpcg
/eJxqahNTEqDmGC1SgRANwb8QgR1r1Foy2ck1kUFVuIBO6Vtjj8/T2hOl2yfp6oV
JJ7JcoJb1PZRmAYVbSSdExeUBB2INRh7pnZveWtv9u0M1LeluZy7biE8uFkUq9Js
mWnV9E56BqLeSmzdlbV+4XV6jgXjAnE6LHEkSv+6HV57DYqMtC1Yt4phpF93ysVE
7hk9d+/iv6gDY+HCx0vbwl4PbtA9Ld0s9K6WJR8PDgfB0Dc10fBADBBwDnnZ//AW
mAXWSmrYM1MUBZyONITI0ogOe/7fmqDaGeuRAGHFdFMJDatGJmcrM63ijEoQdBb9
LiWxJb7EufVrcSsLbgIzcjLUF5txgu2MAs1kHHPHaCJFGkHF3hNg7u+DaES3eI43
VoJJAARhsobQScWE6aj8WsXL4qIB75pXVzu14w0+cCuZwzdgixibJoN5rptDjhpi
dtQVUtSUB1XlHWWjbkLyg+K2zKaW5X39FhkvtZy/mi6ExWjqmpiE/sw3ngGS/LGW
laEf4w+rHU9JWfqn/yx81w7ZprYW+G7MMQKZgJlHF7Nmae87HFnZgzKr1frfLz0J
DeA7ryOVJJGY0NtGpBCRDwSo0NEE8bhJEm7er0RcNz/+Vvg0NbwRK4KdLwDlh//A
8JJ+U+rHdUcQD4KLBxgPbYslfwWoFC0O9O2UjihpMd8709/N5DXjjPmNK4eX+Rzl
0Uni/p3tuQlNv9VYcnV1+w3wlgQ2WOjj48TdayAue9AKumenh9POW3Fb1TZn/pAG
GqEKeUgaXQrnLbc+gioKZTBOPPBBfdzTXays2NkVU9yYzBhh/9VBvDWNIN7N6gUl
81borxtk7j8zC6XoMfQ2h5PL0V9sQ5skKu+9dBvx09yeYKctu2/+41Axjpx2fLZp
N10R9hDT6wpchS2wY25QjTSkFpMrlXsyb2uu6pNxsTJzGxsZK4tyZPDhQ44CAq89
23Gw+Mx0HMWeC+5wJyyQPJLElHPKJYJBK8fQ1Zb24Hz2H+6JRJqaxfbEU1q6cyZz
6J907AM6u9mIy1QYy9KMM0lApxx5dOgxHsntvmbNaX4tTEDhT6rNJ4GtXfFSw9u2
ovBexFkbm0QDhJp9FWMDP01U8B9HxP7X4E4pmbsCwU7JoQbbB4kkeILwJhIgeG+G
dzOl6QH/1FIopDSxhFWMRrsqxdAgfz/omy47FICAFopTmRsH0T/vHkQoBs2nMAto
QHPq6CEhJJpvyhboejAY0/LXYPf20DNVbL5Mj0GBsj5oWAfpO5U+buWIZbXwncqZ
b3J8G1vWDpTljUPEi0Fi6eLhTKurHRTfJErfHvoCzmeW4BkCtoid7cxPVAxTRSwY
fUpCjvaLhDlUL3GlnAK3hBHszP1mkaGPXU8KznvoblMMaLDFYDID4EawxySLD2f2
z4bGI1KSyTJKKPP9wEWv2SccX7LF8cBd66KKFQr8bMJjpgsV1MDVud6JZk8UCWTa
fb4P4GNX5HUul2WIXApbC8l5xi4GrTv8feneMD8lNb1zuodre8KlVE2w1uRgyOcm
OI1jzRl2xfbiLeUrQ+zGMxGOQTS+Sf9nWBeO77hCOsLOUZezz5iC9wsqY8TjH9xB
mFytCKIHUk3lo892RBOKAd+jWBcZxZc8Vvys1ztdOEQH7zGoRnvbTzHZCpOGSvmD
D3sx+yA1VGCn8k5pR28wT0zhNis5HDHjS9sxSrhMGms7NvOoZZirQHWBlMGa3/g8
DRSjTMffmXEO5Ougn0idNgxCAtWA57R9EHMVT0D+AwZ8IeQhc3JwzsjkoG2ku0tt
Y7IxqUbOdTTwJknKUZRe4zECU06FLNuy1bizIWlz2Rb9KxeXLK15uiQzUmpe3wnj
TCdDUq6l3gtAe/jyVwFPM480mEw7QmXSjBSZFxFLFB/Y/JZV0hA0AWrLHc9IU5RF
ciubPiN6uuG2ZPYOIP8iyV505yYJEMDgWobbZf+f638nJtMGCetHTRBQWNIhRIt+
oFmrsPJB6lkE5avB6PQ4x1D86fHJpC69qpf6til/4bfOgj2FeZOFNKxcJ1K8SW6a
NRCAleh0BPgWNY7FELSaIYteuJO5WD54DgKjrE5SXX2gIhNeK6A9gCgdAhMCzcdT
t48cRb+VvgWGyMh7/hcEg5IbynV0MUgMKyTEh+QKoirOR1hCCNRqUKxPuOOtqhFj
6xj4ioXgbB2dKiq9/Bf8Mwcj8fOshw7P/Day/LDcl5dYwpVOgspBrtLNx2aYbiJ6
HNmgtwsPpS15yTJVyt8ppGelRfJJAXJxbVi3OFjr93xlHMSZGaT7fg+3NPNQ4OF7
hPy2SNWCy4AOsALEG31MdFcuStG1BkMP5dCRXm277MIYp2aOvCFcWRKGteUaSWVw
VZLZYMQ20Cam5p70nDTw8/HLb6qu4KxSpJETz7Be5OZn3XFPL5fldiDhLmLoOpBv
nB5J7v7iL9B2yiyMRDSGT6LbOhgtH59y8ZVPUEfw+7+UazMza1iSYArwC829lwvz
tn5G9TzjuZ8CGAJKZyOGggZ0pzdXe+YUC2zg8V8nSV6q9OSxtYcFeTUsqtmB0RTO
SqKS7O8RSk0gs7dnoU95IQgfhKdNzwTEEjk32jhD1SYVpl+HvJKUaemFSym+4tse
xm7L7xAjsS3ybkJFCSMkOuO3xBjy7Dprj8G1wNTksQI2MYH6j1qX0GFOLTGMiI79
Ebp0OYvCh6BKUqmOif6YzwjxTDBFUwMv4FZ44j2FYjoykG+LDqrwTgCR7UucQQ5E
IXJ1KS76Rwv3jqHFzXaaZK5HzNBVNa64w+oyX4kF/8Sumdh04R+UWaeVEU2bIcki
HNDKJbqcl1hcEPYKa2e6d8tRzp2zqUVISvZccj8YSaZG7GAJ7EZCpSHuXa8rKSA2
kN2cxdPJyQyDOaLVFdiGwj4kJM52Y0jM1W28x5ckOZHMpAXQRd6Y8pRBuxZ/DLEx
qyhHblfKq2HIHVnL6586p+44tZDpimEdFYiZOvELEtw7QsqZf0iSxYHCoUwCYQw9
gKTGQlvzlnR67JVMBw7HL5LBTi2rToaEzW7VzIVMBYLHu0W+m9NTA/D9u5mxohCT
Ksx7Lfnua/qkw9cAxrGVx1DjTngR05hiQT2AnMi1GX9lQQwDb/VnkInB/RoxCf2r
2qf1+YQyydnCtyY/azB9b8xEhHYDdx53bgGqNqVcOOZfw5s+iGmWDmCT/ps+ESz7
RmnWNuNI116G6Hq0RVT0HKx5e42uAKx2RUw3+0Jnl3ZpOxUcv+Bknb/ZRUCB/Cw8
zxL3mAtHj45UGNlJshHySJWSYW4T7nCzHYYCa6aBouLHDo4Iq4vSqMBVSSRp2iWu
MVcZ0+FKSxK1sb2eFS+F4WYKUTdZQDfxn5ZnEKehuCCV95tb0wQw0z2LnZqwx91A
XKp7D4WNpCdcgS1O0XLF/Fu0bDh2LTZ2kH9PUhnuHLbv3vfyzwvd6lnR+rp22v9x
6vrFUu0k6mmieJKcvS03CqIi/hsnzgKllayJ1tdavGISp1GdqwxDRjeYeSVwlfjV
0zhvhn0OmYnX7qaUCPiJGKyUf65GRHr0WzB16zEwaopBx8K+LrOfR8tH+EAusnue
ZmyXSAE+3VU7Gyd8TPzj3QSOD8eOQh+3JSnbJHVrCgpyYa9Nc5MfzVOeuX4+FLgA
7pqMG2Xz9uKQgQ0QvIfdaOE8Ec5tIIwiYvwm6CbhE0TFC4SSj8g5uwIxl7nXwd5H
1w92wJlrVweEY3kbAdt8DoosTiP1T4xj2MeJx1Qw+UB3n5/8QZp9kMcPlR6e6iwx
fx57kbGLe4eIaXQ9P6TQWuAS8lvLIX1R1yZ41Oy/jPYwBHbfnIBjG5wvygl25yCW
FA+NN0uTRS8Wo4vtnk+Y4bbai32RcKl1eAer6LJAaprDyinPmOAQMtTSSnBNzqMl
yMRZLbwHo8uPx/mLTu7gPkDlb8pR4/4OVcdNAnEletEEK1bwU/UnYJTA8pG671/i
JvAEXUQ4QNaOyr29Rj5nbs856TCNGECI99YDYGHvOAnXvwGHakCfc4Jqpj2Caouj
RGcnFf6QEHRiY5EUHkEk0xJJHvFItoWec1dBYMryNNgmefHVcgB4chJ0EBEkxjZ3
IGPBkcUz2+O32wgIRu5nVtu5fScKZDdeKnFk3d7DcsFXfH2yYZb3WbsymM26e+aL
wmI+XX6e3ShBSc35baJT+V8/KVFM/L9uHvYSQJA/jULbEjUPTPzsD3BWLWgFFf0A
bvWCIN7v//LAmStvb373Mpo6veJfnDauRpg3ZBPvucuanlpsoKqf3UKebwy6jRPF
20BnlDvGQ0HkmCCL+Mc3tMUAgt/dzOViuJ/i8zZX6yi4d7zZDTcljr5lUiTD2HyV
ERjX4dKiSHokqSOpnQLpUkkSSXICuVx5Q45qqA/cgCvsboQoRLYuLNopf01nH4o1
IgPa8zit/VyZbp0TKnhJQrW/jyYl58cynsj9tzelo8Xn4Q10EXCn2a6s136YO+p/
454WgtvU7vHm83zdCyMrU+6+6Y4VGJRBOgoVi9bd6FNvt/BCa8V0GRFCs/4Iw3u0
0bwH9V9n+pi1lXqZFWqZa5fRbW9Zz+TT3toX4TXllYkFZkJMdyHv7C2n55s4mwx3
6sN6qsn7OpNPudUDHh84HcLUYbsfRtQd0Xv74/nNnW2KuvyAssFhkLClIQAXhnX8
ZfbGUVs8mPK4n4DQHnoc4B/CPGy06yJmB6z1VRm1W9YtIcJN0+P02lHL1rQ3B1Dw
9vPz97qJr2q6DIFRE0fTsVYnoeETC2atrl4R6gcj9Ur1uOekFnDfpUnXOUx7jxyI
m65evIzGh+2LFL/ug/txst7mPuuu3TNF8RSc9+Ez72cJKB6e4KktUYKBVKStgbxA
JSlH+Gb9mzCeIs2lsiYiPF2ENrBJxlZ/XQfkeDqQ2BEl1knQAJOqWmST0ebe9GfN
R6b6kGTiaBBYGzj6+vqlt6rVpOj6aM7WuvxvwxZdeQyIApftuL3UW2FGpgLqXSET
Ss7lPPdyrOejgUfJM4eNykA9+qKYTI0/Wr27mJ9e0sNdkzRE9HkNxJPkcVfFj29y
ic6g2E8E6wgAOEMIsCO2bT/Cid6w+u4dvBIYjzcztOaQY5esR/5V6L8WPoUtUon1
SHgzZubwyFv4OWpJpIKWopL81GZsRaT6crLn9yq0/0quKvUwEKV8Z/tYJTpfuaSN
K2rj71gM6RYbwRiIHnULJRmVV+TYbLhBs7eXkBAJZ/HwhuVS2qbOzFnQlJcMHBcZ
uKlP2z21loqNUVgIB2ph1w5Aup0WUgpbootdMbfzFhPIGIPMLLjQ60dkxZME0wGx
AhEhXdw1P/J9p/4Hl4fddUucLkDimfVHgnhw730sn1SHTS8sw1EpFoGPRNrf2vmp
o26qAIQOvhCdLJDBIsHYIqzB5zjitgLik5VG7peVrDcfLZYERKi6x1hJl08Y/qcY
fn7JvvOlZAEdPNlJQKuVpB4jW5TGWOCT2ch1njswydhHydo9lwJnb8CVko0ORC6p
wvAaonsSeDvZT+Lb4+x6ud5SLPqT6C7P8SRk7H+QsT6hFhuaRmNNBjeAtgj44ylV
QHXWuPIXS0Oa0OWEA2IxpUF6ls7RHU0RSFKBvWEFuWbZmKkp7022jfuQaHPPv1wP
lNG2Yk1QX7ZQwrmOvdXUlvrOLOmG1Hvgdsb8iGtbKkaxdXp2BG1s3Q5kUQUDao4G
IzGYT1kj5OgtwE+mD4qILFjadqO2buNLdrKdpIRRVbTmiJUskAAzF6GN4JL91+zz
m7cEMV/gT2Q+701fTM4yW3mS1tKH7vMs8H0mgXOBEXycniWr7255/JHypruWJ8pq
VCM+eYu5zFC6Ef7+thukU3oVmAWUAZt1uNUOp0kONhkP7DCwXHSuRlI0v7oXyz21
o/tUPgZqmOwCf3DyOxFo4ajgiqWHabwgAicQvHBdhJ7H0lS5YFynU0z9GW4N6H/g
7jSvcPE7HwCP9bIOZuC+oVoYi9m5eN2whDDL8HMOwcqBaoIOtm+h2lQr6SWzOEn4
TinzpYo4P6VvfwbP7KGu9NYh7eXwes1XUP6kTXaxbg+/pLBdas2y8n9BmuVgo+41
5uvAL0Wr0iIuVXwCdLnTP7b8+KXbVcrRM5bQe8SQJGcpjv+yi3fY6txnHwBx2Zag
QzdHTxVXZ+q9F+HzaIyoNohqNmF/AYSnQ3CrkxL9RT6sb5Cr9qziS+qhki+f8KOJ
QU7JLixvbedbs0DXXaZXnPUJHJYbfSB56X5bl9vQl6q07kTBnalRIc5vMBDoJ5Z8
m3Z3iHcxlqf9JcrDg9fn3HD4GnlWD2P42/qw2tNn5xsOon3pC4eI4sYFUJCZqQz+
v+wbboj7h0/TtlhfxYs1Ad4EoaSofzbVy1GB9ZZPjAxDJgOJsZc3DvLHCExaPO9P
SwlIaKca1Yqn5UIIBwVFFXbqPbJ1SL+1hXzJuXr9S+yqOLHuki+xgMm3uZWM6Rmo
ILeCcUW20+toj5fIM5RXQiNXUAxt51lQBCkhxoI9HJumRWNz2RY8wE7eK52FbPGz
Y5v8jOfrNqS3B+gcRD638yHo5vUChbdft/OetZkvExBYfBDaStf3AlKAvadZxtTo
S4gmwPXEsCVrkszJAmOKih0skiahSudWF8VJ5Fgys6XDeG334kbpdPj4o6GHNUF7
2civ2yCpKZMy4J4CQ+q60J4CNrGH/JsNqGOdAMGydpIMVEaTcNZDp2mBtf3cDKvF
0RhE9Gv1CaGCVAMzNsEJcep7QVSxdxkx3+Equ3VgI1R/KLNPoT1YbLYDktENDv1P
GLbF6RIo0ws5cNI/5AL+uzSDYm2mQ5WfIxyRRLDz+Z08KpxLaNCEMamUsUgwSDiQ
KXQyrPxohNydVEFdya/Gh0PT37nQDbxCSJSDAeiYj5W/JBcG5XcJuLEMLPQx9bgY
iIaTKG5HiEIi8XJzeDiEE3E6s5eM1kwQgfiC9xtdNx5bBliVG5bJ3ETkAy48/zta
cqbxBbxvptkp9sz9jfKpl3RSmxoYlMCl246GioOxopzyO20eKUf23BDJ3gZ+UY41
HEIz5G2Tb6Rx00C8oQrn16mPvkHnpvil6ZV5gyA8l0YSE8KrISjl2TvsgWZ11XF9
/2JYUiDaowDYnpYH+xFjoJyL+6iYsQ3iadjvxDifQZWLFvuFV9d7qJwBG0TLSPmb
pFAU6oo7iBNANtmlKr1m8++Ym8PNMgu3ck+MChleZf65FTVHlPVMZbLQGE4tdluY
5pTQXHceU6tAZmba1lOiHKbFiOzsH9zP2Ce/laPLDjf2WtLeWk4LAg9TZqnCDDtB
NPAXcpdkLIuKjQAjy6DH4m0h5xIIW7zaPNX/I2XuESvNblGkYY/NrisWHvPI+BgR
AdpgDAHVSM+3cmUmajF/LQlMAFPz1amRlDVm39FADvR+70zOo5/zxC07X2MngVzJ
GIDC1nV3+drOG9QszFFXO8KOcx7gD+QJUwRqBplK6xtCh/vWEF2Kqg+0gZUr+ywY
x1AIAcwSYrHcsXnJDWXd8IQrB0IJIlJTb4vfv8Djia1qGAXHntAniEt1AmvfM9sX
l7EDS1meWo3RCVHyvKVLZUe0nwkO3qBjDa/s2Uwy42w3b+CS0ynAK7pSxGBe4MAO
eG/tiBeoEQyYtgykCzBvwNUHGApOpuMJvhr4Fne9qKB+1gC9kbhR18cEw7LOnBmi
ZljlNnx66rorqXufiMVn0mf+CCmdlCG+7a9cDiUfvGOPkkZz4sBIp4rXvtBEnbpD
gKAr73onomRErxO6fCxiyxCyazhBm5bAGhEUqRaOdIFl+Hdp8+UejhYofyt2JEAn
TsqqTfxphmJUlAFa4XNJgQH12Mh9oN/qzRlZXTRLTn24cKgKmhXoBaESrlf0BBnx
3Tr+5JEkWQJVUjl7uQCOiaZ432/OSwO4XItH0Fb/dhzPZAQEP0ILnZRttFOlWsjG
zQ0DDfx1pz+85pgCfbDGywqG7OCIM9m06Z64vkxUs1yueYgRh6tGxvV2Lzz+B95P
tUUkGQeYz9uZ1dEj0vGOMf2JW2S8XeAVsHDm4ZZg7oc1tcWJHwEtZm2n5lejGC4k
2SG1WNfZizcXKfu+SQyj8/a5CMh0yhvNqtIYEDZ0Pf/cC4NVVgpy9cSznkVDhdIc
ajtotxiYn+uudzAcxTKTmnqLiQt8hcuQiD/jJ2EXgfOZajypgvL7nRSYAdY+DQjO
EqgaetT3JMkSbJUjAK6AXbHMceajiTcJ6dxrdRnFWps8j4ObQobl7Xq/VO0cvrJ9
ppjOkf6/GsDH5/H7/r+CUEh5EDRDErSwBtJHNo4o2sNWNDhHt6W446X5mOL7juEf
wUOR0UpFOMa+NzhH4S0a7j5MZ7lZiT2lNxDRE+mhdUZ41xpmJJszfObZUkNmVOme
XoakBizhETFL7bgmWzjmjB3XHZOIdlXZnNEVDnWjxMlxG8C/WwtuFgk9gV8L/0PT
+b1g08bs68McVknWkehgsTSLeIdxZSOJvNKRSIzI1208i05wSsEyK3XTfZ5rI08X
eGZJSb2znADKPaYrr+3t5AXK3CQUbk308t3QYzDtLS7XaHyWdtbvVSS18bilHPJE
eGqM1lmLoy/5vRCxX604g20a9LbSTxnBIikDFgSiiLn4LNIyzsDbHOLzUlk30S9I
TWgzVY0cZZMCupWXIeiZxeubePF77TqvFxf9TMAZIQ1VJ+Xin+yKuveBd4G1QI77
4zUABD66JM2/co25m+7nwzUdLY4KA7+gYyYCwvgClkIlZrAqoWHnCKhemBfqA17f
wcdN1gGR5USJjN6Ku9EfxwtKTMrUclwYz7w6lXE2a57hUUnQstHesncKoN1WrOdY
HEzJE3HJ7juermAF68/OxRaiIaQ+BJaPvh4aCBEebNvyn3oNZ7mhJ8aOxhSw7wUJ
HjdJ/vO97QcnpL9TYDVHfsT0sP9PcqoT5cCGCdwez0yfbBafE2RQHjG0RgAtYaDQ
nLKgPk0Voz2k1IozyUqIGIWiwoCWWSXMqnFTBWxf7tRivtopYJgeqx+3wqYYaSwO
ifppXofDhI/o6w2RI+R6B7d04idcB00Y+ytinNH8s6AE/olLgUaHYZEYmpErr/r/
0UT1wR88lHB3gD51v9bqA3suo4GLVmSrOTMENcT1s34mEzgBx7n4BzSX4Z4Lruz1
OXgiVuA/gwTsKGNLgmXDomt+F7g0lFhgYROG2N+G46T+VjL4sdDHIUBEmlHczjhO
G7hXstEJMb3SnyDBr20b5Nmx5zZF86RqmCW0UU/nI0jEJZ77UZPnnfjZ/fb5RSRF
R4Q/3YeWTfDTqcTcn0xcZM8Sko9wHqUPhIq9vnpM6568aUXNglvVy1birPTmuinj
/kTwOIqwrLuV3sryr1aEWlimrZO3bvHb+t8dwFNrbvRaKsVgarE4X8zD8OmRVxmP
TMSY35yjzspdKHA/I2XidPYC4PemlOqez9eTJv+BKw13PFoh1Uo+Jbho3CTGsx4l
/Y8MUsjTZ8AHodX73pWWjF+Jrr+rOPGSoSKcllpl4SuQVsvN6xvGoK51w1BD/6tF
UrGuEHJhbxy4jLHFplZt3tJ6LauGF9ZUVZllFgP9HncdrEF+1j1aRunZYNNEWltA
WdJIy7KfEKzLn3KqC4F95AUnW9Be8ZBPYdFo2fQb7AmYook+0OkSjjBKHV6eU0yq
UNYwhC6d8ez0TItg1FryemYElkcG9r7Z56zz7JMWwQZ8ZKuGhXlHMLj9YV8fEb7x
QkUVNe9RidUGh9slTgcfC/Pj+iZQzzKxNx645IR5GkIy33rGx8kUc9ed7teaCoSd
98G+DHXQhxpgexjhPO+gqUoONFh/K3gG+4d44ZE9ojMLB3gufqEo1xJPF5Smxoes
wMgArOWpmdlRnsj8ISaUDfkZyMr0yigJ/rmH316hBnOLueqk1DRXdcFxMl6rRmLE
ROWSvuuw406/pvyS0QEMj0gTf9KPggi7BQONgBdnMM0TRn71Zc/xsw9+meK41aq/
jZnQ1TM8s64psz2CjqPwrHSLtiXM20aokasNfEjoNsPwb23lcAl0Mu4tOBdRwKsx
xF/cC70srO0fx7pEA3iIBQ1QY8IOVuUtoOCCqZVoKHHN4AawNM4JVJjXjuXwRs2p
Pat3QyRCyu+P9ocJ2VILmcaZLQMtcVqShM6g0l7SbiYmJ5hpS/pYfhul8iClS0aI
UMzNzYUk6YFnZ4HFg4iiixYKOHkyCrc2K77KuLq0pBfJQxG2wxUIxuMZ+e/AyJvm
rRk5E23lYYg+GawDbMIc6JPWDna6aHTKhW54b4+cJL/K3fsZ3B2x3lS2znvZttx3
mtEG6PhhOANBc54gsZlJmAife4epSXXe6mv+CpeGDTXxlIxfZp1jI+xUrTXGb7p8
BPjTnW/JRCOPmUNDq402389wBqkyZRNttpyHT+XC4ezFVhuvS/Ctftw8xOp+8IAZ
tXCLgAXkgbA56oIVStkQBReyJhknW1XdDmwyyzs/Bta+NEYWrQrRuv4+RtQ7CHzY
ow/CQa0/UTDktrI+j3gH+Bv/7Oq2z1hj11OF7wo+aND/goEPuuIg56lGlWddKcMv
1STD1Z6xGCAfvOmOQ7VPfSMyAlQjNPW6B9i0VjU/NneojHSfWTdgndELruyei+yM
GFZVmvJWS8VcMHIVokZI3Qo7+TYmc5A9A7hxjdb6zfI19DGOHIs6sfbMXsY0zmm9
ArTxLyVq8JwBxqlUQgErCURpgBah4VMHkE+TgWqHfty0HlANO5SDQdGqbqNvKwwP
w56BXivndEne7gDII3ISDBaNpMU+qyyZdOHLL4EddP/p2NLdz64Mp2JbDfYszoSw
bsz3mBHnWwdSU71KmIDrxvHlyUBulNmAilyzXZYLqjfGQ1yy6rk0Zx07YQL7W1gm
34yldveTIMS8xnvq7j6FJM1CHopPm5KMXmfDgmvQD4JGBudpBS+OMrh45hPHqV3f
+Vj59yPNj+f7C6SBvGVIcqnsE9qBc1XQZs9vXXCDFIqsu6hu+NBknAhe1waY/yYu
7ZUM//tOHjZw6KI9rJzIYOAwFn4tI7St+tC8P5L10uHHoMMz2UdN0TCn2I5ppiwX
ID8TLEyaMtVhonv6jmo4P66jD9LbqWt0eT2HzgYX1UFJPr8h/65camfZuvoLjWcF
edaPgPEg4EhcpIqBdhJz3vPU9Ld4e0xeaRpypo08N90mQ2AYsqq42RopEmyq+Eio
gX3S7bg4wGE1X3kqfi0O4F8RUO6vBwnr/iPETy4X6nt1I3s212ZgvuMVLp2Q35Qb
4WXFLjb4yRo5TLC5EDOHmqY30FYx73fBEICwUWoF4rCPnI0IJMhX87kXYhekdkTh
jrwyt+fqEN4k/cIzk/ioLIMAFo+vDY+Y6qppdM3W2ezp8YRVM14FSWr3YqG4fYde
23Bt9DjnGbe4rKvIz5trDlAu4BxilF8Sp0ZcRK8y3X2aHZbEQaizbsIn3+ME+mIn
DBayoDiBeBZiXUkCOdCfMDo7zb2nfrimlqvw/OSlPX36xFtEfXt6fgtEzeqvtd8m
9vfrgElo5lejx0oFpcStIHFNOjnu2LvvhcT05h3pYMZFW/LDdhhZgPOra+DmRMfe
dqZfutVA9FW5j/xzGvyebJhWQAwEanRNz0IMPrPlaHd5rh1zAHe55cfzC0/mOPh/
n90u4FXHAXdUBPau6TiHB2QFuIx6y/iUJ6MK7vSGafnTMZ3NPg066yOmriKDHqUx
3H4pjgj6xkM+u5hN5YkFON1/S4MFyHjgbFfOjn2EyQgfbkjm6ABjUTNCbwjxQjfg
83U6QsBw2NgIYc9g9tvtvsI4FTloERbBDJ+BHl8KTmg82WqCHODkYGxaKCE8dRD1
YPUfMFBM/AgXKCIglR4YlmLlX7EjKgA8716yfAq2fszU07H2Lka+pgxRltzxTKgy
BaauikOVHzE2bS0AJAq15tJXHfRQv75+XZzAIFTl2Y9pTMBNHIIgODSDHaEXeOLc
O3XRA8yzta/SWVBpZv/y44KUi6Pb95b53dIZxj65FMHh8nW421RmfAl04EhMk0Bm
aLQIROq009FcgLvkrwUMCGrUTkB6/wmJFN+2TZlm1ySxzjOq7VSUeeLp9n/dMK2S
Y1ONsmJbSnkQopx1FDM/I5DKtlbA4M7xFTNrutaxlaviDicOxeIZc9yAuKUAdpZI
lkseDAkK49bkXc10ZWSulXvwfZfCHOcvHwz2ZwVU/xtJxy62vzVjP0st0WNKzlid
Yd+GmeTq9FRchwBW9LJPdZdLr1EuNHe6ETM9tsUknDwBK4e+B7Cuh7qA+c1MqxnD
Gsa7VeKGXEuQu8z6tEWjoP8A5g5Sb+EsV0hwy0cUvi9HRcDcmDx0FiHpx0b8jRGO
wP0RtI+nPcDAXeXDV7SndoqBKKWX0OloiNW2fVQqlHJr2Ar3wQh0dUxO9Ss920gL
reXrwAA1WhBr35CksP2a8ORc2hUeAt66ay5js/SAN7It77vWLJdjpqjfgcJt18+8
F3+v29qC10vr9JxF+/MfETuJNmInqv6KRH67qvyCACwLxFYO1xSCmnYea+1R3H7d
vpU0tJI4Rlm1SwkBdcUPMNVx4JYa7NMH5hnzide42p5LboBLKicYHGNuLfsSKC7U
KZOuf2gkvv/riBiIb9IhsY3Re96is1JpTRiGCuPA7hKsAOVaEMcKpBDbD+WdAQ7c
XKWEfXtRXQ7R7UXs2hQyZ2s8jAgXCp7CufAAXsu1AmxE4QGrjH1tSwOoB13/OtHy
MMhtogyao4vYcDT5AKfTpyF78zlp92GxZjy8QEA34ZicubuYGf0R/GKG6er1hVKf
Ic4g7jMJzA9/LnilyxP05BvWUJTioDtlK4dOUNtUi4NqAWj6bbcJItagtDcFFgdr
cZ+GSHa7N3szEQv3SXKGNpcgdT/W5+lrxaIfMAzXtmtFRta2p7k2W1SEWQz/Ga3H
ucw1UwX5V0STflpXHAtpvk0qv7gHFEWuN7C3cE0hJPZmxWpRHlw75pvKZwtHp1MJ
GXK6yFLVzDIK/ThOJ22rxG1/hGCEoIIz+PkP4i62Z/P6TjnTyDfU01PA1XBLkNHH
pJBeH5fcrsJUaQdN2XSE+dVuh7TkCXvmivHT1a4amO/XjP3W12VelOhamzNi5GY1
NHANxPQ1TTFbAGTGq4LLO5zaDqwXUNbTWCLMznimp123ZX3NEh+BNrlAcyxHpmig
M7K5qWyl3SFHH2dkVgSfEl67ru6yylxRcBK+dsSpCnRNi/WfbziAGZ2PFNvCHOMG
XeoZcYLjNJsN4erp0AViMKANLI5D4XW40bpBstAn9ChP862nD4Wpmt7TAUJ6F9e6
JdB3jpAkpmL5agBnQ3ayFfEoaeTdXG2/UQjPv9W/pIiCB43TTdllpCatpO8ylB3F
eoPFoDq/2MTbgDlGVblRKe4Cux0hfuiGhxwqgfUS7F5PfFJH2GoCGCSl6NmXXj/J
jn2WE5/elT1PZI7UCChXPDiXStSI2rXGcWg+wsAh/YuVHW+pUUKnc1i1+UQR6j57
pJFoqMIIaiJEF9bhndcxJJvLeoxK0C2TgFC+giUbjVdaf+J6tLpZgkpKYQG1qpaF
WmWTgY+vgpVpl8n/BRmgQP6gTynnuldxRDEBbRTugR8bAoU6iopnwBt9sA8bvAXI
oECWMS1/IL2xfN7Rwmm+BjQuFYIkJAEOMywIZ2R92GM2RFqyMBeFi5GOOhcKAgbq
Ty18qgQAOJ0bfARaoQcWfPsGS2JdRIc8AsVz759nzGoeDUt/ZevmToQc5QZES6zV
4yXava5O5ycVfpkbrS/mxy0anRPV+Rb+719EBXdZ7WdNaNTtZgLX+/i8Fh8Cl+YY
ruhu7HbnZ/MyrrhncQz5hJox6eFcMXaZM8m31cY4guyk6uaQM8vA4rkHeLQpIZD1
WuHhwgP+7jpFJVbiHfq4x8zGH1AqvbA8Nb5yZXs4ZmRvCV2kzwws55rJcTGfZOnn
y+Jfl2qwzBrALjaSQUtcza4tpiZYiGOz82VP592acJQgaTLj+qmujstsPZAASNUm
7ttcyZGZQFcCumYy82lXunyxtTvr48JJv9/un66o2YXuQn1sbuEsGF1U/Jtry84D
QfZfyYVFJ4T+IvX6iqDGJeAYfznDVyosPxMDxo/26KM4MTLeNbhlEfMGhe0+mfMn
Ip5hfRYtWXTSfaoxDIWu8qzgsYAe5GRbybEnwqo8RB7h4cikWEg1HWh7WF4TdfDu
ZHyZ8mlgYl5HD1+mT7aMVQ5RMyUkrBFtc5St5vXpYeDqr1gKOks4wigB98nrNl2w
hL/MRbKb3c06QwLjnw8/MoGC+BXGiPTPPbQ76/h0zOslKsyQ0Ig5cY5lpBICNH1D
iA3+KME5OfQwfmG0bXGIH53b/+HYP9mlxuFVoiwHsPsDaRvNbmkCwovvmEUmrhCi
kec2TbkPY0ygnSDvvIFcmWuywxWveOyudbaDnFGPxOWTidKwHPHRcLXIJ8RQGWPj
CzsRt10U4JJ23aQk2esCLagpV+VebZSgDzJ6wRTd4mIEpaJpbdnrBJXakzvBP3Cp
oNkS1BwF+rrvgauBWO+lfZUnPGR6PoyR4e2RS1F25qMDbsDM0dCVwKb2jyDLGnBX
vh8ptHahbIY5N/04gBzMrRelMtEl7IWyFEUiX9sAkm6p9L8tKeP5nU2I8T/d1e8X
1lbbyMom5cA3unb2CN2fbv8iHwYe/LsCwflf3EwUM09D7fZ4H1NBZFtmL3scsOc/
4awUaDh62vcwY8yEJxOlBBZIyQq8sQebiXgD46sCBNV+wocFqfHePfu8CWQqgJjm
7VuL8Jtt0i99z0G4lPvGiVTL536cju0yKIaGUn6GKurGIBqwfqp+ep2azMrL+G/o
l+1Srvb9vIPGKaH7/gQ/8S7+GGcGEc6FJffq+TmWWjU9fdkLldyBQ7zMoruNeaTN
3Ks+NSBWd0t0PH7xnrPBQYgMX7KK5aesNM1eWYv3k5oKfG7EEOdc4r4PrjRx/aTj
jY9SQt8jIsKuKUgjJJGC95mCnguMki4jMeDzy+KRy3awyI5XUo68RP0kjNT83iT4
+JAa4H5AsIE+Le9p/YdhGIsD3Dd5f08eCVAE6mu5/gKjJLyjE8gJd/gXFbPMXqTD
zaxGNTzf4yKXHHWIa1HYfo78KYjaFB00+zUuzbf5Xd04sqh0RSDkUN31DEZ1izin
+r/DSBTPtDx3D0msovOOnvallazH+/lO6Dm2rA6Q9ADobeysL0RYgAh+cbtqIZRF
E/L+Fi8kv0VkZGE/cLwLbelmk4X90zYky1aOqAslzj+ZhxadFbGdoG2CsHcVQlr4
O67K/C/wtKl5OxhYXbZJ1xREvXjcxJmFHfeAKkCb2qGrv1F293RJ7xyjHQ1b4iSA
JAdbAyAiUYR9rC2DWvBp7wRBPR/+Uizf9kl25dSe4jsKbJFUH35qVkrKS0YwAZis
ESBAy8eYx+u4EOeq3A0JEC+H+NYOpcuGMQjAl7jM8gUHPiEiP2BMG0ZqSTxL5idM
F/uYIWNuCcAP6pPT5slOQ9+J3XhCZ/ajlMfYa/u50jIJUwgbqXljlyGvuOuz3PUo
Y0Yyu+RN8bgY7FHUawWi1btwWK2t6mbAU531fT3Pjijiw8ce6CGaHj1/QshEpxyn
toGhTsLIs5fzYjaHWCzI8A7zqLtvg4tElNyFfrjjm6ge8qvjCzsXELYc3ZTbzdfN
Va+OCvIR7pmUX3FIubiQHn0UDoexmwflXKDrZaX4AG6xKSXtFhJa/WWatiq4/jBC
lcSrcmTCPstXQu4QOD3ab1mFhiUuB72Xivu6cU7Mnn/t4TJHzy9aYZ7KVsXHy3Fi
Nk7UcVYZvvtgYLhVKSQi6HtfLEpdpa9ez4uLPby8S45emBRcJ7qWaHlmDKCTjLiv
qf+y4Qf0OyJUHf50yFvEORwaArJC1Anah4utk5pektbnVLRElOzVRxuP+qVo4HEX
Qv2xEwjthLEJ7YWWX6da3d00MZ+eoyv/D64cGWIkCNqzO6OMsIgopZR6fgmON9VA
RqmJUTuP29TJBWf6hd4S7MVpjvrnPnggENANXjh5w7x1H0s5TfRZrsgi3gj+MGgu
BWm/j8xeVSV2wbvJEMgo+MV0LcxrVRqU/EEjh95aLGvdIbfRB8Q40T+LUAD39Y/P
vkCFkfVSjtSpgX5ucEJYhXLggHJXkjhVsXAZNlA8H1G+dl6lm3Ll411YXNwZMMPc
SVUcPKMfew9eXbYR4gJ0jqHUHRgUpUqdDsiTitr67fOnhh97SoAlR4jE3c8UBYqK
2ZEcvwqMPL4wOmt8DaBnc+431y2sWYEeKExqUgAhrAWe+tGGmX61OWE/Yz/qFVzJ
huA4Ol1dW/1+HwHKQWGdwwwQh1zvFfJnAZNuR5No7iJV/u/pQl63Ry0x5VAfD+P+
51J9FiVHAbJwqhy6zxyGx0/luClK7UBY2CgD0V9UnxaPaEQv5uO98d5UaD3pDVkP
EpuqEKT+5JOapdY8SEHN1nL3CX0EA02SUXQGIabaHyZXJsqYrncprdBKJ2omax1z
PAL+1zNPhHv7mJxbFK4RJkSMDP2xod7UJVdAKK1aKttLRKqM3/ml0CIiWkblreey
70Yv8qNzicKvVY54/yMqlYji9m1FjtZrT2jL5EoeIhg8GPdFqbAlt+Y1yhsoB928
g8hhOhFdwe6G+AWSmneZwH3NQR0l3iYyUQPWctOVNoFpbcCzpnyTbv4qoNscrCuY
ZjVtOBsy/LRmGh7CX7kXaGwQaskmzCdZhBJnusJTE5CUkErdXrBcCFXYBIQETR7N
WASnSUATyOQ6MWcxWVDnT8umhlCj6EfHWvOMNl9fwJ4Ed1PG3kcZfijvk/ClAK/h
IKIo/jCcCwhN7V4zb/Yu3yRpRiNnbiAfcAb9WiHYGBpOxoaHLO1vK/2bgfaB0S/n
xNScqQwm2b8bHCHXZGI3gxT9qVewCEsNW3vidypvr9iXtNG1Z/0VWDYAixHmjM12
Blt9cnYRj1vj4zha+SJIHFp0HmWebrGU7nmf438X1D4ELtN/qeVvrTn0livkRPSI
M0pXk9QM7O/WdAsseytCRD8EdWEICfitckabkzGN1v25TflBw+rDFiRViHkY1wL5
vwIAG0rTxwCrppmdRGgpvSLkr78sJRvKU7N4GzqjqJmX5PwaKgIzIjNLDiE6t4wS
CPsHfNVC9hrF2UQf88NOtqFL2b4952hMe74LAJnKCjODjvy7Z0nSi5ecNNBoMBNu
KFskFUOeOZwJydQhckgiWSVCZl558lgYz1mk7GThjVmzsJCba3m8lBG22wNAKQ0c
K26fJO0rmtKdaRsj7fGwjtd803YQwhG4l2JhF+36qgHezi/ONhElLYjbnuEC8mtk
Fj4a8y9oKTI0Pe3roSZst50ujSyI6u3CPWKFR5mUOTPe2M1ILWjl3L9d70lR5GWl
9pcEcA2fgEjhfQBu1cL8iqUaeaWYyMniDhaOMJSGXdvQ0kOzWghtBBM/FOEbBXEJ
PIrJK606o9P+iA8W8FAbtwC3SxKhzYvpK2mLblrsRonj0r0uHoO+IUbrLm6U643W
AlwTuPHLpmWz9Z32lwdp4zJGeg3iqFKWNRyvJ/ghNmfWhgP1tzpoOtWkzcnKBAwL
IHwdwhJClrMvUL395Lz0bZI6QB0gVcDKwRn1BHkZd6571p/pfsPwmSK5hhzVqpTp
YOz1M7xMog3Yh+gpyMxiF6Pgy+Oc4PJ8MgJFGaQw+iPYeKeY/jbvh+seILp8/M3Y
v8GhMi+FVQHBprX03x20QVg3Pq8LI4Xq1GExpeGemrq/kEvulULlqjszx/BdGC+0
+2t6ZtYKI5dKeAU8jGcecIvN6cnFpZpHzmh2PBx/ptG9SQoAOtQAFtZByUB2s5g3
nlADjC6trCRlfD+y5N/rujwQ2dn8S6wpefK8iCAgrzBnmPzkOJvPGvJTKM2c/Tok
E57nQC5hoacJ5uScMYA49ymetS6LwsLLZCMSG7+lsLPz9XYrRxzike8NWtticDGp
QgK4ym0aob3u6HjcB64ja+vmDktuLbrQyaQvSe1ByUVtVNllVWgb7YI1eh5fDPvJ
8+Ymss5dJv6fsXT0vSHc1c2IOEGsxaKuqJH1TmZABX4Jw6YgYvsXGYVHZLEHKy6W
engUmHnITtSiVBO9K0Xe1qapZwb/+zwLhLJDENeNNXaiFaaGrzBX0V1Ht3CdSQ3B
y8SX6ypuoubP9HXOve7aPw1KR9PLaFPGgaOd5trCexR0p9rk3YpaWE9xFCqvj8Xh
iZThn/fz1jBruOiNy48NjlZxwv3DKwewo5zNan40ctwI7h+hdkZtj98HiTZxoRSs
C4jxQtPyslL6hF7cZVaRwUMT2a8E7w/ZFTHLBBN2tBnXx7sVcwPAFLbxIVFVfTV1
+p9VzZAqiFo2/229+23yKegxfiwpGMMBEitlXkWmNGnbKX5RJJuvNoLZYBR0Da/k
aDtsNxuiFl0lFeZUh81kCSy87N5aCeeAeg646QBbr+DBo84tpSyr5pIF7xQVsd72
HZ9c5aAm9KMHbdhq0FSPvgcaKKFcI7i+utDvh7i/aaG4k4CCnntfw0TKFtMUydz1
zqI+oeZ8ZdLrKUL821Sm6yEG1yvJ66qnZaMTc7/C3TjawnxsZbvbOjbNLvvrc4sd
tQkOk0Ob3EMSjdc++YvuzVvT1pDQJsZde9B+q/MSFLKJzV7ap2DcgOa6fVMd/Bqy
yQ3uVypvMmfr3GVW3k0pZtaE3S9I14eX9h46h8lnAP57RhpXsqIHgE7Lh2r6xh/0
fpMvFHkUp7NOCbc5xoLx5CYs9aIKkABms5J5/N0pWhRcvEkkMwyQUbcqYWW/HvaB
ZBFBoEEaPLj9kLjLtFYYRkEulR0BKr9dsxyKoEId/zbym510sEphlGI566cAB1a4
UZV3oUCVdaZ7EAPX/QK9wGLjbVuMlkqooFmiFyrSgW2p8sokejBqrQOlmpt32fM3
AU8XQ7na1PiyOVkeocqUJwZ7xpfpp27v0SWVIAeb8dV9qMHuldPhq+5kOznn9OTE
9vMXGkIW1iz0nsl2pCko2BuHDnbmVOLjIGEjknJ8QWY3U89BTo0x921K1tioefS5
FgpcmMKfqS9jZsK9QpShlDNdF2HpShpxfBQ4kFmgfMjAlkj1CIl3dS8Z7UWJjx+L
MoiEapqZJbtli5fUr0rpY6KHnqJdHaFGiVkeOrIAR+sRezF0seY3GX83q011zD7j
Z+QtNQjnBjoVfhAM3NmvS4E4jeRspyPgk0eLdqcZCQPmk0kbaPUwk5qy2xKxqoFk
SpD5GwDY4gW7i38Dlg3uKHuIG/uijhmkj7r6UwMnlEgLKsC3DHxHZUjc+419Cewu
uBkVgF/BPMKfpJY8lFg6C/FgM48HP4Gx8cRvQ0qS8lGoDsfttlzj8JzE7ZEAHBxR
qPZ0e492HUgSj890OabkR61iIhSDRycIufiNp48Dy7MFFMDb4+F/JJ/yRWnLyL4D
m5L/UFSi4NIqe3agLhKW0qd/pBmAkxyIygIGvCQ6uYno8YUqkLlOIjbDHW8Q/Kb+
u/LNN9WZi8SJBaFSADzCOTbepqwMZVd1D977hykbIrVy8700C9i1F4ZiZZNhFuAB
iIRwv2+h9VaRAn4/7tv9migUpFAeYQRwbr1r19KUWZB1l6hOR79bmUjnKLcUkpuH
QwD6CQ/IArm+GBa4jGgZjupsWBvEg/PUGh+6x/FeSQMYODAiFk7m53Jv+iEIkFM7
VXRcbzpJ2lr1Xj4kbwNSzEdA5QkGEndm3TWxR8i77Nl8hzWWv8H01YkPm3MGjg++
uwhQ111BOVL2fRFQu63YLjy08jpv0tBT6FGBztLZzZ5rcyhzwdTzuDFmBp6lz/X3
ZDCo2a5fUSpP+4sZLeU4GpONNyPfIMB2Q3eTdWS3xVGHeF73pG8JXP5g5XY9OcY2
aw+iySxYTE5DHCF5gURSbnvqD+hMqrXIJA3c71PD07pdpZ0Xk+Gzp0eaH2TVFk68
/5Wm0kdX8q9gtEeHHeAyIHPtSD8se7ghhpThbxIP3hRB4QMgahMDiH6uNuBiPDnz
05cUBg+XNXwjZjX+bajfRQaj5/Xy8klzUAuMHFytmEPICBSNgagjoNZ/HPDFNwB7
08yOgMePj9eC8uYvTDaKh04Gtf0oCrkQfb68V1n0412vd7vRcweweIgaO5RPMTVB
R04xcKGBPIdJF4Q+8aOjwai3CLRooy5jLlP8ppudqOK3udpWI3mXLgUi9IHx1Hdu
XNcI70HZ4LZ5twfaO3ikJZR276INcQGnF8RcFdHU9xS9M6DGFKnzUCjqVuE227px
JRInnuxYIOnlfBq1WI/Mclbp4qb6tlHN0lmpQ0bty8Z1yWSDoo6aI6h9NvWoaWzX
KJzZAYfBYF+bStcLBxyk65KJG1N7Lbno2yVoPEaOqSiL8uzlYhXPXLRlRdcpWPhz
VCK3Qx5Xk1+MWhpsCmasaZ/UFocoow2hiuUy/JjHBGXr+fWI9JF4gCtJ4pt+R0R9
Pu8zV7Z3L7W+GKqbcxy/7+MzTXaLneOO19AnKsvfQY/4WBw1xIZ4vK2I0fh9e3FU
+puCLEg93itKKWW0gLPE1TIaA3lObaGD6CGcHxmMz5ya8ghlS7ediFJCXO6O/7J5
bH9QwDdGdDjX/MGQD00arWjhWzRdlvXBgs873PNIg0/YOpHOTOafIfpLMFolmpPH
6IgW2ORRHKs27zQPTsBQvElPa7m4wNCXqylthtiIoAmGY4VVYZeqtR1A7urDb/P2
y4lDuqsrj0R/L9A8YA65bDXJhR/McaAcMCIn/0C7aVaPdA6KDT5ZBAsoyJQOPxq6
KJ0E7Phrz2AJwT1pCJQ6PHBq44Y+s87h9qhOgx6/7LRe4XAaShNOHLt9vZ7T6Wjx
m50EviTVeBuY124fay3wNgXrALzugsuou8VPStarJhSd+ZpQPM7JqWTM1VEO6OUs
tQIC3wIewUutGkI4SIToOrEMux1lrLjD9UxGNcgcJlLxZFMdx/lzxhGlBghOtyLX
uopqRcgXBA7QEGala5M5ib4pG56qbC9XuSJxzPjaPxxRmeq2QDrbKCRUsCi5uhQG
eldxA5gMcJRQMl3PFipolAZCeJdsnc3OpT7fcupSz7ispMAreQ2Zn5gBHIcDAFG0
kud3S24xko2qc2E+aKN1uJnhei03HILTft2+qJ0UBPgCR/0GdM3EGYfos6iC2GFS
zyoG6pI5aYvyZLDFGyx/wPR/mdX375cmSAD7XXzMPD1D/OM3OMvhlxB1hkFshLiy
jcOm+PeK3SpJunzTqx7saJI2FUJu2xhMNkKAopg1Xg5UAVpnQG5DJWDXf2vvlhKI
3whSTuwlBmhjxjasWcDuqUcUhUsKD4gO7z2jvuk5wWVnahCf1CTrSanHesRzwt/G
CeHTv/UFOJ5o91lyBaEcXYY2T0ENRTf65ttLK/9SYp8Y9/cbG7esEW8MtgCp7WYW
SRFa1B3Fvrn/VQFm66JfZqs6aZ23TRn8JB7Se3pn11Y0+qFoCof2QslUvLC6M9je
nuUKjjCQYMAUIqkDnxBDW4dveyu46Rh3dS+dJeECl8NVzOyPK6lvswUio+4sZHy1
W7lWoOugke/jnb6l5V1DVowydXzgoX9GEk80/TVETvuhRx5NGFlVBGNfrQy+K0qS
M7i08iuY4WgIdnnHdXa2Tk46nFwJjrFz/gZ4ovHSkDcZQ8LVvNPvfrAhKJm4fCWD
a5W5ke5SaDiS0RDRhttrVwf+r1Ivw8KeAkDGQmMUbpC3IM4LVYUAEe7IKqsBrFlC
psA3pl3ZFt1h3isYqOdiY2nODkUzstx+LsA/AZbGkgTlBYENr4UPdGeWfWFivIPm
d/UKHVQjjQhsoj0SjGJJLuTadFpOKCJijHm/ajcc1O3Tg02PqQ3QXAvZ11Sa+QCP
c1lK4Kq9CTtW1jZYUysbSzaAo4b7CWdvm2NSRa4DQVm6996pVNjW2rxVhqcoodvf
yZGkUtvgbOxpom+3IiVrytKPTM9rnRSnu8aIRTiq8I3Pqra7gMMlw4dJMpYMJaRg
rKOCvUSu63h9FYc9Emiay8ij42ZHOZ3+hSaNIhYSOJV89SlRNrLWcSqSprqqKsRG
ZN8d14YWgBZDmKXrtHRcgbczMzlUR0xtom6sOFOncmNJlj7xzzAHWUs/EiAu+J6U
oZ/MLiNfXoe4lPQVoe7TpPJDk/hcaivuUipsn39MrZM+LRMBsGwWzVTE1TBQ6q4u
+7hHQjhNVcCwlHPNw+CuqA5F5R3pxCqYUcxSgDZwXbxDN3BbrrHG7RJKaZyMaSYN
6kXbIS46vNp1YNGM/af5qRGeJFbsLi7nz+G2BOq00j318tlh2CO8GeapmFOELztL
y19ntsSIjIBqcnWHzOcbT+KUWgtbxL207+FDIQ18sFQwD8VqLsncyaFyX6icUtmL
dnsd7GcvPZLgzqVRllYsnk46bvswnHUW0H/cHnBAxJEgHn3ZJG0w0Vd5gzTSNyix
shy1m9M2mBENtmnXi/b5FXaG1YlhVDdbXgXfxpKxb48DYsvfLiCe8TnF4eNjMkkx
8u69o2TeU7Meg+ANw1sqoSQ0xxtquND0Y5eWETWPujs3u1XgsgtRBvNcrgTjpaSn
Ec77/Xi87SIfPDffheWbrPBAoNbgwcR/bk1ZuiZjbDOxHTlgnz+meuUmZL82n0up
yP/oR+v2TIqF45VZqaYWroKPbL9vZ+FfR5M5lDR3UYM3FHscyGbQIaKmtgJURu2g
JVAGCDSnVAr11lAA7x8PpOgUv7aY9kQd2QoFEPJx/P0WKTh5qa3jCjOijh/XBbnL
xZHt7/EJM6Wp8t2r6QdESquBz7xQaxj5nzkro5sr7j3GJk85YihxaNfmKF2Soi0L
N127ke6er08uoRciaCNE1xO1tnZxcXDVxDjsZ4udrhF5xVAAyC19LsX2vOSku8bq
njlr4bsKWcaRqekSCSTIPErgB08WZUN1gZKy4cLCZgk2MoSg167/uigp42g5pT3+
n9ROmYMxJvHGd/dio8tghJ6jrPx2B3PRYAuJEMoD3phw2w8Wbf61CUKEP7kEki5l
saZahvpVb9H0wMTAvpi6Pjs6K6ViLoXZdDrDSeaX9xGvcpcfYCcgGrbFI1R6/Uzm
1FcWOkOx8JusevymVN0OLDfE/FQwm3MRs7qHRbkbmVk3T+/WtSg/laU1PVt+pYvK
+8tQXnjZL6FuTvKdHw9wss//5WeJyPM+qvtpCLM3uYo9nQune8ShMfB6YDNAr3v5
SJHhcwH+ePV7LUEaVVg2dQoftnDL/b4DyjaAs9uE/6yyiYPezDANdQbTC5bCKu92
kybNkRuqLlg1+VoHfLLjsaHalq8tVXdRwbZdnTUznudcpRdEqzZQ2FTVj9X3CUdO
iu+6MoVLgNqCuwD0NiR/dWAi9JrLFblC6qra1V4ed0hUZs+6QvKS2ZM8egdR+vYR
na72Tb+vAuSmDd78iezguAKcz9THZ+JTY5I2yLSc9z/Ml0m2/pD07lgRySAoBRzH
kASP905PCx5yENHrzVMGkeJZZIvJo7EbcIYvdkMDhJ3vnpCgiP2MJC7CpEOxLbDm
MywMJxU4sO2Cc8/NCiErXi9O+QOHvLXmKP5HOa+iTSlacjH4YNkfhH1OxTW3I03B
vPvS1EQtizGaYgHryrPE9ZKvHjZV6g/9nDxrvun4Ch0rQCU0lz5iU00yzcZiR4sc
TtwdUaQISrQbieIPEBJs4HbZXZgicL+HOFx0alDQocvryxZBGrpbTaPjVzNXNfwh
jskBJt6KksV9eTtLdqGuHGp4YOuj/plJ9KiNj2IM9e1ejQKhn5TqyY4g1AX8HJFS
Uzno+txIsYAV4TffX3ANJ4aT0jJE8+vUHE/4JNGe0cmS1ZRFg4ikI6s+4EubMbdj
sC0sCTclyUYBP185FOLpd/FuT0SE+T85u10hvkthnTdyXDXX8WCLu0CFb5BsBzSs
+KZ5DYafMVQw/Uq4mTX9jl9g8WnrfnCyAMImPFvrZcjnYcPA9enecQTpHZRsM/a5
knt+kxxfm/LH0DPrJP3oVgFKdmwnsz/6szpuEkUzlxJJU/jf0Q9fPM0UtDISyWxh
jvoZPjzRxo457IqhhPI9QS/QOsqMu//esyZa8OED6M0W8oWiZch0OaG6ZpBOlemb
zJMPzfqH3c2tGY/lolm+EvrBTz3Fk0HNj/G4upS20Zq2tlpVj2SNgX5M/dO7tMSf
czScVo3l8JeO1Mx2REo9f2CEiOXDWQP0GXS8tMDWOccp/I8AdTkUldp/0tSi5HGA
+wkxYGXEiLh+FXAXskOwcHRfx9rsouCLpjX8mCLPUeFTFljFM9p/SW7hAOO3PnXl
17UMfgGGOW+UV0QCF+OeRJQNaerwAHS2mL+3f8RNMPN5V/s33NTVRXKGk77SX9xk
eciqOKCiHr69KJoHhod4HuYalKPq3vPnqn9O32Yux/CPWqLzPpDSNkQoBjJvsSkx
535N6fef0VbBBzvU4vrrsp1QzCuWFLBKnP8LYF9ju+QtDMpBW0AULxp6yvsyrYbu
rRGgH9ozHnVVV9t8B8sibLdO1nsUEpWKLVjdayoyqjAb6PMwCMmySGYthdiM8TLy
iBWMAl3HLw28oUthxEteU/IrDXh6+RGi31/0Hhc3FMG8siquW8MGLSPs5s43Tp8b
6de1VvSkjCV1Og+oBU3lgl2XIoqkzZyzVMV4nmRDg0PQoUBFZGhtu7pKqgOXZnkw
22iRTfFmnJdAvBh3XYFAWkOmARgL68QDpjVFMP+dwva4KcTADlpJwKAOVgat4jD8
hUvXtutni63gRBBBXCM8NvW1TEir3Uf1uyNivIvwNycJ+CKeF04JbElEOGP6eGep
J618rJf1r4WD/sMW12Ah5cco3kxTnURjfwZfXXiSkWOSBjNTW/G8M9YLp1KIxez+
yWKnU6dGvW4LeTwRtRNvRHwZB+cgXoUTNY2hiT4cfFJvXlwjhYgAcbWATV8VTQLW
17d07b0iMnGoYXoacLunH1NUsT/zQnQMqfp1Lp9oPqpd0MHR0AMxiTv2LMg24D04
Wmfr0Q7StUu5LGiYXyVu/w2/khHpRVopC0yrbldjl44Js+b7diDglf6d9ReksyUv
9fO3KyjkULBee78bGN7tOlj6qSqTa3IaDnwxwuYlHrDUnZ0/6GaypMhkC3+Ocxgf
O7er1bhrrLd8V2Z2F/iTMAIL2Z7NSuQRNuUp0pYcQoPOpW3MYf2NvM3AvKqatA9g
8VhFzRA9HpAUgfqllKsaF/jF6fxVURvBM/ZiO1SufnLXHRqR8gI3Yp8F9fUk4S9n
umKUn8U+7NBtHgdU/UZvO9H79nrdGNQ5SovJUDCkzythsTeW02Gsag4QmcqP9yff
PcWrKfhsiy6fxAywhreZR0wMu5NZb3YrS1YxGLX9RwEFaIMDmLrRDhYpELDjwi2z
D1K2ityox2j2QRc3r83t264Vh8Ln6JmsavL/Y2ZvqGrrceX5pk8PSaO3XJqAaPXi
7Z6zMajGAPXRR1S3xOrpYfmhLMDriT0Lm8hku8aD4Wixi4En7PEIJVnfTXFRl7uJ
NeVJfkSfoTx1PdlVeYwt8kUBkMV+TsWZ9WUJ1aPQydkIg65eG4iczEB+1YqKrRj5
Qi0wsw/F0h4yC1VFFoxsWUW77Nnvkftg5n26+OQjpdqK9vBGIpW4AaEVaRYlprE3
IfPTtvtCMAfFIgzXr7fceq5W+hN6U8ZJnK56RQ35l8arMjOBwZOCxzgVJ/+WEuIf
iGmIoyXg0hRlfdk4ZEi+k9gDFFD/7kmJRjpgLSP0UTSAhWT92n1gIVytANNggaV2
XGj93YmQj/TdOkACZiXOhkFlxbQRXyrqzNbLZBVYzfYNsb0JvesWoHmi3lz54EMx
VkkSNLJrcZ1iSPkFjvTRd2OVcADyJLO5Aj98g40dUYgB2V9nit8QhWMvoT8NR6Z8
ouqhxUQGXEn1e0r35+cmRhJsA2q3//K1eUzUaAku2DTjVxjVSVF+tJFD/pgonRfb
1tsd6N0AZfxk73GkoaVUXendXvEYo1xqXfQ5MHDdgNrFMT4oe5OHqs23MB5Z3Aff
ahcC4Xlsga9dc9LHUMG0suBGP/wC5N8OYCAQFb5V/as/hrdfiftxegwHlzUVENha
JJXhQ7t69PRfjz7AdcGVTSVploHz6e8ayyIeRRYrt3YxEk6JEB6nrI5DqkZL+YNX
fJ6ji3NImhOjhQLKZElTcGKQKwxajLfo3bbkgeSoX8cmQaxWmBQhSorLtFOk5vzF
BQH5upVLS7NH18Gi2Jxvg5udq8LBLonPbPhBDEUV27hBKr+akhVxh3UNl/kand2U
H1RzbnRXimn5R92uniBwbml60uSJkCaGZAkjPhHZ5eynsG3KVmyPuar72JJ67GY2
0sArNpFIgByNXsSU1zovsSpO33+lXt30Dy3RS25uh1vuGu+BVMKi9yVXzOwnqokc
eNK8CZWdiU8j0snnSa+U9vagSiBb+EXalems8qj7dVH8MDMbI2xHYEJgC6f6kxB8
/CoV+JPAxxetLOEkurw3DSH0WYy8wBQYFjowzZ/wbJtvI61ipk54t8pKdIuAgt4O
T2E39a3fetyFMjdM44kvn5qO592QT062/8QYPSou7EfCoCF1pFczxCuszMShet6c
kbMUMpm6azc9/O876FxWtyVKYAM/Jc+cu2p+CDkKn3rLqw0iAJws16h3kI35d5WC
wdom89xgWWZTS40IsrDVIlE+urA8Myhe3d8LElEke+z/5X8uy0U4SMIZuurKs5OW
XtTfg+pboQeeJ7aNxFKm4bDDA7FhirC58bzvLNmtuTfh7CbLAu7cScA2K+dLJ/nT
7CJ+WwSEKllMv+KFe+gzm+eVJ8tO1tJSAF+xYaTmNH2SP65E3n7eKs8fKxnEKUeL
Mn07PnxLvYfNIiipXn6jahch7DQi2KHJPwiaUdHDSBzcFXoMo6MJZzpxmyNDw9KA
8afnIl+MRMLJlTa489Vq1fLilwIuLoUDSvnIYEugzEEh4s37G9tRSD9K0N/0iZsC
aeqkpc5m49nw25JV94hJyGEklH7UmT/pKzdB61J6/wtKHUSG45Fc7bY31bXnaVmX
YWaTJSHYchN6fFv6SmDyyUokXpfBRjl/HzTuzu2+pliZU+L0mPIjIT0626n8QHaI
GbdiZVJXd2D+pj/Oxxru3x9e8KDnyXYTXNTtAVsti7xkvCSAkORteF7RVf3mz23+
pItHavcCqO1UKEGc/3uHI8owxfCfzAXMy4KiJd5VP/et6CX/ZUSwdpLy5Qj5ESan
fUu0/b/7D9T6tUSzfK8ZwEHiTpLImZHOPm6gJH76aZYI1W30yQNnHMnL/YZk3a87
UsjOLDa/wKOJH+ZZn7LDfUBnb0APQ3WyrUodMRixKAqFRQQRBQqMNqJ9/R4ViR7L
LpXMacDT6eMhr5we6fcvzbYw+GRy2KR3QAEJCaDsZdDU1MwJrpW1yHO9E6Ch0Pbx
I0FTpSfVvXBGnrsqZz7byxj1BbHMOqJ6PsSRTSqVyzs+X/xeL3MhdSbUmQQGzU5G
uJeVkEkkbzcF9erx2Z8u31W5n6UePr0BG3894eWszPmaS155eDiBk/0zk2fKs3sn
xCYcIFHJm5VD0gPR7x3dbJ76T9Y5F9BM/VjTKlCcTMgyURWQrT5UbKWFzmeLvFcT
WhaAaIvFqcUQdG/PVsx3PQ06a7eutPqE3i4UOcbZ6gKPLBpH619MHlsmQTzdZBG3
fFvyKmYMYsgW7r24dRodV8Nhf1T61EMbsH7fSQPyicw3fhdhD5gw/BegZYbi3xLL
Jh9xZNLPz42k93ekc8118Xqh2kBUSuar2w07h3Z6llS6GzrUzMuJjW4IL2IKyGP7
M7Oc6qDeOAGdKwBtBJWs/mTlzrYIDGaqf+PoD3s/g137HOAoe3tSW7ivH4WQdPeC
Sa2ri5wbUp25WWtGAi6SqW2Try2iRtqjBKhe+RgtT3aicZPeGy+JUAOi4gOYcike
6Jnj7eZuFli32IjAEKEixAjkN6ZK2J8Wj91y5EDuMUL2TyGUTfxJfk2FABmTfJo7
LmhEPL1nsr9PJu2/s0yNqroqWhiQ3K+p29J0PiQAvAT7VsVM7f1Rj3zCAolSzU+Y
G9gTwBKHNWJVLPur2goiUWO3lhW3Td4wpKSzE9MtxKqpATzW7PnyuGhd4dtOxqu1
IFu26nBkVyNSfbSJl8zIWoWZPYVRpzY+FE+KMyOuXHdnKo2VVkJootS3KFzELbzm
muP9x0HJLbwepTMb0XUYLck3Ca1irVVTERwinRhlkQTOfOYaKuaxCApF+7fpgj1g
1oAyUYeJe6pzzcLYwNYhMToLE80Q44Xh21xljraRtaWZd/P4tB2byH0vd6Z8InsR
3cofQEI8XJmzdbfnj0L/2XPHwbvsQ1pxHIuRtIqCI0ftrOSNZ4QXmZha4YzW8Yz4
iaeAMg49ru5Ygy1d+G8poB8271y2WcasZur6Qv7QAWhIp1evCY/4AukTmfaKlYF6
VcU6dc5UeoyPoDU7LlvDhPrAzem8u3MWnc8iQC/Y1k4CMqqOR3gXuRuMbv0S6yxQ
/WwaJ45pjt0sTYrIY6k2BAXaT6CdsAvxsBQZUVBEHptGZSx0WPqs1m+Fv8LGZKAX
QwFRTqxgjZ+pB+UNhjZaGqttr7Iuk2QmhH3kVYyUZNcGFAezt0vC8Mox83DCbfyz
7qaqIWaQRTmc6uIU2GsBohKw8FBMGwbuZ7vlqwF7h4z7c0IUj7/VX2I0w7gxiSgz
5GS/rswtS3x50cYxejiDMyy628heciKjFL8mV9ejfU8SGr4XhlC3pdhJlSAsBDRZ
KjuFRhwfL4jhD6jwmQ+0Lc9+hPDqQKo9mb8K46yteuVZfdOGxMeaECGoPabCtSED
/8phVZDqkW1v9w4mr0LvtXQU93fyKmDcvqXegXMB75Kz1dQjfOL4v3MBr5EyMKcY
fURM3FN5v9BfL3p0BeXg2jYkv1NMfV1mrxSWyN5TwarbM/l6nKgCA/f9jTFW3L4I
/oa/JLlup0XtnDzFWCYj9Dfoa+VX2yjP55KQ4nlGFhVxDVKK/isfGNMK6YXE3fxe
6oxe5vjnBHEtG3jHy1ggNlh1sLOLe0GG1x3PaYe7gQhxuCR7yeu3QOcRa71yoTlg
cpmXGzYpt/yntB7Wc5+7Y4jSrWNuOd2VJI1CSh3DhWnRZf4ksfOiNZyxH0So0kWt
BtPVtaPOmBOmVIUCOs47lseFG9Ray6c9WyFfs2TTxwBtQERmRPi7Ks3Cv5jp0Uq3
hrqbu+1Q0o6F+K9cnJUq3j1CPseaFzI7gURAT+7BBm+4hfKYf/Qp4x5AD8r9cxo/
1lxsjIglIckLdsceCm0RdYu1h0a/YsqAIK7oF7x3xyz2EO8dJzFPkaeoSgNb2QXL
0Ip8vMUQfq1T9rQdZuudOKmyuisDUj0HmISeybjSewepsAU2yisE/xRQW0PXIZaP
g796NYRQOVTzU4BBm1aoVE/CZvC0VdI1BR1cgIU749+Lur7VzTg5U+ndyy6CCPXq
CCxiIItH7DzMcRkdj5VmjI21qTs9nCYJf/nhT6REzIPUNJZu9cVWomfvHUAfePpe
PLdhmbTYtpcw8Bel9Rx3s4OoYt48e1s+ZzhJX+K3qS5w1aPaBZJxRY0lc6i2wQnN
d4K+L8dJEGvZO+yh1QxqzJ/UIZ8T1p6awqKylrjkQuprWZSwWKPirWaSnuaESGOi
/4S75qa2Jgcvuy4yJDq5972/fx8717Ta09zWU3p3od//sxw/sFHINVwYTAm/S2Nu
c3RVypXWvkhHLIV+AO3DMIaFkzgx/IeKoFHK1q5Xmw8/65GsFhbsBdwFTgYL8f/z
5JrJlCjAP7BObZVRtyio9WVD9WjMVoKRxSYvOmilaN6nAsVx+KEuG8/CFr+b6J+7
kQpy+OuwLEZheiEmcmVN4gmWUwpooFwVK/5ncSEKwwgwSpGguOglym+MQOnzIUEz
pThI7HjRkmZ08wY+YLU4mqK+foa9kyrLKJrOYeM0E+jxUNKyNeTp50xS5ViCx6En
at2/rkgxZanAr3foyJotu5rVgAxXx61Kj3upWUN48jIUU7Q0/8LRSzLU9RJ0hcx0
2Wo/eIQqxwrNxmp30YZ2Vi/kLaE5Y+YvfCLP0uDCRRvfln44QYrxoGpsXXOWjXa8
g10aJdGFe6djAXZsT3JqHdxf5IuVl5Ejzcq5BmU9SB79ZZFV3dLCkBY202dGLfDx
oCtqkeNPK8NtDBAyG4looLjwjkutgXWFJmY8/K+jAps3tQCJkH/4g0gvmZB4lnCz
jkZ8vGk/lzm2ygVMRt8vmD4ZMHgyPzG2nhw0k0FffMaZemZmCdKn8XealwUNYbyz
LrY0ROroigXrAC0q4/oBB5FlI4qLrh0YnDmchGT/UmxQcqbhlDPghMWj5i9nz4Gy
TUR6a457jNx1iuc1xPYbu7bsGAJf+ZmYM3EeKjOpRhz/edMBOSxyXYKPP6nbSIsr
aPsVsDwoLc8hYwIAQLt3+RWBAp9K23D3am/YWrnOAp02svCioMyofYHE/JpJzg9T
PaBmcoOQzZL7w7RZ0BBupmGeicWejso1fX1NPg5E984UB309jvFyycEIu2y/TJHr
M1xyjLXm28kT+ysKGmF4YIeDikQoCI8f+tU9Scw5UYAApMK/DX0Vqs8+eRZWZNnh
mp/IbjQsR8mZI61BF4Dhev+bu83VCJRyfjQPEIyMNUk/0yP/aEHTQuKU3zfg1Mw7
QiZmnw1hjyKZCkN+z41hWfft7KxPUZGLbxlxmGKaN9nHh1aUIwNUMLicBilH1vsZ
zHITzX67KbYbDR8DVWyFif+65pmQfnwuz0+FkO3JM4Rb39UpJ34g4gYfija0chew
5FhokQLQqjAA/+4f6AJVjCzzpe4mBdOZaB+gsAIMpySc4YbABan8pfF1NiFCpDtx
cGdkVysq/H5GVJ/rBfMecb9AvK1dNg8E9tot4+4DI8UPJJ9AjR48lYiM5Ex8W29U
pdULy61pEE+n4sjVFgG5RtEr44tKs0Db8Ti51rhGpdph+bufUGQCnoVkGHbnHRzH
rACwraEpIz/3Q0TW06G1luKrCMGrjgfqz5sjf6JV+VZXCe1Q/Kja61HMACLlr01K
jsgkuHWvzrIZXcLf7GG4ccDVHb70kiIANSlWcYL/FS4BHC8pIvwhXwPCftRihcr+
gzM6rQos/y4HQPtLaWr/gaQLmj34bS9JzraMKRylrULiJRJYXFslz0Otq7+aumB1
YXYr3lGEb/zQJCRGkDgfvAdFrFn41+LFNGEoYNxozW3Yv8XtEbzJYMICt5Ra68bQ
vr9MerLYJfLWXdEn67nCw0XX0MJNw+KKo8b/F6g98ARg9BBQidohoGf1GsVGoStl
XS9NdYOqMqQZDq/EWX8i0mNNoHE2oYnPIG50Cp1iRwCnukW+2rRI8pisNOOnZOmM
eeUzROyzS+IL44qQaQRNOWnkX0YHrIFGp2HOKPX4n86hLlQpXNsZiy9vzDDYN/rX
XPH6rZXYM7fGGI+qtmE3YgSWh0EZw6hJnsjFnvTveILQQpTCdJgFJGXCKS9gPGzp
Q+95zuj4ZKUYT+54nT4cqcE9y6OTnFvgkkhssUHfBpzuyNOkHWvN5GEfM8dDigtM
dLR2Us6Z2R5qflkr36gY/ZA++yYulGfY7+pXuaT0tCmp1Dt+3eBPnZkQ5j4p1S+8
L95onGVRbV77nxeRd4oR45JYHwFZ1ZDbruSXud5asiJr+AJBZsivl0pIKgkSoa+d
h5jWiH1em7I9IpyudEgSOCPxgY33nLugU89YESr8E9rbCPpPI3cz6RELDL4NpoV+
+jA4geD+mMY0z0kmrSIXKKNODoxGwt69HVrTi5CdHE+7ElhZxxKSpKh3TM/Fs8qm
brEEw5P2Jd0CB8anuJSL8TjXsn6uA+b+ZwbC3p63cMcwgYRtyRJHZV/YVKS16izf
0AtYgcJY3DENjjXOJENBpBB4738h+4qe0gWarG3BtnQ2ZBK+e0ZjALZ7Zoir8L4n
DaucPrNObDFkPwulC0r8TZdgI2IZpkO14dS+TEe+3trZj+1Qy5VB8nSoBv7u7pJj
8Vodn7v/ayFnZhkFq1SB6/uJa24n1+AsG510N8WygEaDYs7KAD6vJ2AoY0KZ7qzG
V0eH/bPKFRT6vtcZBGP9wXCuxWzVLIPZNTLCkBQ1dPDJ39E3Is0q+N6M+VhMTSfZ
vpul9F0GDnHpkM9VNBiIfVkuYmwiBj5Mq7L0Cg4xn+w1GdmS/AI7AysDlHeUbLCU
PZXk355BSQ26rGnuFDtZl2TRDjWO08Kg8RAKqJQpSIkozxTbt4YErsRZn00vZk3N
no9IUg9HjIU6e77wo8X4LlFBlPkD08+bHvjVQvRqNCMKaP3lAVO13tvphY4XCnro
3FEwlgCHu4ZiOyqh8zxRR583ptFl8WaTlqHBTNocgeCAE2/TpOppnxiLYtvR3Ihh
6jfuJEOHU4M2sPqELx7OVXjHptro0IjQuXSNZFJimFLf5ZNPna8tfEPq0iJHuAVJ
LU3siBQssaqVs97fSkRAvh717pihSnyUqNoBsZ/eTl+nBmjy2/XEq6doUibGtdEP
wO8jVvklj4YIBUfLIUPmG/5Upo0wAsOgbgJRvD7AaV4/oOsvZLLRk1S1HKvAxT4i
Whbrfkc31lY2Z2x8IUCaWse+l5q+dOll4v0gK14wQQz5EINKM6RuqTLIqs1LS+HF
hqmsWbh2MP3DfV9IB9MVy+UK73B6bwOx/If72WivICmzfJipYh40xHLMTueHA3r7
A/WYEmPD7cKBjpybVIczgC9+OHRUFc+YduwAmi1OUzLuGvaGPQGF3oR21mfA1vSU
FzTS/btkmGx9bE08XgQz1docppEjn5lgf87d4di22t4R3Ja2DGDEoN07FnkcrTgr
IHA2UTdI+6wBaP325WFf0++9HomXJrrdJbUcx46tSH7rSUAmLag/1S1R6YS7Rmy4
nOyyFoZTyLlLVHjnmBYX6Q3PrSt8mzExiAi2tTfHHVFJp9CfVITUa1DkbjnesCl1
Akx6rkrj6wxctieE2kiPpb3ZPySFnRz/bT9O+gOAr2ZfxfESPE9YdgrnheYJYggx
XG8NkR1GvooMsArngCjy/VAgWSZ6BNR6T2lrKfzpjKaI2rlQ989TUHhctHsZ6e61
w3yN31bjsKG4fjMmsVhqimka8H7fU9/p8Tnfg+uqFGKYCFdBp1iu7rCdmsXAJ3ZB
7nQF1dk75aNNCAOhjDqPzZ8EThXVYnCt9hPUvWsD9eZQrKipBGhRYdDLbVJlxv/H
3gq23hAlRZBdSn/uCV5aaOatDvlH5QmKWLidyZKFPD2xjAq0sSmKzWxItDOkm+jC
5Cq7V9H8QrI55wGyHK/WA0tFKuZQREk82wIaWfikfxPqqYZRHV5h1Y5oidwD29f0
JCYpNNIFkq1naAZ8Pkq2i0935LaPPP3AIpeeGC8a0iPfll0/I8CQ52PKxPoThEt7
2SMUGTqHhJfpDslGtIaRHibLkJ6uzulRnzCPPPV+mptiUUUTOeXxVbtPrYPoA40J
KDb/4VI1pMisLQLfBm7+u5SqRsm+RNA2Exzl72EP2QZiKdhyAMGZVKUS1hbz2vAN
husFK9qIpYNFfv3Jvc0vUd2qJ65Ykhw9Z7VxL36JYs03SKGZ/C+G5ICwt2EPQO5L
uR6JdQUeDTBYYSWAocjlxnuLIL9w/kCukdQX7hUkG4lrA60vl+T8CIXiiV3XkPoE
1T6g6qEXdkytkcVTriJNjScTI6Cbw5uX9FxXbYGiWzETkd+Op/HqEy680iVHBtCM
P45Y/b7QQrF/KG3cR2pzdEpQNp4aBI27X3irGV8gx7b6cx4SZYPMCk7o92heIfDF
vLdIM0gGIBMFUe4WWU9UcIa4aFJNV4LZMzvVmspj7vprw5SD+D9bBzjvIYKzyYZL
MztgqE1yBdICIb3hmwTr69J3Jogm8d+6tQmKDF+Vesat9Rd3YyCmyM3JWC6ue/8y
zjK8w0OCVrTEe0e9vwuQPkU6eYNQ2zapqJF44nXvHIgNeNAN1Jp9agVlTcgeNNl4
uUhts+Q1xIHvqGrZ/ywzfHw8CB2Vh2OH04exk/AkW5PCVAlmVLrvAFJ2Dxo2tnF1
4xNlCY3nro9J1ltjOzw9nCGiq/tL2/+ui2buZq6QZ7/ID5EgGbx020MukDvkBaWL
xCIcPAXsmes4fSjL7uoXEWSoadglBV3cRFG+ZT8kesOJ9qzVnlRFg1faeL6Q0PdC
6/9JowpCpRzNmx4JV4WZ/BxvS/y7Owp6OEQI1Llkxva7WrTIibO+1K2pEkdnke44
8wwR75uVYWS2L6RHGDMnXtI6/Utl01wDaXjK6rqVJAFMfHnCEpp7rS61B+oWnxlQ
jipcI0hIffQyr8tAqZ2+OaIRxzBl9xolhdaQ/d+Ui0y4gdoMC2lRmgK7vTvC9A+8
S4MVYFX/6Z6SdCd3aCy15um3JmhtAa0Hmf5RtNzVkY+7aR/cVlN5dDOFuN2DQaIL
9sAeWEE+9fjQMPoyRIn5xvXOA0NT5eR4qXMq218pvu7NTF4IbMhfbciHUCefD7Ps
vOArobAEaz3CloZ8bTUSVmSQVLHw92fWOT6AheMyIaTy8pMCpEoDta9k6nhIN8lW
o0cbfLHftQhP/mBHCtRLDncoVq3phokIbJ6ybcxwp3BBjRaiUXfczLLfboZUOCxO
EQ7ptO4cmae9Y+DkJtZbLeD4qN8y3jWTI4n/oDtbkR8N9p7s4EWpesbWminhGfN/
/o2ZFioko3rIhTepwJCFLr0MqhvJDdM1r2WAEL5CO211zVlCo9HvfvtRLlhzcEm4
yGO7jAqgQPF1KwJOinCn3e+gDB2yKzQv+AIM7mMfFE7eKtEsPpaCfSMDPTNEKBCB
DeM5XPlFFam/Bl1Scb2QZNyMpSNpyO+pxzMbFroLUB6ZVXldVCLXVftcVY3haxtu
qQBgeAClCgrq+zOJ3ehCQwOkq57NRmNur35pfviTiUoPZqV3tojEuU4T7eV9mGZm
iGJD90BjomTGrv3ZSHa9xXqh8bvTfzN0+WAfUuUP6Czxw/xQ9YXxZdukurBOFzu+
sycFwH826TyPgK2lsv/b9MvklUGMqz8DIviV98wbfJhsq10j5xNV9pCfe8ueAxrs
ETTDlwSIpsi3qpnkS9QxQjVQVtPGsG9dgEk2uqlwrwnXOI/vBRntI7KLvlzAG2WV
j04xy/9JsG0jtuvhwli0+jGDuc/npHemKk5h3FH4BlDmMG3ijrFWKQD3iZ9Gl0Y8
/NaHwUoz5yxTc+R7bHXb3A21XVRQXSVm+GHbinrIxdl9HkunwcaxGESNqLfh9bU0
4jG9VsfmrODUv3lA9qVJxwBjbjCpUrjnwa89/g0FqNimMdVWQi7hSX3DSBBSPXvk
pUjfEqeoj0KUflLGe81evVeDo1k4RWsK37/eUj/b+8ynpEpt/6f8WhFuwUcM8Clm
B8rcmkJhb5K2+46SBQPr2N50WuS9NzAQC7AP/zuzm+hxSXnvYzaaSHHTTiM+yv8b
Qm22QsWEgwtuP8di+K+wTyFJWGb9xBCnQWYQ1dklRjkWU6rlPhLqjUwkzXuoJVng
FXE9vMp/FFG3J+7aFwqOueBxqw2eHYqYFu0o0+fL5jvWkRQfJ5OGU5ijpLkx+buM
3kNdsZnbRJubQauyhzcauiYP4vj5OWMTSE/Tm85UHdXpwih4WcFmhDWvlFPqrrUf
CQv1arngNMLIXWbtxny0qBPwa6NJoyyTN1G01T1OhBph5RzvehQ8iIP4T6JgR7uL
yKw83PNI8Fo+oI320rjcKlRCTb/jGV4wdHLZEsE4RILVLf9hqQfzpFBfT7cf3eal
M8L6DVIuAIdkBjqwlWgNgicdh/x5cs2qdfpvL6WAND0HZIxHoEtfs92mAByc1LYP
CxwJ+6HwS1cLOpK+TmR6l4GhZu2sRnxMadqaggTLMO5rVxecDmzw0mamwO32d7Ja
kKR+cF3ed96kF6qCpQPmjrL2yBr3LClBzhQej7U1FpvfVT/X32WxiT7nxaMwWFw/
o3NtrwReIgAHwTyrIrx7FTePfnx0xJZoXv5UzOyq4oLpEqxaN/xZ0WsbYrMTB5Wx
st3OrnnFWaSTeZei86qjRd1trAu2u1/C+DA/hgvZLMkPGYutTXxIDPh9xg16jeuR
Ye2ifX4t1vTAnL2P045J16q10wroExHPlbW6hgw0qQQjd0bJDZeJsPNe3yhLKJg+
OltuD7yDeWEN3Idq4ADJMRCgqUVmXNkyf8ICt95PO2SIhJ4xYPWnXXfHbl2k/VcC
QAMqDlGY8Dqlozpln2pO6bKHU+YpM6Sbff4ZtrQHwD+Ns+shZHKpocaKWyxtyrAG
Zj4oIwD7A6GjOIVRlPfIPn+y3mMJC65LAW3ZUEXukZt6Eq/yP678Ye+JePlz0k7J
yP4hWS1RlTUGr1VmfnpD1UGKPd2QhXfHPaU7WKes7d8qYesy3MsP3pYxLsEjCONj
STrtKvhx7FxoH+Xex9VOe0Y5KV9eVJid80gzX1y6T+ahMSAgVga06WHxRCBwbYw3
TK+Ao4itmPRP1IGZMh2AB76J/F7G1xC8WJS1YGz9W5mJ46T1PBLSD2JJZazAAt3h
8b9LGut11Gaddpv/FIzjLaap9s1dj7FlbZC6Bj3j8mawl6UUqDE3FROukLPRrNHD
yleb8YvDYLZoaqcIIvqvLTltcM5RdEkp2eiXzFdFkf5zYaKA9cJp93mEraGmxvCW
n39k1yYSvpWaVhu+cU0ClYPq+qK70QWYWtcFMTYe2RQotN1LOjF8SbtVf6sTzIPg
6QsFj37elbti0M6ZR81R37+Epy+EXG/q2HRLZkq+1YB1XE+GUSYuIZTeWoL0sKiC
x4c3bAH24V2gSdPk9NDnQkdcOLIZokMO9sfwatKLYv11Mk7a+qqV16Gz7MnFTfjv
dleQtlynen1JQfzUCJAmpHWBntG049NklpDpY1iZbmh5o7tTGwHkW7PtZm8qKC8G
l8fNpnhKRuT+2Uq34/uuRW9t4qWTmjfYEwPrIDz1ktHXhEvMKBYJp/AIUI25NAFB
RQK7qn/ZuiLKUyKKTyMWsf3+aaGqli5hFmbO6TJB5FEpfJaEjiE2U+dVr99f+YwS
kf4fV6BpLuPoH8WrZztKu5gBRktxAHxSi29hC/ZsUP/i4J7UwX25/g1adjCp6wUb
Xz4qjFAbPH5H25bI4M3E6stB3w5TgMJwFyZbKeB16K++1Ngj9zWNJlKQDEXhhrA+
Vx8Qv21x41expD/QZ2EscgxGuMyg9iEjV9Q4inPS6mdT2o3I6x6FOhVjfic2pfDr
iFYHC+kSS/JlJVFYdubMJ4W7c+6NLTwtv6kd6WP84eWFvcebl+P+AVkzEi9//V8C
veKb1B4JhAlE3+b6isl2f8PTfvAW48PESFP2ZMnqOLvrYONGwJ8sJF7gVI8saVku
k8GdfyuSlekgqJjwIw594xPtjeJ4MqiaSj9e2S4ybZzeVSm3j3UUUozV/n0jVliX
jP5Rv3rYOcdYLCBUsGpXw7pBvmAxkMZ/62b5TjUuzuB99gq1eYY75UqxDdRuXuER
yoKQKAaQ1RaXX3yoiQGqmI0Gj8i4K4+fzYshnHq4LMv8DqlRnLPcNh72jPMsRf6i
cjV95ZGMJAmXcBbG0z5p3QaNOpbAjMa2rq5c1wrkm60Qw7PYCbV2KFGrCyPnaTbl
31GAIvSc61GshmD35sk6L//W/JsaLEFJwVUZRszLyvHM1GJTjSto7jgMC57CAF3l
vfnI+e2dHvioynS7eeXyObT3X2ZDXycSby+TXnq/NRcLqCHq5xE0P4RW0/16PHdW
4O7MJLbF0DvXeaZqLZV1Yuc59p6KD5lE86cfOQyHpSfhNItkuRwIdL/LV4tp21J/
QOqPzJuFzgLaRy+MSe4EP0F2BDITKuV8WISxMTYSkQfzsqp0OviOwkvyIZjBB9AX
iIxivI+e6N4y9q0Q/v/kyeGECizeSrkTPBQ6zEec7/TLzBcWiacuj0e7Cyzaudtr
tkZz1oYcJrpmsmnh9MI5D+ox8T92jPDVH3E62eiqeRaQxM2qgDc3RWFlTIGvOqvO
1K8S8J04CZK1DgFaykdT0K+0tlyQSXIvucTwcz79mPhUWJCR33cyXxmRKgy9D81a
9z+/OLSHvbUaPDhJISNMkTjuJxaZws6eE5XLVbRcz3LMyKcRdphPCNauD5nBfzEG
pZ9bEc8ML2VQmmSClI6+oOmJQ4COO1XyJBnAQZFHNnEGCL4kYu/vuIATDZLzGDeX
ylDq0w1kwuAEv+RMUd3q0i8c/GKsIhIjRVkRM73nwnvmQk6/l+r0N0iy/DTGHOET
6/jQmNfK3D+U4c8D/E1EJwNEy+/ZJGqjgTv0qckOTX2kuMdBigJzSyKYHSHLEn7A
oqeDxfnpEdrliUj6f9qmAF8dODXjiAXF1IlXVQ3LVD2PEyhibKXh1NdJ3S9s84SX
OpEJRSUYK6BA+K+GxpG0tbV4fb6kVjR1kBAzQV/ZyBY5NcSv9EstRP3BDEOAiOjC
a98ulm7vg4vGCJ84FOxaX0ndpP6vwHYWa/y9OLxNmeoRFs6nCD8BckFSgy5yDbkK
mgYeta1UfQVYl/THayVSUjfbXhK3XDmegQ5SlIQpppzRY1ScTNwNr0239LGfXM1c
XjiPrAFjcZSQbC8xiBpw8nG6Pil2MzU8s1tpxwcMm/zO///EwBbqA+206S3gTXG0
ErKFkZxqG56g50Jcamllsxp/r8ZvC9QsZIFiEjL7c++tBUKwIUMaslGLETWPeCFQ
D75x/N434DdsIZbpg15Ktl+jfHHVc8a14MzmQFOPFQ1sWKpBbOIT40XBlDFp/NzK
+a/FiZmAQO8M9T5nGyHYsKZuoDhdy+4JVxM3FTZehAlyzjm12/1uDgBBLqF5LjFV
dkDCwQr5sLCYlylDiBri3D2pJPwVtjimI3IgkW17WcA994TEfwfWYaBqZ5Ycbjoo
xpr7Ogd6rSRdffSbn9YpF7yofPyVofal7WaByK+1nBfAER4ss58flFsxg4YlSujN
fgl22MSUS5Eckguf71xTh9MsXM0DD0KpjoFCg8UTJwyp/OqhhMJS7r8RMxWl31qj
v2ZnMFVQDsbodMiqS53CPToj9g4MUG0z0ajQqNfATXuVk17D1veQ3fM3cSneOhEb
rEwemKA4UKp06weI4DRT2JNZOr9iDKE94PgUWN+84XXGx3SKt+WxpcvCtc4TTw+l
GyGvsVn3g00hY4utgMx35sd5+V0tZyjj6AdDVfcPVnxOMKwpT2BanWe0mko4Hpb4
pVCB18Z/NJ0WtQibbxclgRwS3VUKypG8PggM6GqtpfTniwcI7AdOzoY0JDmQkVuj
T8qtB/8ay4Rg1E23TuP9p71Nav1Dqd8twFUvrvo3wymLRFldyqKYWNyEzceUsXIb
SG2+76N/b5ZAkOvgtMXvb8VzZe4X8z1GjLOonQfNLgON0+gtmIWOz4y/8P9VXqhy
xRYHPSNEfW93RY9HI30Q9Z01odFZWW3vWw2xFKhNX3XPhAnmCA3qTFN+9AZWQZpx
ps0D/Dv2HVdxgys72Gnf2K3eGRoPRmoftrUcVFnT3L6MALly+O1HPYmx0eikpYwb
wuHTzHgvZ69U4DZcIhvo4nLCBTlEUvQs6CQgMr4QO7GitJcu6+7wXW//f9N4yzGw
5dx8eSW9Y5RX4vDKg+NlQHoVWeLLXShYBX7hgscISdS1Nr5jfCppzmYyLrV/dz1B
xpRXakjvfLzvp4g1mdjwKAVsLW4NWpScKesxmrfv+QmUrFNFVNOI4c2N0+B/Z2QQ
sr6pYxgYj1UG273/AeOXfC8b7BnQFueVMEwv+/PRD9mIDKvZUzi+X4uNH1P/9Fo8
WeOwzWWgpfFSnQmnSaVT+qag6/wzTL2zmKcpxSQHwQTqr8tYYXw3uwqgZbK6NK7V
UuavW3ATNH7vBpRcuCIy+rwc1qOROgBBFXYcefV09ubRLFuEFaaHBFnKnTjjIz4h
ITZApLqNHvFzMa4lEVi5uL+ot1p0pQwGwSCJJahI5QCQKsQGhsch4vq02Y1MWvnw
u4Me9OPsogw8Z73VOT2Q2C9IwldOD7fW8wh0gZwohleAoL9A+AkaN4t0Ez0A36qJ
mo245FuJc7U2AqGasFS0JYyU1FjMaVoyCyjSABcq/TA6a/Adtfdz2X5U8Nd88f/e
7rRoaJC2HRyIGdFCPQGx3yoGeAY0Jn5EJQU2HLVQmCgz1MMRi6eyF3v6xiOj3exR
YM0ZGd65oOQZxSBb3BQ+si/DpBaTw4BkK0BE3KWe/7xNYlRZg4GezlJBclyxrJe/
tv0ZOrYNqpWMJr2ji3xL6WPeigvQatY9Nkg5jj3XEorTNylfHt4IebJAUNkNmPAs
ceWW0JbUZBqJNA/ou9HZlZFw35ybzmHc8uXXTzomVdn8uqJUQgOv98GY75fAO6mX
BM+tXOGKKwJjzCAHBnAeQGGQrN/BG5eW+s7EB4R7/o5GWUWgOq8NXhqLSB4ZfjkY
FOqla7dSM1iw3wTYcbK5yWSr/uI02YfYnK2VU6rCkH5QwMnUZwL+S9PDwn7xpre7
Sg1vt062nkLdGx5g4FpjsPp51BrwCvOzUTDTGELvBFZQJSTGn67M485WWS4Jy8+d
nWjpsSxUUUqojzoKKv2qgGu7h9fln30S8bjbF0c47hON8nt9biGv3D8D4PI6P0wW
mIGn8LIJsmrRriY+53tkR9JQBxIpotesf7rAw44X8AA/dUaEX9lSQDFCraBLar8O
p0RIOaiVP3F+HKsW2U0/I6yanGQDwAq/P2vV/XKEgQ+7eqkk7qgKBAUFkBxZ5n3d
J3a58vSpvH7Po2DKqI6WaNOhkKyPV9zemE2NqjI+BJ3tD7RPc42uEojiZyRinXlq
DyIpjufBFi9JoxDqeoBROm2lVvc38ppO+uIQgnJGoeY54hClg9C/5RuosRE12NxI
mxqvwGm3L5JjBmFivI0ybaHiBYnaD0zpzuxnhHB7rXPaWB8KXE/wze6bpLxryMjD
PeC/EnHXpNV9hiekzCZmhgdmptIkXS6B+aaexB+rDhVEotbxWP2nt13DdlG9iJFQ
8btAjjRGVKx3xOKJDd0XuY9nnd+Z9XpCFM48F5IXj4JSE5M5c+iOfV1mOXjrA0Ic
ic42gd/AHEgXL7CB8otuBHqhhna1kBHYuXXUOkqtJpEhy7GXFTxWFXwXcl0zPns/
`pragma protect end_protected
