-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
Fi89jsPgrEWQiVr/0WbTZvcuVW5AHBzN3obZr4+EUiDEeYbowxXzzuy5uvbDZ21RuUlp2JOpF5XJ
ue7yRzMkQ1QqKfB+mGQd9rDmG1ZXRK9QtrGhKAvvHb9MnblxyXVMbIwlkJijBJomt0aIumG5Jytp
MUryLB81HIWzJuXS74/NS3yL/cjgA2UlAnVGPan5sL+CzQxt+apR9xJcY8yZxwGavL7+n67PhmGL
RIV0Ssm0qXK0AcxQa3Av/5svClu7mAYcLaZq5wA5mI58CUSuA7Tyu4bdZaFeRqg2SaOmq4nwxZpy
joi0KjvQmziNOmtn4HirhWO6cbvHwnP3FzrdCQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 8560)
`protect data_block
uEnG5IQ66uVKpiuim95D1SKOM04lQwhXrg/m6fuyinl2pZHj7Fj9yCfIiAxUTRTRbrqOxg5pT8UK
xcBcf/uQVoFtdOzypC7MG9nkEeYy0O1hRiXnp7nvEhVjXIGAO0kAgk0fWJ2sfQc3zInpxUziqWtg
2cSzspivQs9zBRIyfsINQEHEwuHWIN21UmOykApa0TS8SYLxwxMJ7EtZhkg/s7Hsvl3TlPdczo+f
ERH3lg10/6Q1laF8Cyozxk28mmyRk7GVlmVATtSVDsqnwG9q1tgtMbH5rDsLnagrHN5A3/HtCtqw
nKur2cuZd3yUIFJR323m4BW/gsG+ZQjoziHAbE9/y9Ulpktt7fqmDG4u1h2lBUDZIv8HeoxcAK69
g7NCLpz8nQonHPC7yX7U1yL/wCf+4Ues8gzZiKGwxEb2Vbkt0/HyXQ9mneGwqIG8m2KKr4xVaxA0
Br3RLK4XiwvpNQUH6d5y5swGBpTlyyALUA5ENy/LbrAmhXKlTZUG8SYnvJs/EMR2OmZhh6hF+er0
5Ev1SgQeY4HO52/V2HBLPPcHwLDoNKAmh612hvMCHCVnfbHvKoKZrx48mbSrgcVO5sQ3qnbSKkeZ
Z1LG77SPZ/hQdt8/I1JRLlInebAXG8aDW7PWPmENVa6vwzJ2cfZZSxW4YAz8X/BjY2JhmQEQ0ElD
7K5tExHwQy4HRSr8UgXNRB5uQuY1Ew9Uo25Hzu49wrubB422/S281ltR6C7WAWxOS7x8H1vQpmVz
T0EQjXg8Noo+sNmaQy8AkXMQvUdIptpCa60BydxwIWOid4ueDxsqj8iqH8iVqVzQuA4gBiK2R+1E
YLDG6uPeTzj8h0pF6OqdTwHuDz2im5bNfqXO1cJpmdnkum5AFbvtQcMXjE0SLuODIVodoF1cTqZv
8mpVQMixXkKb85Bqa593Y6xVf6r+F0VuGHD8SAmKvVbekk4QXtZZBMdzQOsvSKc6FNOsSz+StLba
XcOTnCdOTNoYy+D1DO++BF3unh1WZkzRzUX1eBpI7DkcNE1s+K8Qrs7RXomgvxo2wCbIGq6FAas9
Q2g8iaQVCrZ8QCFth3UlnNcxaolJmq4JSsYntzPXJ8QOfRlnSL8p34UWxGbWFL2mNQ2X4Ovnm+uv
YEMgFKkAh/YIGGmHh52DdKIMBnA8hGvJfbYKglngxUVo5qADTIJN4Tzn2mwNKkVarx2StwCHdfWZ
URdz+qZJAif2t09dSpzZ8vteC7LeZND/o0Wt5vc+yWanj+ylsgCASzCqyaaEJJv5XvHrjkNygt63
hP1UukbsAYlkdMplY4DWCso+BMiVmGHwOT0AIE/l7/DiQkGHH+zwJhAzPKZ1o7xw62Vx0OJzYnhX
EIly4HDIvKiAQ8lcfBS3l2L/GKtPDCy4hF/o+NFi622wTzhAjQ6bqHPUatEBXcSnAxTS79kDbqjt
xmKYCMXPOMx6GHpqOq+aoeXDx3Lz+6z6r/YRzv7qv56vKWeEOt71rz+yp+lIrThwT1Va5xMyDpMa
Bx0kuBkHrCkOCEd2AZMatkaihklB02A8ktsDr57plh4y/QuhkzMgv3u/ZFyGMImkSVkbs12oBNo4
3tPfiUr15hG6SAsoMVmXQhDiffyTrdiVUKFtZ0LtftDSwFtJ5d4LXObxR3/zxAuKkfFqZh/ScdNB
T3SeekfTYA45xRxptwbCD1ZgZvkLIEwn80bAGtz+7Ms000zkyNgMv8L6NgqAHhaQQU68v6kJUXYW
XcAG8xKPcEL2s2eNwZHJoHoZO6jNqvwWWThWIkcmtuhA6WMNnnPCUPZ/APwSlgbOPsrr+j157d2j
BSxzkq1rxUx/gzy5qfAe+tFtfG9TDrDBThBPLIrr7xcoN0aztkvKw3R2DDj74BtnudEa8sdxxvbm
F7Gyk0SJgPmE4zf5SdmwlqZFo1A82MWvVbwpt5Aev3QI0twvz2Ba9ECnZdW+DPv+KEQ+OwbSEuqQ
1ZC1LcOz1+1usk/V6PBxSrVhXiS0a1/MhAXguZN4dIRMs2im2BGD0jZkBFpe5pNJ+6Ha8Jfdon05
ya5n/xUVwyEp5FyKUdnGlipoe0VWgtc4uoeBmNusTaODhMdDV/26Zt4imEkgWJnz+d3R4HHiwEHq
TvG5bqHAH6D9yuuKdBaCB+V+uLWNGz/RQeLv/oyUnKxKlMFGRkt5fTqlpTGDXjcVAcrV1yVBXZ3j
pNKrPhWKIz2+nBGG14SEX8TibErE5Ud4mYEbxbCEfApiAsjVxFRYWSE11lbpkLLRkVJ2HILo/4Ry
UEd9E+H+lyPoL5B6q25faTXvAUHI9pr1z86+egZwg5o3xGItsye4EhhHqK+Dt5dsbSs9Jx9rLuBd
+JLd8PiXJotwXGlYT2IuuLsCE09zJH1+UdO37UbL/Pa1+UpZF15sym8uqdyRG/eWR92RYS4Hfp5K
fstnc3Ohdca8BFwtHCZ1WZ1OSHg417XqybTpPUj2HAy2vwMmC4yr4JwuZQSHXFRg/d7NAqj551t6
XOc9qGKdcCFtLwk3hfQyY/BBT51xBLNlLRzZ1hTRzNtu5h3GkoTDG+mHJ3dMFU98F39CpEKrNJC6
5ynESnZDTdhD0m2kB8toERtCwVz6bOGns3RysLnsGddd3sRl+HqX1bAPYJhSY8oEOcu9FfHHqdgR
1JMGjjy2RlhX6KLSPkPhxVPC1Pei/StGnCFKsXZXS4PzXU97g6ymvPEo4+8baWTXCmxoSKNbm9tS
oUtEbOQp7HNWgCj1xJfjMg5pyN1eV5Tc2Ov19BJuXq/tiA5X0CG+puIPpGco8jKCWftv6UXZdVD2
4OmRvHWKQKZZrVY5Dl9ygPVA9Zfl5JcqBbbl6vBJsmHdNdbQ7jsW5t4DBNZQuvJFBXgv+sffe+7l
oXxxU3FY3LkTAA3AJN+kEqaPJukayLFVQXAWLfxO0cnEzfDVdzOmSv6AJ2dDoZfSzAEqwIQdCS9D
StIa3RLfkfgK2pc+PBlkdrK25vEWYwFF79FyJSDcVo+z+GYJGuPHcSEb5CazV0T2KlFJiallxbtc
0uLYTsIzmA9s/EWePff+ms76y8yZNrEHxsJdPn39e3gL4Jq2CENu7VwWvUGhb0c6LuJzoyoxVRmp
DEsTAh9d1ScitJUrD6fILovIDbADcXXVHuaqeV90FPZr1q+rmiB+VZ7mrozj0XfjdeUnJFF2wlyP
WEsiNY6T4RTcJF46Ji6Re4v536flmAxMZ7FWUET9PbZrQP/5tljgua7EhfMyrNa1Rb5MahYKkSyQ
VUkvi1N1cgsiNTKBsPNS6E/XfbDORny9vkGkDGE+LsAr+5YMsouO4Rj0krGFATyGKsEYbCtQi4w1
sikbYHLsiTdtJ0I5vWA0YY9KNHrQmHihdd4nnp+51U9vHYEWR/r7lHvF1glonUlzkExT39/D4yyv
s7sT9UilioMMfp+xyVruao0v4hvFUWhdFGlFW/NEvZ1b0XO/o4iE1d//Up7qvvQYuQmTU6p+3/9P
jpw+PZODi2SGXkjPVMeSJaa+AY8GJ+Rhr/HsaGcXTWHUKLqu3TA+anSd6sg9ctXJrbGJ3o9w33Bv
ppw9EVGL0hUveZmona7hlCl/aZFm70IEX3o0Q8dFdtBOmPOwL//fBICoVIP2LDqAJykkhegczBHW
RX1EAeRkdmARIMlXcOOEbdMqDzPbsGLRGG16cVHB2vQ95IGUU7/Unx8yxIzmvamTTPV6mrRv9iIn
2P9wM4Amux0VceaA4KlOH1BAOsaGjIQIedKO9YvC1jX5sTfCRE9L3kik00/M4Jfi9dkV0MdRcY8M
fjbmguEkd81GVySlZXRTYcxOjedpB36B4MFd2YquItIXiXPbMx6pNLxEBjB4zI4R3Ls9E0DqlGpU
OXE5oDJvEfVSB4SGQ8HWxNdDIjxxBWwMo7itd08WPO29daOy9qw24+jAkq6aCE6z6c89mKQ3ulo+
IAabGsNgT6wcVbE3wrpd69ahXQow1OeyyoymlaSRWsdz1DMeq/ETPjUhm4c6oSlUwgtDE7PnitVF
VGNb2pvlT5ajDaSUOpy6XUjZdBdBH9V2T7TBsKTqXu8iUIwMViE2sKO06o7+wPIV5N3qACTtXtzT
rAJkpDXklpRr2UjIa5ztU/UOOx5WSqEmjEeGlfeQH7DOLMLe4bR7rWAwWBJOF2EiMUsdtVkbAKiJ
cwtsq0dH/G9dG5QnOVP+7K7P+SNKFdrocMxktC0d8+kPrsGFurBMsXwtyDNSl6rP+P+GmlEsv5TZ
taDRBXo7eQiPnQ6EJCXfcIefn+T3KUkKZxcU1wiHatGfrp6nVr7HEqhOXekKW6GbJr7eqS80w7ax
9PMRlYM2831Dbkt7Na2TaCD8npsd0+HeB2fO+jaQPUB8cNMeeqyXKoUoGDVee/qs3ikzHJ/VDW0Z
9rUuOtlqj+C+JQGmZM6TciBfucY73FNheLOvGHwKKg2Z9GMfZuS9u2B+O7GQefqXkCMNEFr/G4kG
9Rtt3Q6dArhHZkXK84pzgQ1GEjS6CIUFsj1PTO++2aA97nvwhw3MZOwkMbKUTrFQJdYsUiHGd492
29gZMug3TJth8S7WO4V2K8iE9Su+KDFhkAksGTPOQ4+KyjaDpcuXtJ5Xn2Or4wreWE3NJ/6DD4s8
/UN75ydWSnLG28UtTDq/3EramB+vVL4r6qIhd/Qd2qqSIFuHCkWibidcuyCz3PcPvARnwHGytvBR
jo71rif3s5rHKpMQb+Xdc7166SBC/W4lqtoSkghRX5n60rHI+Lgz/O3VZrP6qAhbPoHqDtFoXsJK
URFO0jhGCWP2VJqMIVcIVuQpuT5QfF7rlRbYCfKW+OZhtWYRtK+RyLTKCxawIJl6AU7y3KCt6Ds8
7lihyJD6rrz2MjO0nvI7VjtVnC+UY67cmrv5SBAtjV48xT9vjQUYoTQeCyEuYTmVXKtJexgyTor1
4drkmoX8BzVV3+iDB6eixEgOD8RAaMswYX/htjj5LB+RBRYYsf17B/Gsg0T/xJGvSU52dNYrC1Qz
DGJWeOla/od6sOsRdP3fjSOhtaZ63H1f3vuwiyziDlS7OCPWboTWMQlXs76hHlbBjhDLB4zsuyS1
o3MoPXHY9OOGho2boK3iD7lEY8wap0NbaelunGyGK3oyViXcW4GLP1RbuK3/z8VJmngCwHU9ntRC
isn6uSGQquGIxLgRaswSJz9w2xAAl/ye65Q6DShh7+1W3SvISV5UXsg3mJ1Qs5jX30UBR83dGy1k
muSO1cvz3cMlTkdtGMwG1fC/qPX9qPR9ebhwrvpuxDsFOtwJRVAC0f+V7gP2KgvLe6C2lsIuIpoR
WMA9zbv49ITJJw6GDA5pVbLKvKtcIE7skULlwc+VQI/lL/3V+Kv05zBHK3UvAtzYHTr41+dJt6Xq
vpYepz+89MoeZmQuSVVqE7RJ2zJ1b2lqgzwYZSP+gtmHMEp2jJFP55AckUysjI5g6HxvgbklENJX
u3d7f1K0TXF8vBII3OROBqsXBIU1k7lTOmrTi4NjJjbh2Qo/0vcAMw37m1SkmfKc9bfpWhZ7s4IM
TYx7FUtKFG+vW34pcIMxGVRVV9+fssKe4HpjiSEr17RU5JnzrXIixYMfGxDb1piUE9bRszBFybHo
yuGHwv43zTE0Wzm/m5QzWBLCLKg88YTrU3PvC4Yvu0EMA+e4Mdq9dP+xKSscVP25HGrM9Ml8JKxn
lhL6gyUhJq8meEyXdh5Km60thyTIu2532wyE8akjkg+ssx66gjD8NcLaGKzN2I4dw+s/BoKcBxtt
Q59WhrrDM0WgN5+ZMYprAxZaQZkW0qsNXypOGXcciLCAXIbnLt9umtRaDq6VLrLIxmctOjBwo3pi
nMWsOJYQ3FhGcMHTIW8LLyTx37NDHrRi+XCr2cyLGL9ZScwkXq7mufzhr1gmpt6WIV6rC6wEQOIb
9HQB4+P+kjjZdLvNlDEW6vtc9MfeuQg/w8aypVjI5+GbSgKxqWIWl67OC5NNy+t/M8pPt4qAEa8D
HqkU6lz4FC8tC6zNJDtbikIKrE2RZOqIJOT7cinK7UI+u8fawmUaUvD07Abuj6UJJ73BFytxq4/t
nSQaYyI1hP04LbZ3oD/4/asYYvca39ZSwcZAwLdiWqChVYdHPCabnDAYtFbYgQur4HJG1ini+6yq
JagCfJZVj6GIhvQXuRPbyUnuIFP6MpfVpdC3G2QbQCzQZDd+UjNeu47eoEJyns7RxavOA1+clJBU
yoKBUxN3HsD1JvVnlbFvVZDmIy7K2fFHtwq3lTlYBRgujsO6Bsbf+cvtyeFX5ZGX1C4nizFlktSS
TIy/mut5NjV8DYVJLE8VBxQBagq2ibVNviviYiF0456RX8/oG4CUSgPmdno6Vrqqh3lQKydfdWnp
Uwtklr7O8Uj6MLmSlB0rkcQwf/l9qfzwFfPz3dHslF4svEL7UenaGdk8M12PeArpaZU6+ARdJXFB
y059BgmUF/WgShWWeHaWB6ZM0MHc+fHKPpYcoLRAPeSfv9NZKBSQWQ4PgTBpUxxK9P915zYonKu2
DbKGM4FLLd1hkrxHZwqzXEAitMVP5N+Nmn6dULQFhXx2L1kCVvkqgepku2g70/GXxC3LQCNNlOgy
uCdU2YYrVtLjL5mQ3ItNyebRNHPeU4Ip9wrsY8SUguGPLoNMUMNlDGazw6tdy6YLD2YkZrG7syl+
EF6ScwVIQ50HW2M8Ifz/IjJrY/7zYV63vFy5YXPQclQWWNIIm3wyGmRc0I8fvIfmHZm053rYXM1+
5rSIfVhA9snDuUy70J0CYqrSQ2YhvRr3YQWcZR8t9fiHgM7MBHOXa9U8TzkT4MRIwfrhxe7DCmYv
SdxKp9ch+a3XyrOh37PEKzdKE4XMILi0XxfheTryaBWkgFEbDps7Qo5kwpwT5rVk7WUOF+W/6uYe
TET2i7D2ZXRZZMzr3bo1Th0vZgIgpy/rHzbIJk+9tuzVJR6nxLfnGBWr4EGXyTF8x/sSvF4Hqx+b
V98ePj9zqEBtMsuvyTrS8fwIWjxCTUvBDnvWwlJyttBJFMkkh9mOkA/EsULcyN1p/0FP/ymBLz6j
Xh1zk4yCo2ZOq34G8Z+Ano7biWd8Y9GyCN9NESdu+7KZjAllaHGfVTJagalrjw+N7/R9BMRwNArJ
2VpyiTuZdHQ1R4XGh9PcgoI7EYZ/1CL8lQscCIKd88GzmyxVOAOgCP6erM1RS9pNLb/1AavfrKEW
gZrDjHeGgsfSYEpOD1+ahzT/M/Qy1u5pK/ZCarIJ+g3gVxXx8KLf3t8Su5+IweKZuDFkTpEfe2/r
9Nfij9spkWqWdv3jNgnK5r1Lnfujh4r5mNyXEAdekpsPbrv2OYjHsGGT5ZTQvccUpW4bjztDPYxO
HOSX9BUFPtflOX/3y+HzQoZqg4wB9oeR74CwMVzz5VJ40dCAFzx/HUHDO5g/NUjtSvU6qadYjE8L
xytdRN6CR+EIJRBJaZqMBlmj038EcbVRwj+Jkt6EF6G11FIUnKHCiRoG7/8zIYJSSnxvDJGavPRH
Vo+YcGgc+cwfZM5MKvyKryrlX2z9G21dzeqa+VnmUjndjfby3sPVmgALv89T2HxGqsbQArXNPXK/
BtHpd6kw9YOCVFlLhGW2FHrEhtXK7BldbSqUrtAWg+VLza3IHZt9Omee2XohgKW81hjNFmeC4c7k
W5vcyIC74URU9szsUhbkj6wqSsFUYKfHp/z4gBv2vaOMOx71H2k9SFQlxVIKteDdMRhfgIXtYnbx
aCNxpjWBzXwQ5N0dEdOcPg/gAXiEPsaWbAT2bPTfEw+CtlB5BD3A4cuAHbqEysK/RK8+5XN1vPZU
774lQa4yb1Crq64PVGyw++q136lvRPJPp2rmyGxxv3xDwZv6mIkgUhMv7Qu6m4kzc17+C6XtI6FD
cwpJbue+QLb/P6zTDtjPr7jFub3B/4YDR5k+IxKNA7Wieb88oLIoq+E3CxrGwo8i1JGCuq/pJKp/
Hqw0dpoE4wAHwQpJtTMicpKLwf38VfsInPDyKZROa9H+qERlrvCVqkUeziWIapNXF1InikOc1hO4
1S/gQTuKKRGYBeszraLnLq+brtlUVy1VobO3jtx2Dix7AFwrigWYjcBklTKe57A2yTu2bv6MdB+D
xDxggHbTXGYJ+AMixchO4XIKMceXzDexycueE0Xc4wDpF+nTIXeMWAGVEfXWZQZSq2028yk5EAsM
ibd2tM3gCPZ6I7llDqXbsMh6DAj/eRG5oMUuB8m//NueQ5a6ywrRCdPz40dou9kgCqfrPtTLi9VY
qVWgfKpEBVZO7N+2L8NZ1J3YirQYPOD9HIiL/d/XQOwM1hRcYzh0Jg7VUhSd0DRSKmMg2/8nqHQz
Jp9fN2mOjN45WShQE3hKg9Qcjsn3mz1Je4UK1M2bwVVeQ8dJOUOhROaHyhlbThaddvJatSYZ60xP
76oNZOGUNJfBOsTTBmEY889yMF6grdOmQz7SuutTM7Eq3yPmybYwC0DWbk3SxGg4XjbVG8ZTc+GG
9xR/c/s0KxAAfgoClMkMfE1ktZCoYyDeoMGA7+5PajsQClTnnSCZPOm6sBNMG4cN6gLippkeYfzd
yN6dt45YlIkAIj3efbNlwV9VrUL6zBzkdptoAoY0y/Qv1zkjXJpu2nOmeiIUDbVy1nBZGd/00vnf
K55nJ6xWm6qTx3jC+oTJjb1y+P67V2X+4NlodIrvKSjw+tmRvPqle7XvQkDCdgTHYhYbiQa3ih8X
DY7fgKIJ/hlvEc4blNBJ3ch07OeGIPY4wOTBx4vcLNHbfQrbdmZXSvJo0Nwei8II2cvYycM/KRAl
N5COIcYJpxNN1GqecH8SyXAj6JsNYBQmXhJW2URD0Ymmy/Fe2M7IU3nj5qz2nUF6f2hb0nNwbWUb
wrDosP3GDjUQVHabhN1Ff017Iwwz9KiGygnT6LzCUTyK+4PeDONrGTHPRnSHC7RsCgEN3tlf9VLb
2F+q72NDE/f3bLe8NcIZDkebbHj0PowSuTRuIrbRZ5PvAef7u+In8V/xd72yEJKTLwMCmupZL/Ug
DQND3HPmOw+i4GklYpW/zQuWs/uLe3vOukdhA1HVpblCCDLx+3ps0VxyADZxFEQGozZE/arzcf/I
ETAylH6MDQQ65b/vvZ1k1eR0A1oYplk3z5ucmn1zbyDsUcsTQ510kreGMH5fzpSNnruYVMR+XpcQ
adi+8lvWvI72OpowTthsJnuervP4jUnjg4wsdgPxIEG/0nR5FENCkLIAR+uUg0vVqOgN4NJ+lrlm
DJRxaxumUb8w36I1LJ5KtojdOVFCEGGAbDK7TJIIUOgwYTE4ZplEjXmr1a+zbxp3anZVEJ4SGslX
Hc2pxn9fwFjEklW7lwJrK2s8JBeKzWC2g9AKSnAADJnIK8QiYLX+NVcuy0yrhXJoUeP7PQOKVr3x
t05F85zNWlhHUBMJmI6z012sptSGClH5ih0Bv9ZT0hiT6gNZKL9Dm/XoLBdEh+zghLHb1ivB+IKs
kwLDvp8DdL4y3OESg07XTT/QBYIn/K1kCb0VzJKR2LbL+6RoF1F8Mxky5GxyxY/cDPflUGuFxLb0
x3VAEY8FFhyElGHRSj1Tob1Uek7m9aVK0GG4HkBm7MBImjAfT/00hPHdoS8nOg6LCmsw91lyQWwN
XEchtci+E2OoZ8ke5Z28MNBVOU0e7dRBFSI4OOHVAbceMR8xGPrQnt1FIF6oDjmESqOxgUT8z4sl
5+p+OX+32dWras4xzzrshayU80SXZ3iwSuEL1SoQJ52idbcv5gIj36JbVsGxwb7GC3Qy4gYSLFqf
s1/00hj30mcmT6Z7OSONi/P0B9nez8q3CjVUkMN4umAX/aJ8Oq89LtUAt83y9kuXuXU58KqURirp
x4VXtn2vSlV8hMriCdSQM+jw6X6RbF7gTHL+VhOVle+zuulaPpslzL1nXEvSOFBy8BOdVP58e/q9
ywptSCx00+xAsPxDoKXr321GmJs4tR5rdcE8fjoiQNwIlcMIhNC4+aenCdfMzAqogb+KMqBM8tV1
/hCxjDGmnvhTrDurp/mBKtWEmzX5XHd/Ock6Xq4wBZhAEvx+P6n8qzJbPdPxtz00GvYNK0+14mW4
r9MOG9AkAniN8RX5mcB3C7otSTNkxQfkRyhRh7ZrviSo+shIlZyAHsdT6iyVjt0T73/yEB1RxPxX
QRGS7qBlFI68q9ATiMY+DLqJflTxEkbDLwU7t3wSXGchjGgkIDRfm+OWVAnj9wKI2+3ABhhIOLYC
6J+TCld4Hdm/n9I9cY8KttLppGogH59ElQ6xEt90TC8cZzZldBRhQj9slbpGnIETHae7dJOBsEmh
7u4M1c60xIUGAM5htc/tXsSso4QJ5kpSGRCvjk7+ZP1EE+bM8X4GPkjnLkobMHmhJjaKZpJims+H
U6hFipzR3SKvm6Xtb7Dy84Bxjp5E7XQTF8PbtB7XODY2KTJzVDQbVYmGOq3rFStCEO+Rf/2WaV05
37U/hFlfMA/wLGCUlhgTkhN436q4hgodh944WsticUUcabGgKrAtqUV7NXgCwgHoT33mK8w5S5Sp
IRPZp1+MYJkWK/DT0+mghbixW0c0uQeO7tLiQwh3HAO+9py+UEwN/sfRGx6Xkm2U7EAJfgbKj7tI
QgIFsXuG0O609J20LsjXrz/Z0JY87tGfw+3OEJ44IS5A/iKPAmYA7kjRvUdlc5ckX2JOwssTOiUr
KohAD6T4+z7EGy+GWQZ2gw9JmFXR7PJxAx2qO6CJit+Idw4xBKzahIBhOofvlqP3Yr+vzBZntG0p
v2xP7qPhUqM3GPPqXHHzwI0w0JLqmLlJ7lJn+UxUGQv/vnvON4GnDZVTgfoELEs1bwRGquPuG98j
rpXn3CzdZonKhFNTdVybEQsbGf/kZNCadnWWd93qb5J5cqxuPHEC1a/E/dub+z9mTWGH8Z3ooNCc
stzO8VcqkB4s1YbaZaM4HkzgHd80XtfDlZMd+x0wont84TxchUW+/mNQgewqI9xDhwYrkbndZ3V7
6PzMpAvFwFpn84aSHAScQUYg6ig9qNg63sfSQ2lbbozbvQ8zu8Zj+mgGF6oQQWVhqb6RK1R7ntnl
MCX2iZKcP1rSVuIfseZcHBoxuxLzWIitTLIEHo7gs7KCkDhmc9app3SSwFwVJM+M6xU/rzwQngJI
A6ZysykAyBldBLHBk8YRvSmfEC7rBC58tFbnvMW8kUQj340N6JNIhRBOEoERnIGtp/T5EAx+9OeT
XHCjofi1ZJ5hkQD/1WyH761nQagferzxcYL1MKXpTipQSCf+K6sQR65GOsCC4D1WvOGKirGJ+hmT
qamYfa9DYQPquFQe6OAl1agfU7LcA1nt1eSIP9Rrk+Kk30PkMQZQJKQ5lMqLXyJ5aCR6H+WdiGQE
BlH2+a6hdf/qXA==
`protect end_protected
