// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.0std
// ALTERA_TIMESTAMP:Wed Apr 26 13:33:39 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
G8HA9qZQ6YRAY1TkO4USudYM0LGSFJFqbupP7BUEnRFAiaAe9/TxtSKMiDZMss2X
n+g0G62QwIck+uXepm/Sac1q2o2gU9nnSsVZz5vqmFluMq2GFmL6aVKw5/DhQKEp
r4OQADO1tCYQBaUoLsKMoKVGyYOe0wtZXUaPXZ5YuK0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 28224)
Wf6O1NteaqDwbSUQorCYeW3Hn5XYIk3J7kfwTquqijyhpcJP+AsCYrjvo0j8DFny
Sui8F5H70KoZqUJ0YQ6805yQ9SxTnOKL1ux7CtNuIeLq0+f8pYOt1yTheFeJe8Zf
3uHbdj1cJ4sI8DPJSW+EP2xA5ztCkDjMlqoXsv58ktMEGH8kr82cu3A8rh4eeXlD
R39urJS7H+KorQ6Yn/qgirobiPKMvdXvYRU2KxhWbyNljw5e/WzGQYjyHLA4Yvbi
ZtaHoKG0laPEN/Dq0qDgXZinOAvvEPzuI0baFsTZtYLnvLCURDyRiVxmIOglP2mc
seXxXrtWYPeMY3PdA1bN/gPvTFxzh2si4Evd9BSCgdQLEOwIiWu0qtd2XhqTsmqt
gZkS3ut9SaUYmJn7Ilt3qIvqna7vYnbRqqNS+CqHaLcJV34IDeJe3RW9JS+sTD4K
qq6J8r6M1n4C9zov9LhGIMYvUqZeTzTY5Qc5iMfmcDAH8sJomVINq2KzTTBiFWmL
jdcm3/DEuZC83YLA68/ogE+FcsZguZR/UR4hr4g/yyov7O0oePz9tYzJ350kL0E1
d64aQLKpI2g/jewqKvr2fasPMhK1fLqS68m0Wb6XXNwaMIyMlAToajpoHqxjsFze
h2ET1FdYQwRvfxT4f0On9vh6haWRdMKKm96Yq60ru/1v3KlHtxR9E1Rwhhg6SAil
QCtiOb8hFmDJof3uL7HwcPKIBe5vPKFAv4qZzZdcZlgjkdPdxSdCOfMVo1KwSuM9
CGltzVvNelEan7r6N7+/+Ei3J9+wItGrAcWYndOrmPQmijEuRv3Guo9Jas8B6pMP
bYe9OpYr91fYpn/h37YAbV7qsXJpl0/dPwzuMRjZruY9xOfx1ffKbxa2xpluI7+V
wzdTkIS1YFYh16FPqzQgqGovupk0A7InQz7sa0xaCC3yE50CHoOpNuYotqhtxtaA
e/JEbJdMTO1co1lU22L6eD/AtXDcjujd8b4NAllA2eYskjIy3yOl2xtPjRHbP3d1
6h0f45+IjSqw4LDDLzupujYSJH0/PnL5rFAL0d8wU2omBqo9QGEtBO+y9UJG2X8T
o4K4ToydnUNWVzhRU3hhtYReTyjlei5JhkikyLFkxcaK8zvpujS9Ph5uPVkVk/jA
CWbQeZ2kbPWXQh0tGkAWLGmCJLSu9gSFGAT6+lK/QAMjMi78OZ1TSa4INPYmbemD
Jcq2TDo5H+F2y7vxTUoSltzKeFtwl7zpMYqRexBwWfDtS7iHg/JBCMn5ebHO7nWY
wMYQOsUZgE94687PkWoaDGejipBZVlI2ZL0tjhWYmm7DijH2EhaPjwPPoNOI8HMo
xrXcxdnbwSa63BxVyKeZ/TheFfK3NBdqNsXQan4H3IYLaoA8JI/jZfE0VMBowleg
JrDlQDx4sNJmzb1PTb6GWksNaZcw2LLDxffVbDSbuA40tMBWfSspmXbShXdpT4Ke
Ae/JLNJsyX0+3BrbEwASYFUAEfYlFrrD+BNF/ncwCPuAKSJqw/R+OTc09qqXn4bt
9EHg9WVLZWwHclZi4cRlBo7n0DAUcGqCBY8jV4c6ljUmG/3mBQdK3H+coc85W9aj
uTb6mq0N4cYspNa4NXkcsNFxEMhfjSgeaccbYa1Wb0EV6S9gC9Mn/0BuY72/KJB9
RroujrR4rGOtgpRu2/CIaWrM8B1WmlfhXgZnbZBaxi5TJ99xkfpisnkEmCMxOY8I
/LKjdtlGKfJCPqEeO1RLkjN8gmulYl6qIUTL68Jz4lYDaSLfEM1vBGM9UASZyudV
Jwm6Wtw3A3UHQ868TYyhIUW6aPrEMbF27Ja+3Py5hDMYMIF+H6fcdTeka2aSLpDl
6bBT7DCPVdF3rdT6p6t1A9AX8+jex/iWSQysK/7h8TxaebmqUkKoBm2ue9rnmtFI
6t6LIbBRf+kFgKDCw8jwoS3/dYhPh/X/VAIMZtUxhJIFuQ2wmcUjl2qJQWjstFU5
sbNInapp2UEYo5h+rrknkvXbjK7/Ro2LGlcfF4VX4dhu+DWKOyxcjby5BmazqQiJ
9BpKdt9IjZHoYMHPdCY22dEjWNRNw9ayK5UBUc/rA7xY8DX0SVuz+M83fy1zjhtY
QuM7DbocaL4vnFvXgrsxbYuCJPuBOMMkGodhlcmDnzGlcs73JNG/4UvWF9vLbMQR
30kAGK9IOnReUhFWQuYG+jBO41PLUPY/yK4Sq8EjpJhyQkXNvlliV9CYQuz1DbEU
sHhJlnart1m9UH6HqxbeX+MeplQS2xV7dhomCLNdS1vWbzlVL4Y+zzRlku9uP1hw
Kt7U+yRrFkO76nUu5gkZAn45jRawmJD5wDzv6vhndMBEHLCvKt7TUmpCvaj5ldlz
4HgCmT8RClN0v3xdo1QUkYqLveTcv4QMIXRffv3p7gu0UcHxi8F+G2RVYOXBr3Gu
+d+aJcQkmQJpMufFZE0/DMf868oqAxVhj65B2X642q7tkWvjULHkSewPrdazEUuh
1EblvS9TItH2diG2lOvk8v99hM8jVvvvy5k+a33SHxSq6T7fuDYNIE4aearnzLGw
kDBRNMwQYnifaY9JvZDxiR1ItVvBE+iS7OqDMfvPaDeiZQF7snB1n5+gsn5B4Ipx
JlVdUp0Z0v7L6t1NNSzgHxR+awF5Ff0XkFIlux+umDT9SIBaLjnedDr8KFRmpdMO
qwmGb+cVNzqr/haoLTheVYb+mx5CGm3Q9qHkIFRzHHYw8FQ+vUCYsdHKiKdo66E3
LckVj98z7xtGYnhJsV4xi8z6JMnMOl8zJxuyzUHABSzDDRTngiiyp6EtVYWQJKdb
Hplr/J+ZQEgbmoq7GSBC9eLdnoqHwsdk+DmuIlIRLQCRZtP+kD51ppSMhZTPrMJ1
Tskkd7oBZIw/f+q8NeQ9LYk5U47SrM2VMwG8P8T3fNzS6qxobkQhMMYLInE/CEIy
o5wLm8FMsZMmOZxq3dZFcorbetJsWTua2f2ZzefKaOeXhM9ggmRHWKypoSoRDqRB
7Yd8qfCIiWpFjvlbYV7knxiESdJdBBgSivi6nl6sllfJyo3axTjNDziai5QVtOpn
c8Po/N0VYDjQttsJYJAfXeM3sSlnoWFZ1SNDwdb68s/5mBW9JMt1SlX8cz1rnKUF
PoVEZIw1IxE52E22LF1A6fPr4+9qzgnbQHaNq5WqNhwra4XJZqS6eFQVDNrL7pJ9
IbYDPObE09dRJuOqpdHIldtUcmEeU2osETNP6f8jJ8oOGNrtAblZiwzFQ6BeVBLF
WPPnCw08bMfuGW8RcVwjyl6B6qH4n/sE9mpD0aXI2Ge7oiaO81JSGY1hq4kn2e/5
qZ7PooxEyHFYziREpAO3jTpRBBFtgPcU6rGNqKm4KJVVWX/EtHIwrWR9veIILXkz
JKflpB1A7mSOuPeon3La2F7/HPg4fytPeYeU0YyuT1UerH8oRjmyXb/UC4xrdQvn
jT7gwAwf9ONQiM8feS9MD5TX/X58hNjJkbP0WZaYCPLv7XSm6EVNQ+muja5nS0tq
N9uKpV8b2LuBcpXliZT3yc6zjejJIJ8D8362MFt8Ve2K4IAkqmulFG8xunfddFGd
iZSAcYqaRfVCts6p9EU6W9OmsRoq5U4UZcIsJgYciOAa7DKrVoKqKFwIwU6MIbzy
kgZEoI4XoDYO4UT5SJv7wW7a4QapJ4Z9VENjxJWaDlG66eXFKv7tum4SJeVJXT90
WWDY1vlFbHaxYN2oF+PmkD2XsfdFhcA6DUuV4kCv+vnaGFGzpwjAy8RBA5t8+GwA
qFMNM8DE5klKNvEEYju+Fy7VxG6QhOxAC0ki3VJWoVFvRAENMAUcQ57L2vc2SWVH
UwOXGC2SaacBFOllp9mfbgYS/UbdXltiitU7zWPU/OAnWnEmTaTaP0jr3g4Anr2g
IBJEKk8QMUrvEmF4sw6ofvGoRTRg/gs0zWwkKRGFCjOXisqseCvlBkgw3hwEYTn3
/CjcLvz53uS3Rag1Ix6of+zfy9FMhQonnVjiIB3tMbyhcxBuNpUbbh9bBAyLzBbu
1b8tc09xhB4fHXHKfo7pH3YsWJF6/b3vHSzOFcr0S/8rewzG9xnm3WBHnpx+pKFq
DxVWt2jiiXatPRZMOFIv1MFIfJ5CKZm7x+2s0X4kqKv5YSOGPg6kMAQPPSWsBXCw
VIQyL8tFD2Gskeq+6OVz0ybw3ywVVNK7DiOt0Y0n2sTg9oGqWWdOeTbbjSq27OcG
/Ku83ZNtTjx41dGYKiVAQ90Q6SX8MrXIkTiAnUskOzFEr6EjR3cLorTK3x+Yc+xE
8eja3gDiMZQHVfB1sogg0gJlvJQK+UqCZ/39K2vnMgek822FhhgJ16BulqSvs3D/
OiJARsR2FCdZvYMXHTweik0URLMEPpEbsQU7snhYcmLtbmvokd/CcZNy2+3oKmJx
PHIFnfGmBlQMx9bWiwOvrEOAk7jPgi81qt2t/kasUijgnws6Lr2uHPgwVQYTI3Fy
WgI048Q1clPwzQzsaWIyJoeetbkqKW3HIk4raEPgkk7leIEf2mYO75HwusT80rFq
Teg5Ck+dAfbN8ih46ThqpCfSXZHbSKPNxyNXHYIiyKP8b23PbJR2mfYIM8f3ylMF
bK6N95MUHtFWljaoTMV7KM8psIWoW0bQ7GiSULcbH0QXfOIbncuWnJq0Td9IzudK
WLIcmUwCyrp8OITyJmAsScpA7VenFdhO1Unk+7AW6Kn8Fe7BDjEgXewXtdY4Ixi8
4XtInAlNqVle/Ev9kn3UIS6+pFMBJYhVdBkYF6vuF7YIF1HS7zTma1ksK7W+Fphw
DHWhrARZBHst1YDjlU0LjWzhpMLtAr55DIDQV13d0lH3W7SRh/6VR8r76unhf9G6
hG+1GhXYL2z84RvGnaU+rkXRef9PYKf371GBwjooDi6brvTKmzpt7dX2EocwpZ0y
kj5Od48XpfaaAnm9qlN9cB8Acg9wQVzFKI9WCEP5vNPipMmnXV2doom56e/lBGxU
qjgSPlrxqYSvUDatLCVZuabyC85W+ymyat9VQVV94iOHkE9AnEt6557OsoGFN7yy
pVJPM6BLIw0HvDw+MTUsDojumQwilxK6MljJY8y+fVq0gw6MK5yxm1UBEijubAD7
6wUQRK5SOG3XU3ndDtpSvk9EXw7zI5yq577mou2hGAeqzwcwBj8/iRjC2WmmYLYF
amqQ8mlPhUv0vRlEYuShXb+dDIg4DzmKf4gLE2oZE89AUu6jSEHYfKDnZkxe4n6I
5mrmOegD7EMCX7B/2AFF9wGBTLsraT0RnS7WQ8I3XDh8QQ0b0nQJgm4Dcx7fQBIE
+0PctDuGNLpmESn/C2E6qSW05jeSqs9fwMbSwtJ8aXMlz8LqnfELH3Ohoy4ORFR+
zOo8ei4uywvKzNm8lxD/rwSygsk9x+FC3I+WwtyUnF/q1k/w3gV6og4npchAdm2L
EUJeehn9fTCItT6df3zlsf0c48gVBXtEp7iO4GmSlTx7xLQoizJ4jKB81h4nz+T0
vwv0ToVuoQzg8T/W6E0rcFDcDxtQ4Fph7doUdvR7BW4/vEA3YdNY2U6RsL+mF0dh
atYJV8IDh+HMg4dypWNr/QVnBGqWWuryLDmwyh8AxHXaRJ5PXk21TgWMxvZuQaFe
iNUe1VZ/M7ST0rlG38LM2gSMItGE9PNRVgGyhMOw/Xq48Gi/hOu57Y14ajvHvgDu
pVp0hGMBRSFiw12jlfIfiM1TyJYzHbaWUuefjgt1Du5ZW9nuuhxvH40MbAo7MYFE
YnI3YUn9uhjEX1pHe5YgxUaeAMdO0g+sqSRx1UWqhMXnU0mhGF8s0tfdAViuUBwl
TtXgSO7//kx4o/bkuy+V9K4y3BjfUs5D6OAunzhqjsZ7TSqHVBMP6id7Dqyl/Z/G
JMAptpJ6kud+qZj0fc67o+CVw+3wAuJKIbowp4ebiwMPG3Yyr1r7vC7RtngWae4V
REUl9WFJtCP21wBvkv4QClZXAeqxBSHY2ZEOJIyidQTk8YIqugXlT786suYiRRVF
nJfPcSMBdeevIa7sanhhE0+U3PxOFCsj8RDn5zponMgOyvWVa3Cy8n8lfeThBySK
mbLMDa7C0ByFP0NGtseYI6iAvE9w0un2itwisD+MmzXfN/U7vc2hPlXyIQ9+fbrB
JRxWFPziCc6QKjqIL8SojLrSsPnsBxTCAYmra9ep2OKFVTsLmZ18Mk0CUUmXrIUF
cCjowQO5iR7ePftrEXQ6DROWe8DidO8RZr0UqPUhQqDzoc5IgZiitzW17MUOX+aw
jhWMPhvJiQ1zevZwamm7/wa4nAfb0olfF262DAQgSZPyzrv3F2QAW14TifJE2AP8
6fvIGaI8qii46KwRSRQjp+jMDVwmWdGFcdmsYdyTqYkMoHQu4P1iwvP38hA+mIWA
Dk+rd2BUNT8VITpXD5umaCT3dlN+89DuzhjMMfF2Yr0YRzOxIo8HQno1TuvdfTSa
R+ltSOcv/R3BgCt8cgyZMR3KYNhzoLUqMecvJHsCnKYSM1KiYzKSqIORzEsqjd/4
tF77JKbbtZJ2RAaZLqGg2sZ6ck4DsHbEW/61YueVm95bh9O8pQJP2bzOqYcDhM9D
v2ck6GEa+pFN1R+NtoAtdNIKCJQJVpgVoB4GqFPI1msSWDknNiOrv9wdXUk8WQ6v
5eiyz2IZf7M7jAxGcQobOozqWgau/vrkQCyRtgyKSiqiAa08yMnt1TK9PJ348dFw
D0pvfZMKVHTa9UmQEdV7M+I0xE8oc7Lv+AGxgK4gdPrSk2g1oqWwkQfn1Jh3IRZx
dkpt/naJVNnw9Wa8zjMXvYL9KuCH0rYnftxUkVSp1/+GdwoCtEGJGEZjFlffzqzG
uAlLmRRWRXwCa8wU41rdo9DyeTEBvw6sd6PzMx3Zp8TWPHKcoEBdAjoUaxBb2w0t
WpSyOjHZD+eQdxFIxJ1ERFQG42UZQAWkXWljo6s/fJ368QXjlRRuxFFf0uY+CqWL
hIZ7bWouv2uO1JbT7/u215UnzOUruBKta0nGsA0ktqai3c/smNrSWQaG62U2DM1G
ISd3h535Senpw7CGGVGgIuKenM5gtawXBX4+ENj2DBZNS+L5SSNHHhv82ab9w2vJ
9nLJTrtmu9aI5wPxyDx43iLviu+GwnHEL99NQAeIAsI3BU/YAPpeETLl+eGROYUp
ZqDIXLIvYU73dCwKtLMrrL8LHgRpLxhj4OKP7kBO8vCh+YW3QsdCqwzBKWAzcPSg
Ddn3xd0xdfIqnqMpx23wqw0LsajggN+L53DfHAqwnMwbNRLZr3vOFWh7NjRmCyUG
sM9t/bqYHjmwYNJc9l+Nm73b8dKtRcmAjuSd39zJMDtPOfgZzQ0TZBoAL9eGdf3o
YsBpctQZfxnqSqvkvI1BK8q1O+obxOA4H8G4CqAs6MQ7ubKAJ5Jd83RQIQ6urTDs
CbCTiHz4WDk9G6mDetEkT/UPJKwF41wQYyZbJos2uaKjflrfg4/2e1dJQf+No8FR
U/q+Fjrx+yDdXV1JgqfEHTUXveeQXHRNpQwAFYerUeN1C1oFWuPOWoZB399taHZT
g6okeNIH5qC29QdZhmrXycMYdL3xGvOoX6k3INhoJHHbCC7tG8XLtwUla2aD2Vab
OvMkApmrE2y9IdOIv0I2DZF1PYvZ9VbnPlLuWp+yiC9E3ClM9XYt60zXWDxmcjHe
Wo5iNlb39lhqPa0sIFhA5bvb6YFl0sB/ZoJwI7OkTCozb1pKoZ4cnBd32V80zpet
vhGBdFMtFWLW6f15duyQSFw3b5gscAdxDkvtoNrHKjEDUK+N4x0ip/aZYjgYvNyl
IDw8ymJbdejT0CvuF7s5MIRWjHnYeoOFxv58qUImk9L+XZoul/tc7e4rZkfQ+2YX
GzXNInnQjEFJ8hpWUOj5NY96yMqsOnRDrKwWny8JW6n8cOO3VVKOOxqNHMr6GDZU
xu7fAXypmyrOjV30UD/DsBE/qwc/dzjiRetabKZCA4GYgd2FC+sXZWE15iYC7QTe
mFCNwwipQ6durkTLXxElEJg7W/rx0KSs0+qkSCndfvHzwzvwVIUgFY8pcxzV3gNO
TdGGhPfpH5NQMRspJnrDa/YEkCO1EjJFBxs5BTO/fAaecedFoad3bO75h/8CwmHt
ERVcAIa74whiRD4fzH0HLXnLbh9ljCbYAnPyMNxcpjfugiJwrAm1LHk3LhmBWNXN
apDhPg/O4gznlofOwpLwtwSWdhdh5nVz/qVxcpmOIXgaWbZQJ0kDAdbfNLNBLFYX
sURsohzLVrpdyv4cLlbhWFslJz5HEFTbjnLQqmP690fmzkWoqTVw7KD6k/AWIRPT
X0OPTX0lar02ZRKUYrDls8R5BcoggkMQQkxfu5hEuoUJGGUKwq1+OgAisAKTe+hZ
PV+4koIZ9X2Z7nKaoBoP7kLUzOgagPkLf6n1Qu6B8R1/sScyN7/ocDkQR63DYjtc
oxnkzenq0UJ7a4Ffaf8XGTPpiZbEsivR1jSSB2flaa3se4QJw7oVX1FXIbL8AsRf
ZEX1g3me1APzals77AwgWS9jpH+5HxPXoIxXDNQLS+TyrzAcWZXuKxa811KtwXDS
DD/+xcL79HxONne5C6ppJ3lbFVkkYkGpRG8EJGPZZ7t98e2eGlROoFVrtlbKBE2I
WZF2qzbYh8URj6P+CoEGuUx6HXaY0qrlfD/9WY3MQ36EbW72L2WUTullDk2STSMM
v8xc96gkmikN4iWkSaAmBHOFsFm0hVkQ8X3NGCQFyZlPmgK7/wrg3f1DMQUnbFnv
ixI+DL/qCwDcKS+o1yNjraaVdYZSUmDzovDLqYrfr5sB8nQHkab2iBjSfrYsnCMy
bNh7O6LU6QQsdKh8Ezy2EjDSRo+3PnWaC5YXXV0BUPJgbSoPPhQJ8wO0steP22Vx
hZ+2dgff35gbjJMYGaG5ToaOy1t8k2eoP1dhl1621PWiivzrf4lt6FewAPFMgviV
ircCTMSyOv5zmrxg5fepV+j8rTgN1vuGgNbXPQ3QAWJ8t9Cr8iFk4hWdgVkCT/9l
I5cJhfGFeyGx5K9P43XeuK5pYaDUj1n3vfxHmrN6mKpaXmc5As8cZdy+7uM4y/v1
N33fzoMVTck2WrbNGzTetWma7Ln+DPFHf52GQogjfycrGPr3BzQLW5pPKA4DM90V
X4Ql9Yui1uEOQ1u8C5EDLeSRpNCXtFx5djL52wjSqC0Ebc2mfrPHNG76vuRhygUj
x75wQooL7X4re2C8OvgngIbiHdBXQz8TNrf8lT3EErPxubZ/WowZvugtwBesdqE0
vUAFAvN7yk0Sy6Ii2juMOsXkUoPNYI8R/bj00KZg8Mo8EfutkvYRlvyvOFuk8HWj
/eP3i4iX+dUoV2v/7LNRdnRchUtH3yUyoTgNgsrlog4sMUDHm4V055B9gPLs5Fcn
jCI+4RM4tq/lALBOT6KjwsYKSIVc3HSBY3h7ZZjybTDLhyswjgw8NjSGMZF6Ux6w
67R6WfBRaClPCEIDX9/0HMtabPv4908hyI7P3fzKQL8BqRSU1619Moj5vXWfFy2k
eDxDftqh55tytFbpfHiFUL6f48Fvwf3IsvzJpx5DLNI4Eda7ME8uFLYu1cpq88Vd
ZQDzRkptMY4zWWchLKB5OY8Qnv3x+KamC8ukLuIcDh6580eZ6uaRdy+bUO0y0dPh
icm4W6j8PvnDk8jmG+wob+6gZatzRqnQuwrHVjCSqejUiioNP8qw045YBxeFMHkB
gVOmVzUpUhhNigtKJepGGbcbClMs5p5CItaDBFTWS0awZqih2jvpHgDW+kJOsJ7F
oAKztwyHpsCU7IsukivqrOSVSU/9hc/31XZK6HG8lZPCAt0KbQrObO2O59uMd0Sd
J1Pm0Y9RtHNTbmsUR836hYVmGQsW7sDgigKnG1TDslQwAwrRxLkwywsLDGFYMDif
Bz+4tBDIObldnWEycD9vVx06foeD6kwhzep8UNP07Gnp7r7QRopbvdwwm/Yf55Ao
S0UPBGwIZW1qd7c9NvvJp/WTjlmozjv0o5qYOnw+ZZyJmqJV0sjFoHcUSrYvMSoE
zlwOmPT0Yu6s7kJDoFX9YZb5L+A26I0r6adIR2+zrPIPhtlT39gUPQUrPcmHIe2Z
rUkIMhu2BbNbTjFxoBK7tZ6cN1wwCPQ1Q79Wz27IYzJ2CA/1W4IS8x4ZRmNhDqdE
CRmF4j2CSoZDyNyxsqC7xc/RY+qDqCbbuenwd79HRQx+tQscJlnAS/tPRHaOqBNE
NAxL/pgk3TCa2QHcnl/aCJps0mDSdj+x5sHnHJMFNQn1nMjl6ObzFsgNGNNkEjr+
kgkaVfhtlWcSXkPhFhCThXeLOLKitb0fjSxfqKWKAOR6+jo+cu/p6G1PcINJkHZx
gu92a7IWxGthvBu/1HtraO9WoyHOFFr9MhF2IQw/CHmBv4T0uyfAOgs+Fj/GFP+o
7hvDq57BNP1hXf1Ge2FFZRMb4ptgvtHT1004SCdOanBy06PnLy/UqX7gy+RpZ50q
aIWDPRK8x1/M5d2SZ5hG+ssE0TBX3ufirf8ZcxuXccYvk/+qB0eOcLhiI+DNU6YF
q/jzps4gW/2nhCRdUz4zdeuQvtWSbK7hKIxN9RAo5ssqmBG2moXtKV0VBqeittc4
G0bOTKSSniRmEoTVE9XcSdGn8DYlMkvU7uuQs/ThMirLCKQiXPdAz9UGrNUbt+HV
jeopXJkqO7d1T77w3r2PjuxWdR3cuzwStMvY1ek0L4IIyNLD29uKZb0bzOmnEZDr
tK3JZkiGEzM9kUGt5v9be/nD/hirewZGTo+dg5Ef7+5gE8PWHpo5Rzg/Qoby828X
2C1hwnHe39pfkmznv6/Z/435BgTeB2jvUl/rhBa8NvhHClOidC4PUkXFZf2BQtVy
qdUQ77S4Edn1QK25bCKF2182ysAVKZsOaI1OQgAJ9hIXRV/yPmPYiZq3YyvSh9fu
gC/+j3V/N2Npj7IuQwSXPZPC+/fMibUWzcbVtM6f13XC62uO7Y+mDn017C3OeNu4
e0EBg/zzGy9ZJX/ixHHLUg4e+5Zcwgfl/PPn1d0empnqtRE1qs1XIdQd5UMB+y51
/Q0cgBoMsB7CFMN7kOWxtwH0kLmnpT+SaTqTjtY2ZHKmZjmRredOyvfAkudtqqob
qr3Do++2epHX2l3CzKStIQwZ9eK+xgIpgpcBlqkhAI6lhewbCUbbTIoIvEBGno4g
lqIC5OMizdqks0o/4WX6vkUvTRPsKOnZJgKiFp0mzSNbuWIAjYX2CP5JVugHppYi
uzS/qY9/qYKIg4B2HhuXwMifS41KGyM1sbCTmyD/MCx9nWPLdmeFo1tLO4sN1Ea7
Q19omQS8Ex7dY++JmMMaznqyKJiPPLPVUXtIVc7HORDmRgdQGIPdyrWC15oL5wS0
x0Ec8gMQcQNk7UcheUnRtocOSj1F7tajztCOzFklxboluMONX81QCZXM5wj61UNd
/rtKjn9WQuNcxoAnKLBgADKSmjUTqy4gxfAWza3uz/DHAeV6ACnuqWjPuMEn4Upv
UXCWPPu2TEo6DSk/YeI0ml41muHvZGCh+S7XIjnhDSgU+WXmiherRRchFT36nYHm
UTbtN6E2nPjuGTcoYgdcy0p7p3sL1a41y6TtIdBtMvH/FzuN7VmusigeawHScKSm
m0yr9a46slc/XlAEj1wfyFrFNoEwpviDBQjO3IDpyVqSUo0U7seXdhcPA90T+OlX
4jtYjVl/fdDogXZqT4QIjjBITJRtH2RE2v7omdtjyER24ayP8cVxAnpWdlpe4nZQ
HPj8eUloKOQmSoJNmsjGYR/S4gwGwCnCzg+9h+TLRhkJI9tqjqIfbEbyhapjmFcX
cBo1oL29h5OjHPtg4uU4Ny7lRSAR41nhTLJWczb1KPJITpGsGurbVanZqEb5THkv
bgM7VMA+GQChCq3rloCR2PCcT1WKtUDnqXSuBE4FEOyFVzc78DPT5xo4LsT66IXl
rnr94YhjUTNdgOAHjURgjTManEh0EP+0ZV2/SzhnSAinYBSLRoDSGLvpL1imyEH1
w12DaNFH/Vy2aoCAkC+hHDyMbpTg8p2lKqxC8oOKe9fpQeSfPmjpHPuw7VbJ8uE8
z0fFvW1l5vLQbCTA+iCPOaMVL4s0+QVHD07sSm36Y9wFrXRXspqAfwIJ73X3dqQS
r05HlzF609FHh21DS1xCVDjnSg9PET3VPvZAGyw7SrwBdq7rp8BlJd5WqaFBvrSL
/OgHVV8nrMseVw1D3MaJjY7MpA3IgWvuSz0wWZdDFLkn3GVHpy2+d3bzxXDthsqk
52W0J2wfY6K+LRMfx3XwY/WbF5uG2wiTQzLJEUgng34gKvAkNnaOWzBV5THm70gb
rLDfj+Wjp0/uVVpIXxIGVyl1VWE7mExoXJ6B4/i5CDIhNM01ZuAtLv5+utQxhPIJ
a9u2UvqOwGi1hueXCb71YKtzaKWYX818prnixcdZulTjGCk1bpWHQ+JbMSmAlQSp
zkS0bAnCLbtZTzTPC2cPPLDiW93th5Ylj3dbv61X2M/KBdjws9FECiNlLxWb3FU5
CJw6/9osox5e8dxOlPst+ytRWgHg4URkMNWUnXWSWopSns2o471O0923qPdr+Qkk
P3gSOUm2591ZdvQk0XQUGVclEyPp7tXWox0vZXlTUSJhtqmdq4cWMKnBOlIX65SK
4BvQC4yPs4zEgWVpSiqaZa/XTYhtLXkNnwhoQa/7YAaOb87iVxgHNXRFOnD3OX6K
wkdYOqUpIbLNXSVjlOZqqCEAzamRRz9DOKlCwKwXRakY5WbZZDeAUCeZCnAEClJX
urJzy+wXi6za91wcqnVqmhluHHuo7uAU0nyUZrQ4tVPiK5pG/LHVwo5Ev3f23Wm/
TzH6Kqgj77OTIzHpTtilbOQTkpASLf8IHMVuweFkxC48F9n+G6QBWYQSsQ2B202m
HWn3O3PypyHRFiQ/O/f7ipRhWDAg7BGz03ELSjuLhv5WjUZqLLBNgurhLS4St5cW
JlYlmxcQpLVnYzULYOD/tjORia4CI/w1aArOUGD1bRGBCQTg6JepVxkzJRdPP7R/
wJvbJEc9N+VxRbWs4WZSjzwghhZYDqYa/88xTBZXB5MgBCGEZ3FQtUj2gtIF81N9
HgZcN3oLWND1r5h41WLpp1VzZLkB1h1uuZFksrnGVE2tSUD9hV+br6G2eR2MjYz+
iLV26j7JY+D2NRrlyIORZ2TymmWCa+LKbs9oJcCGbBs6s/vsq1/x5iOZ75TKFuhf
lxSVqVrA71w5YvvVzSCs60NemgW3XSdgdSfSRCAJB0wdJIbO2biOD1taOcCnbX7Y
KyaOyj32mO/b6FyhUexwNbVtXJmn3sWe27h6Vdf/T+ZDfIlO4/17x+rDrU0p67Xw
0yD++9rCLJ2lsCrBuAScgwK516PsiNKsWX10mIGfD533o730YYoHDn9JHjtYtrUi
kBuutmSvj3XiXxyzfG6nrWezg3UuNjBa9XefUBxSX0ff84nftQMjvQiWs8q/ImyP
i0rIhsaiCN2jXv3FP3+rOw5DDlug8cTvA6jx7d1ZdEQUG2Yq6FCIH4gqaS5ZeidN
eZduKG49ELJYrc+HwLdMSdGY5TPovpYWAm6Vx9A9lRQac5DXDDSRSHHgsCt95Sxb
fyl5uYKLbbhAgzAyiQfdFK3BeVRjwRmj4Ghdl13P9MSLkCbdbVSfnylog3bqRYSm
wq4qUtZ9hG5PeUfbHY/mnxrsbzofeYBM6wLOD35yrsnDToFjoSvn17j2F1IFo7v8
AyYSQGNQlal7bVxNajBtifuEOOjoQpFBn/35Wejb+S0wGq2OeIGpZ2TXha+fFo9N
elve9dFrhW4O3cwyC3IZ+MHkq1Br3NxC2IV8h+6+bhOqYu19mlDFYsKc5A7zQDFw
0ewzrN7EDmhevqKsIeUwaBGF/i3wY8zTHt05GYn6/sRS4s19/pgxIM5BJONQ/Xyo
a28fWuN/FDHJfvAEra+4oKEIyWEepv0ezxxGphb33d27aS3rUwxI3mTeya48ioJk
nLl7MdPc14D84O7I+Rp1dICdVyNpuLCrcWhRF8s/KeNDquODZmr4br6s2yTPo7rH
BUHKuXPg5AJczmNWmIfTETMaq4kjcbckIVQvjTAM2cLCskPCRz8LOMHE90tE32kz
oF7lwTCGP6DuOQCsVzSQW9OeeQ/kNIsPbZMRtt80QVseG0z9wVr9nNmD0uDb5zrD
MgPdq1Q+N2EX4o0Jxkhu84NsYsP1OLW+dkqmF3tO6QASep3/GxamAKwqWV78EPVN
YXY3XhJJsA7paAFCaxoQrvPpsnr82DZdQxYs0n7Klz5CV3bJssocQZghA6LNarjP
3F9UMeu8iCXFHtC8YWblEPpP27iJYc8iRlJ8stzzW5P/kMz8mmquG/TeXDJaSfZA
6fxgFeJNDFKxPS97fEd1B/Gj8fAtnnslUDRvrvh1ImumzVH4POy7+L7rg1vu0zAf
/mS74PM86u7itFYOP/6NY6s6p7IDnyiMbr22BxcnJeMPXVEKNQNAWycED9Tsd2/h
7gbwuhpdFP49smV9KoHB1B20Cs6kVIcbxv0RAO1Uc64gzooOGdo+5hav2m+h6W5s
cMnjy1rbfh5t9fyfiF6jWQ7uM6sOdNjRcamFwYVI9LE3MkpmZIlvZ3/z6jB/h/Lj
Dfe9lgLbxr/lmcozQGvF4H6h3dzAKayXUiYwOzSRLhXiU3c6WYIeHmtGubnRJ1io
n0odhoI2mLKOZH1+vnAR4yj60QbpLdgzzv/CczmzRt/7TtcwB5W2AEtyVM1iHWJo
l0wdzybvTf35OEYmyAiLk7JrLQG6d/pRD3yfFUplyoLxqcl6EoOkKZP5I++e6Mdi
a/Zqdlj6OoZoJCRbDGK1xSCxo3CBvBYyKsN+KsOiLt44n6hvAhMRyCV98VzwKOmv
9Lu/UvkdeLFBuPZ55rAocH8BvLtj2oFqjPLAfO85jD6VBQEyK5rjYCFQ4WmqVEze
+I1puQX5Au9fM3EKK1I8I4MN/we5txP8jLisWAf6y4C9HSghoevduzZuhCai1vCK
xd6cd+/Rr2V0aEtYmbjdOckjbnJn/BMaB5Ol3XD/TQBZrxD9ulfmUARK8YcsZVmG
qxtIb2GqG9SgW7PMwjrfUjRe8DWCO0WmmsDkXYCfgqOuEH/OfrORfSJkGk1LY5L7
T61ALt9I7UldK9t7511SmNxTXY27DEntkDAIl5YAEPjcw4+OW8s45BHxsGSNh/yT
/CT2BMFemOeYyGQ5+P7Dxfghu70AQGwE68q0NoEJFlTTQsQ1vK8ih38aGVfP21QE
kiEBfeJOLKiEn67ii9CDZMB1UnyRYQWHSCuK80yutMgB/vIlO9yIk+fTtL1tRpyx
mD/BjuFFRwMUKQAOoed5ZyOMeeNWHZ581zQWGY9SuBRij7OL/XGTTAii6Dqjkg+g
sHZw2ozQZ+xaUpUEJCCaaL/LPoi0vSqS6WYhnbVWlvlfjA13uOkyaRBRYa82y21A
JjuFtJ5dpDPmEJHJ2w3+asy3Li0vBkUqDGHPpmFWWsGvjr1lisQOlnJhtJ/gsYXP
CJ8lqFSWtnr/MdHw4WQ0wmxtM7x2UJViV9mIMjQWS1Dk6f8qJlvGYFUMjNhaIwGY
P2GDDVMhUYLlAr/JOj6C2m6bltq0xpVTVEb35iieddOx+1u+HEL/wkIm5MsynAib
SyrweT32rb/9VPQ4MgjQFcuXo0Ji7i5zyYkSkxVNZ7DJZ+kC7jeKWdNhj0dxzZG0
69B8UYZGbG7WLt5aBa55XBa+Xo/6rLG88WDYTmW70qPirObEVbvF2N6xvR06JH6g
LS0g66JQl7hiIfPXXaZP4nhOI0Ck3DfD6rJY9CEfCCP6KP2TkdHYN52uOygEZGUn
v9EOPdbGFBq47UDuQNpFMAEojBNmxnmkEWPws2HcYDYmaFNiLHgZR+PAIFMmlpzD
H3iJxaBlFFRVRYloGtRzCg3PFAUFLYieV1b0CM7JE+pydvteSPpKPqpsV81ZT2op
jQ7Mb6YsbGCb1wTDH1iq3ACYjCcHu/QVzqmmQuZWEObDqrNb1oDAOUGs8Zu+m+Lz
cXX3ekC7U0IamQ/wwUb8jXMzg1AlgyxTRB52gTKz2/mz16H3QCUOmZ67G79Q9K1n
dbnTMpAPIVKkfeFgKRmLn3b1dJJx0vVnyx+xMfVtIEBzHJIz/sSrqDYZskVxx/sH
zpa8Szuyz5+cLzODI6k7ddOanA6b/9ZwZr189XTBr1EPiTi2lBN897HFL/ftHAlE
CtFjYYqJ2W/eeLg/yIAZG0qI8XtDu9cJgGGTk9z279rYFB+Aq2DTwjeIK3lMdUTv
+tW2rj0l8FQAoabrYkmavkhF6Mch+E7bxY1XOYForavx+iLwH8yZItQ4KVW2F4x1
fIo+ogv6hnj6lLnxko79SfP+c8eIqVy57Y4E+0JCExXComCp5XXZ0QA5bjSfb9Cw
S2vJcyrTo+AIk1Zvnq+KpYVORhYANIovQfLB7c8boFvYTWzH2EAcFTww45puP7yt
rCy+kW/0maoBI24lpj+sydfEB73bbdnBN9tkt+fUmpRLuf2DauR15Yan3F3Wd9/f
QwEJR3xIeu4IJptcNaHrSCV5y94bI/CRf01GHRB2++Y1lMFLccCsBnHqLnaohWLA
gLifd037mlCpLD3U4SgbN6rl62TmkwRUliYmSCNvo+vGtJv5MV+Ys/R7u7XRdNBj
CgKT9VIOqBMROOsLhhEkCC8sPxibGNlIXQKFT8DZybQYaeeGBLAqwGIi26H1g2r+
b0Uj8TwI3Q6/4HjW4zxGkIckgmRaRSrSZi47i9EDePWfzf5FBsJDsLyj9qmfEgqH
AyZl7xiMtO/ZpDKU1fHOsHE7efGFgxQ08qhURV+KQkwjsa7xXi7D0JTPnM5ZDW0Q
EcwgVQfz40cHlH3k6RNgLU3hM6XQ37bvTPSS15tesLBE5KUiawOOmZQvc89PnGDc
IQtj+nxeh+5CtNPF/enoRt0ZgcZld4ppnuwPElcgbLsYmPcQZxgwlQl08FNrbW1Y
D4YW0XhOBoGrmvx9ePNQTtiMDrM43V/g2kG9ORZqT0ISCNXvCYzZEc/PlVew7SHb
Ve9PbJziwbemszcb/HadHft6fP0ST2UPj8vzRNBDUEa0xD+/ORzAdb9r+IJqdcEr
lkd4AFtnDaUVwgG/JWQxdtdViwV8YRwb5xcsZ7Rm/KiXhZ1H5JLXCstxOiAgTKeN
5QJ8rgp6aYa0eknzNB8Qt3kQJq9OVPKN7JcCdlre+GwZ2d0EZRGXEEhfKUROoAQR
0IGes4whLjFsM7x1VZCQ9FBH1dmQpFsx6W7R4e28RGerIEwf4/YLCpX464C5saEb
axhzHi0hPxhbokIwtuj872sw6msPNlMmIsgBV8xwjGGp8+09dkM1ARP+msvtfSTv
9E9FEVCS20TJr0c/8MjRFzhOeEb5ScyiRv2gU4RYKElx4EroPervSQerdjb1jFyg
fMfdKj1mLixHREYVOMa76Y29xjxsJ3P18vwxGebpnR/K6+1o+DMwWEMcISkAyenC
evYdiP3uNsgRjEU8myxg5vgsJxLyeH+Hebi2zfg5Gdo65sR+eQ9fGPfPREWGq9Pr
Swpjndv21KuMsom274dF6RmG8Og58ZGZ9mbxrvEEyA1eivvd9fwb8Kf+kxtPxt1S
Ag5sfeIFHs/32vrztdhEtXs6VPPtpK3lYe1XP4LtbXdff5yItskF8iuD/Xn5jjPM
MuDssvmyGVGuZFAgs1yfEq6rsY5ZusBlfJgZlCB7LYszoLkhULdUzvOz3vCj+XiM
tS3BgneRSVg8D+z2GWhKA6NQCaGenVPmrWtCVw4/mKDzBgrNgwiWB3javMlZVmHM
w4YBaN2uRHXvsnymM0ogymh3F9LOkhvddWGopIXn3M/eRoUb4506gvxt4WFacBLd
zN4qz3bn0m/eGCy+GhCLFIdqMF2S8trGrQ8OWdaCliwIYPH+ULWz0sy3xo5op+14
n7955esRvL9Mc9qSMHgdmzemgzWRjd69+dkksEpc3fQIO8VlfUtGFYP20VSiK9MW
MCoql0lAENp+guCdZuBjLcVztoH4ofQ49q0K+6VRA3ZoFMR15bD8CnpO9Vzo0qBK
CD3eKYRLc0r8xGY7Uv/MxvZ3PMERXrRveBMg1CTc0WktlURb1d6/3cwCs2waNFxs
JHtW6++i0ItZJC/2kw1vkp1NBL1s3Ukva5UM25XtWPWr23tp7YM3wzJNGniNASSf
qLb9UR1rsMzDfe8F6r5C/gIkCjyjBEX5JCMpYNWWk8CuTq/AzH5D9yfG7kPlSxv7
k+8Hf+8MUSDWLZQlqUwvH9uHg1NB5mrqjox7NWj4fTUkNO0w6Qe9PWiSIB9k/d0h
ZmJKcyuBjm+JqUxrDZR+xqnceA9xVon2Ahfoiwt5kI9w4U2PTJ9eXyLUl7qxDN2Z
W8npALFR/R7mqEjeuCuBKYna6JtQ4bdmTcLoyjIbdhTfJvFTx+1+ijiFBi1E0f5f
C+kZsm+XkKWpsQlYLp/EZR+fnTRAC/aVYhE+DlI1UtXNkByQB5iAW8KtWiv9QIif
wje9kEHGLDI/0h/Jk4o5j/PtIzpW5OcG87bnRWiuvPYAp2TqS5+mqUkoeWXngKdm
d2rH6RK53R/RSs4Hj1HsVNhnuO2Hr1v9ipsWbV7bMtg12W/4kQeGl/mKmMPJWX3V
RpGlKX/RISmugmeOY3L7O0/gmCDUjBAbd3mc7YW7vabTdJB17dnCg3ovR8kWAB17
OVNwcXqH/uPaJXCgOxw9SjGY+pkvqudQ1khgy6y3J04mAgoXqaLI2stzRygtMFtc
WnKhmPU6HzLuYAcyaxwcbj9K3KlIJ/8WON2zwV88H8SSOpkZ3qKQKkN0ODoiGrFL
EgNKhp9JF8h+Sbpsu+egG41i0udq5521yCZLfz2GYGEwACM8jF2sqLunSQ+jfGSw
C6xTrrk/1is0PEovGer5u3uSplwXHxsPfAGOaK5BIS3+ZVFPixA8cjAe06g1vis8
Ro5wjMyAsmN7adEA6QMJyOiUsPo2yR8JPU/7eg0SbmHJbF7s+ImTtqS8PtAmd1AD
tDg+lMW3hXR4/t26wymOVCDGHMb3NfE7pHYRrkZwVPpkohs1vSJ6NmlmNweVuxH4
1FHKuJs1wdT/9EWEpVJNYnSfTW/1nXhGP9hO7F3l+E7DKmDlT4iahC7+6zFcyWtF
RzqJoDLzq1ZkESZ8876vErsw4oHX5gmxsQ/i8IuBTR96T8pnR9Pk1gPU/vpjI6/Z
QlKmQ7gEvYKRv3fNE/r3JZ+F5aGslJsrs1LkaQJ13GQZblKE4/I3G8XDwrZkmtX1
K6R/Xo0lBJX/OQt/eC7+9b908155mqZeWN3ktmjO/vk7KIsxw+BrQjgcq1Ja86La
ga8crMmhN+2gKrbJVdMpgcE2ZQ1d6/77KFQbCmMh8Z29EseWYQniOmkcriD2i7Js
oZpTtw7YAXWHn1uGkzxfaCW/qx5PTvrYuFzwlkes/nCTRw1qsRgdmBWCUSIuVNnX
Stz+uPqmwqvbkSjE9oeC3iNMM2gisQLsMaCuJ6FwwHaAA7K6hUl32vLAL16jl1Ch
R5Mak6u+VrrzmvV+QMlN1OTxhPTxrBZEm4seJG3EeHME0xpOSN3enj6ZFG5Z+IVM
pOC5CVCF36XrSmp3R8YUS89T0bgUy/jEuEYcf5gZswgGo6yAT+w1x/DCa8Svv7ed
cULqPFVe8lFjTYTIvz/JKb0sDF5AuH5Aczju/zrItVwnCp0ZspIuf03clBZC9Ezw
4vDaZ7HKPxQNSYI1esDxgZ2mLtlLirVC/rGYnLjraAL1wf0Imyb4NJ8mP5a+UbAl
/BQj+ZtwuCb7Q9jsGTKSOZZql+D1GZPhZNdV8W9TO6xSYb8koR48pbwGe4YW7NAR
IZuiRlB/E8uqdtXUguVOUkk+FgGYDNRMT5zRJXyTaSeyiefe2iTSV/gOhL3KvVER
/1ogw10aDOVGnXtNmrAte48RelLNshaMplsYubNTbZcVpHSucoh9iQM/4RUe3oFc
zxQATTQnkto1pjkdsHiFGbRPfnVtnnY0IhkBxJ7Oo9HOqpv0wjynspRqxsLD/kjB
pvV7GzGepo2DeNhXhUN2EfFkkcaa4DvYb2+8cKctgsghfrsPXzVYTgbq61KdEfNW
3kNQr4LmsExhy2/uAIisFNr31+ioPRp0DIi52KreV9Tl1K+43U800u4bdokjqdLc
KL/ECa3/SDzWNXiKp+vcb4T0MAQUSvzn2f5O+VzSeO/xyXJHanX0V8EUerBFHdKF
zOnUoePBajUelhMtaPsz1aGfZcJNfxr+mNAfSVUn/wyQ/q0CLhqm/vjA8eXf4/iE
rXkgT0jZN/RlXfdXx7oLI7L2yzOHmTQL+in38VSf+Psj57irYW1tSFeqe/1DAF7Y
sF5ZpPhKSAFywQHZ2hpqwso7PaolFqEoD0pZyL66rHsLxE0UzcgfdEMkUsYzXEgM
k2SjjynUFVgiesyW6mPjpLOnTeVpv8+e0UHbcSMngYuLas10dGuavex8KzGYkiJ8
4eXnuf98d/5LhUvDOmAfo//mUHHug0/YKr3Jm2JqW07DuJEvqT0Cyh3/bpoMzpeN
XJMMAZcgvWSgkEEIMwWxi8UpYKhmdFaNIXs1MMcWozq/pEswZHnUNx5UWR8g+F+Z
1msvPv8PJzmORd3qwvzqt8HGDsYKZ4HcCs7XcEq+w94N5VqJOkRkojFQDaB45ARS
VhtS9P15g1amxw30x4e5z5OAdoxrSEMUl8EsAEj0nwoozqr1q1iGSVR6vQhphf0n
qG3ePDiO+yylU2Vkc27u73fxlaGXmKCHEQlxgwir2ERJBdbvspwagblyY+bUTuDK
/aMqhMeqb6HViwBKotGNF6IIklRz6ehXdxcKLdiYDFLZnJ3RVdx0jAGwfeDCN/K8
IWzKPFjn7SHPaghFAIsLJj4uWTrJ2Su3J2pz3WzFobhRTD3KF0Ny51AdWCny/Y8V
eDkktmr5eIP2MZgQoamgFRHpY1oioy2Hg1rkt1ugp0JiZhBeSAGfhzrSy45ZEVIE
xTBakiEbayKNnBFN1dMKljyZ2hiZERn1OxTAJZTwebCO48Y0qmyNIdg4uWp8z6DE
pI//nATFX0K0CA3RlG/MQeEoprshZG9RHDmtmphdrSjPZWFIoDyhGX2C9sGlb8+l
wpY4FZ2NUslAN19dFOI2zibzgRpp6MuJxR0W+EMZywjCOGsAf0cN30SI3KGJZZCw
zXppCMYLRLVvBkYJ6Qjc4Up7ST8YqwDpu4X1XQ7YyZrL0Nvjxrvwe/XpDzqRL14V
djRhKPNELZaR0J81r1i1nkokrZuzKoWyE73tQpL/Bp8hwACf8jLBnkcOXrvIX5RJ
fXRi3GLwk6mq0D0yJvo7su3LxVRgpFwxr4oJeNvuDEDuF8t1I87PsP+H8kuAEZGg
yLhF4rHApx4St4UA2Xb9hd5oszUx5WIB72KqNVELkRaDS2NjfsT2OWox+5sE8K42
U6L+tFpdBqkd5RNYNhz/K9riJJzEycF2nDSVhKmedn6Z+nay1MpDk4ipBnix59Uu
7FZsJ6ygKe7tOnwsI5pVmDHTtJV/4oCPyqZtyQDfO1y9qAtZLSxyOCYEcA4K65Ki
uM+ZRvlkXNqo6GbFuJ+Kqugq2X+IM1QFTr6y+GZ9HOpyLR4xg9VuUTOACIDKdbeY
/Pm2Alh0pQ7+99g/AW0Fl7Kc8ktHSMIUBWBB0G1YMLXH7fMCwv8KHq5hinRsBHfa
o7U8McKM9C2HUXTzuzFXn9g0mOuvtB83EKUwD1ePeZy3AL48T009NLyc5elvsfN1
az83TJKZJ0xxTI/Zj0pfrm7jpQ4l7FxIUEykioeijpyGUKByfAkI94zpXb3RXrgt
mwvS9/rTrsEAhyhJPNbxTuEe0twUoEzzRBdQl5/IY7u/tSkj7netdRWrxrlghtbZ
nVdPPlSR3fG5iexoV/sGg6CAzs/44TR5yJOUPWZHZS6xJNN+pZUQWKWXeZx4Rxxx
5fVkLTwGB+jrJX6c9uYh0iJhPK1a8KIQMe5yJaeVLBiVGL4rZC1pnkewV6LslJPK
G8QKx3dGDqqM4DdmijmoTmTnVr6ykFe31XFRWWpZOMSc8N25DpuhcO1L7irTPqUq
yvD2R5UzoJDLujrO9gwOveBefeRTBzSAz7N7GpPHonvvXmrMyVtsFnqVDG9HiITy
jjy5i6wyeG1ban6mvnMsRmgF6FKWfYabaANCUClfmH28hWiOF4VbL/dCiKfjihfR
t3r4KYF5TvNhN0RcryBD+BlvxUuYThYFJbHI4bbEzmNYGjqj3OQTcsEcyI6EEFPp
uRqn9sfEbOdBugNabnqkaB2xX1TTDu7Unb1bVclgXk4yXmf4UmlkX1ZJoB7xwW3S
Z2b+LMQ3U1wThSfDVp0P3GBJkWRPo7ev/yMgcLiClhjN34Nd9L0tCKo5SZogeLON
D+9cTS8IYa4+TJ75V6pSj7PygCGhCLUjd8TumehAZ4UeWErh0kjvRiLd87ZZPnnS
h5SB0x65DCGeZX4MXFSSOZ75OIp8CCn13cNiwfCd2AyhryE0SRRJjbZbi7i0dEGu
6FzSib3kTxXn/CDseOuVzmEawVY9VwzLBn63hARru5lxL2boUzfAeRO6GjOjPp8I
V/aCILW+otfGpjbkSTYMKpNi3V3uyN7r7z2lg2wnnnsoNS3Bxj6hLcPt5L0YNUqF
f6Hkg/fctEDG/7nbdQeFHOvgxr7VqIaVVSYEB64C52Sq1UPZMq+A2mYvLVen1gLO
9L+zmyh9IFx1WQhINxuPJz28lyAoQdXvg0rMd0YPLXNxE9sxbOLYtkFvnQOuuKbn
jTEQ7yT86ke+ddCUwp91waOzAJGwMcHkVlBX7iHQQE1EN0AxGZ7x75UFw0mk2STw
pH8MoEuFQysY1Lyn2iEo/0ak05blTsJcH7Il4KLTkjIsFbQv5kT9EJWU7rDfzUzk
P1/TZsjuqZwUB+v8rQ2q0Npt47A9GGIZRJZP88IUGCFw3nefLmNKtGEMqPtatoig
KkEywB78BPXtlkA/aFpDGxoFcmOu54iGIiyPqKRRTE3NSP0eDR2xVjgRLbRmHBLD
OCWyJgS5LO9uX3Xo2TOOVDWJxMFTnJxUlaS/hBKQwLdWq6Q/MSLz4UN5kEWjITIl
Jn4pj8sA9I1dA1ugZ9FTqCbgOS50uSxDfTtoBODfiw7+OjphdRfaXzZyax+0hXSm
0/lbsjHrwRvhUiLfS6Rec6jLQACpww30J2GiXD61zOKiatnFpb7afHRN554FuCXN
RmrkDV+R3tO7h3PECzf6yQiDwYCnL88Tcc3N1y08YCzGA/Ub6XDk1QiAJGNEuWI5
jpLNsOiIf68T9i4EKxr7kOU9ViCuR4sT4Drrk+734XaTMRGuSVvKL2SxjycYoH8w
d0bDoBA8OFXyGL4VL+3qnGF/lzKx1kSoSrZwoV9B4EaanRO8SvCQOBbQh6F8aIh7
wNUWGQUXFOGOCI76VTSv1vZHl3HxHqgLBsK/Fi/0VD9+q8LQ3BpEpVzqrB+prUkY
2RjmjBDvYY+7cl4eZ8OcK3mxDEIEe2QSgLjl0bR0DbGzRJe00tksJbDqy8vLBFol
eOJiRF94MFHSQMm0La6/IAYXuMM/cS50YXcEHsRv58jsETnrgaYmDHMpt5zaEdzi
ltNjC4VkMdBPyjb3dGKz04FX7xNlI/Gdlq9uGK1bioWi4EMolKg2h9+lUHwk5a7B
++Dzy29UPIJChiKI4Norj6xY38UuqFywbiJ73Kxilhxq6isd0y++5kRI4dUfUqCA
d4zbZJc1DhY3Vg9rCpdMYL3Nv/hqSQVQjbCeZTHTbS7hPuCDfDk772kEl2io/+Gk
z0VondeCbS/r+gAWqIIE+Bd5hbrWHtWgcR9uT9+daV8h86Ew2aOYs3aHjfvN5XEE
QZByIHY35BBTpUvgsJMSj4J7gr1GUA5vAEuY+ccDz89h8GFtwYcKJJSjZpS1IKhW
dk9JHfYBTkOwemiz6fP8gD0Wifn2R1MAnGo/pBUVOz5JAmZ9YH/+HuiiKbo9LHX+
AyVEBXzQxj/ij/suR7KmSMkm3sZqOY3URv6h629pWMfC3TZbaYSZAHbMdQJlVdy6
R3YpSm64EV7U/lpiCSibegsa4mKWjq3fgHy0I6nV5svGZMSGKcJxi/vrRqY9E0Nx
7jSPyrI3L4Rml1dl26YLnjTVZQvdZ0flVWa8P90guUc1FgmueGytDNQru8fMdkEI
QbQ5G4OIwO+Lu1f3+jG+ste0erOHjDgA4I/pDG6Q64xS1WbzWWaw4vLVQEfcPkj3
jYVlxFI2k96zQe2WsNN8pTut5FGSIObcDmqLE5dacgdaFI8fhdvZpRnXhCirWML5
fxdL4zQ7XWYo/FVdwDjtiF8PnKbV61mWh07AI7tkJ3wwwR/yTSUvIVUEoChuVL2F
sBx3QQIFQz11BiMrcRgmTtV6uE955JijEmuZUt5p8+qCMk3nBidfdNrytLfOyK43
SaW3u116E2tQAKDBCOZ28Sus7/n+1V70Sqb7wHnldMx8kTvgwf7ySfX/iH5HFpHQ
2YlxxJR04Z8nwLtZbLlid2vpsRqH2nmQSGmf8au9luiBxxU0PS1BIXgZ8Uk3wQ/8
/WiS9KDxhddinnLglpKa59pD5RksoWF6V3s/hOqk+cnRj7ZTJvGoeUVjRdWqifMq
0zIjuf2J73QdpFnFmh8lU0LyVDb/zChfTSZG9Y1EDTFaLAW0ReKY13T/ASiH3Nq3
XhgZoHB49j85nmGmIcYLFKIKSoTzXsOaS970Mr8tS6w9STelyG7A6WGUAruKfCuJ
GKiugPzb9zjcwVZdsRS+mseDb1a0geUcjHz7olQVG04TaBz3xgaM/V458GoUZ82U
sf4D9jgDjD14MZrCjo1ZMElsuyNR3e61qNAvQZ8TgUdtrRo2dmxIFzxMhjWgMRwH
KZ/PXUYvkwYFFA9ufsiasrlOIq85+KBYt+cf/NQCGdTV36J47yRNdw1j5m8qDZ4m
pbqLl5Aa0JA/3IC5lUpl8eq9rEl1zgHeqDZqeFen2XBCkc5+aajTM1pQXbY13HN8
mh8KnWdU5UDzJDnk0Dm9NeMR8WnKO0f5rrQCGISun7UmPHEhyMLfpx7V/eTgwLjx
n3QhtMIyr85nKe+wTKas8J+kNfEBgTfd1ZOGx2cCRYv+z5Nm1u6TrSVDWcXiJbYP
AxqK0IS+x2hBictFXYRaUeYj3GrnmXLZQY3Z4x/WY7kNEKFrpztWeqUWDal0LeMK
Y26BIMN7UXPQbo2aHeGFA7Xcp1R0EsoKopFsr5EDOPAn1JB6ilvzhX/oydCzWFb0
TtDYWiwdOg2E6hH3sIhEZAXnCPGMGuXAHnhewlAFQkeb60gLo9+s02RaLxbp0vAG
E6xYfkxk/9QKSU0evg8ISqJQtzs3t6bn+3nHcQnfPNg7L3/sUizvMDhK/ydFfn/A
/ROy4CcizQtpZuQamtylFXUbZpoK3kSgQ6o3nSgBA46zMqZPQDkPERsbRdHbnpHp
iJaJCb4MdLTUg7Urz9VL2OG+hCuQUGQbIGSO3tBEiCr39e3CxmeK8p8MDRmxrHEC
7oXxiwAltHll/Tug/Ro+BQ0DBkeJsOdYQKZtRfxTF6AciRA+C5YdzG8U5FzNJv3g
dykqpI+OIcOKZC0yopNgahX8qPpUr1Pz3Mckq/h3gRXFrIbE1Z095B4hYNvwi/8t
VyWBnYSps9FlYhe5wgDgJczDAp/vw3FAdviAMpVXCBIWsH96jceufSZLRorGz253
Et54VGweL9uGzEHZwNeo4KWYMda9JtXfCh16uZScJZsFSC9toN/vpVsjDPtVorO+
qu+5izSJs3ajEJKBnkVb3wZ0BozThRCnwn5wGVSarru+mC2ToiOtAPGzPa21EHTt
3QfD0WUleNsJZkRtuEbNbtBXD8YSePX33b6nSzL0tcMzr6kjO2KMyCZvhlZzVFMR
EcsReve3uvcrm/nF0QKC5sktg9W7aPtB6RW5idUMWvvN8nK54941S7VdyehCbFFY
X+9EG1Gz53eZr1wvUwpqCNV7ryx2sr3sotqFvG4Cs7ySthsrJescpp/cVAQZJpFp
Km4l7H6prROYPoN8ye3em3jHt7znxEeYbJUIoWVjadxao0puPQ/pa70bsLU9Eav/
KGGEnfIdfas0Wgdt4Njd813JfWur1nt8G8TT3YyFk4DgLZXB4rvUt+MXmTJ3f/Pp
xKDK8viPnTNZlrP6azco4o/Xq/idBCzMo9xwzcA13a/F0uVKu8v8JV43xIE8ZPpf
IrapJyNX8fUtv3/FR8SLLcH05K5+MJyuSdSD3riEq5YOs5OPQOBbvk9J3oRjKyld
BiG+jSlW8PmK9SxP3s0IQEmK6Q3z5oZgG2hPWI6V5wCJA3/5kYNwYg8S7GQwO2hH
j1SY6VDhz1iIp9uR6/7Eqe2QLnEGGs9LBKJWUJsJTVsI7Lt+k8zYGfMsLoLoc7jg
InhEgqVpqJCCjQLEXbneDYUs1oi2SqmN4OBBfpQKAs7kH5F0DBs9ugEsTAz0BdSS
3BDEj/qP3XyHdUPQaLWp5HRMFyJ3UaW9wPPmhBZwmgVphq3aG/dSMBjR/RDdTD0E
2LfKznQsETZcGy/n1WFtKRTyeM8cKTHYOgFiBQ2IR1p+QB02rNw7fvL5Mc6zaRpF
dH3Os1rOhIeCXQWCDfMhVa4RB2xCsRTZoBeK3FyBKKSgQHyByII8N/CH2iZNvEGw
sQ54w0sK/OzDmdvorB9pttPnxYM7p4PD6KG74RyWIoEvWoavKyfvjESc6fBCaQMn
92VfYng8nZcrn/ZC+WcLhh4raXkHz5ikmz8LdFy1HPdkkcuUZ1Sw/ssRzN0EgG0T
tGXjpKNdkd6rTptuVma4Acx2CBKJIO4tGOcHhQDgFNjoBDyHGH9K9Ra3tUnFOFf2
jco5ZNjgUjKO0l31fva85lXuqfDwT/EmyvztXb3YRGLUzzdTPs/iscqn8gNK1ZhM
CqBtfdqf8hyTpqgZhKU2cJt6B8xHS7UiSoP/FtUQmTnNbeNtXIlKJlLrzjx6h7K6
7IiIJYDtZWSD+gqVtULFroTwI7I2gE/P+JKmkk+JyHn2amj1RR9cWecMPcNqzwnL
ylcM7+f8BLJ4U+mn1gDaLUea2/zcFthgSdTLZkHwHDI/qs8gcbHLKhqpruCtsYoE
zXfFCZOye0PD5W2xWSm91U64iq6W/mLtyhf+jkMAXbDVU7lyh8ciT6vD8O9UEcOS
If5uB+TE0PZC0bNZ1fAV7Tv67U5KZHJosAiDj1SI1F8f7452OCnHflnh96Duqqic
zBR3DpTrXfZ0Otda0DtIfWr88n+/h/XkTnBlLEHRFATwEwnFdyZmnIxKTKyeVQv7
ZTI8bhy56cDB3N+5WrPLVX5OFZCOfBb7F6H7WbZvpYjCarqzjuDA8HVy6mWIl3/Q
IWLEdvB9gS0rE3j/vtas46TSAC5GOCkOM5x1TaWDjHdwhLcwbagHtX9fCot/YtEQ
ElDoxkB/f9WpzVPJJxTY8x+gMkIOHzrnRu/SUMCgxQoMvuEdaMeY8y3XLIFcrhUh
a2cosjBG3smNK0IIYE20j7QJS/jU9Ns9ZGKbcsu14b13tuKEv3txgfbEBaaBbc9r
GCfzlu/9bZo1DvZfytkyLYPPKg5qwbwRn4RVS+JPz7maFi7SCia1fPaOYD4dIUEk
TWYxNC9E0dfEsZcqPVbJsWeJmgfoUgE+dUxO4GJKZyOH1e3ttkmSSXWxxbOPueEj
E+5G72mmJKW2HzsUC4/egdnEZSxl62D+wLzTRhKKYib0XKqg/wP5J9x1tqOOEkZ0
nYTN0EKICjuuCky0oWsFFTfS7zru/Xdjrdr0jjO+PLpAFpXe5YDM06C0UI+VUq1e
fAJx7cCy8yrZ9GOVbSI4k5HORqRbG3JQ18vJGAlGZ1Gd0KSceHHALXollJ9O/9HD
ZWvKAoinr/qtclWz9p4Tcr8QEQ3QN1PI+/N1eT7UUqwbq7AUHCeYYH0iX5NRVK+C
5jWxPDHOz56/qVUdCxWeF2rMvZMCAkbNO8I+xVJG2gSdrVNDmKgMgcgqp5hHi5iU
OMJVuQ8MNYZdiFh/S9aCixYNanXXWLyxF1Z6Jay+T+snALsOOtk4hzRJ8oBjDzLg
94iMyu/bJ+sqMU959xQnvct2wg9rwte0V8qdPQ+TkOS99Rx1q4g6h3l/046CujYw
/VDfhxlczomdonEQ1KNvbGdbG5Q0Dk8rnjbUfLoDdpqcr0dXaG7Q1EGTmG5L0EDe
bcD9LkktUcmiznVN9Xa1W7ZKYRzQWxYpxahh0pJFjZKGd2at3E4iT89OV0mRDnu4
rMRYjd4HlutYwiw56NB9G8QJepkD20t7N4Ese5OPQ7fUw71m5Ka/Rotg9yemuOug
l4jo7g/Vds7n6m3CYoIhfuP++PAPKsiEPUcyD8TfNrUQOESuda6006/dRhtrb5Dw
7XtIYMbn79hj5UwHKwM+Itbu3zKBDn9IP2j4gOKwOrT7ZM1/fRQwyUcKn+4aFJ2n
u87JGA+IaNvFVTNceL/974e8uDuN0+1/k4CNXeDHY3aVkUFi/bk7ksheY6o2kuP/
rsRW6Z/V7QPCBBjCTzMqgg3jeNhoqJyZF8MSTD3zrS+aXVyXtGIHlJIh3b1CPwgq
ZU38XUe+mSUwjQXMRqcqHC9muIU8YGMCthwZKB93795N4wrdeqeVMuOOIUVazeIS
oidcoK+eQXqjq6RfEQ9z5W4ch5xbE5HDurB2BItZk2h8y/MrejD2c4wOh53NqbtZ
1Zk5jmo2ZoOAXkO1fxExwwKb3+DPZpg2HaPdDvDs7RqFlEQPAGPPr804Y4K523iM
jXLsfeGsl58/T9binf0VQE5hh0gm2rxusdPM+i1GSYyNqom3M/0WBU9Ev89cr+nI
R019p8DHS8Xw6p51IJjwo/cvdft5TuE/XMRDYaZDF0AnMMH/vKrUe8nzg0lvoqhi
YQZfQMkYLS81lmi/5CNaFrfDGFVhEfIR8W/UbCasQIqFfke40qEKmWp//meYKeOT
zGwIKtL+7Papc+VYUz0XPmaar2fP/8DfEALyRJbS1A57nzaIabHrdmNA5QviNkOY
sXKBCbmIaVVo0uLHSepphdo9EivqXUNxkSsu1D1KHtMGJoVoqGqdQVUQ/Rx4D3R1
yZ2AivVpcoa+HVEm8XewBp+xBt7Yh4Dci0JLEtzJTPiHDbOeiSflw720m+AxAIE7
Q8GcR/Y1Ov1x2YeZlTXlmUzHuLa70DOfPKcF2ZjRBN18AiZX3S47KA6RRtIdeyjH
szH81NRjFknEyLmb22PZ6pWyqemm0zFYt3SNcW3Ve4AbAOUl9481aFSTwQxq4xgJ
CT1gdnwwMgWsBAjSb+VrgrytPZyN7It94zYCSMLtKg6AQMx4CZYRW1W0AukR3UD3
5JszWkWlWQUxs47VyM+Y85GfbZ8AHIGUoWmvZc+fPeUjybH+bHVROvE7C4guJ+KR
EuDi6TeeDxE98ybdxyjk1wzQpczCBSznwC/t8kyyxe4vH6XCf5/Frx03Bmeo769A
3rXuRfZIH7/3QIWe+hNGSAEPpBt71n2RbftKBm1zqN6GqAjxfU+7LVSBkAoB0t50
KmWj+Da+UbcSgtZkZ3/MU2Fw/FG/YREG25UFEcopu+itv5HddIHsC6+FBNY76HXl
ilF79lKBvIx/7Kwiq3c7RB/y7IQV/LwmmeEqoYVuTBFv/FKKR6MOsd/ucQVIUB43
371D3T0Kxp+bzav+xuCmq8CqBcZoddsAMgtevHWQuBKkjl8kmm8SN358pU/MqiD1
RXxnfGzVQo2rKpVdQgCwF7fQiXDoPZHZZ0iN9iclJUvQzPblZxgEIsvrCIvQqcto
LcZY9ky6VAJDFW7nAGQvfqBh+mIErHuBHNtJ7pUTkxBfb5s9zqyZljabqKbj4b4X
VyS7e/HgetdhRgCwSZwYPcFVw5ep95OMoNPyAxMoQJrEdeKhxHyKgMPviUGd1Olm
4EAUaXYgY8NbZunJlC5GAZ9NrYsbVWPnKPta+lcJWbGrKRK1m8MF3JiThctbLUzV
QKuD3+tEp+FPPgTFvm1BC6iDwKFegm5ggB1eF/B3JICp9dWkmkwvgD9PPj94EZ2e
DFN9BNhNwLTes7lZ//yreXaKY/xapYPXOlJhZw+6/Htfe8PhSMW5P+K4I7SbDfpi
RdmZoa/TFUUR5VWPO6SbM8SQFZXGoRE/E580wxueQ6MsrToz8ZuLGyHDTqO2vkHI
hjFXJIy4FMpC2D21T971/KD6zub9bMFd0h4+LLFNUSpRi9yC+5UAg9ckmX0r7mO0
7uKBZvYVgPTe47LVlBjvg9BA476ErW13A+OvOyjGIMuIt6wmCp77QU7hQKJ9Y0F0
obGik+xJJqMC7h43VZlijGrVaJgB9LqTzNDGpkYVis+ABCwI3cU7DZnLZp4DGpK7
LQSnQ63/shuuRa+vNwAWdL5OvNKvssZb0DIoZAd3tGlnpoa40goFkIlqkhrOd9fF
9BpHcreFNkVl3xhzBzqEIgt6LbkyAtjQj+lir/2OuglGuTUKIVsXEjOKEfMx8elV
0oVFXx5NPGSxzimg4xw/AQB0DlfL6lRaUrJFsDARGuc5kq91Cxyo8OUrXlB6oN+T
RiCF56DwcS11hWScE34gg8z5vyydib5QXfkg/y9q7wvR5gawy2l3fjAh9E4lUMzP
oZyAiM3PE4Z7LwaCcFQZBHk9EvzMVo7RDTCF0HktiO2TSCaE5+g5vHJ6BQtSEr4G
gJ44jwKmEF7y0x7bTD6LTXyz0x+ixN/9hMIto32K/q31YvhY9u7oZZBMn86WyLMg
HctjBZUoXRSqKYPyL1XHyuXsHD0/BsjuugLdXmGsjmGguGf/X6njxxTCEMVyZHUI
cfvFwN1pN25umjEcAzhLRJGw4exA+eYQzuGLHO3QcWsBxw7DQtmUX2m7aX4sPQ5M
WT0Cl5K0O0sHJdZO8KwrybZaiUHQ7s9c/iUiXlfMVRrfwkKmpFWAltMyMfurYzdr
QzrJuFGgGam5cpWoxdzO7SkTA3Xvv7Ndae9T3cYc8LbPBUhbUeXT7EPbGh8tRi8i
T+jxxYmXhPrmF0rRbIpIZdO8I8sOPgHCz9HlIqsS0QeVnBLbTTuwt+WnL9t1Ligi
6YD8ePauaiQZJ8kRuCw4kz/FW8tznIeI7gvTjhB9uOZDnlyZSl2HLh1nH/hiuynQ
qlQdcOkyFyATMaCK5jCNuS25IBxYrjm78S+3QkrrVXZBvaK6POAY7+wnhXw32TsJ
V56GZBrxTRX2S95iFnCArG1NdoNbYPs/nzliwjAspTsBdO4rMF4+3aVgjzWI/xiD
rPSIoX7AwYAjFJ/lD2kYch0oQHEkV9HKyA50mYwD/TeXRIzpUReYNs0XkwSRETfM
Db6g+8XGmw+B2U6Uw3DuZEnXnjOzRvpRhlG31+W6P0sLXfKW5eBK8AR0Isj1xzFt
aku/JzmAOdqcsJJVXYleEsNApWJ7jmsjujXuMGqEoT/CngUK0SSBwzJHt+aOKDUV
Df4FsARxay2Yuo3D+SItObiglAnIKuoMJxZLB/Rv4GTcxUxzzZwnsFc1niQx5p3x
8Ugj1lKeqp3W3Z/27xWvi38N227i4CEZk5AnHMI8e4B1ssReALxhiQfYgZnmodVi
sRBlsx0XnxowngUZ2eWi9cFNG2ilOd5NEVa4cprMXR58QWsq+Cen5RvaxSokVWIK
ovG7LP8rAdsuporDMmFEXUJEtl7JWkdy86epAEUPMUbv170Wx3bDIfOtVGKtKkRc
RONomZAMb52RowkGS6pi8I59W5K8PHRfyuw+URVIqi64kHAEZRZ0y4L00J/yJDCI
nKt2cSsuZAWnZRrDItu4oHWeSSvH9lx4dOvId4uW8r6r2ghUP8AI+l5TgWcIxbE0
98mCEpZRbQiozCMDmCCkuUDD+pl520ScGt/ef0aHo29KNUiccl8BNAAcawoaIwcO
jj078hie4c6eP+UX4hraSKVXZbRbDrkX/dwAHrX8eI4BvItqUPrcpxPrnnygExRO
KZAXlj2Y7ADky0NbUUPU32AGTe4Zh5GCJaY5q9NjyWB60eWFOJi+vtZRQ5QwGVuo
nuMrkRMjqdyQJSFEuOU79Wdw9v+afhi0yuIJ0QtWn327b8L9nchNFYJmBmeduw8/
HEoF3go9bvjAwRUyHSPBRtXQvTmvatPCzppYOWn9SSdnIvSRZgvTb/MrQyYn37Ro
lvKX5A4U8lnTVxIOmdnWYL2jRgMdIA3XWh4ZIF67EA3QthPRB4oHk1dH2/hN87kb
rOvZ5JaSZjXZ/OGY0f+RXBEvRGZcNMlgHBRDHLJcud1aQDAXZjXiOn7LAc33+jGh
IdqNJtmFBm4dkdq+h3ZEoj+p1HYNaBLDDpIsm0W/UK4SWUlH+yZoQMjJAl3p7Zqj
ql5xMUjs/leZOtA6qqPahQkgzDxBoEHgAFAHPqWvGRNKpCLGEPWBiO8Jvkl+rd2D
BU+9H2HE7yUu61UWuWzhKeiI3HqtRiRi7exBF4vXRyaqxQOMTn8AlDT3J5c380GZ
81BQ5mBjh5ooSYH7u25JnqVBZ6xGD/EN1T0u4lKc4uzQHVVDvEFXUDpOURh4d/TB
9XBiTH6xBBlespY3kTVpp5YpPJM4dCyKNQJBXP4SI0OEMOL7OkdYtmppAIpmdBa6
ed5ty9V2UbB40wVZd02Fvjut+ueJj9JERrdns3JJhfhOsiaWxUtStpHpXf2d73xT
iPS6Ri6pKjFGR0xj0Lz4FG74DyjA8Wez+UU6yCR1zqmL9KHGV93ahc2FEfKSrdb1
scECKz2C9UChanwlQUI6KgV3+5MYG79hz+itqZbgaGN9/JFe9Pfvx3JB3KI4hsjc
MvXx/OUGi86G46S58oYROjFZSIWJE4Jm9hrhvTTmPO2ZZbASqFnmnz/T9g/xeXfy
5RFerm1y12yeB0Mv8UkJoDW6vr+d3dLE6Kx6h9oVh33w9fmOJ9qigumaC3LXj4so
weHDDrJEMrvu3+efpzVvyTb8DhFKaad1leRLr+pZskilMePg7gvvGZwT2/wXVLtW
7wKg1GtqTw5LhYf7R+ntGWv9q9sty0eM//OwywwCIdDEwM3EHuP8jSTdEW5sXsBh
w0WnuW3Ieoq8Vto5/n/+aPQOxEFw2X6UOjkSHezCU33rB3j6Z62IEtcNl4bwjbBs
ocGbRsuNYxp3OqIucBUYesdTC5lcEYSuEiycHz7i7LNeqNhRs0snmafO36PsqzF4
7yiDuxrniD2sF5dykDFY8PWxIpiGICBuABekYbGmwXvr+xPPyoAKNG68yVX+LHuY
IQt9P+Hh9zf/NuAiQqqTU/Fn4i9uIEfgpafHA/7LOeZqAB4m33A1tLmXvKidBJts
lo1VXb9flHu/6M1Jc/H4nt+n5T25WnYtg7/jMCOnFVQp5yY833LPp+LxB+7LYtEQ
0eJNpnuVG7XePmHcf0Xma/1fJy2UGzbTA1NL5Vqbi8r6khAcbtprVIoTbk2XrZk2
D0OfeA4qJQuCiWAziO61V+zr5Fp8bnIHqcBddQYFHUmIIwbOEuVTH36JH9gPYu1J
tLPrpncmwy6de0RVXpokf2HXhZaoDyN4e/cUapZEq7XYmyla0g8ustg5+p20RjD6
8Tiy2H+8yTtUQRibUi9+p67i0NL1ShH0DHdT5e1j9IkuXKfc40mNlsjTdil/krda
xGH3z1VF7jTBvB1+5FKzAwe5f23q34vCqB7Ro3ZqmrpoakQD/hfnGV/23+d2ICso
D5fKCPSUdr/E1T3xIUqLQLzKvBK7SZ8TxD4PTpKSZTeRtnmbQYnRT7i1ly0SAVak
Qi2gyaRnQpwvlCl7FtYDFjFauzEY9KPJIfP+p0b2pklglaCFvieWM9eTdXD4lRR+
NhU/p4qt7ZMfO6LvjhMoTsbXrCZ+UfhYocp+RwdDiFalAoy2BClxA4EDwbNTo9OX
MqPhiZFvAXBIv46bgXVSRA8rFfy7wQ7wnxO24wO75bvt725bxAqn/+BFV9rbBk5N
rPeX39fr9UujoH49AkIV+UV3vWN/+lCJolOnn8U2tbNJypoc+ZXuKzYz+KA4KW7M
Cc2hXWQS+PqvB02P82Yc2bZ+wOBSKEdKaWUsfMIbPdPcxUZ4a56TDQPaNh9wnerP
l1jLxS51V9GGMaGTtJNgiK3B/i5cwT8ddrSL0LEnXeG1z3Spyi7HkJCr6McsNFuf
okaHpTLFch2ZYWGAfxIVEAk+63wqySOfHLmhddTLTZgWo8WdPGWThwqDCgjBwzGF
iAEEmrfWEzvByHsqEqG6n7gfZFz2b9MJKLeatgGw5iFiG2bpYXAHFy8RvRPVmQAq
SyM/yNs7pq1LDnJ1xFDQt7rINpd3UEj7W/6Z3F8QlZkt+DbiyKF8AiO3WwYeMdXr
QSRAlqwfbdPvODlifmIW6gSVCxmwIWKR+oeT0Y10ax8bPwSVhKn2WUo1xrWQvMEQ
8a4+ttRQM3Xlfs7E9+1JPCK+auzI/QHPHtBNroMpLy3JZ2ZuL6BV4s2xwFhs0LGA
KbfKrs74FhFuDLLxI8JFGzvR/6RQnLVAPQ1OfG45ouimOt3URutmem8LzmrXJhX4
NQAK6n/N8wT+nish1VHNPSfv3dooaCxusPGKKnfrqQ/Pwxery4D/sVwq+qCj8o3B
9uY6Pt3V+6omZPQV7OgTkS3HZKaYsJVib38AgWNpoNXvGgfVePInkIHDdljPopos
4XaB0kg6GsBllxNg/OlDg2Y8uhU6pDK3bwbCZX/MT9tEFMxRvtMn7Vm0GTmoawoP
cp3ghZpGiWS5d2bNNL4Utxg9Qkh1P35X5S5EMDJw8S6ciNtz5fkkJbNZ5+1pmoyS
FZN0mAb+RLeKYZxi2sVcfjx8p7XZpdgutZE5ynLd6kCKTZUUjzadmFYaV/dGLswa
HPmH//0k5a6osaWDJF6+p4cK/CijlFuAhOgwj5FP7BUSsFLL0zCXhp2OHKEg8LwS
jKieSMkBiD/346ta19bCty5NBti53lOUERmNT0fYKESrWlFyp3gjIpZ0dfZQ9vnI
yUm4KKqxt2Rf4y9Nr21/TRKdwI+XufRGAZYfAOu/+AU4dIgDLle/XV8miHHxvW1E
JCJOX8Tf2z25LjY+cu6C9hEZC0L23STEAIZzJqePy3aO/l2ayuBdvbVTB3yTQlw2
SaLd9LjmMZ4RE1nJqJ5ym+sapeyi/6VEoC62pUk3YlA+5sRmf5vKkpAAag8rb57R
nYUK02im+Fij4x2M2IfISSplIRA8FLi2t+GAHzUt/Y56q604KM41H/o6Q1/A4uqw
ZR8ve2SnzzAvwAETku72qmtqgBnPTtMlY+G/xZffpehimCjmIDUSg15KaKEtaz23
wmSVM9N7OYv9eDYd9OClP5mZdAsdmZuOJ252/ZxtnBC/eNAVCh/LFuFb3hm98Lva
JqFVCEPpTHBo61xaaaNblU61pap53XrnzjrkgUuEHrk5A01vssxyuWqaIlvBKNT+
ne5S6M5EMrgqsWDq2p6Xpq42+7a72paQ1B5VB/zbS6SAfnRrh1xYJ+owjTBZmbUk
689Oa87v/3KZ3cLOxEJggNCF710NXWiKGqMFcEitU3rFIeAB9+uU62U4nhUUkHSb
wDbdDytlxEXwbHaUuu63RsEXK7pHa3esIuDOnAQxfbAR++CY7Xg+0jDo67KZ97xN
ywZz7il8Tsx4an4tDIvHzQe0YisQIVKUpop0qOt8dE0QY+yUNcZsDlNFbN8VS4OX
AGE5fAk+D94Z3rbkDBWFIzYQcNcH9MEp2295SeLcq/wfMzwYT43+rhCjyrHCbJKf
MEDulDS3B+fYCOuk0JYG1JgU7DEZC+j57TSzXyW/jHVKB7R++wxS9ToXcXRuUG1W
pXpcMM0Y9Sho08BiOzNHvwgWg+pLe3Yfw4WEvNlwoHfgFjfv/ue+x4RCJLp2sGHk
LBqN97A43BNjtFPHVA995dnMI32KbZDrvwrKutcjg3fOGW1cQDwEsYP+B7I6XL+B
Bacj8ak5a6wDqMvst7ZcYphtdiXsMUupTHjprGqPtxtNq0Bp9H1RUlVGXBiJa5yW
CtBkAvWrtLPEKXCJAsLI6WMXUYNbgQxnXGFlFXM24ouKEuDFh1GINCHr7HOFwqGh
maHuwdHrtgd0zpIDmc45eRbC2ldkvlbT0RvNI7FQrYM4FjNQIpQ1T3jY4kfXSp5b
PeM6YIkWl8IG7shmlsb3rl7Pr8+CKuq1ora66e7BTi194nDi+VDHJ2PoulVEt9Y3
P9MjkI3QM/YhqzU63s4cvTLLm5UYukxuJWKPbsQC76HyMksMJkm729hZpPj+VIIC
DtyjaiJpN8bVGdJYtiA8e+s34QFZj9lhZAuxIpwh90ZkOnY/wnOdTcPPPUTOU7L0
rKmG8JsxBxP2FOP9kbC7JUR4QkGoOWU3vcHmnFAuL0SgtTVxU1aiFG3Itvur2squ
GernHFKEEap/R32BxyHG7xwXc7+BFgLT0LRHilc4xpzU8+W5OhGZzeW3pcES+/5j
yLvPbM79SRGp+CF8xwuUzDNuqpm2ze81ouc2JwKjybUbs7U2p8GcgbpCAiWQRbGD
12CTdJMdEp0XBh8T966OhIDeOMOkLoAM+pWVrX1mvQb0xvsvRlqjddYHH9q8/0Ro
/nA9Z9mhF491rYB0srgvkNKylSyGKLnTSGX3RTHYUyqKus0U0Kveg/L8ovHK3ObL
h05m1oI+mKLrAxRTBRPel/BgjEISB+Zw6dwK+3UHyA9KACZEiJAm6Kxez4DjckQO
rZVbJZo3VPstkfaJgN1XhJkBlVGVrK976r/aYG2vEQQObvvFRyf/c4Qvcr7afuki
rOHBJEIf0Ez4vIIeCo4OaraWBt8iaKiH84axZkWKNYFg5fiiNCukQ9sbL4bzA8Nk
baBBd5SJQggTYPNEHe9rb57wYNJU1niJPP6H5zfOGYQ/5FXyUNGRW/D+cNJl9Um6
JYfyvkWIWxpPpF2Api6ol6dLSj5oaCOjFI7mJCOdSQDgOTagSMkfwYzJlocU67pb
8aQ0lgLoR5NJ8StRAzysY9EGP0ur7P9hv9IcdyASGD2SVY+2BKXEsR1Ruy5DvTiS
a547gfs2uLOwfOCE/NlelE49WHlg4xv8olowkMH5csqsVeDG6TKF/NebynKqtxac
tDGIt3CPreWtEYYrnU7ynAm1yUnLNfoY8N41XJIlB7BNTkYggQTpSV5UrJgjI/xy
ciLS7TGe2lGOZLYH6hp6zpr2rd0MdxTrMJEs1op0bLnxtxQFtXAjVFaGcstaOmPo
v6VIfUiO0wqqRT8JoP4WOHRsAeTXuNaiWiPXfc2q7pQHoVztDjBUk47wrBBHCzmG
RdnZ87NlTz7o3rrUn12UfKj7nA9OgYCwoWaNEDIIcaDUpsFpNniRtXmpIEOeitxz
OyhN8+OVjxVaJW7kYlQi/xyIyAvZ2MgLUwiGE4omZFF0q1aCDZxOtV35VnQnTrq0
1QvAcd0vQXxoCLYK1rFPJCKKTGyRVWTAIKDgnVykYYQkYltlsN42XCUKarpCmXs4
mrEZ7KkxbkV0h9tTrbs/oNf0JdmP5gUDzfWCFVuymE2wdOfaO50KvRLSi9B2wVWd
`pragma protect end_protected
