// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:36:46 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
i9hKlUc/4LevIox7MNckfJ0V1Hr5rjjQv7Vkwnpx6S9h+VRC+L2NM5+GUdknR+xm
w4/VeDULXHA8io/s7EDJWt4X7O1lEUCnIHxduMChO9TVIHPZVD3UveryluVE0mY3
GOAUqrcT9YXHFoLYjc0Xens2Myw3m2bJv5Wnyw7qLNI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 19616)
qA/620CoTJVjnWF0rTNY9DQUk/bEQ0EwkDNsoZX+OejG6GwtlSN4kfEtbYPV9lVa
JqLAfYWrLM8S2W+rALgzilqGAghj7a0UQGmnCudZbELMl2IWKGJKtdvl4zRhJGP8
qcb8EuwrLTCRbobBtb0gY12tSFT68WIq6ROzwKzuHHYRF2iLvrGqdrpec0q26Vx/
2aMOt/gQvRLZfA1PspTTtt8v8sprPRtxCdVH+B/aDsUVdfpuZqyDhV3TZ51GCCw6
FI1g4JQORfB93lbA/zVC2iCQsSknpbkubxl2camOqMacGCYXQw6FDeWOazv7GSU+
BVXXPD6HCw91NItK+Uu8ZxH6tXUGRFRKfatetbZwrTUOOGCvoQzwwfk93iRjoPUp
Tv6DlAiYwLXnNM5FwIon/CNHi1UkGvB5ZAsxDUQL71DNRDFMoxIfDnIuzeC1KVyY
lJ5oapjJEKWaODHEA59MeElj/BhIXJQK28dvIq9/YKSseRQCNvrfbgpeZuvEky+Y
q6bsrqu2NJoK3xMmKBn9dclWAVfpPikNGRXD9Fqs4ZIroarAt1/3UJvo6rM+TprO
ADfAsstkGoN97Z5cHimrm7v1j1VYYALwyRGdqapNJ6lxmkUF8DU59N9WgAQ2vFf4
aj2WwfuEEsDi71W0a9k3pLY6EfwAWcgl9GDLO7em9mksN26BguHoqLnRY73m+iJy
+IIFuLeulrwGJgBqMZ3w1fmXkOyOJcO2Y7eBr67FBgka9Z+/Dbq5SIUjX8VEPV/C
LOlH9fxPS3DctsP8AY/L3BHfNFJ/yy7iAperwYN680K7RyBBMTvSN1If63NQAu8Z
76qZX1e9Axjem9XUtW2rJQXpdJ4UHxh2V6eyMSZgPZRZhMRPSsCmtW0zpS/xkexv
O95y+59Ofhz1Ju2TadfcGO3GoO7djeouG16qJCCKiTR16WMIror1U3GPcE9Ucipg
aFk9XlM3e2zTeWnGzDIhZUu3Bh4GZ0VdcSJOUujCvJqZ0loAOgFKu8L6zUOiKnBH
18l+HAWPtH6Fox1BwN7T3IhiXLZi9NjTjTZ0xRkdH2u1fWTuzGq6mElTEsc8pnDo
NarJ/zejIf5lkWfqP53v6GPG+MnA0QvNry8GBjZixSypv7LDeY3ItToWvbt/yhWE
65obPa3hTd4LJK1rD/G83vf8iEdUXdv5yjbWZc/vuUqyJmYCCV4ac40lAP+Fwt36
1qTgiMWj5e0kyv2zBNsC45AoT/3aYZIB/uBkuqOF0uPcc0n0uqHCPDe8HBfyTt7j
07UoaYO+SORmwXpFwn0MD3SLR+tTUNbQvRrwiIMShSc0k/qcHN2VMamwO2rZzeWe
gDfi4rQldCEhkPIMQygyC9jDmkLOBQPth1FIvgJ+ci1ZhU2UWOnATIKYkMnyrOen
HumlZJWEpTWNO3UOkcoRvqKqvgnhViuYy0Jh4yVo+l9dZbSfAGoAmVqGg5dxIeIW
BR7CQdNJxdqLvft1F56m8SaXIQ/YMJjfSn834hdAUW2H3XJI6TIDVtGefHewrPAl
3YLR01gHzJdbQQUXvvFCwnvRQg0sWEc629u98376FA+SUxqzRwOOdHWgsJeb3PhI
8LBAUHpkihbM8O9EZCP/F4L7Bfen4w2n8naScNnkjgVcpl3J9jy/hrqBOGg323+T
bghZJ4F7idFiywjFRLjGfzxUjL3X20SsVSGB8RDCdKlrW21BldD3WPVcyjA4+hyw
S4SwzYX8Edyo2jrFLh/aGBwtNaTaXxwqxASqfPb+UbSK6iKLP9dNcGf0R9D+9u9p
3bhdD+gZfo+C7mbeqR4HSDPQgfDU6ZQ42hiiMsuicd+CU2xEEjElLMGGYPvc02tq
fNC5BGXExpH8k/3NaniirrUyPmk1KmnP+leU7mzlaQaziEKPPNLRtOYQeDl21FIb
TJ2cvoPA6FpkgI2Izo9BNKOQnUMZIlsU7hS6pKbowW3RvndV3UxIrAsXqpBN7wUV
0FOvkCQsyptrEbLAggTo4nRG0gxk1gzC4ONX8sVBXLjSrxvqtj1UTLkuxt1535hg
vNZn6eSJYhBjH56oupOGAikBCeR1c0qdnHdmukfqGHxlArGeJ8JK2kM2UE3Wcxzk
9VMKKzVcKPmdscRhLsVvC1hBH0z4h8ewNphKu1eJILhmlfL+9rKI/ewCwI4YJluZ
5kI8F4CwCqmFr01+p5Y60saugS2lvVwOQ3gD2+jZpSP/73uK24GlGNF1mmjdu+Lj
Z5JYplUjRMlZReM1xAMtYOXv4bZQVD5dZ0+YZG/gBxohTrUUJ+Evlsgn/2NGejia
KxER66CRhY+3XrJBymR4aRyM2nFE7vk7cqaVDSuwoEp3uSEN2OWCLi4pB+pKsfCc
cEOYOaYXkTonNo+G1/uHTxpjvUpMLTPCRmR9opoDA3GAII40A7S4zGXbcCLdPsWv
7RPcKxG2qK1bSKpCvlQy1PcFnZniEiscbS3cH2q67XhsWkRAB4pFZ6Vo4gruYmKX
0lk6QPv+Bd9TI1b6a24eAiH+XwZKHGrDJ5pKBchSPkFs5JM1FyS8ZWi/Z1Fq06r3
OGx6V72+fdXYXgnL6K/nUSr5FMsK3RgQ6BUGd+kQJ7U4+/SzYjORUdvDz37b2YYL
Q9Zt4M1h6UYOfwooQdbRYK6kgykVUPRYEiQVY2NfugZW9mdj9lVs7MM6E69G2bry
/IObW+5JWwnP4Irc6eLmOFG+zecwa4E6X9Clg9hhHKoGAywdgt5VFK8jSQ2VAyDQ
vQ029OYyJf1XpDLsMlnjjnk52W3N+5T0XAY00wqKtcSQKUO52qhQ0do3OHpL6VDk
IIUc9OsoD3NWwC4vljmLpPqbbOnuaM8XulsHtdc7qUuHzf8kANu/gybN9nRFeY5u
r4WZSgnA5ZY4RH6DHBp51RU4oF0ZV8LlzhI7E9xat+ssyL4hZtIO4eTqOPsMegDa
PmT4gQDWS78BH3iy6b8+/tPmNJoDEmt227sz2penCeDgi1r3WIUqowg+lwrb+aEV
upYS8UPI2ZSnmq3sOlZoHEvVO1SIyoy1ODwnsl9s2iBltkcup62XcxcdClBnharu
6uYK0vksyAzVLTHTx4ihgu3J/T3Y9QkC/40r6+sil/GKBuntGL+fH9g8gKk2J8M/
gCI8NecwarkHTjc6uPRFdNd8fOTpYUkNJISzExYdLZ/Mzx3kBE/bCpVUBbF14fUw
YgjoIGMa/DSzSA8vJ8+a7ogBDmDlukm56SjuOW/Av+PQL589Tj6MtM/48CPpD5/Y
U59na2u/Vhlci3GQ7r8bfZOxki8zzwcL8rxPOkdZSWfHfPPlpLSmPuIHvmuPyDyY
i2G8gQLg/y0u2Fxnj7BZ873Xvy1LiDVSVRcMPGi4A3/CQqtz13KuoyT8HCDxou/g
uRVM4AYTj/ePycMWJn7yQqGy7//UyV1X1JHfI34wbigl5SfMLe7Un+LaPKw27H21
+xQ0ynhuq6fA7rmXSEVXN6bD32LAeKdts8RS37SNSd7qee74sEuosYL54I0vVhMt
1h4pZrSzBkes5qGEJbFjNPEC0IVvrZRzGADYWE8LcVgsq8ANH61qjckg99rDVvdc
6JF/GIxwC5HJ2OnDeGzISEeVwRWF2TjKYIxWgiQMnnpXWlgbeArg/D1mm2dq9hry
ECd8WB2E+fapkJSCW77RItfXvfZzg6hb4ZEdam+XyigwFNVooNV315Tw/R7Qv4vP
S1wV3GpxDsbeJccyqyYSolJccTvY3UdX8kFW7oFUc15wQKuXm/yGxaxo80msfHW3
YwCJlbKdAXstrUWexZSsm3rmiZgnakzQ/s5u7Tw2Yf01WEWZi2g4RwBcSN9t9ccJ
5H4J3kBtdmOFP1sxJdKcftYmqDN155aEH1TV4S/YfnWOkbb+yJ9BPKmqUzthPCAC
91X4DlxylU3rglaOKbOjYY+U/d5zNFGNf5YzOgudhflRJFziBpO39WwJpBEbARe4
gNsod2Bo1nugDKN7ioe0689oo0I954e55o85HRNqYE3oD9wHh/LaPQz6vV56jCa4
isr6ig23WP2C/edGVTL+HPOKf/t8b4K+1ld3g29Wlos8Nuw4xZe87aBUCjjlYeZu
JkmT4O5vq+P5l5sN5MBQd80KIKxtNI38Syc+J2qqNwuh54gnTlnN1loowSvzy7bR
wn8ii/DNrih09ss2neQNC36XwKkObNKHZkcF6dhwd/VLn/RbNQZbltAVs6XMxAql
wMd3qicOXtGmvfBwTYghtvjvk3YM9YFToE248TYLb6as//rEQ/Zjo3JCkEkHq1IZ
pEIdbhrftkrIKX4Wf9Q+w+gD/AYCoRqo+EY0FQ4ctcYGGOU9g3yrPC0BGmBX5h0K
qC6Fv9KlOaVOzBNx04V7lwbXrbRKrnzgipa/zgGSc8YEOvKKeaLtHslY1qxSmLos
QF7uD1xPhmTyPcd6Qxi7ymCgWeoXvlJypimzRfPHRgTQmDPdpPkhHzZdNEXyAlR3
lZU15MUvWHOYpCIMzALkxaIEwR+edlG5gLq+RLTK0eogFtU5Qby4rkODrts1lswX
qSdQGMFilRUh+OAvhVyZSUJoi00GXes06Yzr3aRYio4Gk5enAZAxFAP5+EpJkHx6
s9ynsEs2s93MsnEHTXQn4Gxc2tP8GjpZWNov+kIetcXw1P8au3tQ4QVCAHZm5fuN
42LWVtqukTQ+KkpSZtoqXyar9JI+q57JUy6mMsLVJQ7/Y1beqXgEoRrbFzKRDzUY
5QM85ZBMJmO9D13IfYsTxCe01d5uFiD8UxmV2OA8IAP14VWJqrQXAhNwlbtVyf5N
+9nnmAP8I+BgukK6IqHl0IpAdBY7Dhjdt2pFmqY1I1TxCGvWYRibp652/Sqss6qT
4Hg8LfSczAZAA9MkAAZ74T3mQ6Psgbd1zPvX321R0irDeO6SUhCpPFu08xO4hJh7
J74CLXJfLKOJUCcvSlGOMcdMzf2IVMSJqF6Z+Q4nJ42FletYYb+hF6gfLkle2KkN
A6PK2B+6eCncnOl0E+MXBejEnpSTe0wWIJowa6HjQlOFV7TwRlmq1FxyXCVhaOrM
EU+cZntSUuCXZRSgQbfn5jem62PsOmGgswp6/yU2et8ndcPv0/GXT+iTP3fl3L0G
iXFjAyGEwnIzbUuLnIrZwmwWqSufDJlGEKR7fag0I+hBARTdKIut7mNqDk9G/cc+
KAHxBeQHoUKoJCXAYAhh9DqZ3NDmrDyzFiFDMfxLx9KmjC+K/QxnuITx05lOEwMZ
F+oCRgy9flGpnqFAeK9VisiH7OJloLfAWix16j6z7o/u7rwYlOvxY2+0jvY44KOU
TEKKOzx22cLvijFkLOBF4buvufPai4F5mAy+HyjPwcu6qZVyadcKzB+NDnfpR6Js
1zCRcQkQ0vJ4KKpFUvg5ZXTG+kkdp+PT1+bDFTJoo6/6zPfKSdx0XulNU8jTO479
ZXxGww8FVvn4DQe9VRiyHcFmdBRYbPRdkNEOc0aLUeAGTEZo7COJUYm4uQ5AYwkH
m049BnW+3yYDAhOYHpx7VWxxGJ2q+9ZJrXu4QxJz4EypH8GBNZbwSVc817yeF7OK
FbYTTzUuAC0fg3EYSDP/ZhVqowJKNBafBVKqytivhwpFI/XGFqNxslt3V+cri6uc
UPHOcQTe80/GhxgEqw+3HS86NpsrQ0hIpvhaVpC9f1J8Z0ZFjyyOLgvUgw5+Xp1u
UIQ4CWA3/f0gzG8g6vyH3PoK4/u9XAr54NsBqAW1oGFp9OfOAgshyQDtSYtZagGj
1lntfnPn5c/cFq5Dh9GFBqo7xDCggXHmVWb9LAi1zVVgiz8BNP3JLbnLCp5PLM1b
wJO+X9wzX9Zbcx5XlUqx994flcLNoEfac72bB5eV3blldHOSUjivT3w/Zea4mqjU
YCF1TnjNxXOOfJ2asr08F8KK4CCK88FK+TwF3ZfMvlo88/4bpKkRQ857iVR2kReO
iOG8iECOCHSYjmvjaTjeGjo8bjPFLaEorgW1vDUGWvUPNUqzDT+ZhzJHjnSi5Q8E
OVeqr3J5lXRd1w3UdEUuhPWmLkC3kMMPEKkAvzeVMztSMFmIMtCw4ikte1bcD68I
oO/fJr/LeSTvXmMCX5HEHJkWrEiTBzRgetd8rkc64D0vAkf5FSHuimHzV+hpRnoS
zHfpdQletlfN9rIFXs3xAsGQ7ir/OJYBlffnNX+GfWa9S3dd9TOu/Z/QIhquJRxq
rC+QUr6zVt8PBQx0IFY4cnC9wgRz9mOpZjV22Zrh5TMW++OamhMCYDl00h55pGD8
8CX1IG1Y8vtjNKSNCt2/JyFSlutcb52IESnq68wshLKhdQY04AvSw3b9IhxF9z9y
TWOgjRC/XbvQWfkKVdaiNLNxYlPUH0FxCd/IvXuDoQ6bjQePlEHS0oXemNi8vkMZ
D1dFjEcn8zGXujzg3uUVVBjX+G47F5bDmZzgS4DUIWV4g3Lta4mJqm0izCaqkEJJ
eTlz/xLZ/q5uEDLFus4GnlcZNTXwpVJBM4SnSse/fl1zoT8CV59uE2NGQ/pvh1VH
02RDREf3WJRBdvkOXoqTZBOGLAJhvwfpafPlPXeeKHuZDHeaZuFpgK9yfK0lajSo
W6TEq4xFV41U/SHUifSTcWHbh75VMxzR4S8yQDSzBLPt7QXM0zpUkJ7mqqg0O4Dg
Qlw8xnxpQ/X9O7UfC6sv/rhMl58J5hoJ4yAKQyJX3SxsMfcKFsIUvKQg3fuJpmZU
uaFVV1o6Kt72IerOTb5yq8hektCi077iyZBSlHB+T0QLagdIwIcuhgGDvfc+gHMJ
dEOYT4Qec4cuqbSPtarBd85lf8wR2np5kgJy9FzVn+DOU0YoAq21/oTkkeu5Rsn5
Y/IS7k/ZP2q82MizoV1opoqMqBO3yi448digwAJQze+lEQ66/yk0e3mfxor7jZ+6
UJLeJmBljesoM0tvJcce6qOTIF+orqUOR4HBvuNvNBTjH/nfemZKveoUIOp2TzzD
8MzO6Yh91mk0FCgsmPqBSE/389+HtZel8FjA7ijjpSTryAgslPr4e0sXuOU+4weu
oiKYNu3dFHgNBji+pkuqK6jczh8GAslyRTrdmKk7u41aRf62Efu1/EPBSxGinWq5
XEtGoYY9BfrXKBRPX2SfJMDn9zLsktnJygCDvsLAs1LpTQruP4j82lRXoqkJeE/W
+J8MixtWlckTP6Lr99dSdZCdaxcK4Huk2oWC2aXuFCPTQf0DRyxzT3QQFY1cQIzj
OwrGtZyvcT6CsWFxO9JZoEsU/WUpyrIDFVJC/P4JGIvpyOKBd+xVpcSvQJ4+DrL1
9etaDwmHgYMYMNh1HWk4v6ueAraYGU3n/efPdHjhGUbXlRKV0La2+8PbIau7RJ6f
zz64Kd4bJqsHEpV1L0G7Yls4XpNjFFr+6SGQpUNlAucvx/Za/1LfNY0z3ByIWrb7
H5XEHnUiEzBzRlm27+e06XM61SmyQX0Hb1y/5qoOjsvSF8RQOVUOFGr0gjGuMajA
XmF7g8nfHMQlivXzI8qOug7dUVtDVwS56dWsiCuCS/2qHu2jHyxOXKey5hbpdJ5U
FQWuBKyhGShb0lJY80gQQPXicKJDZ7PXa94aIY6MbHLIEoAITNdXCLgv3e4S8Dmm
LIAyh+Xr4Vwpvuz6IYUEzj1qHD6/Q27c7eQfquMYq0ucnDOBg4WRogb8ocwrfi5D
DOI/UFquqiXFXd54kt8NFmSUje4TT44PCda9Z7mBVbOZJXnRPe3XSbWM4xydDZHO
GjAr+cvAlGLfOxdAUTiyiV68nif/LO9NXKEwFCi/yJcjm8BFv6dOLuJ2EIQzXzAf
8KgDsA3QIAs+Jrfy72vN5yLk4gKuqyQOfx1HXONMIWUpgW1a5Jo+5DGHnaV+E5dg
zr46EwONlROx7rMDkWUtNhCwEi5OAQlWn14tz8cTnrFvin++3k+s1L4CKTN0aw0Z
6yvsYMosQnLUI1fzhZgpWr7bTPg1M3qEfE2sbPiOHZYcj7L6W8ydwOf0e020CIYc
xZwjXHzdC5/yzShIzTduYBiIT91KxzI7bfxOSXEJGtehiajuWNAyAtI4mhZorJBP
sTNIaj8V1syvXwZwtJheRi4KYTwKd0+6wv9u5n4QWy5BhW/FqWlwzx60jgs1xRZ4
8HUP9KWS3enlCW/FSw9Afa9xTafNmDwE/ojueNmrd47wcFiKr6zHYRd29tb0+q0C
872YpG+pmRCF0Fc3aPuTybKYyIyXFWWNAn3GOonqW3NZUJT+nnSNXeJeLUWO6fXN
BMruepQZdQ+KKVOQc0LD4feeXWRKTw8uwhIGpbnM2qelwKOp28yjepFjR2KVnk2v
SRszDbZvEuckSdcVYOpVraiWhPWNixK2ptLA6FOeP/6XwPMKwKNhnHRLNBF3GNST
ecVoAsDwAdzgwvpbaV1zPMax8lai7f+foz58qCgOTBIPEOx92GMQaT00lXbK3OS3
5v+I7ngAKw1gJxifg5xN2yr1fWfyffLLu5Ll+rjlbn/A1S2nSvBhN3MQVgVo+2Mk
LTgDI6Q/n57NpidQTGmVxX+bKiiDMIbbNyq8yzHILORbUNfWcFu0NOAvWLzPQot2
5xHDdsAJDMt9yG5HUowJ3sZLs+oswyGkWeohhkudjvrUcMKlmXineKAn+bcf9e6C
Dr+lkj2a0GVANCAJjzxF7YYg0EiZRB19e0Zyoai0c+PxsLNhP7KhWPEKxur0Cjz0
gQ/Yt5jdIrgOBbKdt50QdwKVUnrQuWM0punzMJDkOomsV+JsgieoiAHTs3t5VeQu
tcE/3omrOLVKsz5YHAzV6Sb5FOgDJcRHOHOFP/P9wGDCWYGZDS6ijHq24reX0qwB
w+9eI1rTqQu3KoFH16h9F4TDqLBnAMPh6ohswDfOXMw71umAVexpV0IL2XxCbzgC
P8OVy7XhRiz8fkuL680FopHDowEctXjRfDOM/OPAERWPFEsYGZXoho6kVS9nv5Jd
a22jSJ64X7HtAVzWVF4Du1wT4BWkmaTrb2lyOKWa86RDD8g61aDGz0Z5HkabrFTr
HxRBP6eaBRloZACpYH9h/clGicZ1Q928JOZG2ZxBQG9HtxJ/pAH3C6o11ww9vShJ
eqTOOj9nlrwvehE4FH5MXFFALQYRph0MVL3s74xNWE1a3HXCO4adxZFfFhRFFWwl
bRfOCPh732dxjk3hn0BMD+LIKNEJheBxzE31lDgTUkHMBCgHu0M+zt9OtOrGSQpe
DaXw9UI4dUKHgV14RwCHWEjkz8F7fuyoUcbAcJWkntiGf9nWrcXMK7aGaIy1cTxF
ivn8nmGra6iqEELUfaZmXoFeQbdp/V4/AHHqZTpYOGcy+qsIorUIQNCZBjO0l353
aMzRmpzCPV9jxbRpw6jqD99cD5jv5u76vgH69o4hML7gn/Q4sANZPyD85/5xlRLk
AeaCI4cIWYG3TQkE1IlPn9hDxD8HdnY106GI0sxvuzCIAi1CO+4doSyuOoS/WCgz
KPHhYZt0JhnTUyYJ/7H9twzcsRLfpk5Pjq55pQj89Tz54W+Md9tOk4PGxW7LvRxY
+1Fo8aiTa/Ic40XQ54CY8fRJUvcHFPKN2r+FAmhHKqbAfr0hwrSYswHM0ufSiGSC
109N40KeziaqpxVnSOgOrpR7S4syjdA8C0xWK+/mZWsF7L0sRIYWaXVrsNNsjNkw
JpRR87EwKEGpKyPqIzXNCcshuSIU8Cvorc3ZHgPcdAfp1B0Yk2K2IlPIWDgVt4lZ
PrYNrk8GciJeA1Z06y1JUxY8MFqtB6osHach11EM0jMvvq57sddClxCOsdNERpZA
+g1+c9dPWB5rrNx96gnC/rmZ1+V4bfNrrd8Ym3xF2Tqj/AO7aYeHUh1UrkbSgvyW
wa4t10XyHPoLQ8Vx5esFehD9wMgyUBZLdiB8exYqJlh+EJ6MTsVZm1ZgAB1O0Fr8
Wg+9kD8QiVlDN7MLjdgkw/21iI4ugPOz8bDhdXe1Hef1s2p8xO9xmh3ABXdpXS4N
4ZohhuLIzHX8BbrbkGSc9ZkLzVfU4p6aYbrWYEQ3LURXusBP3/EI1ScQBh7Wc0u/
F1nONg+sA5Sbz2aNeXIX/g3bINzPBQo36wPx2bCFxT+mxqkvwVd506hHGl68Tdio
NBzrrYQb51pVrJ/+34eE/O/3TbFPLCzBNyapEjGoOylDOPs8p6oGThvd54cAUZRj
BfuWOMjhzyStPRW9/2daSu+NR03XE2sNj04nkmwGdE3x4EIMxfTcf6DWScVV2LQv
xSx0gV0TyVMGXSCvMeIxIn4iD+PdOUvzIar/KCq2dIdUXCtWt2StACZ4yFMc/j9U
iR33M4AVmHMhxkkXiJrXR3A9hUQ1swYvI43XHkj6w2X2d1rbZaZ6cfhtju6HVoP/
8iE7KuKmILBkqHc1ynL7l7uzv+hYdsB/+8P1mGwLDooUvxmi1s3BvzFK6+b+wLhI
uiu1vmJEzWYSruFSUzDRcswn+HyfON5MeRV2oCfQPTjKNVF2Nt9UgMCnyHA9iTsp
4APY0NrrLF2RkSFZVdwC0HqZRrpnIA4InJIJiksF8Pmg0m7MotD7tjidt/MoQC1+
k5498niB3i9botH6XFLvLuLzz9eTOJFNlGgjYT2qQ7OTYdga4k0KZAWqSiDepImG
u6fb+vkQzUfxfRLEgKS21j6uwvcbROWa+jGCTz1Z4k4SaW2kdFNNHr7vQFIqYaYR
woQseq4JAc5xPTnAWyBfJD1GbqVBGErFf9ZYijfxw3JNZvccgmZN1rkwpCgO3Hf/
PUP+sOAtgqMV4S+Sz3gQDiYRqx25eaLtYvKlZ5NxMyPiOSh+bbeBF0OaQUiEYmMB
pFCOy1ByfVWDdlEuE9X6+T0icBUlksxkr9SB7TIX9lU7zCL6cXs6v7hCBMDvrYd7
RgGVGCUlt0YxPHY7XpW0b2Ovv/LKE93Jqqq1TGTG8IGS2hlrzcjc6Hn1uxTCab5w
ZOoYwJz5K+NA09lpgJWwdhK0dEmbs/FF6CLVKMv3EEYkwZvXktp2oCSVtso6KEy0
9gtk0WbGr7jZo8T2GQKu1jDj8ImzhlAKyiwUm21vfe7Phkay6o9o6LrK/th1OPmx
yDyDY8dLshRzJJZKGk4iQXu8rn5A0/TTnglMLRBDJqwmFse9YyFOrJfC2ofHYSpk
vCIu5VhSTvGyZTu3QeK6kHHXD5VHo/wA5jvv0D3RjeiUDZ9+FJzwvoRdsNQYkE1N
SEdtGCh+Ot4sA1HQSnKVDS/OK0357X+1BXxNWKf1Q5EjxqHBofSySS/8AZBj5m9m
gjD696fw9kZYBfxrGTYolZWjAv4wpAGhQEulrUWHOB2tGD3sz/plVXATiD7+RuDn
8s0Mt7sZJM1Vp8c+X0Fpv2K0BjPJK77NNOrKF4oCkgjGlkl+3jaVPuJe5l/e5fkR
Mav+YpphUZDXP8foyWlTRn3THMtHJQZocqRNkquAYajPuL/wFLql5lR+yXXL3abm
aDGTAtYveRZXcAfB5PQ3Agrr0zwmCIq8QitQMOsk0k0mPQADpFe5N8wq0OtwOffU
TukFRhwKms9fPCpdxAxsvmvXJe1pw2BdBtp9J5CL9aU1DZbKlgA2fzgNqiemdnSe
LYqNmig1Timn54Hmz/cIuly5MNvhXqC0RSPb2OWoPSeT2+0LBcOtKK81SmvbHbJA
Lno1BGEx7kIy1QqySgTszvVCHmoBTjejyOB0VrcHoAgedEgG2Z7jGI/aNh+uVRmM
qhFzPyOCkjNI0P02Gy2V/NdGYCnmPPsbnWDtDq93iH1zR3dqRIARLdzAqAeqU0D5
Hm0G+9hFtc/qMbD3oEvoPxCayB1Cc023soZBth09MmgDNs0nSFDIS7yy57HcO13x
DL8BY9QNf6kpf5LdhbH2PexFWuTZTR+zx1EfvwX0DsiWrT0qC64spj4Y7B4JuKc4
IFBpebvQjRvWvGtFiInlElhVRXfxmjuYoODpOO5B01d6kwI9J1L++T6jm532gbkL
Nf/32Q51LvneViNLNXeS1njkKw/bTI6Pgsg8K8sSzdg00Z3eKG1FzGw9eXZUKSkY
4bECAAh7RUIIFflBtBfZs+jngqte/kQxRobzfGrSWi1WsJuGckLSlA9K74vW6Qre
OQQ2qPX6kMnymRPQGyTX6E/VU/H1pnX5cBQfZHryo4rBNR0MOVqubDDj+KzvDTjd
C7XBsvHV1w7RuzySy/N1r2bCjy/euBKGPKBdP8bCFLgBRu5u/XNfrP6JRVELYpoY
AXPBD90oGCHUYwU6ZUiQTuVHEA6IS2De89lo1AdxJ8qacg8Vl/Xwn1KU/4+YQDEz
ZdedSQ6LxhYLHeMf/IlmWZrjIitBU4/fqo9B5idE3UnRwy7FBZiQ6yqI7ztGD7yO
YXY2+VHSO77zvC+2mL3tT2BmGUUZJnRiy6vko0UUA9IoIhBQnrLvZCZyNCEfGlXJ
8cPodkrlyRLlL/oxppaI5E1OuthUuk/3d83vyaqyz4f1elbAfqElE8BtRa7wUzFw
y14zWhr6hVPuHHTdgFBDNSSqUDoLb8gRx24XivaJIZ/UJKC8/TMMlN9bB8C+DIAi
TJn1GsGorTR6HZTVzUStFXZ6/pzU4J38F9JYhxd00uBcpHcT/afh+40DTtFzRBVW
JyoUPcS0OJrMU2Zh7zKdIOHRFuNvqU/+8oQzmfCZ9OxtPX5SapT4UGEo8uoAwrE0
v6cvmivt+eUHY9kYJBOmmbhtR37GoI05R690LwZ/T/DUsAFxxHAUJYLu+C/kmK9A
QGWaYPl7TTqqC3EqPmy+d5wE0wMdM2tK4ioLmQOTrL3xhN4VZXE/eHCOzaWHUsKp
dAt6uSbiVgPlgbOpCFPlgm0YLOz/OJ6Vz+GS0K3vldzGqLfeUqs2711Y1MJ4mTzX
DXIoTfzm/182/VAzUoWhDD2BUw9uOtfO4gc+Xmhk3cIc9Qn42eTJr23ixU10uzUp
JWNApBsE3FCYu2jBMFnLHQBGqT8JOrtLSiqfVsH0BIet8oiXGtkn97W8oHhM3OG/
25A3cFu2Rj7rxwfCVfFC+ZNk+VRsk+VCvTImjndtHJDPrbxCH+K+prheqW1WR/V0
7gXlLiUlxP6KWVsuMqe7gEDUarh3lJA6If2VcKXWyhmZyWyXKDX38zFaPTy9Ovoq
GzLebkzuf4xhA8rkFQVvCUIOqC4YBoyng50ZLfvmWJwayqYdP/xb479M4AJMQU0N
2D4QZkRXa/61TVq/XtXC29HCMfSwhcdcUB7/95CZk0H3j0K7eKZLRiGKmk/4R9Rv
FToxMItudEqmVMFvMJOwSfzvXQZ1oyxDT+YREqhuxjuQDod3OfGakzin9sktCqoG
Z+j+JW3HCGJKb1NS6sVASwNHEam1xgXUXaIrOB6Q/PazZ361PD2DvF/RkX7kCX2i
8FzgQ9uiMhdxyioECGoW8sz/c5lwqW6Ig+Q7ALopLG6xYeoW6huPqub0aLebCZzu
XrZB8rD3PCvMKR6xRb7s8i6dxiDsUld5y3qu548q3wDvJQ2eqO8vVHWU75v2G3fP
D+g8WhIBcL3fbUzdl3TlSgszO6EtanKb8HpfBJlKYz22NCm89e5tNa3Ni9Ss8ccL
6VqSGCcYVYhbOw71mlSh10sLKs+m+FE4icp+Fd8yoN6Y2ch+vrogtNPbSMZCyGgf
Mr0NGoLkELPdthvO+hNteHBtgDGEtDjJufYR6LHzik5EJnW2dhbU7vsvaQP5SSle
D09fTCRZFEkuMl8G3Vpy1YrsB0vFthBFqyqmXU1ST+cO12XNyr4kK4A/BMZgvzdB
aqSeOn5vSA9evp7krOUkcYhuMUHOlgT6WgVDcFWXFf1H5J9sMyFyUeCXHLcKEQ5f
L1NwJN6xlNTSUbygLBMbaJKRqDy5l1AlYaiRuet9l14eKr3Kf41lVB/niZkSxohv
vhkoHrEl8+fbCrLkvVSTxzryV39wY88djqH6mrrULuijUOUPVTXTd+Tr9x96qneg
JJtu0wUSBdsClEpeDgGbXMK0iM5QOnnSa9lUuCZ4xC1d83O7P74Iiylmr40Uv8uB
2h+Wm258b41+01gNpq6I6Q8JJ99omeaaCyoTUT7a4xpnGs8mT/Ud5UFUSoKfmTZq
n4tkFCGLOyGKAff/ify75G6hKGUqz7JDu6ENxgfAMX4pgPSf9P7HXe+9hOIifu/g
/5fCkRhXZus8IWacU5FNtrFeZu4klsvq752V6InGHoCoXSbX2JIv+hGxmJnUZshV
4bnPjLR1T4GPlGRBh0cvfjOZ51b7YBZ/G2krohIlE4viIzoGA7Wy334QsPNWF9Zu
fxW6iYDExnKxT+rm30f9tJXWHk291dP64hs/DVbkpe5eZq1F91IfmT6gHgCZJe8E
dR+zz/VNhyo+WXpR5AMqTF7gYA2PGzMPsEQVXkKqOqG8icqKpuay+8SoTDglNAXI
akGe+eYcoarWSNan2GivZz0vDdVUzT7LCUvMXdPwVnlas92ABJ65bqzI2PDOuMoi
LeRjlxd5fdP6KPSCsw/Z/YJCnVeyOeWXBlTNYmTD0vAMTT5qL9cDgqxt9WFYsyF0
UCwzOZrfWb833feMfrn6sMBubkVKlAn2qUknDQPFGhoXlg19l87NZRwABftwSctX
Gz38BqPpJeeefbm8/F2I5vTiX+8RfEDnrnq4RBkMp71i6GqJiy37MtcseqFm/9ez
E526xi8oOVxJo4+X1qUge+7hGSp9DTPe3V7FFoEcSe3F5MEjXb74mRmWqUNRycTz
sJWY7wC65BGVuRRcMisXmKsgx7aTF35y6OJtrLnuunhiqyFYMvIdqM8ecX79kJvv
YECWxax/EYJCfA8hefsapkhUg809g++F9Jg0ztdW34zSDijT3g2a8KodXrPcHQNL
xrG5DzIgZsujsOXDzOmZrGGDOAVXvUaOqLXiVTNfiYYBEtmkmqTJl2IeHsgGAjuI
dNmob6VRk1m4eKr6zrZt8YiUXmneiMyAPbLmrtOZX7LQb9Hy/YlAtx+nrzaCXnQu
KD0OLQnoWCOTauaKGSv+MMK1l789gfgzRNXQJzjQaMylQGiD+r5n1C08RN0E4t6V
1eJLScUfUeYqisBaD62RlDVZbwLC514N2hJ/PJpU9BtTVssmRb4LaP38r1VxOZ/X
8T42yygwp3pxW+E5+BbfobO+J4FYHdAG5eGMgsBi+Ys3vlTncDHMnM9qajS313qi
burxLK3A8TCuaGZoW38Nd7h1d/enU4FhZaOdBPmoAwcxmurBKyEbd+15Xtj3x7HV
O3QXYouecPhouzXA4NjJ5xpd9tnsPX+vkgeZD9Uu4j/Yt/znwlyHhEFAtory6bEz
uXcWZp5ESvaIWXDE6B0MCL8oIHlMywWborG4zbm/+ZpeMHZv6ZScNJF7/ONB4X3U
OqoVS66Ydp7KmNSxzrjWXbeb1ozuHwUFT9UCnTKgeDf0CS5kdSoKatvsg3XBSvd6
H3Hpu/pKTZ8s2Olg5/jdBg7YKy1EPJQQ8rS/aWZy4BZttFiP6rQioDHJi+zQJNmc
jVub2FP8XZg+Ypv0gQ9gxlgi/1aEY4OBsXakLUmy99AH54q/NsmknFP2ErtXZQpQ
WIYmVNhuxUHRvyU5ATmouwv0eJb/leFkP5Ve2riV1SE59howc8o9lp3gXVby70Wx
R9Tgm/2Esub/jSmwwYWgAiK74BVdsGQ7/pOpYExR8VSN+FnPJL3NSNPZRave1/4O
tSxbVWsOQ+0jykNpj/UVmSzBiMmQuO8ZigNsHsXpfhqkRSsTwyF4d5CUF4qFRa0V
UQRclGUQ7dJzdju+B785O5QIFVR5XB2BpUnZ6E2GdsD42nKTgYcH2NyS00wZGyGv
pYr7GS57wWMJRc9617Xq6MLY1GF7s4F0kOcmJl2Y1xF9I1/nJLG7tsU8IG01BQiO
GwR1Y9IKlV8+SjgWc/rntxGRmGo+lodsHypXnfCk4JxQolaWdiQU3Rq2JoELBf5A
DCs/e4n4zU47ZUbwamIfdfWccP0/Vg8KB+MBzGhAHaJ5QeZrz1gQKPsfimjTSBZW
4KjCd+hFqDTXmiZXazDqmi+U6hGE1s5EzxfcxWBBpanrBVCyYw1Zneq/ppKlbyUU
ptUWO36gy1wXICjxgGAEYypqYymE1s3/VtXaOq52d+zfI/LkjTS+/bwBboj7OVPY
l18Z3mclAIp3jhPedMWyA4RVEyPoHWiHNkJBzB7x+yYrVzv5VCLroNfGOo9La++e
5nVGxHj3PemWBiPRyq6MSeCf0h1yrosHCZJg/RqOoQ0od8HOg5eAlrU7SIudV14g
9+oWgXQGvlrmUnhDJyjSPb87svqR1rFfuw99ZisXNYmDB78oW/+ydiqsGXK3WPVK
DceSiE+vtv61oPWqCVB2QoGoaWcU2xYo4qABvuAFyQjsgcqdnVbsJe5Ms5K/x+g2
jDas4rga3mQkGfmxnF/YwDBp+RD4Y7rHDJjdOb3DPaqxn74+nP5zE1XcZ/Ibho+6
IrM8NGRG14/CU6Yu8zTQ8QpnCqrUI5jTVS/7syk4KaxAf9/4hNexzU4nZ7aqT5b+
kJHGFpNC5z8LklbBQWeQZmX2UQEMWlJvre18vto2fQhkLG3BmzBGOJWaXIRonDaW
v3QZH4Ay7qCAUg5+bGHHAE0G76LdRM4ziWx5KSMMHACEgxE81Ce2+U6KQyjXd/Kh
AoPQzB/3UClqOclqYTNazNvloMpRjRFqWZiYcVSXsN1zcfyaScej9J/I1xH2QXnG
mS1WzVT/w8erZ94e5TQIqA9LylBB65tnmYI1dbWpT1h3FQXs2QUmklfabTuSgo5P
8ArnGTF/kH1B5HG8kV7gJEHeCLp6VzbOu5sdE72/LaELQVUdGiKg2GH26NqhhYZ+
Lft0QQZu7dkd3jKk8nlrMy7IWlc29CoVH9NyJjQ8Ai2xKxMpESwWcmES2x3NVb/R
OU0Ue6vP0tBoWqRJPNNXik8XC52hxcfzLcZCF/pB67H3HC1Ye7WM/szh1cElx3X7
XsEvUZo3449TT9vpgEsD72RqC114GEGO3ZD7BCJZ315jNC6Sy9kJpHLyYrjyecCp
tCP3S8tPJhwO8SPmMIBhlghFl6TVrXOohX8F2Ji/0GNj9EpF4LYl8cJ2FrCqsulW
XFULPMf+RO0Tdw4fBgTfZkQKbFPQhyCD4ksVb1po9v6sM28xi1aeBh0d+1Oi4+vx
K5cyhtlR7ru+v9R1IzkMJK/cELCABO/bC63vU/iupDUsNIcOmSN6qFOksHcNj0j3
dj7dBSwXOWdSGxLH1YDuHTz4CoQUyPh2gGYGct0eGVL3Hl4ObtHjlpT2tHbAeBGK
SAPosmuHgkYRPh4JYb/6868wO9w3HqPr9htfrZzrG4kCK6d5+lDPnQDPyArb7u8g
j939SflLw36yCydU62d5gblcTELGi7eMovP3Fas7bcoOk0fUBL0HpiEczuJcb0pE
9TR766jc87xEUqBQnqtFTZoJoTFW7ITfTmM/PU8/j0Dz16Rn3mSrCRyrWfx4Qqp6
CBI2A0hAMEkCoZuMfYustMTckJE2Yp4qKWcX4nZpOzS6e57on7NG2c/INYkU6LRc
wb9usdQzJMX/ZOVAoVvK2+4DfNycmk/ncleU6bYQkaYf+YWbxtRe7NKpcy52ZtHh
dVgNLGfwalreqdNI2wN5znIs6IfeDKgVTlB5yiuCQWFUcr3n1dCr1TbRtl+UQHA6
bwtUh1p4mr6Zd3itbY1BKQVNIw10Y7ntnvfXmdoJNkkvgV3jpGVebZqSs17n+XKB
LM44PUZiWHlfyQ7Ob3XcfvkvnAFP78A/h4vbQ0LoRxdqxQOi1YU4zPpNyQE6VDCU
nWe6doGXTm+YxCOFK7G4pkiYebdksjqn4cJDlIyIBE8+n/JIbiLoLAtiPlstvPp4
OOtwjCw1zEepsBTtFQWyFSOP6xJpZXfZfsWYKJesU+3I1wFi72BKiulq/B6+N7m/
LBX4qdgqO+W1cAkMoK1vUQT8SgJhJnoo4dZBMDEKJYByHtrMoixPsnEfihqM/Yyq
ZuOUc5N9n01WRZJi/QVNLj4tIGrJeQO2Tl76lsHAgTV09jQ09uoZcY5L6OJZnLRa
MTzf1xJ70D3ZJ1ld4a2I5OEnyZ7gLsnCHx7LfXllqmTI8DFurul8m0QqJTjo0AH6
omOPnaXHaU7gKjcz5MZISsxMqqfJdKL9j/mFbBtv41P1WkTTpsSWVAF4VBRjZXwA
F7bV+JQwqlKff/5xwkCrlEkCkiL6qDsal03SQNgPCKLFLdaBgFk6Jt/4jodsoEU5
TKd0eaeZUP1IwoZ/OAH+qU0q/z7FgG+seIOR6O3ViKSlFdTiPY+C/Ko2pBDQDuYI
AelHGyABl7FVLyIl6CAmXFFJsdlPCIzWg00nMJj98SIjzRB7mtqWzxPCdMNc+cg3
4DBxAzekbisgCMjdMrA4B6zTauNTUtxJAOVjiWNE8RwztYeGYiegJd7BA3rzOKUT
5VAcvzAXADfAAS4YLx+9tEAccocmMzKBSMF1FqgmAFZDrXl1OcMLrKhOeBnRpFaD
y67DJzOOMiCXwN14vb1gJHIx6UXs/YYtkbQDm/o8KouCEOVMbO/w3Axgv/4QhWmT
xSiTZaFksauE+mg0rZoe8mpb3tx6Re0JCSGtaIOmOGqstdhgsYedrMebDRHDoZD0
QZcu3io4jV7VfnKVtn0n4N0HlPSCDoZYVvFGHhGqswEnImEM9kH3EWbE1QdY1cYn
nxhk+wNhHX5YhnbVWtz20AbfxKb66kp0KFT/Y4IXfesuGreduBpNhK8vlhhUX8nb
hpsHqK2oAMCOBHWA/QMfuuBUgCcV26ZTQmpddySIyjBD5rfQp2AiQqwZGQ937uLw
KmwQShtEJbAquJpCRKExHdPf25uZk4RUxgRGvr2s14xHZYzEvJIyvzSY6jGbRBkr
+EGM/tpZXUvFK5fCVSWGZbBoP6ZW+ah/H4B78oXA6p69qbGz5bcyQo/Vc24C3Jqh
/N6AhWz4mRn0v/UTGjhe8+/avxnfNfY6uz8diIp9WptCPru1M3/R8MYZbFKgN2js
Op6ZSlHeKcjMwOK9givSugazmeQJGGottc4NAdr8OSpLjxhZSkQjqVy2QDbfaxMT
zoPuOYXaL1j978TxCSqY+7JPVumBozydj4GFtMwkNjROxkTMfHizW6xPx1SJkjz8
0E6KSz+EldUmtLR+gfsGS6ondEgsrxoJcMHIPvH5yyPoNSNTBHuIQlP/YXfKXisU
XYdPMebpotz4o1uMbvcandvJgeDZBiLncydq1kJGBOFaufN7q2GH24NlpPhyGAeR
pMABfEh85MwEq9b9QCEl5sIudByq8cC+g4AQm06xHv65u11vYCHzPBmK3CSUotrm
yALOGhA4f7q7UcyaocI8se5u4BFt+Qbqa0sf/MA2eCvWl5dwfofrtv1Fzi+8644a
FnO47eTow+y6Xyp5UblgcroM29M/NDL8+UWVdyXS5nhjzrUnNDBIPkXmH71Bi+zV
OeJ1jLjxlGXO1bcCH4vu2dBONgAycO7yQSCl6uwwWGPRLN7o1pFaHE1rDww6xWOQ
t//UcWGiyRv/9LL9lPP1qvSEH43bdaOq99/31jezoSClrI8odhVLdR7bnp2+Q+71
J+BhhgIFLl9ceMxjvYr4OSVO1qr48yYNnruJTa2z1vxILKNQOtp7Lh6Z3ClSSwpA
R3f4LCITOJNj3VIGdmPmfkz+6qc70wnny5ghkg6/WRbaV6oaNK8l+quePuDdIyCJ
aUJmT3kqdT9rY/BUD9cvUA0AUr/hj4qs1fC5a+DTgNYcZ9c0TtZwabKrF6jufDXj
bl0LXAUgaic1YNPl3OCgwFb1ipN2uMNT93Kf9lnDiGlqrEsx0UHR5T66i5FxeM1r
ZK/tw+DXyxjEE1NxSPKyYa/CtN92+tm5CuA5MDAOwuZsFgg6n7l9Z/tH9GNZt7Ev
C2bzWM8Fu8+KfYMXr3M/SYbu3Gz8QBo/i1xdkRAmCqSy3Y733PuXPSAj4fx7WYLz
+gfG53bJlueVqT/3Az5HA3Kf/bnQPWFIcvYKobLEtMIi9ebwE3ylBBf7BLTi4qsg
o6S+8UosGL1uMIPYWam1MeV/pkocVYWCbnqISKrgMrn5+73eQQoyNhKTZRARPTJc
7tPqrpld4cfILb/OF09au0/S+tTcVp4Qj2ITRE3195PCS1O+sz6RsV+QoWaUxJzO
f9WDql37GUUoRD04260gjIPcUe0lYQtYbZUrO8Cz47ld1zKlX53p6KAPzYyET0s7
V8n0+jAgRgIL5C+fe6gIj/a/KnXSeS5wBHAOM7F1w0zUxyK37/M38YbWWWz0/xVA
Z6YPmdW+7VBWH/zd3AyMiesNqsl2j56MUReqad+qkH39Kx6evRcEmGDqGAndbpW6
Kp6PMDg2KZYwbKcTuDKzAqA8Q5tnI28No1YT5/iuWO7VPNMiq3h6whEjTF87VzdA
kNsZnGEUP9sM4B6Z5406175cLISfGhDuOVDT1UbH7GRcC0ptXRSsR/fV66ZcnRlT
1AhHdev9rFlygw/+WvLgUJ9f6jFQQHCUL5t0sN4oPDu6v0eGt64V2JjlsO1UBUhD
WGOxZrxP8jvADMTwt4mVk2klnlpJPc0edbxItqicJjby+eparBH0Bc7OwOgcya4F
AeNmWTvIth0FsX6/zQmzeOzvydWDUl4ihcu4tJ679D3VJa1ERnW8a6JuCX2jqsmk
TP2rYjnYqNjKmZVtzCkJsw7s7ZmqlMeP8j0NJzMpXC8FDsCI71ZOe3vTW166/BIh
xj7npKdvCZwtKYTvvFoWph7ILwNLu1UstG3EM5sQvzj5U8aT3KwNnWlOLPWsjoz6
qeSYR0vwbBetZeYzrhzoYSoNDTWlczkGOE9C3ExGBVPLvJF9QS/tH7UhWnT64gQ2
sk/Ze0LNOKWDe4qqRmqph9wntD92aH8ZnfISndKX6qE+LIBxR34i7tAWTocl9Ziv
7OlhSGLXGMws1PYUAAj0U5+fJFAp3nTD1gPgalOMgdyGoN7jwxj9b3/6B/oHE1xT
73ByNe9WmZKnlp5r9bw6twdiAGU+g5pWekEY5LfKzYrWTK62ocTXMhMN704x3fM5
qlxE5qdZwVqwQ63nwRZ3trBNLPO7ZxSXhkNiVfKFLHslhsRrob09QDIKRpRjdiq2
TxpSLx7f+mXZ5EAK0KmhhpalOMab9rKtwjD8h/yPpehoix7GdBDq8qFMAUEuLUpY
GpWxNwtpFJNC6E04G584ingKjjk3G6OzcUBSxtK9doCwwaH2qN2Xsk/4Ntla3lzf
IIs4EQh2N/DUGITCy7NrqUuoakuIdd3a2XLcaXtjjUmElSs4bnkmAtwcZEeGdlZY
BW/VPHWuqNQQ7ogJZcokytu7KGs1QhO6xTYerSe+ebfoOL8Q00Vmu1HPJVgIWo7G
cbPZV4Ni+0J/aVlbprePvODiAEayWDtJuqn4zmpnqaDkQpvehKgPvI24PMhKMAwD
cgceOL61TwLWIGgiXHdjXEdgMEH/Q0FNgzDaJoTwri/qTo2EMWeDgJDfo66ugj09
L/7qRM9gip1RrAzZqn6vYDSJLrKrL80Lqt6fnm5kd2yrH5GpgaZBcQRGkcIdEYxM
mWwFutRZZ82+4CNpBkxx/uTemeuki9mTtZXnmAc5yYpSDLOcXlrx9xHbxNhbUXnS
IMb+o/QP2Ow3DARbU191WFY9RT4YhQbhqJrBJSaLHSJNf1RqvVr6Kf24uV5z122H
s/CEuyVmkaM8RzsQ50rq73SU9V9//UBRqicSVtzVX7zoaPacAY15/YWHmCcZL20f
2irXIE7UKjeVI00YN0Tk5u+tri+ExnMFc5js5OUBEvfd4CvaeENyYqhK/4sbC43Y
r4cdd/8EAJEArGwFfzPbLovZDDDB3n3K0Lr3ezoIEL5IYCDv6B6U4zjAnqrk5I9t
7AEzZQbXVHpvO9KW2xB5g42gvxZwDoUrmj5id2LDkUxhPvZWAYiJgwaVDYmVmo64
1Ye0iv2CQ7qBVaHwKFbGr3umpNmm3XvFuazBfhbFm3Qy5hSwhuywo9Epsz9fN6+D
eVZAabt2He46+JtlU8mSVWv/OINttfgKKxdCyZcOLZZlWBWqoAF9RD6+ODIBRgd2
ttxNaK3QuDnPgQVtlfbsInq55/Magq4kT2DKnNXOU3hBjlM0yTvzbq5AXyveX8uH
gFe0p8849IMtOeiHOMaMvgIdR1rsGsfIYVggJWu81o+oZwddwyGOCiSo8E+xa7Rx
TgiuuhlSWUMNmTW1K4SCwBgXmAyFSxTZNfCOEGE2s9NfIe1G7VosVT+VG/xb4kzA
31wmMH14mkG1AGtZgkD8jsYLF1S6KqmUehOxRUp9Zn5ryezAQQ0KRbdDcqR/8hkb
kyJ5UZ2Z6yz+hI703SCVBFy3bwt8vzhPpm/nQ6DpZAIkIQAP0ELMVo1X2cPhY6va
NHKCJUTIEz9fADttcdNVOHh7o9x2VUWuPg0BnQhWOI/ef6TX0WH5Rs69wvQZJvly
2zqHGnagDBX11l8KDCkaTL5L4kI45gmdYf2WkowxudhoKLF241QBdMkz5hhOs7Mx
XEgyk3NXkV3X81B8PMW0HJqNjfM1fHJBa31cIfB1hRnLsuhYvfLBa0QBNh57Enkj
7MhWh6dlb42XVvDBrCc/b6SonyBnA+vt0/zH8ECivtd5cmc6Rp171D3kWPJ7TRmp
tGVht6ae5KqEIO1XaA2EvrovMwuQkzJCdt1Q3XRDUTKqIlWozEkfmUtDl5+PFAMY
V7o0XcpPU/RQ6/hssrYPW4644URtr3slN2XnUaBdPKOLlQEpY6qMwLSt1Jbe5tVZ
9cmY5G/x8/U3thORO5SSu/PH6TC6lckT0WTq806Btbf4PoOcpeWFzhzkVIO3x+Is
IUm9/0M8WMsxhMJxr5jizQiUi4r0V45qbtIDxz7f2XviV9jkPD2znAoCC/o2a4+f
CrxIGDsIVGfFwJRAd4d/8C5x6kLTZjEEvRwDOs8vWTF6pApuij45hsCpq6hp2lgT
v8pNLvmnFxlBoWnxX5jpYmyz/Tpy6w1LB9x+tE3Kbnz8eM/bnw07QP8glX92SdS4
q9Fr7pNW6bN3EBrzSCSgjnuAtQBiSft3GHnkoNZ8THv6lycb1i/5D4GxnXs83RiM
YBHT3/lT7pIHEioEIVEFdX1OL7M795D7jOpEqaFfiKueBfslwyt8qvWe07f9ddm9
g40ecI2GG3s4gYVhSfCLjrJvfYJdfnOYHXNzwBTq0m7/OUsmj8QndTJaZIqwrBuU
QiL5zpdV66z/1wQb5bnSyodyla7Tr9dT87LjwgHhQMNVXxg8gPeEnkB10CZFh+1t
4cd2K5V7ioejX0jwWmsroEWfiUBwwa/7nx1ZKwt6TWDUx5QD0V+BVGCH0zz9jkO6
NOS+hu0Z4Qnl27Zlix/qTtuVo3Y56gBGHKdOpoVBU3BtGIQ02+00SMfsN7UYDjoX
eLPvIVb0eLBX9QUZLDFqWZE2NPaiPn3yzY3TrHf0nvTioCJ5o3tn/tjRI/y+IXgX
URPWWyaKwXdL79GBalCGnNzzS9HtKcZh9fyx8IETn9RmfEl0acC9mjC+INUoKBla
E7PLD/uB07/3dksqtoNYlFBXwgXVml4j5SCKcNg+7Zt29ggdVaCFjWAVrGI27Dus
Qo8SHH1kcN29/S+82VtBCQOSc5zeYM2V2frxecNl5m/NgZZ0VwAOEDBk+7Arm09e
Wsr/WhbZU4Od6cTof7jZyeuDbQ8bZZgo195bLZQ+ei6mMClULRMtjKJ62IfkbuJo
eMhlK6eRQZ+yh/Q3sXRSBsJQsxmoID5CyhhyB8BSPzLRGAynia+vay3y3DveSuTo
IGKIAZzKRCWj/PfmpjXpo1eqk9naCIUkoOcZ+40WJkSbNubZGOhKhPNfGwXdf5gE
aWINS7BuiVXmWbpFBKIq5i0mSo/oUooW055ZKKVInwQ+lwUqoRJys9EUlWtSqe3A
nrhgAlgQpw3h9Ta9bTLYLmsWC+g+f/9zyFPpR6LpTxBuGZYadpYv2m/x/+gtKVic
Yz/8Fa3LAlEd0vG4FEI8LQJmO14z2XNZQw13TAGSnEGXtoqP9dCAGTspVwMCDqtL
giujfrYeU/rdVcznlBAtvMrNFqEpbmHvupEAjwvPDApbXn9vbvBAbSgpX0JBYUCJ
l4UWws8HfN/rhNG+LxA2GJcCbxXlOzBhsC58mD71ojlt+iYr5KMZlpxZgT27g2qB
gvxCWqtp97bWdgjhAoHalcz1ClKRjjU4WH1DYt47g+3K4RRErwdtd5bfU644gAh1
oS5R0K/eSF6KRkmPRW8SyXSsbfoBIbdj2iZS2+nfH+Gw1LQfgWtcqQLydIYQNNyw
iuE9J9sclqCSG/KmSSxkCt8v9BFsLVQ1qi3uDG4tCjQZ167otoAWTXoxOEwoiHe6
8iPN1JABGxyRANIAadCNvQoXk40ez9DaroA40dEj0i6coc5tuezJQKGVJR+CIF8o
bipctig6BNQCFVqCgw+VbjD40CUZR10JpziAsVJEgMgrHITnf3dw13TTFxT+DDaF
G4sMO1hp3p8i0/Bi8VqD2Velns6Hu182P+ozlB/+Qy2Z0C8wdOzwkLAbCWtuiO4K
SCZim/6L9pjsPMGeZMku9d1zBRUktrZioDfmK+kVwF59Pf1y9YpkMqggAzHMCDb+
CO2uYhj1Of/6RKfiNUbRQfXC26Ic7tdR/orWzfWEdfHEPY2b1oIf6GD8SfQx+P2B
kgUlYSMyC+Q3Yr7Zya53mjO8dcEcJ/s/nRgjtURZbcrlP8qpPrUzSEwSoaRhPyF2
MS3ScGIROpt0Mcq+CxSfeXIc7XT2hYPuaCn8nSMH6fG7N0PLteNRMATP3LRfsv0k
C9vkwW5PdOLt55Sim/MnheNqX6Abn4UqAkuUKN0bCLH9Y5Bz9mBnbeTYIkS4IVz+
TNfeedCBZ+oJnG0i9KPeeEEEm3vP59+SGru5eXfG60apoQpkBuZ8f/ZhioZ7cVmm
dRsOYWR+1MqLyX6OTmyDxzyyWSLA90Lzsfvf1fPOJB7S86SCp/5Ih1qSucCnr3ir
+XIZCsFmrpHyCLPZ0X1f7abLIUV8OobcdSHkQSsKB6dDslpr9gRFHRCsAcEwvnK0
59l9Q5ZfoEBRTpJab+qiO7gphFJpulBSOZXt4JHtWw/HhNus6UYJRLqmpfB+J5Fm
hOUwAJpG0nf12yNhqEhPvMzS2P8UdjflYRwj63U7eLDKpnBSkiBYe+4260iZzr0B
RVZE2F8BUrNO8oSwMX+8ItD08iSzDH6v5bisoH6yZ84ZOE7KLN6GE/OOsl3LdD0R
2AmyjC5ZVWsv9RwxyHQKdjIFvEySnSJM+GyHcw1i9gNTTNQaImGUm0ykfSYqNASP
OjggEYCqatk6qEkkcoI+PAE5n9/jD2mqmhIetkvnHjolfdpuciupOmDN8x9ydRcv
3MzCnkrDjB/3+wOdttQfjW0aoZFa+KoAaTK0/N1TcNQOuM7KARbaAhk6zL2IBo7Q
WSV2azh5mIQS8jnGr0mKHEl4FkimSJkd1OpCFPlYyYewENUXpqzWRJh8qLQXIqWw
BH/l29kGoRA63lVOBxRb39C2N7r/OXWnE1ZP7u3lIyv8flfyXxv/2GUafaItU7+W
IbfeuolY3IW8S0kMEr054wnzYCFODH4l+HX6KhXX2uk12u67CC7M96QFC3OZEhUG
bK0xhBfovWFvyvbOep9tPQy5PbB08nVDvHmtRIgYHd4/q8OdORmd4vmWFCjrRy4+
xQXoYaBSTb/0XtZLUktGwhgrJPGf3zv5fOTjPOUxgAgqGpgmX6rhtZJ10glUvs0L
6B8rEUK7feCQKb0XWPW2Z4POzpSUV28e6KNfSEg1WeRfJYrR8+kg4x7aZXq8GA61
Wz/6jbp9t4eje+/sR0HjFMbVlGdNGTmZDw9EKyQtvc7DijH4Ty/qDaH2Zw13HOuu
ZvFx8Slw5xNAlRmOuJ090V8x5B/HSdUTZq0KiQRZMXPpiH68uP5XJZOEuDtKhlmN
WkH41hjA3dHDb8Hiz1ri/BKH2aPim7bS5CdXWB9txbcfGGAE3yR0ixbxIUaK4VZY
EvNA6ww9Ppi+1IF4fhTV3kFlrXdTyQTVGv2UuQFFbe3c/yGF1MeHHuWvkZEy/0B6
RTbvRv1Eaq2quCbj1JmGqsMOgB4tmyVfa8MZsm1j5l0=
`pragma protect end_protected
