// (C) 2001-2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
jk0YKhW9iZYK66Rc3mkpAiLh1uBdQ2+gxlo+E3hAF1EHGe7TRXCGXlFAOmnQi2fJQ6idXmXo4WEz
VB/RxG/Ck1w0Q6g62+JxUTpNsTg2pvYZQRXz7Loqirq97LxSkgDdvKF1X+8JstZDK4lpD0Mebp3/
fbHf/8SEQRokVDrDEUnl2fBB2ZeyvJ2PSQQ0E3Q7PKXMPHpEt7HkRrGgJpTAf6h6FjUNPsKdz/HK
6P6nUGufmySqlTz7hFhQdbo60yfqZHhRtghaNt1F52S/Q+gimeEp26B4KQ+PnNfx236fG6MNXP/2
YeE5/+Cq3FRWTxcIZVquaagHmncPR8C17Q+tWQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 14000)
JOjjo8N9O6Jo0D3OpCCrp+cZNF7F950RCldrGNmhZbDQbPsAVc6j4/FQRUK/EgP34a2hmTXSL9ef
W+enSAe9B3uMqUx84goIl0YGLTTpXwZvi+Mb6VCtRjPW4zz8PpTrCFhljBTasCef63kjnRMbAZoU
GTXWmN0v+eAKPMbXkIvQ8bt85/n7pflwAseh2RRWODximPjqDW/mRerLDTodHqdwHG494+SiUPFY
M/i0sG251cIaFJT+tleuYW6AhzBfzV9pvccrjh3AHpVBZp5s6VDcch+cSMaYoupXGNNnamPYNJ/V
jYrZvdCzhkt9A7vboEyjJa+x4G1Rp95ZcqWXK10GnJwcBlgvSe/eXwQvPW4uaAZywL4j1G6LDQBv
7CKgepnfeNMC92a3cI+i7YdNb8rbMhVfASzn8/up3b7KmjWwEqk5vLQGc6AIWEf6dQmKQKJRSVTJ
2MFiDWXTr9coMSmWwBpBYR+Vx85Z3BkGHP0YShxgEJXX7nvG9HKpBym4nNme5g5a228cmM5dtfpX
kRrpqlW7/5c31Z6Bq6ntfMWZCDjx5Uapdhg3M3oxL6Kl8zy6lrpor2/TXH0gRHTrBnznccC8U3SY
9lzEG9XS+7hmCMxA/oLFDuMunki1jaXSFY49DRTX3w7DzbkmrFLErLdSef2OFEehELbw6kpC+dXN
2vb8IMTR1VBsUv9oY5Y0IeehzX2LK8kkW1tYQRjcCctVkpKyCkBw1aJZ0fbKgZmGMRSfgWrVBMSh
4P6oskzddvliDMCXFGJeKS3w7W2KGXDwpJ9BL6hQhYwaMG6EG1c3p4i0Q+ppl0PxcxvbkZRSIWR2
/FtczTTcOtrFe1PpEceVKcXWpNoq82GPkObyzzdq1HlCGbFkRNW7et1kbfWj20o4UlqeZSgVDzTX
TM44nTXgUru4aRAVog0g0kSKjVl3zFFpQ0YwKwfYfcxl/lDiwZNR6pctrk135E+szq2bOpfFG/Dy
mIWwbRA0xexw1YaTXywcqawUNkKX1Jb6iwvuCZA6ZM6xyTXOqfiYFppaO3i2DlKI5CFu7H3Sb1ep
6YLl9X07SF/bJgxn8O7vjWwmT9q7EWrwSJKZeA8MCfeGt5CPmeR+Vbw52tLSOpOVP5/dzpf5DIxN
F6yA8yFFnmmCasqPcxIz2zIWTgM0cHelLpMVmSlxWti1Vrmd1S3NHgeRZ1xlYASIFrEbR4eyeHH4
zEUDY3THK2K9nOJQwG+csvxw5o3Dbh/98AQ0fR4Hs6cUE+3man3I3SeIffIQeCluyXD6BFMtmEmA
tNHO9/ORrRc8lkjFHJxBVrRfpwm++Wc1PqNqDmF9h3bKuqgDdGUTDCRlXw1eHdVfEZnOOSSHSUuV
4s+VnQIV16OCk6LQ474iTUJ31UaWUxY21sS9DSGRi8nLPD29dcevbPnMvNJri63sFM4sqaTqr36N
0SeFtHCKy3UJCdEaQTxe7zZkHpiN1emCEXKDbsCLo7vWtO05fy4GamCWxRm50OsLj1OlllIE4xVR
MagoYlLlPqbBocEHecrqrfm7eLXXs7nNjgw7DLXSBwqPRApruepk4auwYMbURYTJ13Fecm2IsHB8
TN6Ie8AocatKJCj3Rv6EOZ6+hTO4kvvH4Dq/umuzMCpBMObLh+0lxdq3VLiH/03n3aWcChft6BK4
Eu3es7zHc9+u40XXYvh1ex447046wMg2BlX3rbePMTki6qWGew+z0g2FfyFmBz7RilblsUl4EMmv
Lq1+e0XdcViXf7AIbezVa57A6nipLdyd7NB2AHopILj6LV9lDLQ4qHckvTw17Ziq9NdkhiwBF6I3
MnFO1zjM8wmYch6prADJ/2M1eGGQhLw6yBwbGjxXqXnK+aFfeQeFYVkrutn55ppOVOU993ZsghnJ
9+xtZuZd2G+WhLikFhsTQ85QghOus3QwG6dWdiqlvN80Lmmb4YEwNvXkEGs5UDpJ8igtsMWK0/FT
kw3XMAdAuz0POzum0xHLHBswq7Z2MzcaFZ8xHXHzJFWKN+UGUkpYXxBkFY48eiZsGUQJzpC6HxiR
0dBJLH/0vCRKkJbO3t9K5M8n0JMAVt7sUy93ThqNvCRh0XzDr6A6V88aMnen4mQM2EO7xk461QuK
qmN/fLRSXCYqz/zeLEyOuxodVMESAvxUIMnFkAUBPM86ax573P1ECpYxOtJzuukpcdJhCDumdKb7
8dGRCSB+RHSccLDLWgcEOGErPyOd0kywnGYN3YHnMGMBtd39ekb8pubPEscC4doYC2SCCAOzJRVP
RhLdd+g+4ZoU55GFWGkuLfMyagbBL+pTMRhtyve1hCw3gmY3B9xyZuDA9MzeQIE3fPgw6A1HiMzT
RXU7KIFHEh2z8FhWTE9yWAlrKo5r3yOSfDoFR4UFQVhddgtIxupabEbli2V+kugsaXrajVHAMygI
qkWaMHe7W5lgBDP68c5uWu0YTrA2zVWuQwd9REoqlShigZd24SkFIObr5xK87z08ULM5IFMEfa51
bE7E002BpX79Q24RiEWC+Hda73vLNvWK8OM8cLEChmGUBxv2fQv2wqQZ/VBiLcXXhDd0+nS5aprD
9zXr7IHwPTmSqNEE/tmodTIZvZTjQrCXlRjWcdEuwikPWk7Yznry3eKcfajbqijhIk+CXdFNg9D1
UHTAZ19DN/fIqTzTEXVhiwnTLRSOwDqCdELQFh7JXxD/YsFdlzhOPRq1JiSnyenbcL9T+EM7iFgQ
17O/cOQj+TkKMKudOQlui2FOY0yXM+HNpBqZ5fSKL8F+6eMHRkSAbwoYg+Ex1YwZxIws8hE8iDOc
+BFMW/S9tgYK3omb3JSiAVK7r3nbp14rVmFhZZy/cq7Xxj/vDfI31ploSXkamILzwBirO3n+/BYD
uWPA5xQmfXEzjYJoN4VLvUtQsY8rLVtCFjrQZTnJZfNvP60z5OOtWTb3PLf8EYn1qreWpeGjlmwP
mTzZvVmdwMiyzvfD4go5Yeni6vFgkx6yTmBr5hd4wILNbADgo55j5pN5l6KM5igIhAD3KjPuzUqS
7YV3ChL9kfwjMr+uuFoLa7GmXCRsfWu/MAv5xqIsnjX99i9q5Adz48vRWA+08hip4WyZ9SdVYNKb
2+Bui39X4llhSFrAL+jZDy9fLlOwSaRXCAvfjq72hyUQeqSEm5/53W/QpkuMTGirm3O5oMvi5j1n
XKPeO9s0uyloskOMQn9FEPlY2TloHYei2vgYdd51cdmSuzpW3A/xnF+6yewdVl1DdB5D+X+cuSNK
WztPv6W+ZP6ZoMLTNOZOgO0uPmMqL7Bqyv/oiXU8HKy600tbs7pp9t7XhdWieKNDGxbur9FWbH5V
iN2ynZdYWICrY6V3j9u751t/zzoeLXrPnkV9IoQ1fmwro5DraZEk6LOSe75igAOmqYR1ULkU+mag
IItUrZ7Pkf2wdcgPbsHqWl79Mz9AFHXkPqLaCGOHzT4b3OetuHHglzFARNvrDbE0D0pMvrsoZCil
6UPNMrORy7XWrg+yEg588kVk9oDjjmRWzCgczg5YGWYF3xRV4OxPWD6MApR/DMFpEzd2fRJBUGd/
zVJGwsUgOnHOcOAF3qAmeOMo7oxj0+1KjK69H3RfQwnlX6mKKIjfMAOpUfDke1md5Evo32DhYfxs
x36sMCizXuU3iuGp8+6uEdqT5hi09sLbvl5qrbKPBRyjqhHbZ/iaXo/++IGG5HEXWxlxfcgcEyne
7VkklSiNzgf7mTsyudYU17kTtaWS+GFtntsJKh3eV0vcQIyP4Jzy/KM+dhNKgNvDtxa1T6o6lghW
8zYoyO4B+9jBAsAuaslI+WDx2KwEiAptuzrkoPNsUzj+VYnde6Zx0LJE13MTnRN0a6v9HNf/D1DX
kVmWL8gwhoC/+iyUENVdbvsKVZoc8R8Skv7dslydVwDu78zswG7xsDptE3+XIe9iy8xG3hR2gkhz
Fnl9mMPJSn0B6SwPR5d6BA53JCXC9UzcqMnWgnDyCkBOdVwDoMpHYHBXVWJBOo4H3rQGvPCTOU4b
Ronb8R8vyWYk31S/cIzXbQaSAs6m7N84fiIkA2VgPyD/J2we7RW6Wvm8JgtX5KvsSxIUZxfHi0jo
ItJvResgyiUcAqXk2MxHBdcOJc9bOA1eRu6QHUzfPFFeznrLZHH1AXPmekfRhLbFGeZbcxeN/c3T
fBfuCwIRQX3hcy5YE1NMY4tJ7qwqrjMZcQ7jDgD/t11MPOEpuPaxyuc4xx9UkzKRv3CYwFL73e0r
m1SbI5yLMr7eejJutHi4GNJcgcRo5z1UTvBLp5PJgItenEPCANiKApkjJVXNmmXTJbADauCKLm0N
YDmzcQZ+SLpU8DMwgQROlfbQ2a5w2Ark0MMbGwGteYzZoBljlvZUAY2oul+aSabqH7KVVNrtb63F
svG8+Yg4vbnx40hSL+ysQkWBnQp9GvMbcBK0sKbpilkPSGhrycOgce26/YpshJfnQ6HOqsWFG1vx
+NcuQ3QH0IaXW1v8MrijnLLYnO28KX0R2k70rm+vv0K5WEBTCMGr+Dow19hU5FAKECcw2qE6NCoM
HhGNO9ep9Cc6ZCrS9UR9EmRhj515LCbZc2OAMa6880O+55rumqtedECIdIE3chXsP6xWWV/Baa4O
tTOaH7WdgI1bN2sLNalHYVMnuXtdSbzCOzla8TW2/kkYSPnzRPWYL7ImRKO1+WU+6UKNpnJgpfqg
HcaffVe3qMCIcubWs4p2jkG1zHFoZrC7EwFjgg7lWoGMBvWepb+XZqgZXOJsJeW0XQ+YQZF2cs0V
LiFykOo2Obi8Oa/8MnDuyXK3OE4KEStQIXDFIX6RwpY1DDh6fARzU+40uTqTvohSOyoWChBpgXer
S15gMPztZ9KSSsYq1ePRVisfB/s8HDi1ANcecE/bc0E+rw9C6snM2oVmdtVh1HfP6odaxqgID068
v9JPweBc5eZnLh28YRSmrXrQJHDLnJVJVekZedDzbacNUsdLmZ9L2DaFQhsPb+rsf83DEmJ1TlrA
5/rnb1OA4P4rkh6GFA+wdyHY59BIf0DrEaavgNrW46MyAOxs4mnQupyBb3pH+/1G6dangmflB/05
Uzl/bvRPPCS8d2AK+Py1GKzuCz0QTZqacHba/U6z7+MDILtLxaaYXYcxV4YF0jsTjLnlkprmC1tA
xEIa3jrPRxNcPYKzbK3L00H9HE7SQzyjOYs8OFJ36WHjDI2Hpt0iTddVZ1kpgvG6VsCBERlymZVi
EGUcLYBlfzp5QHNCXT/ntXMOcEyLnD9GSVWBJAJF+ZLbkbywut3yZrE8v1tw1QTIYL9wdZ960zBm
7c91ORfgchZCDeH5+0NowGRkLUrzG203mrT6CWgim8UL6IpmTS1vJUKcSkQp2PlpXRMtW6/YnJM1
JVkFAEAMPX/PS+B/ZchQ9p5mvBQqdE3vrNPS4kx3erIXaBN0UlE98u/WVKg5lrnZmo3uQCNYPeRd
lDWbaKPidyoPxh7qtX3RK/J0SJvzzW87Ih58llVOOBVmOFDJOYjwnloqUXe8B9UL2vYKcbW35QNZ
4THn5wBfHY7KhPfNGLhh/s7n4aNB2yK0cZ7eTFMiBiM/J4G/u03eFskfY1VpyI2XQJ7wlPSOgt/P
JcJWL2Dz7dR6U9K7tNXNHY48LoUpUcBcwv9NpUkKsZZTVymAaqEdBLHFUxPU0CFDZp6v9RDfyMtV
6CkR30RppZiNVVowgFGU+bSOhuGdZYJ1v7AvBhActOr1m5tuOktBmwivg2UPHoXA++HYwnMr5sQx
8OMZG60QI/ywGdlc7cgT3oYQLbuBo8kPpd2WoizNy/qdPiuUzClqjlB07DuW7V2ny4p1smJgIlpd
YT14+xWTYpWENoIyAW1KxIZqKmzP6Axn00oBCP6rt4k0+OGf05fJtNrFhR5ZrNgkDYiYzz9Ojn72
iHpLEm539kyUHUZLIskUZwzh+x36hTugg+eUoEoaWwp8Decpqtiso3xHxOwSYfysNi/Opx1GHSG1
VBv3t0Vj6LSUDwkhxSECsNW1rTLADAY2EQqNX19283BAhDeSdBgZPcUTS7pw3dz6noNqUOMS6vOH
tPFJ8nzZK3yMtRER3CZU0Tx5lwJnJJG14nygWDxZ9yKlz2wSd5QAK+wjDFTJ3BLbyjJRkMCm3GV8
Y+/2D5+gsak0L5r5JVj8p3MZGryxlZA4VAvXGzddkARCIFNGkNWbv/MZ0Inqw2B6vSzVcmvEFIiA
60X73WeuZPyYLdQb3XjKZRSlPScWX/mdD3ur7Vo1Ui1ROgIY6u3cwguKuMhcvYVvOGjdNQUq2J06
1U6JOEVFT6Taw2sFjWsdCVDJMCBcKmP+8vEhsLlH991e5xPgPXjTWVt61PZCSY1cnpi8B2GuCkbq
y0Ztm7708OiZkFyjChVUd6/h0Fc6PLdaD5BImRPGecpplx3M0Hwfb3elEfxdtGrQuXRIdvXqmzg9
KqFJ1zdMvlTtSX1+NDelHsbJZQFY7DAvkTcvLKdn14O35KYuP04CSYHW4vqDf5tQkeiV/iGnJhYJ
DSLbuTx5fO2Y40tLz9zi8ZGiycnHxHAbB9wG9Vab8mVj8RDOJR5OoT4XGW3tn+I/7n30Yd9aArFJ
p3yjNhQvvTCAVSZNutl7omBlWagJWy5zuVod3GcQ4KYmuJz0Sd5F5UY+mQ/myDO2UuPRgpI8dYcL
gKZ+7BvZabQJ4JX5rAT6H119fRUf+OOZlTqt5A1n3z4S502kY7TL1BJIn9Bq3au/AHlInB/Rxemr
K3kQE+tUpwCwCkTkGTFriGdwtP5HD637ZncvV1gquK4FlofM1cYgq/Hh6UpSFbeVdndxE+UI3xsV
4qsU3dTQnRV5kog55aGVtOkEtLaKPQhcRLmSMY6Y4SxRldpQr0s8chGv2E+E+3tdYeXANs572ipO
nCRup+v76UTT307bj4AFSEApjdUgwr7XLqpiqSqgTk6DSoGLCD4GgCdgyFE8/F+3n9pQvC6yt50a
BQwshOWyoUAIoxYKQXJF3acs2oYdgqvdHcH8gClMkb952CvvjXAw1AvEPnxqLrEBezQz3UVNf7p2
ws8bFiLJ6xjcrd7grTN1fqRpkW6yjFWeuXcmHpVh/8XX1OMuIRsJlQYf44cCL9BNM4RCszk+vXru
q/zVBCPJWflO6if+Qo25GPAGPlFTDHrpW2eQUecyBxRmswh97bkG4JMe0P3V9KqxlgEBTPVmS0Og
mKma/fQuq001ztyq0BJnw3lOm9KLMoZQvhXSzS5NCcvVAoPN5GriXy+MxGvt4TYj2Dp4LPdmDmJM
mwVNnxjfYVq0a/LRKPBIE8WzLkN/RrR0Pppp8y5Ot+SuasLc+jkCg0z+znmVMTrjvR3aWsmJrBBR
lI/XDIABLRR1mbYp7OMFHHG3UjR5mLmDrMiKf4c218ae528tn0NLINce9G5nkidgnii4/wADGyjE
Rj+Y6naa3oJQqffJj6WbhcQHhIZ/sKDRn5UanEpRiHHCgmESd+TnRAjAVR5HhKcLgW5b4c3Wq6mJ
k1CTPF2dC8v/u844wVuoP7v39cg42zUvYBFYs0NoU2lZveF/EQjPvkt+VeRnnIY3dvtNabjVMuKA
WNe+6oS7HDI8KFCGcKMsk1LygW0BR/tnwooAehsGmcSmZZUtYw+XXbpAsFkRPErma0kDYankFjcE
ObegbLFXKI4wy0peiA1+Glh5oknCTw656lEU5MRICuZFW+VCfyBxjtAfHbTsQmEmox/yvnoxUHnM
EZU00rJOAIEl1aFKSbz6DOPAq9qyR3eSW15wB/7mywqXiCrA8JyoeJUbcLUmdJQDL1QBhWQQxQgb
jocUssh5YhpIJxBsYTAHT1VMIfJDgyyiw28pAKp1FVSdhKP8gfUZ1tcrwtoTRqFnCvLStkim0yEZ
dW/laRnEj8aYy96HYu9BQ1wh2Gnaki0/1YH6Vf06LphQc7hoLSVCLpqyGwk304H0SiPrbufN+7ro
AWnePsz6RXVJFSE99e2gCL4a4QuV3cq7BmDaTS0b128+MaNRb+Z8Trgmu/CoxbDQDpifQMAc3l+/
QIQGz7xkoc4GLKwdznizom728shCPsDoGqAdEbry8WpuiyVFhsPrXtQjf7jsyt1hHPvUiZj5OOQM
IZ7eC6f9RPA8XdRJjVHx1ny9nZnJqXUNfPtl8zZoy1acJ6T5/jv9u1TOCJ3sofF9xx8LnDwBphsx
0bl71pZe/B4rJFyiN4T73ctuOfwZgS3yud8fHZlqQzgg2FByuQkzJGhtuF9jMckpbxzOdIJ04RLn
9j5PHZI2dcYEcttFlqpkVPotlMtWBPOoU4tWaukEENBfbWo9bn+SbgDmU+9Z5tTPPCMcKJgIoSi+
LsZIibvR2BtYG1aiYFl1xKi46GIdQTKqdt7tIDmn+AE8FWD4BvQNZonWIFvygz2jX7XCJ3QD7W13
hYm8Dgt3U2oBkaNhYGYYL8WvHYKUKHmVjN2uPmOzPM1IEiKQm6dFCxkfnYkZEdRgPqeozNtm0f/F
OMOlOk05lWqoZXZIqX65CJFdPFKe8jWPYeJRzTJhiw51W8EyK/jRCusluOlqOAjAnQntuu05ezo7
gf4w3/QJpxaU5c/I9TFhLiksEuw4r/jspuX3/hGubBdGc3Lid06bFyYJqv75SV4dqzvqxt2Qhmld
B+VsrIC1yWV4lHGmG6QG8pBbhf+6e3dr5pcK+u3GT2SQK28qMKjaheVJJjhf7ULt78TBOEUAnlbm
C4ARpked4LykTz2nX0h6KMr8JPxlMC2kqaf0o3zxoOJ0MJHBmcdyHWWFbK8YhEXgwVgTvUZnrXVj
ciNd3zv13Zy1n75i8t1LmxFDxQvVyBITxSn1+AhX2GYP2rFknbfTTDZVjpfMAkdTyOaIALB9ohtn
N8nWkL4nSo93H30JiYQJLhBmvdquyrRcqlyPOlKVoASyX8aREkzvtIV0SjxCgCAJaIk/ds4XHcDs
U5pjvHLWzBtHnHLh57oatSPz+EK4aRRJI4deJTm9dRMjFxF+K/sUHdOuzbyzjivMPF1OQqa2LnJE
9opxN6yeNaHjqfKHLuLZZhaGzC94Ml6vwCIJAUG0IB5ubzSfixh1ovnl5DJk85qWoumN9sYcMRut
2WW++it367tQrc+nWa1mc7b1oBfmaLYMDJr+eR4ywlps5T7oCgl1jZ427+1B/Xeq7QJOK5uEJNRn
e2sntX+3oNanI77dW4JtkBaVGOfFiUIxTnT3GnhBr48aupCI0d4zIicjQUVKPQ1M4XSea/RE5gIF
j2LtQjd6nyObT3tpwtC9zH24IZbzDuXL3s13RtQSitYBj6KwG2g5EIfuJ5qNmbax9SFAUd2S+/1J
mEMw+nV35Y/BWVCh3JB/U/QDkE2yyyTbd+cFQxRx5qGWxVtvezsvUafhDpNkGfJAoltzX0/bfz1C
HdBQnr2OQc+gexPxlwEHYGs4ly3r4bk6HfNgMo3SHBnmnvqQcTzadcdTnm1PxYY33DhG6TvrZ7+R
7dXu4zBcm9hCc5G5Ih+w2lKdNy21wFllR9vWnNW4YXBBEgTxMWeaHGwBR+fNW8bX6FgzoaxvxstQ
OJPCRWxLDdmYixIDSnOC/5tAAwf1JcqhOZzXSoyNlziGXQSypRt/g0cQIGVPc5zGYdSLAxwcYZ1D
k2nATK1n9qaHREaeqtrFegX09DmpY9W3+Glgb7LypPIgk0+TdMEsJt20eqR9N3PeFAKTcMp6gVFu
U+Fm+y1Jw8pG+/wddGYHII8Z3QG4Tadaxr39D7bQ+FctEJWz04/Lu/FvsNKX0V/hFoFETNn1gZFA
+SRhFNIdmfl6CVai8iDqoICsUJEkFmqFy0vo20yAEOol3E1GAZdoVY+uMvUUCWAn/77gbjO2NiUd
8UPUrscPLqzcmVsXgP/+FSEg3UKuMbyFDjgXtWEto0LPCRETYub4BMHR2xh5gQn03O+ySBmjp8ws
UpA6q9UbaA5e1PQQMn36Y2eTYKfpgBBK8iCV/bFppNs/mzSOrW2dQHbbUyI3+epPCV4SpmLI+938
M7ZIzU1p/bPHsDzk1MllK+2/10XuLJxZdsWxy3y84RyMNzmRfHpmB+6QCiDPAg6LNvBOSkV0PFcJ
047t1brelLMKboaygVMCHLH/pkCB6FDMPTKAojN+OgmubVOgKfAhSeH4FVbz16nZkqjAg4AdQK/C
onelNjqGZY4ug+1uv5keB/jZdeCSWEYVigt5hnwAys96p3iSd/frLqIlJDvUcFCG+5B0PKPkmlff
yVveNEIumbZN4Qdw0muK7FryS1C4tNvwC46t8GfEjG2IvADqkVC5oZPHlwRfGZcqF306tuwBua2s
zgajKG7GY0KoNZSHhKsHvUE1cQy/L6IGbInYZftC36vsdHThDzN9YVYmKdKG6ARBB9M7pPdjZJD/
07ySLie7Dn0jaINcmmh4LxkR/o6n8/LKyJTrJpCJAKn2IXEi6Y/9PJKgPpe5tHfuFOy1LKYZNkTB
W/xMpl2EsiRFWuyywIhRb7GodEe6vNMie0a8qMe+egu/g6OeokrE2NkTCJuNJfGTKPlvrAnd5sb/
7Efr2ZBxzFcVeZNn86kKpa/upSnsx+46ARsffLdfPsxdsm32cYLHHbA7qWkswFPUJSbnkqNxerlM
t+VcEkr62dSvFgRWrLYndJcVkz3bsuNWNQGHQQjS+DhT8JiyMWezYeVcjL2JWBfMEWtCxpUxak75
OA/uorEeVYMDGdkewsSbtjlh8EcLlnMU89cZShAeqkcBxUVWxSKLMHJubfPSE0rJbMROYM0Dsts6
0VhCq9t0bC3JpuC7KVaIeKh/EV+j4CdV5JoiDWjIyCcRqW23fsvyLFRNuYfpLlbz1QGqH93ysPVf
x77i2ZkkIZepUzgRGBCIiq6EMb/X+Eh/q8vo72JVdbqUIZmmu+hNMHl9kiEkA+UqytZy2+WcewIp
Vbb0MQH9wa9Cb36gpGAUhF3VaqeyLn2aIhk+RY/jT61uqVvwJNBn8R9NBFYcpRYgc6qdZTd/r519
zQ5OElZUnD1MBRrSIPAFKA0icQDLW6EwZXlHj+KQiqjckKjbhMw5pnGq1trRVINyqlK65QxQ1rEX
kOQ5mPTPcPuPHBJwqmvNObStOwZ2lyns2dflTeo6hLSuHDIII0bPBaLUprP1ihRvzktydvCV26JO
GM0N3cqtIoj2FJEtHTSn4uxfRHOBGEv/7+XQI2q4gRpZJtRH99AnijKC666maErRRMw9Ao6TM6lp
CIL/3mDXD8nUBpULXmLcjLfooKHMdeMnKOqnEnVH62G/0snjDMxui4yTL31uESufLyF3E90sTq8n
tw43WxnSq7SPg0BgkMAg/5AAklUyGgvrhAkSsqPxtWIhgn0lRgQG2oBHIUJ/gZCUlFaqaegmHklT
/4/t2WbsvgGOK5QkVHcuMxhOQCThMTqwpIrwtzOZM43oxWOnYcLSdoL+p9kglZUGKoisMEO0zoeD
jagpNXWzk92YfzoWleu3nmSyFk3Q2bsQ5whQs59vtIcYLqUnV698shBss5hPRsQBsVir2YGMfWQo
U/859oiC4cOtfzqMnmCNAN0YPbfEjzJf2gSUGa8mnk9CeplPylKZOodHTfRR4vdYy4ur2qAunAtf
vymaMvPb0m2MdbT58sfxlvs0eX4GlySbe/jkKhdUjtyM3+Ha+6tR2t22iywoPcnBZAokw+Rj7vuG
EQoFFg1gyJseZQwiubsUioItwDP86JwB/oM4ZoUOdkyC6nBCWb7PYdV6HpH3A4vn26+cnwGJp43U
kEpsSJ6i96i2xfJtF5rvMeRx+XqfvBkCG++Bwix7LL4LDoV2HsIpIfygmX2M/UqaHP8+c6OC6dLe
jTh/HXQqDdUfF56EiyL5AZtoFx1fxvIulo8pBBkOBXskGDXYqXG7vJ+22zPkDBaCYQad1A+1rYgT
HnCWGBvxsKsPsrB1++VK8V2b2L2UrsyZAYOLTKQnvag7yvKw+coAUn07gJvM0B9hdWs60EVo9miK
v4noHrw3Am1vct9kFYlsb9xKerc2g87aRPmJSsL758Qp677tcz+bIUD5BSOj/GIPhlF1Mj9TSc9/
SazqFygawFfdb83BtqTDlGp5EiYN8rt6FQjw/cOwsjrUAAtbGaFF/F/HzX9EV1XJ+yEVc6Kcb+gH
0RTIPyLbbAxCWEcl7XLDqyjXrAP/EuMFFAKIBYE6mfSkk5I4lL20CrYQ2xWqXkJsBFJ8pKMtVbku
mNcyr5R5+/BNP1X/F38dGcu5iLbh5vTmE+y1kaL2hJgFCwxi3lxqRbXguCJln5J2FGUIvDRJoZFJ
DMz8+IU3LgIHCht5TYEDEqIkh551M9E1fiqVlmODvenNcjudo0LKnegt2CiAPzj6OzW0b53PiqGf
4S1UhzUDzLrBtWSkXh+pykQwwEIJhxxul0KoP3Qk6CqoywhfJ/RJEdFDZ0w4lwozz0lCYnAqfTYg
Xzc1Br/PQnkRCNKP9+vSG5zelIg5Bv9MHJE0rNnp7zxa8aTtJwDxKV4lmRQ/6EwtFbzrqUfA/07q
JdKxOcgJlHev1m0cHjqZIYqlRvVOvWwMx8dC5e1in21jFJnFV/wzKLa7npYw7OWycTyyvWx1OEOJ
I1sxRs4IKlafaGE78CUzjrqLBN3PT0SYQAXW07UVjAybAIPvNfcxKvl1KRG3MFjBYTERoSMzNn9n
5sbPCk8INjz5S9BttBg6yvuMkJX5NgC6sl4vcY5hVLgieeZjuw6uFZijS94Tzo2T0JzG7R0MiVYc
zeUhVCekik3b4jMUbpM8VkCo7OUsC8uvtHRtr+Uu/PZkMw0arbZ8Pz2stT+U7Qsi+EZHTF/sctRp
z9/nhio7wz4Pl9906rkrkDZxLCG+CeOjJPExPU/KN+9T5P60ekXjfBNMQjQqNlCXunALKqjU8c5h
HyAdhbs2AetBuTvjIC2xt8eb0Uy/mCFAmpTnOs8yusdM5SJjYSgNj5ACCs8s6Femokb+Q8f/sKWm
G9E/lpG/NTXhjF8yXiZt/lqceVtPpXGSJJIQ1gq33u3HmS9CJMgL4vmdElDxlFQuVTsQPFTa5J9G
KSf2AcPHbxObcz4coeDJxGYwvj973xeX7bsFEs1bteSBR9UzLiWPYifW7960BTHF1h2IM9AFCmYM
worMg3wd6lu87uZJ1bT7R3BRRYzzn0kHo6pbHMYMlghyGP9D5NuXRjvp/A9ak4lJLiFV+vj9KB7P
DjZZ6+hO8VLSEoRyuCFja/Ibh/ZjRWEw4DdF3KVHtWg+0VQLmFYZO18tbbSJJCCr8VmdTtzbQ1d0
6WyGJTXjqGbdH4x4xDU9sAP6wVK/G2d9pW5aIZE4eDmrmbtYlIYvS+GQEXZgp1Ss095SSS8ejzOv
4xRf+GwP1CVoujiQ9mal1DbSPHWR06aRlzbeB9HQiofdQlT4k2wKwxZZODzfhMUEOja/7A2peAts
UtwAJG8EUFzu4gM+mr1beKHkms1MlzWPAJ+k5PE8C++F7vN9WxLFvajPTSJ//PPvhRPrvIIjIKco
5pAhze8rUG2zDO6iGvBiHJWzgakRMgjC9AH8p2ds4ugDz0Xvl+akoF++/NvER3a3Q0h5Ofo9VlU9
xkB5MeFsUYsAq9srzpgcklRZmOUcahgdoVSs5aF2KuX4yrztsfxFyx9bZPxD2JuPyB07K5mrSYP2
qf7BilB02IDb+gg0vAGBy0dDIC5MDJPoo1hKg47v/eeFLjXzu6E3yV6r6gZa/IP6wqA3gVn56M83
1uo4pTS5ivpYdfjpt10FfnmClQOS56s70D7bpSDf1QWNZRSrTMomhlDZgA+F05La6U7PuSCtPHIk
9dBSxlHDtkMbVaBottHxtA79YQadxugchJUmLF8bd6fecxQr1BWWUUaKCTImOfClh+5GM1n0npz8
1pZ0zIZteScxIRVWi7moe1CYTTCYgJ4qy+NZVT5Om8NHk04AqKa9LLMSA75B0k9q6ANGnMg3/+/G
P0P6LfbZqrsGQjpq7z7Kj/sXsacn+Ni8931sAa0RjRDSiM8/FdYwcw31YH1tCK9/+xG370lcjR6p
PQnVhE7kiZ4phTo+pKOgALPxbvJRWcK5H8pk/coG3qrxupIdY1sNUPkWpZa/1czYYW3XClQ+CP6R
7RNeTUdgFq9cGdmIedKkZyJcDF/s227rSK3PxNSiO9Zc2Uts34/tIEBCW7QUeeqqB0yOwII5bbPB
/PRPY74nLfHeflTBvNYh2XB/fAlRUxSCF1jSLo4avSpu8/CmrGSd0HGPbJo4CO+dFa9ewWdh1UPO
R00V+OuLHxJbkS86QgkzlJnYQEPB7MCaBuvOk/7/0vk+7NzNhMsHGwOemr//QGv2DEXQYwtGMsZy
fOpz93uXTj7T9BPM50Gm2HK4rB+SpyB1S1mz2pn3jwiKaRqWS7aIK7BsJ6CZEltvQQUhJY0IdBJn
N2hL2r76b4bWDqtkzTRelvv2Dhpm59DE5/yhjAYBfeDa4xQtev7NFW9nXWIMgXyByJuDKNMWQc6A
wCGQ6dwkpNQonBzodoH+O6vU9xqqzi/lKIRFQfm9VDxWk98DqhEsG3cV5Eozfw8umdL2ZkXk9JIK
Y8yENaOKomaVZSWkbf5Vt2P7iHKo+9qQbQNKwyu2G3bE2xmIEY1I9svwo4mFm/uhUWVEyU9WdUnh
sjpBltPHyWLv63ci93LPud2hSauwfisP6fSgjoLCXMhil7ZX9+n41jeVYt8+Nb21uXPZJ07zUIUE
w7Vjns2i55Ghc9YSrnP8rEBAqIDrWdcVmgHvh1Ngh6RTKLQKGM3KcgJYahprdXSf4WhftPBSHrlg
5EYbvE8yMcYv5xQjoMj4Ilke4ewAxS3XVzFMB/KggCLheysDVEwoWmGADFL4M/IDa4nSZPxY5bbH
Wh0GWCXXBOneJLWge7SABSfDQTKAX3IDsGEn1dCCASgMtLWCtyi1Jm9/qRIvz7BDKqAFDVdq+G5j
scKAGMxT/GUZOoLrjPw3PKg9RnxjOfWRdtD9bKbVO1Dw0zAH82VJUcV+kV/0N+M/othWnN3xTkpN
mRAqyFTsoxsJXAJWCzwu6p1HHUNcSVNPRLlLAqz41gQuhzbyaUWHN4Ww2WW6a1sT9t1mOVG6AWbZ
7EBR0tO73ZrVavBQtgKnsH04PClTA3beipx506n3ew/WEEeCG75vu7Ket0gnjdH9Rv33zJmSseku
fcQ85U4/0qn4CQLAQ/NVjh89aribiH6yTsMyCaVEGsmRo27EpiafcLgTqryrTFShOl+/0kxXDGFx
wqOs94Ev1vCHMKAGc3Z88MB/MSPh3tcb3flImTRMfSGi+OIvl3jrtcLOgM1UAZvsVtY1i/zl+OJp
er9dBToRMvYJLy4K3K8TQV/Gdlgw3SVrpMSzWoJnzFCQm2S+elQkM9bdQeoPoPPPJOLDlLEbjubG
VvnUppiVb3N9V1Z03PJnSlEiCVNvLS9KOUCZ1cbe3YWqyHxIHNCDXFuKhTMzQjp5tRpWDGEETX/b
i+gVBjh0oFmvulH3RTkb1oVEl0O3jnmGuDH4ReSZoCE7CoFU8Uu7YL8emWNGjiyaLix4dSeix1YK
HXiKa3MPqulSgxlLEIb2n8SN32QZD8LARiFfZRXM9LAfYtUC6UXSv55hIqvN0Bb9N9NKD9XYg1ZQ
40Y2dmqU/Oi4bURWmKknKBr7huX2PRxrheVo8Lqcu03FMORayxPgD3pX0+Vjd5jbcO98pjg/b6go
mKPRnFaJUZH0FTW5H5FwbHhn1Khvk983tNpJ8psrHDGTr6EElGnjrDc42O94sAZ/AaaMgFu30LZj
lBbeno+UORfdp984IAd9RvZVzBLzp6dI6yR8Hq/4LcGE7tGT/V+GslCRQvmO8MX2qpzUCmFkihNq
l5Vc7Eq3HYKYJu6ndtU/SkMO12Svrf8a6TGRXdqU/kdeGV1UumqiGDPcwkeTJrVXP1cVddY+GfS/
8JgAolSOS9EV2bYV2EbEzyl+O/rIwqgfuKexUz/T9WTGVV23qwXlK865HvvBgFIaxRc18/XLYiMO
g+Jw6VPxvJZ4JKQ7/hGjeRmw2sQhXWbe/RLV5tAyCzEdDHLOOx2n6vd4vtQn3QFweixfueJ2vky/
Go4IqwqXdHsvBHsHtE+dPm4XtqgbUFaqR0bUUpXHeoEz5PeWJ8hC1XaCl9ChuPN/qodej6u3LmD6
TUkN6NmGpFXk2SOtl5AB7UbnoTGQ/eagIhsPC9XnGjyeZdalcV1f/3aOgdx+xK0Lr5G9ZryhSjnQ
9Qg73zyCzKut3l2iV7vb07h8uZjsMQydikvdp3iyqxYK71WWhzNn/JIkiME69nA37hgkwhCdkYyT
GWrz+stJ3bUUIMa9MN5i17PPfOTDYJTG6hzCi/r5TuPw5i/tPBInZn5tdJyH65FQmEpbQSf+J9nj
9jCfk/KvEykVXyOH0HmkCqIoN9DqmrVLmHs1cXfxZikoG46JmRc6z99ZzBQ4OC0pN7a7tzrX2R+P
PjDXEmfCQVBXjfb8qJfdISJwV6uWfMQZi8gPJwc4JQ+/lyfkfiAPeqmOW8365t11mn9bAjIsaCn5
XpjckAlJtG9jggiM70ZFMl1KnWkS40D3ntnoqYrdyTc0f2CHtJHrOhGtKR/2z4HrDw3qRDWUFvt5
32G9lr/UJHFZCPTTvgQh4PGL5w9sdtXBMm5z9D80pAwboHiDiKlF35Y5BN+Hqio+uGqnK+tCAinF
4l+LEC7AnuPt3hOKQq509KSGiGjN2sSlWAa+Ank0hntcgBZAWDLRDw6Pz75vUUH3Y3GWKjXv8CwO
hg7Trkdcia6sywYv5sJunvfNpx1Tfc824dr2b+pEE7LCc8M2MvCShWSpOd7nLOpgBp9wSWUaxG4V
tK2KeLRbx4cylyJj8E2U56Hfm1OGoQ4eS44LXXiMXkKbiPlN4wZiRP2RiyG9s4Q7vPObOA18jzob
6+sq4fDg05kdEBJyIYx/gFOX9ZN6poV0tRj1exTeN8fIJhX4EQE5bqxIvMZ7hVPucyJ/rlQZxScG
SNaJLuNVeEQrpoC5DLTQRIpfLUMaTnn1vBWSV9sxUdd9iVHKI2xL7xD8pO2f+7q5RA2Wkt+HSQpV
e0c5MWz5ROpOKpqLBSJLmcNJu3/k/ob6smYrt4x+mFCrUQJae4OFQwJ5CNDvHN0g/25dDQKHsJUk
Uee9EjoePy26OujGAGNDqtdBA7HgKJnTX4JeNapC1weWCjwHh+0ar/RTyu96RRwFSH2MwsUO/7QG
Xusg33pUFKxw2z23s+up/oRuauAQDv0L2Ylf8edBT8/So0KRh9tdgcBZx78EnxhlL5+HPHIfb1tc
LcqKbWBaNw7jw+rLrphqUiM+jmkmlUTJ6193rovcn+hJ5iK4v03CwUXOLplVgZJa6IidRAqMwJyq
/1O6nGizSTteTp905eSaFNxSpPnx6bZhLraDCXtgN46qZuZ+K0c7m2TDizitNWwTv6Bput1GcQP6
pHLRLgsC9kDFdRWLf7o98Cyx7t41ya+VKeZoBsX/XB7/hqTqrvA3iPMhn4RHj8Ip+2Zm7up40fBE
9Iw0y1EFtsd5GOfFJdulHmyoTpZ+Xc81/3KUbARLJx7154GJeklIGrkEYJUSt38UwwUg7i4vfFeq
ho5V7E0YEBJQ4XWC9LpLWJdo8a0O54+viu4NzBWm+tdG9DcRC3KFfexTZ/IttfyxL+HXLFj2xYIQ
/4yY8LgVglkw4Vai2HZhje/Eg6j8xrT/pB8uMKh5pSmRupCSR53JtR+ZGfCmcnmVE1RWAsERp+GP
ylbyWB0P024A+p4tZCHh5vEJbh9lSLWl8eg/fjovgHjr6YZIDRgnsBeBK7WD/p1j1X8INAbX1sjl
56r3e6SYSS8j/+CLYUbLhgbZqrjNjyUeGmrPjk+0lNu9zMl4iKxUAUwr1UauO/hK2yYPs55KqZwa
6btO9NJOcAH6p3YPHw7bX65r/kw8T0h9menfLjOcd6WUgS3oGqrd06zU/0k3EDHSga8sdOZR/RH3
ZUQL9sM1IV03M+I7OQyNDZty5c++4iXQRerjPExL2kce8XEl/tRGhnat7SC0PDW8zxSBC1+vaGyk
uNDgdDUcib/jO6qOq5rIYMZQL8ENIY5yuEyK+n+//OLEIySGgswnOfJSKH9Sku9lHYcdBe0jsSaj
kLpVCrQPksXihnHcyKDQyVVa4j9Sp2rAU3qRYjLNuYbyIhz2FfGu5KgwCF56CMHUd5LCN2yiHl67
u9KyZzTAdo5N9/Dsax6+2V+/9hme/tcJEQZqtcQBu9plCmFRPUsG/8/DIKRpZFi0JROLk9iy4K8O
8a+OXgh5YjBH5jZMj9V7t8PJbXsKv5rs+kVT43qiv818aueNGkYStfGHFhWpVVVVT5aPBzAVDMZE
tMhvy+mlOpWaLlfZJREZqzgy4diDr4ra5T0yU3Yaj03fVzDCpC3tXEibnY9/ctegoKtc3cW7MHvG
LJDFdO9bRskpfSkEwkghNUlH6VtXAkUAdMixmpZSlEiqheFnfr5X5NeoyjJ6h265+nocW6tw638v
srsnE7vQP665K97he7SsVR1MbroafT7P/ZLJyxOG2liORfAk5UKvtSBzVziqqADP+qDj05bNJ+rt
ekz7GmiZ9kJFhpVR6WMDI7QshEY/cIYDjpbgRnlM1OACWCk=
`pragma protect end_protected
