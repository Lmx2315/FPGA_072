// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:36:58 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
LP2D8MxAbx4bN9vR0+vrS9JLUynpvkFjbGzIaMLhd7UNfRL+zmTbGeLe1K92c9X9
oEMHY0wnBYEARHgT0hLyKA6yw5trGoh0XG0b7cbIMIk07j59bV8KSgBpp7O/K0dc
Wd34n0oLXlWYtqaUWWMW7u9zvMXiy3tvuQqV8c0NPLs=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11472)
uMg2D3KoC/xqt23xQo7QzNNc5lbrtrYLEIbTo/+FLVFqbKxeQx//9IZJa+iG0PeO
EpyAF7/Q7dj3zZQBeb4FwyTEaSYVl+6j2d37RWCG2e7zCyn3Ca2cKFvF9po0yiP0
8DtD1I35YLV3r6Nc5aSG1qOCglibm95bmoAomtgGzqWiLT8vUglCCJo9+bTi5GIV
lBxf/2mQ/2+nRX7D686DrTvHpVqVeumhT06hpuWiUlH2IYjDwVI70Jf3UW6YrB9i
vuDfv0HUbeNMO00K9fF4M3/oOU32XwnOyJoobM0H+64/BOV9ssPSPhZBr0/1niqz
WbpSnwe8Ut+fohU515ANCDQMgjdTBEgddBduiep0L0UObN94pEzbXdAGQQgRnc1a
N6bEN1+UMew7p8X0zVg+QYRVno6YYVJWpHGnGptfTe7SGbNtHAh8k7YFEftBKewT
v/ftc+FbyNixTThwGY4HwodzOiEBGxV1gJcgOa+GPGe/Mu+CHRMUvNLqcJYj8rl/
bJ9lFBvAsn+YDQ2gW1vNoSnPafLCKMGtLXDpqMhzUgpNPeLdvmnUd4AHWknVuHUh
nwXL5QOuva1a8eny/D6JisZQUTE0rHcx0oPCtT8Ty1BN7c5p34tS3U2xQ2pWh6sg
0C/tl0C3SKAbQ3U8JGnrM1O35QVQDNfExoY/oFmsbQJKnpHEKpGqkxwzPG/uxlfj
XlbjPLgtYqbj1UOoj6BU4CNAAFkc++pMhxdsp/5tqS4xhUQ8PKBI7OfJPjxC6RCH
A6hcVOjLJct/Y67Q387pxFJw/dehBbiRkKqRN5qhdZ1aabgJMDgxdcViq/GA3oW0
9gOabBA0JMdBoFATe4yHRyDcKFjEv51KuVGPPs/sAMY1aw6LHlz2wm1QhtjTc6Ug
IHds2j5BUUZvVwBQbtWJjfFw5qjA1Krmc7ovjT6nkHUWRTChWrU6154vhQeM/v5q
MwouB3VuctNHI74A5m0h9sYXAiFvefca9b1n6vPZxQY9lkUA/o3+6ITbEHJtlveq
DEI3o48/wgc6BWywVcPGxQJisa+8Kl87mKsJcS8Xa/vCd7S2xcEvW7jfbPeMC49o
XIRMxkA4m7rf1wFVtFCepLEEcLRhA4ISMYSHu240kNumuYHWhBOEbUnOaaGmu8s0
2OLpdGZYZsCnW/Zlzt+nYTnddrvcRYa01pG0RSfUeVWsICDNFsLgonbPx1oDEUGz
AQrd/dsJZYncx5xfPLSQM9i6yAAjueI1XsTW5wnPyFECaBSeYANvaJhrctPwrC6B
eIqMvjoP7Sijxe34rOpQb0JgkL+yGZnt/AqjxSk+f/pFvG4g03SDtMjdtk5wuaRT
XJNwG2y9AsSaX7XBNQPs5DIE9Zn6o7kXdlrvIhq+YMlG4x95xrR7mW8H0A4Kcaux
23MvALyLaqRlevSG0kRqyjokVtQ9FrJoCMt8xT5Z9a/p+t1IA4pHGSCJpPpZO8Ah
KuBm+E/pnLaHRryc8tIKWvCYv8sU3XCeSt2teW0XFJha5aoMYC8R1luFEJjW0u56
iw5f4+2kNf5sDqSyp9P57e5iiloUMD4EKYORjtL29YdWI+iLKhwCE2dfWadbYJR7
p+BBaj11mzVgkfG3yc7ADDP5rnwg5I+PUEbr8VlHtzx1PRjHLVixRQ4JZ36HYSow
aApKqNaZUI0D/p5cFJVPtBkokz1ktrsh2C1MUzl37Gk4SkfNa2SanttHalL7RpbK
xalBg2h1gzzz02VLdSb4Qda6y2yZdTRm0UpeOxcEkCuV2YnxHXCJwY2g+4f6no8U
7ed+f5LInoNn92XWBaUVt1lN5nNJTGkSE8n3de/iyKSm8+hl7LRwxrp5CUetrUF6
fsTlG7CurVZ/Jx2oXH9ijOHlOZUvrIL/sEpYfQZvC4Ysm2ghotnumfYeM5MTillb
Ei5eFoW+vVEJJSRDqfiDIW9u23imp2EY9RYQEtzrJCvjGrfN8yf3HnQC8xJ1zsUw
lMw50VI76T81jgCNFMKvRxc5EvBXa9Sy2XBCeN/1Bl44tUZuAiqy2M34HOTL8ANC
rDA0CRMzi7IoM9kPc7PcZ0FebnL3r2dhYy21oQhByapTNzWsN6BrUOsy/EnfIJC6
6h7FMhFjBHXrfduinpXe+fBvkwjlmdnzqRVeNwge1kryejweQCOwK2W7WJutoe8S
jS2AhxAkV2PE60XFqSUfeLNBEyGj3q5XzmiNtYuwshpEzOj46h/+v2JLy9EH8nI5
FFj5LIZP6gWeHgZnTvOwwZwqZ4tC3HVG8Q5JMi2xyeXEuEceq9g0ZZpb9D0xlW+g
UwsGw+BeWjuCIQqUXilgoliNtk+DvHowwOYyKGwZxkUD4+bVlBxKW2EvLU5V3+D0
mTHfAZiwSuTWeJcyeoUMgpXV8PHJfBsDnTmL1fUeUnSVhlI0IzcpwfJsGxXlYlLl
W34H4SwW7yCgQ/sB/PeSuhtj+N6z6JcDHlVbNW9PN37i1V5uWYGaGRGc5mYGejpF
SrSm+vNtQ02wQJ0kvbgRdKpKuJ/fwjafdM6bVIOYbickhC0T5VTMREZWsE4KWcF8
v410iO+LE34NAd+b0CHyzgkje9Y+eTIqidDBU8y38nNFYi/mZJvYginuAlDQNVXp
JsEGVsLPEU8DtjgAXWAzPoQEL2CN9bz5a4/Uuv9VNiJ04x39bBNu5OviMgU0t2nJ
OkN9gAHnyoR6HEK+szet+GsroSYeV3w9JAvTBdQtwAlMCsIpw+8l3jK5lw9b8tIC
9wl/I77kmKpY7uVVpLHQevxLXGvPGNXEmRmuHiZkrycXLjmnBzvnHBljqL489Vpc
PLxBbLHj9+mVFIRUEg1UoFutDgsGWchy6vRbOM11uQZizA4G0g335i5ENcgkBPX+
MKW4nwtOTakzXKea/jwoWi/7lU6Wwt4Oxh9PaHGCNJoxriHq1Nk4rVQJ+TPU6ETs
wbo9X2WTHvwXsuAd6th00jBURhRQmQLSiYe1BPyjvoB9DvkPOiAPer/RaDFP53Ed
bOLnOE8vwEjEdY8UUm/Csw7Z4lRn52y1BcONRBpdeujF79Kb0RY+OOfnpQkSNxBr
rY6JpPVyz2uHH92T18N1ARB6m/anETV238hWSE5wC7/v07Jpat9C9T8rrf7xSJb8
6Dx+VYO1UyLv94yKVz2q49E00iSJe1hvCJvLsZTiNI0CaNdazhlJgNQFEuSrfH4p
tovxIa4EBuXVx4H9nKb/B3QUcjXLWJYOt+oUTzpgTbjUuNcx2fA53O7o29RX0M1V
5r6/PNuCM6LoFW/mAYFwuLkvYcwwdbIRKqne6ZymU7O6h2izJdgBbGD4Ff6vq4T2
tLP57729RV3dV4r2FIjBrQmVzE69xqANxqlSdcP/k6bZ2p+MP0vHFVYQLr84xRuJ
MtF8U85b4aNzWmBndqN3xXfWUT9ZWwy1doTkNbR+LhVh+lpBJqnlZJiZMXjchsw6
IPIzE5C5aT2/vyMBHZavm+PCwWPGhudt1mkUdCUIpHz/YNJzUfLmQLrESMNtgRrS
/bluvPoJJyl/CyIxK8boI9gpMdxEdTVOqRGF5sfL/AaInNPsrh7diST2xXtc3mvO
Tw/2usy7kPcb/wKozfESL0ypzYG42/oH9bu97B4rX6NDZ+y9cXs3nGaTPb+ftts8
VeIeN0LK3Ljo29/nYHweGLkMhpcJPl4FJWpC3ZKprFIkfXHgxFrWEFaNN0ZbrzVV
oY/wcD7DRKKm7Bm1iHP0woHPfqjk6UxCiAzS99h55z1G2TN3W5jDBzgQaYvkU50p
QQzi6wX4goFsEXQlp2MjkRlxJw32BkqHwCSQhkV884PCIb1F9OF+kJ/xR5uI1HLq
c4p3WHMgxjBqbUEumXC5OzQlT/77xZSVBEwM4yu5+9ag/70bxVUxzIMzuUsRQyeH
gf4ZRNxBwjQpTtFL2zQkEvLQXdhR7x9BvxWsLDDE6StGta4NOtwwTGwQqw8ITk4f
gD1RQj3zs0qcK+kPloIBwjaAGa8lfAYYIlsXi8NLFnna7o61uD1FqnjspFdk1m38
XQxlwHyMkgEKGPEj0aJoyeZHNBYsQxLm9XiqRCfWQjght1EmBj/rJ3LX4ZvHQyDq
MqwtnVO00vnnRruEWy6seMWa4XW/zSQxGxIgCk0S9zPD3IISTnAn+HikgUqxI17b
n4NFv046x7fTPA3t0OKd3DmkYBDKHbGECgHU6Ckwz2wqy/I0hCgsh6zg973t0C4f
TMNfflk90QmToKD+ih6Xx1Nygcv5WdfqCltRQ8NrhEHTRzYYY18RJ5BCrSN9rmHg
n1aCsVP/FTN0h07xCpGNb1ozJyNM0rVIgDf1Jb80D25d4Jo9Wq/fbUDzR3KECS8M
1D0ASFV/PRWo8aKdG0gS0QX0LCvKj6y0GQ0cZ6xHg3HQhn9Y52g28R6f9PFE1Ott
h+MCRQP4hKzFEH8fwX+P47aPUba6CwMrvHCDf6XSb8DV4e+IxzV1nEqnqtvX29w/
+R+xHZwnsgyvRneaRCPafq+WhoX43ji194ZGCyDszgipKr1QsIO50IhuqXwyYbao
2NzB3EZfKfBIMax8VSmTmnNTLzJZPRWfcleK7DsNreMVMy2u7nithTfDGHmmd5EE
2JXjXtV+CwugfRqU3Bf/7yXSFs3IHDjFsqVhC4Fdzg2aorAsjfFZQiOaDYw6+qly
8N51OMe2eKAytpN+8pvXCQcRhCY2Xa2ZzfLdCyfi1gb5t9iEbAZMt1/lta7W3S7r
k/Q6n9grYi5WmRWv5vjHlg3AbLxec9y0hRl1iUm7iP9CpI1jHGfistHbQOIArOos
2Xa6DuSZ1amv585i0roc5XrHbJhGvoAzdkZjmnE7DmgVjGS1rnX+9fkSSBMor+TF
Cknh1UCs3bdg3T0HBtLH3BfbMZSjDvUPeBrcfK6OK/Tt6vqRJ7yaDhmHHKBZhTiM
gNRoOeKiLgaiDiiwBx1xN4N+oNKXmYxvmngDcbwlSRcOE73dS1eLBhAejn2/TQg4
EYqULifVYF0MYG138XgjJ0ZEVV7Cw7K6+a9TwCtLXE+I06J++Pp3VE8GxJuw/XIU
EVU6umgCvUHXnRUgFiAsJKaufnRO9OD9LTKK4oQFfSCJnTo8Xi0sjO19mF0kQrJF
9Yr9Lz0rtNT9yI0wFGb2aPDm89wAgy33Cjfe9FIQng32bLGjLWG55HAargFH7hGk
tw+rFB8VqmK2SkzYUW46Eut1/eX0h5SBYHx4WEN0Pd9+4fIVpuRs+ZCTs/R+aZty
R3fvZcedJcckd5mkgSn677yWVG8sd9oBN3k5WsHUJfGC1rTU95Ye63YfpRsrDcax
5r4ZkuF90nqJ9yFvn2hE7BZIN+L+6UAZ1JQk2yw1n6mUm4hX61LEMUR4zFezRSGx
+RyZQaEGEAJpy/Z2ZP0YnV0rJnXtNM9p3692YpK3ngtKj6jOvagWz31Typ+zwaqP
uGFIoWzJqkq6oi8J9pOoTswRUj7hafmjuaiWtP33guUTTwKtWiCfv/vlgefixJus
zZFpsnQLO0xQAjqG0slvjdOhfr/ezqkZDrZDindAbSdDekEuwxh6BRe4SbxgKo/G
IGKGZiUwRlJx3ha1L8CWWJsoZKOHUv+Ur+QmtzREZhTRznxfrNIZnGmqnVRrnIdw
YGSz2qr/oUbKWU7IM4P8O4DciSTkHv2FcHovPRJ+7Mhl7rYzD3sNBEIOckftSONU
tHmUsxDz4mxL951yPkO82EdnDgsHRR7QYfErzmDkPVgBl+Xph9B/4TSR6xE1E7lD
emJSrdYFr++YyOkTNEGNroecrIn4hNx/aYITUspPBrrLtHwapiQeoiDS4wqHiucK
Cv8acsXPRRP1DK249uesuvCaja+jne+sCCopH7+5hweL49cgieosN19SPZzJRjiq
ArsHZu9zXpQ8UVzhFHDqiDM1Z2ApAX8lFAiUx38N3TnG0ZMiC8nc37xrXGovePlz
ep5i+hZXHLnqWuGGY4VVQYuEWgSx7ANvZjiOOPLKmXiL6vELigBpIappsipQtWOP
ply3N2FFKqo9r1zZF2fK+bGRfoMo+9h424ggWhw0V192HmrVzDAaPGFDtZlOtBPs
HO4qI52ezOj4zfGV9K8auocW/06vX7X5br8mMrKlW3KUdZZaMB1SWEv4DWfkMJ1N
vKgYgcmfvQbiOXrmGQE0ich3NVXNeElTfWa//BPryfqbYS6wFaT8ROxCSdiXMinG
njGifRFtugDb9yQdq1LO7/Kbeuwyn2PSuR5TI9IK56hdmpfj3NnEEvn3+R4uAetd
ct83ffSgMQEflakRB+8evrBeTx1VdsA7gzveNDg1d9LeoGbJLNNEyQ6CteM3gbRi
XQgfSFmqLKpPSu1i3asnx7o+Pbf51HN72J0Mim4uUSe272PnXFMYYOPbeqb/hTzC
e+QLmSjpeIz6mRayDYOc5k7nW9qb4F8tUrpJ5yockraJAg7LtTdiGyrVSZSPBTyz
l/LteGM8saWqxCqukYdYcZVyTM3HePW7gysd5hoI2dmi1fkBMXe7ts5AzQ7biW2V
eIucna6XL9/cdM+Sh4/O6wc43m6pC/p9gW0mkFs8arOU436COoyhpBHqQOpoxkZK
u7LRGkhwaZ/rNLNr9PJAXcotAANOnG5C5PlDOYTW6V0rFr63QI8KosrFfmoDDkLL
IxWl6HUAyx8K5errQSqdNG8JqkD015BzbMxl9lsVwpDjfQ29s1N/10uok8g7lO9w
XzyQLPA2+8twKBuHzdBkKEUPt2tjfi4wUt6I86fp1i+VxMhbvEgxDOX1YwvZCX/F
XS+y4K3P0G+915JghEXcHptkYoFiNcyYH6RUdvXdB7NlYyV4RmeDozOAv2egT0h+
NR7wsOaetjir7U/7x9tO/D2ZNQ3XJsX1X1OUR5QUy/B+F7XU0v2i5JhQF0/GWS//
MFsETPqjmpvviM98457barHdxnXuec59dpw+zL2ZmdCrvYrE7amdBAZQjEUPyMSX
xLoFvLEMNQgUXynEcYqm+eoZusrQu1cPBeJYKbWKDJ3uw6hqo08E2F3Cge1yNMKK
PXaagbuyi0q5MpyvVi2PaYE2lWi5dkmRjgl83Wtot5dwUlVdhNEdn0jWN8Qhkwz9
41tLEz5z0nMfLBPyMaL88tZXFgH72WHMk64ndOEH1juvwyDgkaf62xZss7gCyq9F
anovtDOWPdeXxLL0Ln8PcPWo6Ph6UUDaIMXOrq3EHNy/W/hCGubHo/f65ZinQQrt
W2pDiWo7v27TlgEF66YIfGW21iPiBgn1vWSddCYNqIi3yyTW1WOUBcRN6Rbfh8q4
iIiiAowdetQBeRUjj2hK8HOY2jbigyidNGt1hzh6e5nNFTogaGh/ntanxAAcORzF
FrMiEvU4ZrI5ExHYE6N9bsYNGZqQewz676PHSv7/ROTql2lJ8G5PoquQg1SyOBj3
mZfeGOWnroC3GljhAhp4SyInSupYEfD028SewiE3fGbxHNphgjOe6a90s6JMn5aE
AiqOqnzTEFlXajvWcp/g8tteQMlesP6Uk5Yjrhx8YS0FjVlkASTzbNQiQQCk8SaA
RjagqvH9FS25LR96TE46qhjfJBb2eO07QD9MyDng66iEqACOSU+mimpA8jGHehG0
X9E0L7LiAPV2Cnx3xCwXiuatkA5G+aPksVBVJ1RITF0wNlI7GVsZh7cl9CWwLrob
CvxTc7yO7x1VCqDAuMt+nhtIM7V6smiCydQTY/EyVa9kezTUv9srY9ow3g2PYBD6
mn4Pxx4TbnqSRX1ptRXZ9AOqA26UIzTDY0PlyawZ49N7OVYzv2vCuqyPn5/SxoLo
Oikc5FHvuO2JsCdqBggtWZDjTxZMYJlDNG63p3WeqSWxYfYfVyWyhgGhkfysa5L6
OSGjEMusJGLHp8nO5FouYSYLPsfL8G7PQgWpTqO9j3ogs9uEOqLZFDmD4f2yI1a+
rqOMlLtNThoisxz7Pc5ff/herTegqFqwgTZl7OOcxB7suP84BW6vVEtnE34iLL/t
uGg+lVfBBM//CPSsFHq9plIf1zIB8zVyZztAY6OF+iD+nDvOzydo+gOofyS7U1Yh
dYDRmB+wI4eJ76l3rzInZF9PuMv6A2iB5Ea9zChWBW6bZnGubG2WMtXNALmRW9xP
wRcMDXujDWW8sjUwsrKRkgVm3KC5LIr9POzNXtevhDmU8U22zqFzkSz+O+ZFNUFn
PagBOMfEFMpHzrZ/bXLp4R9q0VsN7zr12TIB5EHpDI5hEQV3AjqunHrC4Df4GZo5
81C+PFDYgVvQIgZPisyn4UBotnx3/yHk2rldxjJfBdcUkPB+XjOSM64IR5NzgRdT
FHTVoaEPwM123Xow23hdpRu/iKXlQBhF0k17csCO0u6/MvZlCZ+nzhyEIhBfhndL
fJYU7CyLARP2SSidNDua7KfpVtRmXLpZrQhiFMK5fYpeUt3OnraAC7Px+QKUPfu7
mkwnDlqIZXNofFWd4rX5aYgwNIEsQSbHKQoRHI4+1yc9+VqKWSheSuTdETGy2o1N
4Kf1dh7vG6/Z9gd3XLaVodnVKcjd04jLhXmIOY2uQ5CfA7eI+/TnK8J+vPcvJlO8
dMy/UVSzL3B0ooJkToKsmQrmDR+odD+qup+kpG5GUlGxQl2sLiqbMhLqhq69ctNT
Tqa18NYSIihe5IiGarNLFs+oYHzGBA+xOiiEZ202Ju+enyScRx80QJrrCKtRU3vq
h22NrI2WL6mDXbAVKq+DBxGVeep2N1Mav4VMwVMIkPtOYOjlBgIhEsNSDx9Hb6BV
9sCDIUzblDIU0w0CfHaroD5WCbo70nTZgU3E/c2PN+v+XEv6BR7O8shIZWyMpSVF
unRwHbpGhZYDLo5TWrEBPmpk4OhGwOpDVAANCJZP+siXIFkj3HyNMwNVC7vsav2+
uT68mr7sMj62N0EWso4iv9G8GbYOaimvtv9IBcl7QJ73EtFJ7S/ip2gBcBwhACdg
FTVHeJbuXPKtVMAE2rPC/t18BPTvT3hQ+OEsrdTTpw2mCo//X4nD0FRfE4rqNZuy
jLOJTojweiIJWcP9gtClthrR6mRj58bYEV6s3DghiXrSQBbKPrJdJC5UEl+dkhLE
59BZi0Wbek4sA5G6DE9Bfx0NC82IdEbBDb5ZtVzykkPpYXBUUyw3mydlOTDuMpao
7goqWRPBzCpxBXJerYE2KRCa9s4AeBPfkUN5y0olRXYqdBMKf9ReEni8fx55qrQ0
xOEljY/n0+I6HjfVylRM7hCEJ7obVohTuHKBDLsOQgb8vbvMvbzzhRQJzIaZYqzs
cLHCzKd6HvlK26YZX2+eyje2x3IT9JFrflLzmByZT/PhSHqju3dJo1ZvsdGfb+6f
8+lvO6CQ6q0QtXLaTmxssZoLTu18G06WGRXb1AOI7fMsMQCiCg5DusWj0UKeEzku
b7pl2NOCy1bQEE6MQnCDuDdK3zL/9R340GTVyO0ktAdP+RNvcCT3y9OlvRir+cNS
wsx2FNx4GjwEvZcnXb3RbTKlGOaLiqVgAtBWH45zZMSeAnRbdf61hVodBu2d0pzR
bWtqmiTnY7adE1t0RZVW3CvlmL8+5UNP6McQuy2joY/tAQMJ4vyRZJoj3uk2bjGB
497aZZN9czTluUDKXgdyj6KN+q2fRL/sngnrxUnEn4MqLFMne0GvFq/DpyT+NbYq
Bf3X/br6xSXpZjnWWqzPRz2vVJJPTGBF4OvbLTe8iLmjbWNT/q3wVpfIeSZEzpws
jk3S8yFAKkDX17YEucycbgE9Osj0zvYWcUKd1tnspSURatD6wqLsBCEqt1cIpGE2
DRsWJhavnReA+1g2BBCrMKSKVJD8j2L6cNFyJ9o87Abg+y26PLDK2rWRFVftUQFQ
OSbT1uS6KaNEiTC+terImISCc/fHC+ezrBdzzNOWaQLB5zDm2OnRz3NZ5Fi/+tXk
a/32nsRw/5mimUdWq58lsNn3P1SNA4MJ+b+vKpj9hS0cH4ZcsO0q04i8SmPnY2bq
fF4WUAeas7atvKDE5J+XEuQmQCqIzQ3eeGVgF6n8afaX1Nqcdmc3kPJImXfTwvIp
X9MNom/M1TqeDoj9Ww3jqFdhSIMXg35KF1KV72wYG5leZiqpx9eaVCtaCBSLPpAm
y0+ko+CG56oZx4R6fiODmbjjMDzFLU7zlANzyGYm6uILa1zushyLXLU2Hq5OyjMB
w90cYpV2kc5BJVrbAwjFfTFcNTbBSrhoUKHqv0NEmOek5OZgMYU8ZJtqP0bMbA3H
IftnRdc+5TxcqOKtnahUPL7Rz+uzcpoPkNWUMPpWIz/V9uuy3970aOKot0J91xV7
Q7Idvu1IcIZnAmzVXzJKSRW8ocMJhDXQqGv2festniwmex1LWXU5THj07Uf8iNiI
aTNPb6EqPIidfgTkdhvrDZBPqqhL/G1ZlcEVBsw36QEHba+tPs+2Bv+4DCc0im+u
/e5p5zvzzqH7u0qwhhrP/lfsRJoFSrWF6g8GlLFtI0cLdI9lgHxdNbtCT11PN/er
1hsZcrRd6+lBddAchLgSZoOCRczfTDLJvydG22IhgyVbubJ7zj66Wcrrj9LqW/Wo
fefpLqDrl87md5rIShV6N+RHsey3oSuTAbxSyJQjKmWNv6H9DkoQXnrbEnwa+1ty
AKp3kwj/ITGLcvPgLG8/qyCOnp4zYhVmtgtUAbCONqFqLBOf5Rv9ojcB4NzO6xII
j50+T8Ipt7idepdIQEosRrdEsQsjCIqSAiiHfBBcTp/NjQjQg6kn6YP47BpXlXFh
wMe7V9lRDjpuzxusdYPiVnv8cYHrJ+IN73PUhdQkLOGBpKenFVbGEwo7Fn58kfRQ
2b0SdpTaoKq1e2fEhPVvq+6Abn6Fu8x16N1p8Pfg9fqQLOsrr8yrCoSkDn0w3T2x
KYvAlsA+R+TfNpK3BjXZ1W6JJ4uIOzaSCIpxqfjwWFzrVp/pl5KIgJjtar4OUC3m
5o6O/7vaH6ZO4bgmpkqfDzR73HTQCpRcHfiTZGnggQklGLpXrXgBmgp/S1k9UGSg
Jka2hlHhWbxSkuKAGBb7Nbf8/1losWGaXu5rRD0eLLIugsJkbJ4Yc/n5IAwlw6QN
rtnLmM9Anulo8S7EZiSHzdrQiOG+u0p7LW6iX82OhI+h3wvwx0TPO4u8OIsU9mrP
0TeKfqEhxvavHPI8hzPgJRy6ayuJnE8nyM6R00fx984pUeIqBjKubWgQnFqvFG25
AZ2Hotj895Q/qeChV1W7yk5CjJsIUuWlVApq0ApZrbEjln4iYEhMOYaNmMPUlLMx
n36hDcxaRMqudMSRBACdmcjAYdhOJfSkug6cO82PfmVeFcMbhSx4kOAxIeuWQKAD
8r/ZQ0+zOoNVZNc1pAvG/DdLfYf0+1w3Sc98rFgzw/KhI7bHJCG4T1n9COE0ns56
4QwvoiB7TlxAHTQlqLo8ZTiFDZS9ipN3/CBbiq2gC/RvuKKyVrcBK79fdhXGXImI
PoqGH3IOmDgQCTp2S8dZd6psSkmFYNeF/XcLKAXbGdVd1Ju9EbT+Q3oDvy0qrFan
14Ce9ogU2wWAYcu8bkhF9t4z2/9fJBvQB/tyYh/vDouZOiDCRPFLZ1AU+K0DFrlb
DmOGMjI9QS1oXHVQSepJs9gFkNTs1474o80TSSxHii5snTIUMDonHnq+VJUgtwtY
PVT9nsetCqvcdAe44veH+FqwBltLEsHySoeGVKYFk+F7adNexzNjkanfV0HQ7qXr
bovEhpa/oxn4Cl4b0JcH0cpNccZRUb6JzblQIRbE9slIrJ4z8xAxUwEUvv/9GCQW
/60VlUOuPPFhNX471XXC2rG3asgyPUX1QIVEsABwBGBWCt5wa0J6UnQY6zas5oKn
MY01zxByGeC4crShJUe6aDJtZoG5jMlKNdCL//ezYlXKKiMNnXbV1ibAgimrHXoj
ElLH00V4BbkgwGvm0n7817NQYCABjEZvzlr57abQPs0+XAwmbyvhIRrGJUG8C5GL
tcboR7gr0oe7AJ5Bqw/DinefBl4fLvI6fgOxCpA4lVtGYPfC4/JWOLEP6C0lrgs2
+Yu3isrdFsyeX4ceg/cAEgXTqxFXnwaiM5uhJ0hSrn8VFdUzbb/MCi2x07ABDnjJ
AngxY5kMmaqBKSGlmMjDg5g0yyy/ghqHcf8jhXILXI9qnEJjm8ZhKzFW1uL3Q2zl
wj5ggfoVUwWUTFQBgxj1TGJWFZD4I+ubpwn05T5B51yRxvfihLOk4MVbGbG8mpb2
EUnxkjc97rUc38jbYzn7imIk2fcwjEFm3aJM0X1dWKEKbpCClPFoFtX0B0y08K2c
Cf/NQ4in0kkCrSvtPeXQMk5deuurfOoe8QsVnN5mypyQ1iau26RaJrn+1gg3zi0N
3Q2U7wE2DtGFlWyV4u0vZu3MhH5drQTAiedhX5q996EgSMdtEgioE1nCHz6UWO3o
O/l+QjIHGsLKx8qadN8jA4roPCpm2Xf/h5DbeyGhWxujPjfQP1JM0khXwET+QWZl
6QvtYtcXPji7PqQZU4/KVLgJLdGTnFHb1ZWBVbzt0B6QSMe8LCnsNPgjEIh4dTjj
lqmCBtYZs+RJ6GBK9v5SluGlPP3t0wX28weCmiS/YDqiSbMONBXfGy9PeOrRuta3
qjzX60Cr28cw1A94agKUm6QEMiJnCzK2v1Eh2qF8s8InHJ2LjoYg1dOpDDDISk9H
SxkNNS23Ro+sSkh5ZSHno+5Nn6K4L8nHx4raHEI36dBrN7g2ucYL7v70XF6h0TOh
cAny4IFNJA1cHI3FcpZCZ+JWXqtWsZyvCODyhO8Hv+s9RFkzmPpLTBcJipVrajaV
YeYbUf3zzB5UFT+7UiyCgIiu8FPnEnSDAqUHLBOQU7/spXAN9DuJttALjVmE8XXs
3WVzvgLf6Q9s+m+HXwZaZmWDJuKBMLUXDD4A/+bSjqQydXkN//nwCeaAo01mvhhV
2/pr40k3qqiOUW+3rD3ctvtTKOgslHOJB7C3ClNggFgJ5g9GnvzNCfH2JcswTjPZ
h2pSb1B/xjhU0GEGjBiOAkJvQwEOnZ6nx4lalylYtOCViYfpsWZz98PUFYOy9PgX
MbZac83XdvP+ZjE7ZnYGfkh+QGD2h7bivQk6Pqz3uagaqrXyhBMFwPz2qKdOwbds
4ZFzwhdOhzr68V1D/L22mNvYj6DNs5DGuE6kTKonTF5I8dZCU1iCWxFJCe2IwTX1
c8HlVrm8BOguRczEbVv16yMWHR24A6q5moqoLGfRydeGt7AUZChfu3OYUuDGB3bE
i5Hq+SA+a9174JmNx+Nx5eDXOH7VhyUTu+H1IK/QCSOCaCsWDbPXwQdEPs5ufIHH
GeLV5OEgZgzOL2O1eGgW7YniKvbU23LyD+s4QNG5ckpTm8iMMPjfk6bNUDs853bF
ZwEIRiXWPUzj1jhOW8PDf/miwbTOHOUQk0wgMMssqZvDmD52HyycuOgNTrJVI31B
olXifWNW0f+w51y43rE0X9pNRou1aJIv7K7p4a2mRzV8Kgnxq5XtxUScchhpuEmk
Ksn3R0/miVbT1EYoPfRNtt5KACfnOuz6XBa2sFytAioz2hUIcx24EPqtFtUJWYfy
f90RJ2zqZVUYfa0qopn6Plj0Mft0zkjKxvqZiXdXw2IJFwQNRvpIKVRjYs4C8lbD
V2kS+ndctHdvSojykWwYBISZuWZja9pNkv77nX61W/BGcETB+IiPfmfTc1A0rlEU
9ne7+oLcWqWkPjl7f3RCPvrj426QEOO7Rl2TMZE+lMEK2xdexqILKlwLRJARQFwK
mkMA1vs0cWa+Z5+LfNbXeAjahUEnR6AgbBsQ0uh0E5Yh3Bp0R/SiHZvJ+IAV3Ypa
PZohaYXV4HAXOY8JtpTcpBwPSDgVGYqJXrhnaZ8595Xa4acg0lDzQ3N/HDClH01s
9XA+5A3d0U3hicZLXu4PCMuysQN6vncV8YNAmC9OgE47EqMjzvuoO44Fi/n+QhPN
yVzLMP1YYvQwrUKGEWHADpuj5kQ2RHfdHQo5lFt9jC1r/FXh39PTAvJyXwcO7TMI
+e6YtrlmYSoyOJr2UAN2IVenPV8JXPP5bq5k8aWXTIqzubxFN99ju0yvg6bybrxA
M8VY6FJXG/FNkNbTAR/i443c76jArkV1qsRo56znUY6JJLL0jiiR+LMM8iWHid+j
COKD28IlVsd9n4xc4OLejJ0w30pELOPT5OjssSJTeSZHEYoMGcsOIy3KpPhrTG+S
j/kfDRm5sRaU6IbGezf4hJdvo8o+9ZuppGZs2Jq3mr9p3TMFoP0VDSsjX7lE/Q0m
yvEnNrIEZ/9kUQZofURxfvrqwZCTn7PsO614Xp6QIoM9UBLYT7DS7uvtlFK4Zy8O
i/nNQp5nB6rPjJxdVbSELdKWJ2gX5XsG+DDBRtz0ovt4HxNUkvInklE+eTAr41gg
svUNDVvCyOPGTXsCX0Twv9uxP+PL1iOJoIPyNw1BstadGnE80KZUH6gAejTV20al
ogr3l0E9Yhu/GnVw64jrT5OyEI+m1EvwONWZQF8AmmZm4IQ2LNcR8jJCOiMhNpCE
jupQlq6QHnApv2NUx+tFewBGjo2psZtxz10urdbihg6eZNEJxoqAS7UGa++fdFnI
/p6fuqTlfAAawInOl9dxP4aaunormcyRxH4hvqz92/xJwSnsyOx/JIurmKl7h/Ld
wYJTkG5zmNZHRzn+vaoZX/xPpFPGt3GrhkRr7B6Kk58NQbrqIJ/x/OyrYlkImIjD
DycTlVua+ObFkTjAemCxPBxXBmDzVSgFSYbwBw6vHeBgR6YzSyy77ReN4FaD2c4c
IEennA3QAE6WfDOvTbZ201mG9P+G6lnnY+4gMYqACH7i0H82MDOUHfZb86Oq9qVe
kSd9Hk83F2iGsY5smtyOpgrdH0fYAqpKJqLJSBWRAEyOhQyBopemiFIIt6vFOPeg
fxPUkZByHa365ajzUuvGB+kFe4xd6Sq5XwcMJhjTkVs3HV73HDfIcTnqGIrl2Coy
xM++kNehOvrWwNuamOQURB53I/PXJc1ejdxia3qMlaGVSe/uX3Qk29HYnD1jCTRe
lLfvQXEZRPOOnTEIls5JdRfRmBBMhLz5O5Kw1tYIzPl55MOWqxWOXgJXjX9dTVHZ
AUf/wucVUd0p6oRcpvnLVCbipD6I+VeF5yFBnqiOMwSGLyzAOKH8CsX3rRwRmgQC
O7N0p6h6gTDJ0RHN4NTOkIaFfWknoqR5AFF4CobHCjGh9y7qDIZd7jeTdUfZcDQc
AYNitM35g55aKNHcdANsXVAKqbsxMJZETmoRbVFBgh+CYCI3OgB1s9/5PjOhzJgR
`pragma protect end_protected
