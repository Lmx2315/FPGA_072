// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:37:00 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
r1cpc6wTFhX0MSx3yXcdMjN1lWOjTGBP9O+4Zx9+9Aa8z53wDPegb8iE6YIADD7H
xDuDhczpt2BWfQEeeRIIkar1Nyb3tgcuZkut3gV6FxaoEJE6yghpkCzpV5FrNRRg
X3QVTJBahgZuxWh19PMjNsyY1NsAynUSenPDg64vzds=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6400)
MYptrvOTSqgE9keumGfqSc4NIBTZm8JJTx8/XPoLT8flu5eL19nRt4fPwCb9U7g5
zm/sxMqPdCTNA3TiAsWUA6GBzt146NPx4KLymKL998piQ68PlXk4a7bloApEhXmY
/VZwezmuDEwGsbzTvPART9OeDiO33CQLPwbbv4t80J0g65F9iNw/DPy/i51nlOeQ
4ikgeuHV/VeV6RrQMOu8sVunQWlyj16wf1K4tcKJVUJaXpjXkdtaRKnmbpi8J+Wz
9d/tUXaArjWWC2m3BvpQ2iAo24qI8rM5e6/PuJT6pOW65S//VsvGK/TuoxgevDKV
h6KLQKdrMbI9sFvmGWkGVuvIH0LnU9OQBBSl+5N47fVQWHXixAFaQdDplHevvk+t
mlArxp6EE8YdRNUkkJ+6fDcrbP1ZW7Ztj0dtTzuo+chGTL2WTyWMf5nVbezLCF/8
7ZvsSBk37anLxgZCTssmwC4xrBunq8dn3ErRG1SY2EuGFurBcEPtD7l3IGbojBPb
x9+DAWoWucrkcJ6X1/G+xlmGPuGYJv4nboD/D3YazATbqctGASGktUToumbQecMF
TzRwKXPL1V/u6zxgxZDKSpM7dZMY+3IPmnqsM4DCQQXO9BhqMFYa+AwPNQtoB2NX
UQv0LS7YTlZ5RqbM4aeTqnf8Dl/rKkWzqJsrr429qOuKwGs5/SqmZnrWcBNdldQx
Htad+cPpbzIuouLmy1kgvGjUe8+T1UM+XoH9ZLIkNja1FuOOgeY9aGflNcQE6hPi
NciDy78aCl7qqLvrtzSklE6QFdkOZhrJEq9jmHyLQ+/q56lx6dq3saxFnWw3I2g0
B27RH4LI3i2fJ23GOUVDoZ75bNY58Pvi/TbI2lgzbzckZ810KFdaP1gRuHzdCrxX
RdHutTyn5PMhRhEKYgswz+0Q0NrsXxR3JlN5kZNJshCw97zqAzOVnPkOvEyvMCVP
8z0Rq+qKuguQ+MshtDiYf4xpnVAzaVD/3dOXBouCqTmvwtlBGFocCRZ21TyBEHnu
WqBhyITEa8oaGRMsFFqX6ZZ7YQWP6xkKJC6G4Z3ZbFceODDokZvSDBYGtswqEpAN
Mjgi/rjAryRUvIxzx6SX1dET1bC6KVF68dLItDdk+WbZ0Wk/3fiTLzUsaDI25xba
vtnRjR+CFcndlJvVNWGeNPLnHSQ6v/tCFb8h/jR7hNe+kEVqnhNnGisSWuo4Ehfm
zkhXK8DSbsyVx+02vDW8eJXIxJKTjcOsVNe3YejNwAO48/ooK+vLEvnJCttxlKuZ
jJCfxmxjuheJVcgRt7dsvClXsgmMZmhnsmx8OlyTPZQaXSnboyyPqiagQis2Ddkv
J3w7m/bw9fdC3vLGX5tDqXkjG+g5bbRn7Sv7zjG+Pk8AoaFg2SSQQjNMst94qIIV
mgNJcKI6H6l/j6/+zqYcvFNj/3dMmzH/1hhr7gIpta84fFHdPHnGGslzIj/UIvqK
YFwesXQNGszxH2eI6ZMzdV8f4xueEj+aI+HhD8RJoCIwtuPgyi7VjMwI/ol9Zzr4
YgzfcmJjR5OhwPKPvYT2PxfKh/05hXXpl4Lm+FAhg1WSxCdJnCYkY2hEaohocQW8
zFONOh1nK9BBH7J1RVqO8Y4i9Iyhj1RN7Xgk2qQO0cogjr7x7MiMAO/2pLnlbJm9
5rGojdCU0+niM6MpYbh+PkzrBjoVXk8x+ALOXcS1oT+z6xaEZK/2bPFpzfc2DHY4
ylbxRWAkE1nqkCOUVNIGEdTTk1E5ISxngCUmuLdYlx8kj5FVp/LD5pnhRpDCKPKH
opJMmPN0LqzdClWziWISPz8X8EncFeim8dtGmzs57/B0QJFBQmPCYF8LK/iYsUcq
cHaJ4TfsUADL7T8E9/FHzPs+92puPXu+sZQP5ULOcL4Sb1RJ8f7MJG8P0MpAO9/O
kc98ECel0mW8XgvcvyO72o74zfCgipuewRwi6ZMmcY/PehnRwB4t5Onzl+wS+RpN
aFhhDUsfWUlOHsARp276nSHcQqtMVZCHlyy1Nk9LlLqhq6zcs2bVerF+XvOAZ+bm
d0UYJ85p6xnHhm191eWA5dOi9XYy4+P9Sk54QBrPodzjz9f0h86ne1bZ8147XMD/
XG6ETkr1+PwaZ6HwJqEUfb4E8gTAVWtH0mT1I9PcC1RrDlBRR7fqhIgXzDeVkxOX
Qx8UE346IR4wQIHl7xxBAJdkjA+8P92ACJHsuYWiVffN8P8O9fBevdhIWrpnfz5o
PG8Mwguqy2k0/VzS2g1ld3GNBCNHbHdxkZAlbrg2GzsE9G6UQjBml6yZ3y5ZgoBx
MYlbR9gFXvKPLKXCej/xubgh99+Jl4BigQYGvCa4RBB9JW+jbbE5xXJ0H1BIAZqP
DD0c5/zx3DO2cSZvudaym0J4/UvLAtPuNBV85lmVhaoxJP6mPlRsDs5hv8kOtyGU
cWaXfNJQAnRT0gxKlv+5+wGba7iBCiKxKeXSswWPXiB9Gw88jvEqy/f+Pvi1yiLc
EBo8+SKUXqLclKk7bRBReJoQWUMJl/2lNWyVYcohIacT1CPcmKa93O2wZD3yZkJA
gQmcJVJERR4OiKEualQjaBcJnTBWNGgFTSJN78ekvhmthAjfgpahFKPu/pFETphV
Nrs6iJoBTM5Of9d48KnKzmZ6RR35dYtCy1ejMpFK7FzHkXvmj6fR48IRz/ZAQ0oK
hktHM+oDDG4EeI1nuT2qs8MvlaabU3WqQb0ttRfuWrW5VUUfI57Cdf2XH6izQlJk
HqPAV6AsBbRXmoImeNDzSi1BTqEMM2nxxjgbAwHDXDhono3thnPek0IGYSgES8bO
VOnhPiZp4jJmbQfQiCln0NFwEkml42f8ZveoCBaG3PZIDnKq7KPoub/EYGIyrvuP
lqcZOhtHDzi2ENxBE9LSBs9BrURPXxsv7nvDIO6z9niGU3Yo8InBHVOoh6tmxMTn
2oJCkgykVQbySpO6k/69bekX4/LYTWJwpMhIeERg9/82mWZn9ZbRLxj+xvHPG5it
8fFMVNuUMDPoh5X6fKhAIwo8iLmmy2TNiIOySAd9xQZgfYfWxeZRBWTmDUg+gdVl
bDtZSW77XxN9w8XNvY46DkH0Y6XeyNvoOH83hxnFa00FfAmSrR6qfSL4f2ueApP4
ZsSufFlFkVG3OpO+6PrvoDTQ+2F1nhaA/bgFZgZ654Zmdh7035Xh4sNCDuWydcyz
nhc89lODPLU3PIvdvgmh4zjbwn/8GAupNE0C7zQ1nCEk2yHFq7Iq/uQvtSfn8Crz
pC/TnAOTfTj5G82VVJQf3vmWCdeCEO4k4uraV4Xie/m7y7tlhkbEFPaKW9UMi4aP
7L/dXdzwtO1OqtZUIKvFHr0QkX3JM9GX/dyFLImSyisd/AvVKWnnjO0nUeiKlR4n
qF2BnFayFwmyKa9TCZrVZwh8GMfaA1qweNRRZhizgQDZs792HTXn6/Ws0CclDHkY
8w/4oJXY1REKdkSA6n+iP5U+E/NApJJrDrQOxyLYn3WH7jd9R2DOVlZu03Y/Yt60
4HIZ5F4YHKQctEiFOdmF+qyBf2X3Ve5wPn+LQlPlUIm8DnfZuvh9nULHWmknS0gq
uCHUuKTQeiZ2bAxoaMV56Nk7j00LuzzStAhYiAV9RFPaFkkptTJNqHXeb6tlBNe2
EBl3ybcjxxW1TLDbnk717+i1PpFRkoaJeTP9rd95+L6Hi71qWRIxPqVkw1F/GjIx
/WTXPnWS5bWo8/+GWGBVC8ClHl6Q+8kHZYzpXgDOSm0Q2Jj7xVhwZA8sNaY9Nwn4
DlpghBGtU0WoSmByGXCuROgB/2fLEkn/enLNoAKT5ttxVmfWkW7MKg4ewVzvHoUh
IFsiruRkR/z0JLcJmknCccDwtI9eJEv24R3P1Rm2I87SwPk2KC4v+d/23WhGjIeB
6XJ6GO+ZkRjk6Kye+viKiB+0s5xZHle2+HmaICPBuLZnohPvEwiu+FnvSLBqfGcl
mmEBGRys4DLwfBApKd9XPcAg9CwJcbXL2ZhEFiawWv/jc4HxyumZo/cpRHlAW2Z2
wasRGYEGlHlFA/f1v+RH52qq/RtRRKkdY8bZ7chtnybSLn6T1NVicimmATq7GysW
WPaf6TnldaJgB/Aer3nvzo6tqBTZnZQf5eNZFv+auHiJe7FszI9/V+UDAIjd/iYd
FmKrvKG6X72kDyUkg2qVAIasDBF01K0ufpyvAMnEx/z0Coe4R1Z0VC0PM8S+BZn9
07hb6Oh/hVKMVWa+y9stZdpFSul0u5/mibSd9zIWhzGNdlMfLIvBLhSMCnqVbGWH
AFLZxVsV7X7KZiwemi8PX0BGvI9q4uH/4nJAAkn6HKiQdGC3gpcsEu0boXiRGiQ8
IxnAJl/KTHnldlnvAWTDCSphrMkJoLG0scxhlYoNTF+y7uRuB6uKRZGOnoS1oQOv
EiuHo89FWQsFTQlyxi2D7zm/gSw0ypC0zaExeRR6qTiZ4a7+99Rdje7/59N+z8Lk
H26vV596OtHNtBndPvkBwdYKo+PfoVQtt9sCdpkBHeU+0y8Tc0YZ7mt77skIbUFu
7A9uraqdbxKrpo2v/+uz8/JQlxqTrHsXf1q/xQCF9oCaxiL0I1qdHyCqsU2SiXti
TIsXQhoT8Kt9hJC2bKfBx9XSc3RQdmuHTkGa7ZuJyEU2w4Q3w5YiTsw+IXqWkVxp
ie2cAi0SDy7k2uL9n/x5V5ctQRm4thT9mmAQhoPPCl+kgfW3TkKn9kcc+t8OTFqF
WY6N1CJ8sJzoSsgsgnw90kQFLSXrVl3ZJEAOYDAAkgjoNc7SJcMoNSrgid31x9De
0IEmIPhCq43X4C3AFAUz7Wox33Bde4aaxRVpjIntCdS+mRbzW8MwUfI033JCNTHi
GOl2+FsGr79+hSMPQVRB2uTWOr9qO7Fu1qj+Te0EOgDUqMt6ivd0VqkWMilUI+5e
cMRsqBRZzvKtvTkjzWtgyxlFii3FH3x8GRVpP7uUuUaEtbY+jyBHT5cyugs0a7U6
PFvjsvT4C/V1ORMtE3UU0CSuIxzW6pLLwV6dRKXvM2Oxe3rjqnXPyt3HrrSf4asC
N3ynD0SkNXolhGru2tolSUQ/mLDFwn3FGvuXUWc8CsDOexy2ZwvbSXon7jXt+ADk
qFoQIMdwTEal/Ejpwaql+iE60nnGwoYEiVs6/v3GGp1t4ClLTL6TxtXgr7ezexp8
2V+L414PPDP8Q2MuAPfefBKhbDMRxy78mCuq7ucQv01iGr7VF+ge4sGkNnQ08IG1
S48v3xk8hh28Q2oKlf/boLKb9Bb4txoFLst2S0hY/1rOY7cVwvrvLqAy1y00crcy
ra0QFnikyw677T2YVNUrj1DiWaI9v/UBK5Yan+7B27mNylkL/Dq1Gb4Lrp98hdPv
HoV9bcPGNxpXCoLGVD4pigB75QHuoYCqK4OiQ/v1Y22SY4AN2M6Xb5/vZHCekMnK
4Bc0bp4T7FjdJAzlXhGcC49H+T4eDg8QQeZGq/y1aOrBnf9/BTSuTUKRtnGEWlVI
GwIJgrP0of/06brXLbP6GgDOAEh7tUe+VMtOHbzBv9Eyh09u49hHqAP/Chj/DMSs
Is9LRbmWSUtm7smFcX6ojTQgn8DymuVxbBk+FgOlctpPCQJCPStdUlAJWnuZWX33
lWfKVidOqJ6Wn5S37oZ3R3N+8n+aFUJsH4PKJw0IqIv9fBARtqMPg2puQtXOKE/V
F87a9/dqRfCjfpoKmj6QTFF/oGEfgRprqM2TqE2VFHmaYq3MHcPM46LdGu6jEnZg
G3wI/8PIl/6ow/kPJRG73oVnf1XDG+R+lUekDMph/TxiiGoDLh1TvYi6DWhJODZ9
sm2WnBdD5RqVIVs3s9gBHC1SGRRgFl6FbA/oMpZszg1K/zdIRveA1pUva8KB1PiM
rfdYgNYrfMc3F2jIhxYlA9GqrGpPSyuH0b0dUu4/FDx7aBTVzl3re6KOfdmXHs8L
bCkk5F1iZworxla+q/RKpgwogfVpFxAyru406oR8xKc9VhYKsiB1bjbUhy+80Fwu
0WnI0v/vtWxNLQY5kV9SjGKmAHlshB/oFwKnMmjr/RmyDkx7iL4nsi8s5QR3lo2e
T1f3Fn+cm3qYK61SNiDLL+DSFxaE1MhazGNDEU14xolrKDrpa9dyjr8uuQqYFSBy
Ivj+xYreNca55Ig3OJPGL6CRxWhEHNcdk8SP/Cg/f2NG0L+VDIY842HD7Qd+2AxD
nFyPs05TO+rJozsOXhLLPN/TSdAJLtBjkPektD+xflLHWG0yIsXfXNt8zTEnkC8+
VmQofPF5UrQUsSdzBZn1IT7xPAJZt/e6/58fBmx/bf1cOqbIwUNpKvh9mVrreqIN
xMbMoYgTsHnerZP6xtYafbSvIx3rrFgjoL7ezwzu5UbAceqMBO44pAlYASg/QpoZ
2FJlFhxsaSP/IJNSQHa0JelVppJ4DDFPbfht97CpKTasKkoB4MpamvO0XCu0SWZx
3pmFlXu3OHES2XbhgNp9esDJVHw5jsZ30dt0o/Ntj+T8gtH8Szgqoo5WMeTbBx2G
8bNl8sBlFHqmNPuzTovrHClevLlFVuhcu95tE6Vs0D4Ku8vRLzRK/f1JqVCHGOp+
b7j83LSuj4brvQhrFEkIIbb0lIhsJSLGa+l1geA1gNOg2ZAsCRAWuqyu0uhEeJcf
2a264zpPsYJsyw5athdvFB+o9ELXQN3HewLK8GHQWUVLZ1+zPphJ2KrJGUBXiiRZ
bq9SFWqflblOAxhhfbyxe1Rf10vsdrKAC3MbBRPqns9TBcChb+9QdLWa1aNMyp0E
dDszeWhSnWncOP5cXvH2KBbdTfFlNyB8/nyKqMUEXADJB9FSszqf6A0UGAWBr2BL
nMMpcFM1+JyRfRGQPJE8u1FAR/5oat43jkwwvHa02uZU7cEoZGY8HTjaOD9MbAys
GPESHVfBq/EOprtGxfZAIdi1SEpwzugoRMFL4CAlPKSwlF2k+AwGQvjMzcqY4qjb
F8P6Cv2H2yPueg53qQYk4FyK1Ly3+QNFBZmUh5hUDne9SZpwy5a0t5oQdwm2hjOs
nTu/hY2vqOEE70QPCAVOmffV6BDWqPZXvlds+fhrjE7eRKEOja2aPUDIR+JxsA6w
C2690aWJJsnwR3f6CMzniVdhwjgrLa6AIkNu9S3Jm/s6ju7gv8MEt3oh3/bQ1GPM
h2qc2m3XCzQPxbXbCPKCBfpUWnHCAW0H+XOYpCOXFn+Jz5VbtaTmdPWiz2gBKdsa
yFDhj6om5+UCovV9hiF5N3d8YP7L2javz9ymFQdeKUZJsaOdPxxsetexhIbadPMv
fXLfmv/SsquT/OeBflT6unwXlwM3lHuE+DjYEugmdd9yesu6An5zkj/JFyV76APT
g9jezuQERJnFnSkknHGBt0PIqy5kZB2UEAa40yWg3l4UAZ3xZL2Rtem7HhV4/kBb
A4eXy+pLFvP68YnrkmYbNVs5IPhpFvsQK2HYk1CCOyLR5CTGKXmVKYg8ekI9J/AL
r6RJyT9FFFSZGrKDqk6eW6mSaoqR0MbFMJi2imYCGAEr9W3/XsbWdVforn+1Q4EV
EKTG/or0Vf2y6fZtC5sQ01ZuOXJg96n6gw1Hrif/bLAWTtR/rmP9KgjPXwsvg08e
bcJAJc97Jh301Wxh9B++PoprFVOwCoVA9lzxdRmJFj7W5cKLI44+iJL8zk0znwLy
9d+Rlz6YxSMHRv4mfz9vRJoJL0rfHWTehVs8IaIVHXB5YQlkamge+oVHlCBUsghY
uaPNleXBphQ2uqbuU1PpTNCALrvIEhFUC3aqitPqcNVSVNzRA/ZWO9XVklDwhr4G
uZYsVg9G5oW4lARleSz8oyG2ONWdqHgj07yDhGSwA7e46HPuNmL+c0bGXeDXuH/n
u7Az5MttFxuM5oKeGPopFfkAQQzkku6n8IakxuB7wWhaA16b/RvUYp34jt5sx61e
c6Zw8ttR4EMLGXpsXbPLEVk+9z6Z5TpZ/SbwRmQuRv+tET8EOEWGnQDN+UGcrGf2
IOZ03yBAgtRHpX6K4sL4JiJszEfaJn8waiy6LBY6EPmjUti5ZBPIfjnmdnZLjdTT
eLA2ulYetJKYgN3WYvdq7v3zEmmHQOB0Elq/YU4b5f/aWc1MFdzSOFuiWG05MkSm
ofnU5igGDoUVq8zQbU/Mwxba9OMt7EXqAxLKOmTUHeFW6HwdIHkQUcrixj/DF+sm
JndojF8Vq/K1VvNT4QOkzIKwvA7724kNATRUKBJxnDzrk1BZlcTFdqEq2rX9IulS
yUF0rkHUbKG7Znc4vkqepm8u6ez8UYTtaVKqnuksQnVzAb4CyjpwGpR5j53I4nD3
wEC2mfX3R2FwpmW4f1i5YYZrXltU43lCrHarh2vRlak9a1S3d/uFEwqFxA/M0iBI
0ecd9r9JeXG5Q2xyG9QCRJIf924sj7V14c7EpyU1RpwViZsQBVLaT2pOWxrBGOUH
l11FEzmm2Lz+zYDQckmRF9drAg7M6UsrCdgp86AES7/utb+ljh77OUWVWYIFDBR4
ljP4WDylj6hP9HDwtfu+iA==
`pragma protect end_protected
