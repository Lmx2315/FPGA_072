// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.0std
// ALTERA_TIMESTAMP:Wed Apr 26 13:33:37 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
FRudhlU++2IAfO2NEcMRNaE+aqo5m6n5JfAHELUIW7hYTt3Ky5pQ/53LtVrrRjN3
6E2xrhuLl7CVuWenHQqAV/kqJYKhvgPx4iKcreTfPg0XBrZvXdqS59h8vsPCtUrv
ldFl+hEynB4AWu7+AYXya1AX4vZGk1Y6XfxMxljE1qw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 12432)
Im7EIPcXtcrIL3/pewsrB7ATR8lDssAsMrgJ5bdfP1mz+tmsBHgfMuKXZtjo54m3
VPEqiQmbZswzpfNDFZH1SfLtkpXLQSgYuWf6Mgv3q2/Bpd/LY0TDNeWMAg8upYUH
85jCr945a2hRB1QFfiBA0ZZSeleauLnM05l9q+7cNA3YxNQRm2ACMVBKtH3rZqTl
Srl7s5ZYmP5ZV4rZz1XxPhJBnBXl1fOnRMd2f074odH8l2D+r8s2HP0AI5XFdTMH
DyoR9+L7IQAQgw5SgXpoOYI9yCtQoBu5vOIGIyI1ZGyk5cMsh6MqsFDSZWiwOOFs
EpLJaSv2ptOsBWRwgFHpZipTVJeROByQFb5WarkUaqbS9wevx/GHvFojF6TNR6Ve
0rWfCStoiR3CMk3sZOKvsaJ6ezL03GmwnIb8C3tL/lR2vGIbz+4jB4bfeUw3bDos
XMyJ4Qf7NkQG4OsoxiUhkWbxZG/6fPukJLNsNfvUMH3JNKiloMu/ec6NN+gaurfk
tRfJVSxzugo2gsS4zliODDIGqqE+QwKNaRlnBy74Xha8cDsOpJ7f8wlg4UZlmeHZ
T53pta4K6EQPlV9I5fDDSqP8aL5cFdQpK1vbVRzmvagGXynEYXwCXhbmJaxtbvI3
uQe41h4ThQdPHAKCstfiRugdqvE7AXY+ou1kYrcN321BYxLkdugVrwDXYwXemRRx
S5w63jCmfKotgHz59Ci2vlanf4aXlz7llGehfkN/1Q/fI1sWv00W7ENPDBSoLvXm
XbR98ySilre3YPiArdBa2cel1JhMxsOKy043E2UzbwFQ/vRkVahMGBHwLNQkGrbS
7ITv/234nONHN+huGQWUrYHmxJQ/e5j8F1dYjUa/rL6ebzNEESXwBmxdpZo6lP7J
kZ+V5H/hdzgrI14eRfEjfT04LoRhMSYCqmIAWS3x2dGOc75YvqU5foqC1VdzDo4s
P80PcnqDZ0zEg7d1XmRxfzY4alvIvWb/cs/+h8mrWIF7idGiszVdqBbR637y8n0O
mt1ihVS+Az9Pfirmr4svAxfJapvlce4EJ/jRyMcY9v+DDmpdlTWvv77JZdXlvAbd
FOJ383aB9N9SglJh1NAtnYN3ns+7InBKdgy+pKg4NKaSGqJ0B/716lnLGvLFkfB6
i+iS/ljdtDsaivYyw9V09zaJ6zkWeZ8HSWr4ZU+EjbY4MRjMzGBn2comtA6LTTYN
QHMHnYmPmoP4thzbgbak/sa3tr+8yIoEInbQEo5NB1E3gLQ82h4VBT397s9ZcD++
cThRH/x+uK4VGcHQI2bOG2a1qlSAn1FKF1U40yrDj3uk26REYXzD+oXWan9jG0Uy
fBWU415KCGvnhm9yAD3/xZ+zPYTXFX8rJEzeBmTOKaqMxnKSCpNDLldcvndVSrh6
VHOGAbU4WniVtdlHJ8HHV3w2LGPvyEi07KUliytxwHYunQ7XkVPk/McK4ljw4EsV
RLuKtcMf4kzXTR//XVVtLMoFS1nxLjZA05e4LBQKQAYQ7jNWJKShYOnpU3z2+Ckl
hLGckuA9jP9EcbXgSvApddPEShXKiwHL7336kdWDZ3H/YWgVfvrZ9XaSNbl4joJz
apw+IqO4Dr1wD8EoBztfCwqTXoubAB2qHTZf+WXRLdjl/AzO6m4LHrxbkA6cNTZo
6LkpTVC3UQ1V5pfoKEVcGAqmkV9TtQtdUFAXnYsReL0aqfrVsFenpogjOeGa6LtK
nOu/6a0F3PQ5DLamZbG6o+QNWDiPOL4u9wMwUeXI7JGq01RhT6dQpPc1+NZfGdBl
GaYiS32L0zQ7Qocb7wZ2kH9JU4Lg+A/158p3oQplM74qBQanX25tVONqzXvLVCIN
w3BHQF5PFiy1upXgk/lMC3x0RV08174aZ+FHJ9YzsRfhiweV2dxmt52ypOsNYb/C
FHkKf9kpXJJ1oU1CTrAw/IFZq/uK57f/9r1XpBSTkGoOOLenLxaPWno56lS8tffP
N6o+NnEtJS36I/P2vdBlYIUtR2BQbE9HFF5X8pBlGlTX8jvcxyuJl9BQe+hdXBHi
6eNK5dYklouUNUEI/5JHbF+8tqKu1uy8+3jpuQqOTL6s9Kg41+TKnlFoTyhbrkvi
2pD6neRL9e3k+1G20hEVbMUhIa6IPRtDu4IOtvyabnHuJJ7veXUNIKAv5TuL7Vlv
7xBjCIb98CFfuimaSO2IT6LqsTN60jhey5PqYNzBKTaIjVy7vbriv1pOspGF50Rr
1GhkoHf2Aq1y33u4X7n/+hAqdeApu6Ymz0ydvBf+GWGc0kHqKT0PUDTSiJ2/qPbx
fuB3jwKad5O8hBcgcK5vT2dY01s+fh9bn2/F8TLxC7yxXsx3nS8VjLHjIv5q19Te
wJqShATJDjKr9tIlhbh6Ry2esHolXQyyM3n0S/ImnXn6v2Nw7CEN3BSLR5esBUGv
EB4LN0Vy6i7W8MsI3pxUDTzMghXBSO0LBwILzaDoweC8zmqKfLrkncFlY/fok+J1
yfpd9LOHF2YwserIgylrOUjGWppj3PWb3+Bz/1izfKeZvT95+9mV6sNDpPZ/+IQI
ytcy6oZ6NefC/SiTGfFojI/cC3wsgNnY2u6hCyNijx0OC4zTy+Xno6ocR6j58i04
mc5hzBHdECsIkfRveLXcR3lStAq/pUa05H3oVL5QvpRf28tamq9mIzU9RKtvfptS
2UXJN2uqCE7Geg/jHBQ3mXlgHSWy9YH/T/mA0dpIRUhyoqkieksGdJSV7KftZjP/
KXnxNv26JkEzhE3VTqp3vxbbKte3jqPJMWQIsKXKsnLSi1Hn4wn6lb1M7qmmf1r0
OFzshy00HtJ6AdDUwPgFjryD7LbobQKxq/LlcPqANuPuCvrX0kqtBuDdH2TiLgWS
KNoPCS496qnXGxuU3PFzUx8CUIVbDXJedR1idiNio2mvwi63yoNF/uTw4FGi+yVR
t/slWk51kAq/k1pJGPfXkPRYxlDVKHlnO5NxG0sjRtjSzdpGNKNEp3VqtV+SujtX
S8HcHkWYum7L2022P0LDPeMoy5t6wPgrUwX4iR+tA725EHYWYrJYi5HUsNWCfXXY
jr6pGQLBoqx+BUkDKtxqCD1jq48VXalpHeA2NmvJ5VWtB1leFr+SKwK5BIINbtAU
yJNPV25aZhPo6Ego0tqSA6sfIzOd50/QgsPGqse9GDihgTtQirDkErTAZA8Z7e8z
3qBkdF2A2SkLQsoC90Npv/eFJ6Z8dbxGcINqc+4yJQriPFFokxaQFukplPFm9jlY
8thp2Rkc585a3TUv4z9GtqDIhSLNCIN2R1/PRHxxoIbzD9XXSyKyEPW5Blkd1bWW
3WZn2C7CYZywJ/Zq+SpHk+IZiqSdIZKBwuf5HapYH0F03RCHh5jJs4gVWogO6zjc
bBPzURMgsiMM1OA0ISkR57qahs5nPrdBm8mGz18gQ+P/OTvxrKcKVUexpIvJlK11
ekX9GLBDSks6rubjsR/FiH8IgTVzD1gC1hJDHWZ4T6a7IZCXzNBLlH3Rs+yYpvpT
v88N6hqeJJQKw13cF2dZdGRr0eHmuOskbdt0ES1DzdVxMyqdXnzzZDgtdTG1aEzW
m0JhIqSQUgvk0gY5yUQE9QO/NG18OzQw/eWeWXJxi2PyUfqe0ewOjPXYWbKN8IDa
HNPFbFdolfwfmc2kQPjS99Hlbv8tuoFlgVjcVGJP1aPkA8cKvA2JUgD76pd0onmX
fxA+vdz3FywYvrBHVXhcTi8JIM1u3EdWpFWNRpr0zz1FHzlZr0gHO3MhTkDdKPqZ
dxeQ9gOxl9Mp39Ye0as/6U0AY0w6+CCyW8CSlkhGSVle5OUcuw8qPFpcxTBmKiPm
S8qrpwYyd2dqLssxtI1bpkz+KBVcxBvY9PbeUOYkULEHcqGs6jCfsDl96WiLlkOS
6GfcWOn6hmznvdVbtf9v5YgtE1rjCI4sfAkFE1Itc6/8k+txGY4RoQ46KZgHRMAK
Oz/AfOi9KIsCn+Olj5PRB63LOgZNrF00VdNIEOq7McEBiJKU58rl0GAcOgLaIKa7
sH4s2ifAXdkE+CAQRFQNkM5QTQGo02mdc6KNePBOakCCc6IayUxYbnFE7e3TUtHe
5oaJFud3rdwY816ivrnQbKXeIyuU/ag0HS7jrp7XW7WOFbcgPJVU9mJXiXsS915R
dz7c2cpD6odJflLU3rv6UugCKUmGJL+PtHAqAarVZNZeMRVgnr5BbqZFKIoW6Xq6
fT83RyTd7e+2Wrl3wmOWDeuG2RcWYR6ZQ8XXMRnvpNjlZ2nhlSHZ6dWFzNRiXXNM
t/H6KNOS+yAC8+tQpT4gIGpfPSm/qrjOrICojUT5DwyUbp5Grax6EbLEBD8Ny9sn
Nm/YF+Fthi+D2VhCqy2hq1dnYpQy7JoYqQ1R6yOjFqi6lGg8O2+mzkNTSBOSmzGA
lIZcndsjOKlshMoHSYXK7hbv34pZfpSy1blhQTKCJtTDNcrpiYU+e5MYa8m7aWhq
i97CWV5XfcfevV7bOkkGfbTCC+KxBVSan3Qc7Mz91v1Fey9C4VdgmjDSc9sW8Yay
qTt/OhAxTtF8p+MSVC5jpXHDrTOcZeB92EHCggYEPMbyAH9s2qzvXvy4PDmVRn1U
X+SkoSzg6jrvqCuB3ooghT1rdUjDQpt0hhcsoibwb8ALcRFeIlH5CtLZLUhy9BUn
8G26Hrz3rzGjuvNF1vGlJ90X8unr259XAqPmvSFhRnQxP+DtLuXmyrcC7uZYc1J0
FdlE/9+sgE7MO0DWBTwZlm8zfJioCnO/rBlihr4swt26wkLkYnnP4y0dLg+vf6fn
9KHGebGVLvNrbI0ToAKutnV6iKT+4OX/pTrQlQ13RrlJtxpP4r/GDBiW0p2/siTo
Df+s0uy7ejKM2gwXpQrtl50A6RlfX3wMF98aymWvxQDKMKEZHBt1vSJAioJXvvYM
ebufhCzCxA/nRwR9E/Truf5ypM3Ber2NJCIaB8O/i09vP2QEllvtQiaR+oFGzsBX
21NQynHmbv4vSesa6VbFdBAEAgtvsJtXW5fhQra42hx8p2R/7s0r8qcTmu5NoUhO
aLx5Snr/imBljY68ZwAeHK+9GkYtDzeyRsgUjWthyCskgfyQ9W16+pOM5Y8dBrhj
sj8IqFLD98E0MBQNmsHwkkiGz85mlR/vatGNgiRuXIE5e2evbGQllxvwX8DlA2dg
cVJbcmcX/4YO2oLpt0w+yvhdBLn7ytH6Z7HH0epOSIIvXWtO2ERHfsDHnucNbq4K
cNWuV1XLCmnAGWBuYR/Ar2tFOdSoQfaJ0Vafs/FOIHE2BUMHE5P6XrYOAQ+pZrFr
sa35VTU+EX+YeEeU5Q7LL0v5MJ89bAarAPFS5etg7t07sv3tNJWrNz8EmsVqQx7H
R2DdxtgvZlgXZtWYneaDQE8EaclHPo8LT3tdWZlZCJCGi3eCluX95Hi61hxtT44x
e5z4uqr/UZ+PiYGBhhHn+5LGCYq98JIZphJuv+MmqFYtiEc6dsaRzmiMsjKocTdb
JagEuX/m39hkwOj9hpFyRQvthelDDhjYX/COg6n+qnRka1AvVjZtyGVWZzhgQx0F
uO+gKE5i5GBhe9LpTnMdOeqUKBEHdBe5rR9DdU/juGept3iTi5K7EWjbJB4A7tKb
6gp+FzlCMNv805+xWPTCtyZ7eqXz/lGrLODzNxIcuQqR1vF88Lz2EMkhNq+ddmg8
T7DTotNFI0tCJiNof9DUO+iMpveXIaScQav2AKdh+BElxQ9PxcGnktTzdAelvcCr
cVx3k+LUkMyGQMGOJxGNAbDx0eDcLesUmaKgyzmDXOpEgsA4GxJjW88Z6Uw7X+T5
TeIIDrw214K8xzviwQXJ54n5yBivNLTIpPBM7kNw3H4Y9drUwt7jdONodKa+Ehvk
jjyggxN6zFU5Do05dXdnhWzAJwy5qiZaKCpOJt9sA0+u1aL0t86IHcYXfJ5wrUZO
DCVNLUwo9PsyfpVskiNzVCH9HeSjoRVgas9iatNfFLJUQwpBxXdW6XxbV1PLrWId
wU7790lPpxDHsunFOCr/1pYucqWBz/mEWfgROI3X8Us2R+G8lJ4VZTL5sOB6mUy0
Yjj3x7Xl72xHbhVKxJ2NBzgTXZtTN6fjeDtKpDyNmiDGPEQFjdHzD/9bj5H1WXDH
9z1bIy5594Cw//yEOyLUAR3scXQLhMAbOZXpCOyttNcO/rvsWyRHwIkulEqO1XRE
KPVcllrJjtJODJzpe46xVIMOgyzU3xkEc3zdDDw7rerpEyvPnKH7EuqbBQS3HV5P
CSC40BmhlrNjHPNQH0dHXSC9hBRQdH3mJNcYeRSCYV2fdXW8RuCCub+We2/llf5V
FPiuowVLISQN4bfnJBTekgQcOPxmNfGKcuXXT+WHsNLPt7JtGDZma2OmVeGDu6vG
YgGg6/kzYDYjtuONRhLAD6A598dhX2yrU6gPlOlzcX9b3WqufluV1+AtYlvsILxP
eWDYj8XIVZ5nlZquwaWyuXCIxJesEBzMqFG4a6QhzBuE/mzd3hSkMsiFEOmNk1xF
iClmJGEmG2dUGtC+TrKpoDSNqjthsuJKWIEHdQdxYuzJsZNViwTLlTY5D1mqiUvE
DAFA7FXcsW0oLZH/Xr0TSJVGr+zuJB2fh9oZHSQK77wVWX6qEvKe4+v8HZ5ITsGE
jQSrVoYa/01pimaKsgxFpbd2v4EZs64sUKdlSezmlsrRyOk18wNEJcMMz3Ap/S/T
vLzktRQGiDCGib/MgKpHjPZLzlESQOIKnZnVEiC4zDpXdTndC9i/a69OfSa2kEcy
sUXKxDrj7jwc/Vyunk5d/55UZbaTfzinG0b1xRwk3xjpevMecLoZB8OkkgCIdSDP
GMPGy8RvMZvJpGVIl5t03UK+/iKNPrcASFjqBhjtOz6TV8UGmTACb0hxcRC9z8Qo
Oo7G99XhSOK+8FwHdgPvJPcrk+BaU2GA4T7m24MPdtvz+qQ1qYBXAURE2dUZnEoR
XqZXZdPrtSiOSyTEba6qHPvP8Az6IZ07YKxg+QiY4uR/vJg0xuXrSRHC+6zUpVa0
atfr/zKyFV1bL7iDEjKYQcRYMEqJ4H2bKBlFTLoRnGt0cLWrb8koCBEpSCSyOtj9
cYDowoqOmTxlWHLWEkD0MKYq6lD9TCiZSeCteP6bjCuhX12c4tnW0oLM8K7LY/lL
Wi9OkELGoEIJq3PbOsnrq3Puj0G0WJ2Si9eDxR5ZjhYjWnof7sjBBnr7NLw9b8Jb
QYJ+EhfhvowW/esgJOdZxNwEJZlgH5FkRGAqmX8eaQyzDMt9kUP4dgbMO2ScUG9X
BBLtws4YpBM7WoxfyE1bEYwJmrS/gcUeLk8dple6UbCS5FHbZRXhFEXTpE1hNfDu
PgluefAyYxn8Ffa07+xvSjQrQt7EIBNVIdWjsbOW0mmuS4j8TCpQMXaH7NfwlyVr
2ev1ty5l27KrAylL9kgLad3rLe+lIeqdy4OQ56q8XrZgP7f7td0XxeDe1FsedI73
TUGbOZKTUmAbERD6AUkrW/vllj3nEsfBqgNpdzl/pj68VqzDeJ+OmXnBBCoyB3LR
pICO6lWmMYQA79eGk6lsMvK8ukwFo+xH5mRy8n1AziYeDKZPc601MrAVTkrQ+Xx9
WcvU3IEzb0Mz/nMUSF1tD0Tsy76tKYLdNlQlkcw6MB/aRX9XpRiDo3iwM4voANNV
BVvbcH6ZaJsqkKMLdukUCL2Rrn/j+YQKMTzkxm/0iq6PDs09k6DwOB/rPyp5Ewjf
5SWvLqW7R5umnijkgLIK4yx9bdu5EMlQwKNXbIY4gEpn7ObUDkw6pGfUTL2+BKuF
OHWEDOu3YhF/8JTwhKVg23LIyKtCkSOOJdRN4Hm/VTpeN2qRO/jHEXVDgkAbNQLg
9b9ux1IwCvKN9mJlj2pEyMvWPUWH6KzPj7Bw3kFj59rKG7M4et8mie6w9isbXUUT
fh4z0YGvrWd7Jtc1xK/ItmP/w4CG3bA1H7xNq/PYp/dkrb/gZndVV2efmpbK4DmD
ghb96Qc5Q/3qaHgENg1Alsjw2RJMYAkWM1RMLK2qmFbUexdUkxXz9YDASKfo/q94
Q8OdAAA+OE1pscZslfrvejzawmdz+piIuxKZPXbaaJWlz16WoQN/So/z7AbBO0l1
7bj+8WRlxOtplQ4iugfhMLYqJaoI4HMXcf3Ft8pnJeXZoIKm8tvhjzhBjRLvJejH
5biSEsu2Mcr+TNQ/LoTeXf2OV5ciiW05f7hpgkOC+LMJi87LdQ1+Q+u0RwLI9KYn
aGz0y7QEDFc4kHw4E4ReU3kQ7KeVoku0f+gXvGNAIJeGtcVvG8R54QwlRCk+Jcyl
4+pLqu3kf2uVObMPjD8PgAtrFu97/iT+KufWK53s/Z/PKlTWbedbM4ZlzNOOwK7m
vIuLf2uYyeqKoYrwjH/M8/+DU4j/Xcmi5HEwImo+UwabE/I2unIcGwMpoQgQB/EQ
wN+FQ0T8BNP2AlWi6UBgK63DWXPczXb8SesfgDg99l+bNc9WjeOjKBsophccxXq5
gXq6A6R8Lc+JyfT0iDkjhlGMwi3g4DPLMSZfBhxZQUn+Tw5eeWvaDGVSzIUfdwYS
t87O4diNM8oQRoFpf2y0Oma40j4i/R2uY0nEb9n6aShJAy/rS+oGKrIZNSe75mZk
9RxjVmfewvnj7jCvH50FXF4EMGsuhTikmyb6wqQ2bx5lN6AqsOA22whzy7NJ+qQL
NZRYTtr7GPBNg43kdlC+I8eJP6Qyv6qhwvwYn8ny7H/V8NZnwzglhPYL1F7wQjvU
Eb0zqTiqTUjfwtnZAzlPCvMdFIIWRd6qIxv6hGK50bublgIdbEtr0JQOljQ680Uw
0EjhIy50WtrtjAs8xbeS4VMRmKWwq0XgcJTX0u8kM9f3XffxVveFFNUSIq26As7I
KzB6oyv00IuD+Yzc3CK/r2R4RfFAUTbD/cJSIpecPTvcpHj5OOvK3Yttg9UoP5N8
3vy+gavR1YCrK6aXxgF7WmjEzpS8xV7G807KrCRT0SBvk6m99yTRPp9ro9f/xYxw
D/GlL60FumBtdcdjKspS8U7icGY8gVek6R5SHqc8dP7oevYBVQ9auyWn7syxBiFJ
WghGfgkPeM6n4ahRmX8cRQGf+EzJqn3i5mloqg5WhE1VKcgBi5hgTWQXsp3aZUHf
NaUW1Rr5U6jVfjYDvXpB1JZiF7MiFLPBY7kMWKHGnd6iTkgEbhNbjdh1ZA7mz3IQ
2K22XADqjblX4p2Qt1y6N+/5WadWVbah6Ei5sr5tR+Smzu/c/kTYE3qsieubZy77
JATRLy4eygI28aRffP9Z+fqy3qBe87WXbJc5RmM4chmu474XnJJowh4KHBJG3GT+
akTJG7RWLz7ZevHo9rtvfkL/Dy/TkIOxElLWy0Z/HIdlnUja1r96oRKei0JA6wUh
4zq+PDW7KEBwMXgxTE7N7nTjqOhAtrP5yS8qH1eq8R8m5HJph/WYw7de+ykrz87L
C/XUiaVacyy0YUpxBKV3BEOVPpAHvxH6gWBGPCT+8oR99mgjKXlyuUpvIAahjokh
VJb/eRpbvX0pnkhNFLmIaN51VOyowRit5mjr0NUgHhlrREdKlFyeY65szxGc9K+P
Rr1A8snkQ9dmoZNtlM21pCMhzmbW0llul0fM6fGRM8RxuCuwAITvHKG7oQYSPnrx
T3G4eIGQd/grf3ye3u4/K6rcYqN9Zaqmv1ICsoKB5knaA+llECmL7mDeA5m/oQbM
AbInOqZqWz+vpV2SV2JPGWbrLtcS6Mx3KHI1CA4pE+XSNttrBXMv8a6c6EkhghVk
t/Hdhpwj06TxB+XHfh0TGR2DeaabRgdm8nbjbiJNgEyX8Hjl0D/m+ciZYMFCPL9t
TL9XfQGV11IPCY9TnEN+yVzGAGDAVu2eIWa7TD0//eAIUXC6dg+oEpli5kq51qJ0
ajFobzvOUH7apIl9UCjJORz1tyE4RyL/DHByslKYKfACVWYTKIHO095wPtyn55z1
+F5YtDpJul5Xh4t/wCz/x4wSrdHoI20AwqW16FX41KSQ2jZSdFBGk7FsuGbs5QuW
YG2bpN5c1nVARvL3pPTfesSfLY91IMdusA4SY6HKJOAiFQcBly2INW6h1RPs1BxQ
4ZKkaw4zwfwmrOJccr2sKMpu09Kz/TRcgdyoFujgoC7EYryaU4RvdDPLownh8gkb
PlWKOYlPYHQhgfHm5SRraedoEMSKf5UIDEcesMY5/xbdswEkL4NQpp9+51isGses
xfepe2q4joRjwS1LGo8b6J670VC1qGgBTBynEwRzyWhmdMneBKzTGSRUhzd1/sqT
iSP/r312ra0Es4oCYT+WNmb7QumWhPRQWHBy6zbQZ7QW/oATL05kvtcguRf6UGgI
h33RLWQIaCHxkU9NpSPpnUXgeami6jMvi6Myzk1yutAkcJmZK2qANkoUCQin6WZE
5gJwTkx3HGgjO6l45eyASo6DJQASYrj6CBzFWNC2A6nj1CasWarSUE1BsE+LoOiy
Q8OmCiZO9xM8rERYBl02iEWquFLWVlTNf0sYy3Y91Q+ZXxZeUdIycYIBqzalNwhi
zP/oRvlYJkr/hbmb4QyWEOouS0U6IMEv0lvUhhy3TWQLUvHeSuLCHvLMx4ZZVd1Q
qmkTcL4MAzfge0cwYZPTExKsQA1MlbL2Rj8eGFD/x2Q/BGLEeIh4dOlfoR9Nhaod
IRaQsdcTFUWhnmhPfOIswk0r9rS4ue6rY6tDr9w88OZaV9W7p4fwlnfyI9iQ4BqR
oQlCOl+A+q1FlMSvH1hrmI1CzazSqBuCot3nFBeMylV4fkD0Bb/olBjRw+UmhwVQ
cbGmYv/VR2yPkZ7tNx4W2/X3WwEO2Cr1UabrX6Ergm0ek5U1PciBx4hZvV45ZSQK
9Sm4yA8bOb7my5vSSEVGcnCWBTZORrrj34+ro7N1ozfXSynO2i7n7u7t/V6igd5x
yN9gou3C/JJaDc8bS2gqgYvHrqb16UVwhzttxK24OdsXmCVArruAv19ZtBnSg5El
M7nPZReN8xzdTZ6E2SUIETzxLcQd3SMux6beZce1QczBsV4njQeLsUDJswSDFTAy
3iTzFukZk0eu02lCYv0Ak4KZFnUk2v6lNgMqVCxZzaGA1w23NOckaH0qJdOBshub
llcJ4772RUxgzRZozIlb9Yc/nWs4L4u3P8vzKRV/q6TXpKv4Gr1thX8h+ileVcwD
wbvVeovEBNLyweFfceTXSdWW53Mc6n91w/Yd+OuXiuHRUQw+i7Xt+8Wpg5dUxkgH
zU8Yxm0kOUrITTNPCBtJnlNodRahVnHscwgAI63Do5SRrbLgVIIceNOGQlcyHteT
s9AvPYuPvJckVFXPD4wbbbj7LrkP+aPKog1zP85sIrvG9VEpGuNQtUtdRsFoqvUY
dVzJ8UbIgWoLCCkg1x+pwa5wZRdVUWor6sYvCCKezR7ZLQHGjmjZNSl+VUklJV6I
vjx0EeQwBpQ3pdDA7k9QbVmSaquL1Z5LaC/nXjh/jdHdcicJNxeObqsK+gOzNRvt
JbmqMvxxmSgbEU1LZqIcYC8HNwHJuuED6AvxtqI6RCdVSj9HXHV7SCDWnjnBtW3M
N9TgAQLfifzzuwp4qHW3AleCGUyVWquFU3Jzz7GiPNoR2Ma8aQlSgo/LQPz+Sje4
uTFE3omZYALrMXZbg2IcXTss7iGwGM9siRovKKOl8PTHWkgSJG4v48LK95iuV4cu
U7S8l04AVnKbPR+YVJbNRyyi3T13AUcirRQa8EfHTWuPlgnpzLiNpTfmFwnm6QEx
cCj/tNMLkunVIjguUBv1SZMCrKtNyRhTQuHMfs4abXXSwCzc5HIaTrSPXLxblb71
df+3VmPDIl0TuW4v8mzTiUXn5CG7GAyBZ0w8PmjDyHnhyGn6UiuwhXsIShsQ+Uxd
YVP6Rkk49L6LbwXPqEczqHrkuPdP/JdcUqBbUrS8aFpNABHkrexQmxb+0O9KfCnc
BGljq+ZtP8jY1rhu31KaOXa2KqL9r0W62E6TZfY/NWdpBDAnk4wjcv9w1MZrr5b0
HLAa6JStPhUZcUZ7afiSkq7vg1a6s2UhvnMtaA1odGvTbTKJ/hyv1QP6arnjv+Dc
OOFmrvjlHxTDJJmrHKOZgYuU80HCj2jXN1cZqRluu/G0i9h7IknjXls5HVc9zo+Y
o5J4CPp8w5IxxlJX/crLhXdUwtONBwzG01j3Og0UK7MLgFtEME5bNjij8TAUcJqb
aPzXSGVO2OaGNkN+X1b3eV2qVdlNrYjWYPu1cKHazNQnPSjpK4LT1kn/woKAswms
BbIEG9XBcU+8d0I1WKd1TL/FUSql2UeQ1tyf3DPCJg3whb9yFJkjm5h/1iax6p39
HpqEDFJImE7A8dBsygilRf0mmVm+GklAb6VwEJ6tEi0kqkeViu6RSQlGqtHu8W00
xOzlmZHk2VT55iINR/IOaaUx1sXGW8axaIGXm2nBTI+GxmyxKt6NqYHFPuill6j/
fbhfRyiQqBrF9UfFQn2cm08ZurVNnefDzaq1f4J1l2Nunxmwre683Wucw2lliBqp
4J23C2nz3+BJrKZp16DYvZAkE07c3g7Xj4d3IUaKyNGrTwSTVYFSq71D5kUsWfTX
UPCVQOLpwgstf4w4Xs9RNWq5res9X5orhoawGke4tbkv18WcdtfFMqA87c0IdV9Z
Gzx/pEOb+5GrGmTdCr3I7JB46F0kjqnghygiIfYIuZXQInFuElg3YKjCPJnrheog
iBi5X8TYk2F8VitWLJgSYabcTmCAwpa9cS9U7JL1PuNnk+yoQ9YAj2TIWD27IYXS
Ls/dRcaDvPFPkLYSXlAF9fXPBPv3FZ27bDxeh6uZ5eFTEgWrz+8VuohntFfz9YA0
w5r13WPiPoxm3577Olvh6QNhKkFTP1udamygElOxswm0O2eW6J8HpVsH3YhaA11D
5j/fNAlK92xQ1+duZbNKumB/xrzG5ey4P1dnTGLmaiq0PFBI4kFo2+GHTsA4L/qF
AS2UIyrfCYMhlyo53KMQCqomc1/KYLVg8X7fIHxT7tYyYV+FilaW7f9624cTYcFa
13WIykVk+PPwLNzQfaJ0Xzj/k8MVmaiNZ/jMiwyKR/2Nt/Ds8M8x3ZVg8TkiZlEf
JllmNCKIqhC5tepLlreh+d55hLJZA+9ONwM/RyvEmzNoqwjyebxk/2mMKSSpz5BQ
oLr+fX3HUkh+l7tp4aVhh2v9nfE1dGAOEHMcVTzXCJiDIf0LKrP5gu1Vcq3TUp2A
J7zcy7sBNxse4JBa7V+/qQIYr1p07szKg7W75Zxw7f1GexBExE43Rrt0lM9tXU/S
knbuzpbdZXCvBHImgXYNgoi6nz5aYIX9ey1WVZ3tF6Qzd8cG4qsxdISftS+mKQ0I
aw/NIxi6ZzZ49CBB9hpt6b8eyQGANDQ5+ekwg/do8011A72T5dXv+hMb9/S5nEuw
f7PN0c5HnnaS+WkihK+JGZCfsZtfNLVz0GyxmxfZjvfiDbssTdiK5P3zwJmq7A+8
qrs0m7qC2h0HxzltJIFGE6vM5epM0GPpWAjydSFli2jFI6GVWM5nKD4L//NY4TOM
5xp5Mfx6+bNlRRTrX/qRayVxISb+975DuSl9sE0ndz82qUAmf1pgGr9wg7pvt1Un
9pqrqqD8nFBK2b4te0XdHcsCjp4oySLAR7Ey8u+lBdKXJHW5M8XqhPDqTD2o/oax
gYG008NJFrlvbxYb2gZQJfwZuOzbCe3mEWm1cdrICmJOV5ZjdaRougZGmS592P4E
lRjDo7DVKJuUtmG9VEM8dDlLXpM8lNWXU4mxqzqB16X3LC6sa7F6yK0zSF1I9/J9
BvgNWNwkE+7ZHyMwvsYeGR5akGui+tfTirg97v9zdFF1TIeU1wwF+EVkbXnLc+xF
fQMT+UAiEqjXibyUD6Crzs8tb1ja043zOAZAvK1E5w+1C1kyv4hOpQfgI+82VqyB
ZbdDj1RW7S/BVRt8mCKIHuWfKxIVwYK4FA/3kqCJqz+2wLw5XoyjkEeC0H2fm2Ro
x5YICqQWriN3ABVqfIdc6HVh/B8gWF4WlbJvsNbb82ZwAyTiHbUi6Z+XTYXrvNnc
YBuX7vTXrFz6YDHfNxQbnHh/OG4AacSVXVvf0h5SrOjcQtCzlRB3gydbxqVafQsp
Rr+yOFT7I2fvEcdk8W1aONgZHHdJWKo5u8D2ObaqxzvCxMHdS+bGJ6tyOfcwZ3Dy
VthH4tEzY7tXpREfZ6oC019GLl8UXJIiS2PD+sORJMM4SeWGq9dHJcuA0UMNv633
24D/bW4GjDV5R4/jE3Ryocn3Lh1fkruC45IIOcu/B+bM3lWDxqqK3iqUaeBtknt8
ge17CLeAZ7J4DTVtAKRGyadjMj3FC3jK9h63x0cvABSCLyYbr34AvVzgTLZJ9d6y
NPXPnPg8PWefULlPxbbQ4rNe/q/IWDc46pu8w1rF8yhwEnC1cl7SZc1NmMDH37iB
xc0X0KNjmWE7OLc9XPs4vaAqayTlEPtmBk+xZNBw8J2IOQpc4qSQ8x7H/IsIAmP7
Y9qlRjz7RQW/Ww3fxY9m4XahcPLmAE8pBhcSJFbIxd5uJ0fE7RVUs+MsEewQYsor
dGf4pYFCSWxFUnnNFFij8rTgcMdb4jACLa+cYGatMq+HZjBe2ukATpwmEQ1K4mMN
+P82S66Ewbg8W014qCbo6mJJoT09G41ZHJQekQ1HyWnQrwNGVxzxePcCK2q55m3q
TmFK/e/COhhp4t/sMJyekgz/8TsGhf4h1/z8pZMWhmDDGC9ui6POMiqT5mqk7OHw
bNxJtvazdfWsjP6O0YHJwBmgSeYjBF5LUb6+7rJShG2IytNbS+L1jc7SN473Yy4v
fXjUdPBEEGg2dluEbCEtbX3Z9KWZmuBt+uwjFJksGhRlkm2/2DO3B0O0kBHTcfUP
j79hqoe8Y5z9drPFFV6yOQSsbRh6skRUcxu/9Vy+v4EJWzjzcVSmrvaeDjqzpXn4
2vACKTGXZBmiU9Opi3A6a5RY5BP9+u6Fvoi7mQ8wtwmPC0a7gseLUpTDr/ECJ+Ry
gcMkLl2oI4lXzNcTUF42GwRfKXpqkFoi14HGDe+2B7Y2QDadMJkCWNc9BbV7aFK+
a0X/yEQOWjya0G0fRTLix3iZTiMZTGyPWCTgYr1W5y6+vZsoQaAy9jzWKl/FGvzH
1ILHVBDqCyFCCNRPNLtWzW6mAzTjJHArvhg9lFlJF002nI4HzFYmVanQ3oIaDBBI
ScdZ/bocvIFK2oPMd+ehccbAsH5tyGE0zvQ4UD6STEPSfx/WFaBhLxxtIq7Uf2vl
vahbAdK23Z6y+1oZKFtjcgT7y8BebLim/Dvvv+juOZNiwy1cxCCD+N3cto7cfOdJ
0ovSvjZ7q3AJrPEKeCd057cOUde42hXCEbsTlVVxOM0/5tPFSW9ExCAhvYkqklSh
thJie9vD3dx+i2GmFDrYS4JqBfjkQ5V5q3i+h1xgxx238sP2cdTpipnEBc9ShyDV
RSGVsAl3XTDj57tpYfq536KDm6g20TbZ5mBfE6OHljfIbuqfFI6xT5zADBhl6PFa
HSo9tjYHk6ctvxKUO7FaxjfMOeUb+cq8xwO3dnJ4WcadXelWtFbzjcANm7vHvtrh
G1ol0KL4p0il3Ug2TAGATSX//nT3pyXfTeUxXQlQKBmBD9cjQKWzVa9NrjF+4IqK
SqvyKeV3ugfYEuOVjBCGqJUWuJvHVK1Gu9ojIM2iuHfd0/vYFl266TqxhEK3ZiJM
qemS7pO/B3AmX3ajIfmOZHYCfwQKG0h+do9bbsMrn/Jsxcu0R7uSI3fT//2LDKUZ
fPViB2+CT9AenbyU2aR7Pw/7Bl74h1VxTkPS4BFs7GqN9hgjY+zMSvmIQgjOSmwR
mz9JeAU37m1NISC6YbO+ZgjkQDEm3R6SpbQFVJ+iUepmdbfTK9g5D5n+fny0rhN6
+vBWfdrLINSGsW0JluQiKFwv2jfZQThJsiLf8zjq21mw/EywIQzWlB6S5pkiTEu+
+KThDitPRBMB1m4j3rdgWmF2bUO0QtEgd2YnzMqMNOIrXuLYhIz2G8wq5WEiixim
jNRYCNRJsCEbKplDPklD5GaAbwpfvRocOKJRtpLR0xUMCbxpBFLm6AWQr8zdA3VS
nT20C4Zdd3ih3O7qp/pAzo6dW8E6dl6aWF3d01L3BLpvm57TtY6P4zPb0o7ETmMJ
vrzjKgZKKMVJhr3QHpUCXEe8KHFvLL1f1YKPR3ZiMA8iW1U3ZvMcfoHXH8COy4ts
fgM5ls5UALBSawwl3PH1c9t/uaf6yRRehuPAy8U6DSl16EhVXaTgKIaMW8aGNBw5
6fIPGLYqCJs4y7V0PBvdbCxG5pOgXJtNwjXQIYsCC+DXWgSsRysJ0naicDOICjoc
Com+KsIFrcuq6wtyny0FnaPK5gmhhuy9kMiLK/gda9fuAt7GhcTJXmt+hxEpQLzP
oyjaap8x9ELQR/QGsZURxhAHlZTec3nE3ON09je6XZC+foRKp21GCHxZQK8kyEyF
dRITPMHPRWADl9MY58i+APS14bBBejG6pGkZ5qlr82J6O2YGh7CCCFneSlZ3K0//
`pragma protect end_protected
