// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:36:50 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
YurD831+nJXmZP2V9h1qgega5KxRWAJKmHe3tX8xhnHZ0BlYHqPq05BDEMWAJilq
IFS/Pw8uaVnSoxxOCjs5DDfjMCF+A77v+29KNZlQHT7JJuaS3w0clrwtLMbh2Ejr
4M9B5OXQp7Eds+2xZYsfVJAiN3to9vk6+mI/KakQHKc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5776)
2sqhAplj/Zr2io+Jquk7uQCpw7THt+WcgFMUw4yDJEzqBHqdkVtnpXi3Lj5X1pit
hMA0Yseg8wbMmOdcJlwIg2LnUIoIFOOvcmLGXdoXjGjRjHHKL0xBxxtrnZyLZgOx
holIcugwwxMXnD5IPYRTVmCpqhqncrXJrOi4X5+5r6mJGCEvaULkkoxsG+WcQ628
n7KHwycdTaW18sPOKQSfaM5Yk0GPyQ+0AGqXsyLc113D1CMk0ygnn9MMQalXXFHY
RllbqgTIGEwk2ENlskWwFng55YQQIw0+Njyi4NEUo8RFNka7CmTpOpHynOcH8YI5
m7r20hM7aLcpCxjDRabGbFnzkgt2kJBqG1WVCgwJH6O5x/nhNVXpCXMbyrDEjQpa
hv7p49gLH57m1P4YEt/OT2qDwvjZFDwMNEMnvbAy9vTkguYJ1gFgrofDBEnLX3Oh
8AFij1+Y2n1DPsgR+jMngkSTYIegfH77VgEpGQEKobmc0tQ6o89EqabcaRK2slrY
kNMguHv9mO2cQeReFGSTYwjZ3oEbMyW4zf0de/LgC8tJbiZC0lUU3+OjeeZ0LKNT
eYrYGKS4v3QPAaa06PDxd+LtfyEUp0s5sQzkAfmybo4t3HmSEZowBOGc/S+Q3lBE
k+a2QGUOdVLGcrl2RkBA6zA1ha3JxRr1kcaJqNnEAyJgRrWYi3vZQXzQtlXPhHqX
3Y6KlKakzcmU7uK/NW8dnd8fvMuRZQxIfPWWnP1Nsq9UNlzbZFgzg0utzVT7ccOu
CMSJz3UYcMW6S8s2+bKP1ZsBIVVzHNkJeC6L8UaVR6W8UdtSaJuyOSnMtJE0Vt+m
TvoD8y+ofTYbavBfLbBLHYE1rNJuwiEy2jwS6bioiNWvN5TNngK8PvHR3ZIgwh0M
eorU6wbP9SrEAHmK6w7XdOM7NSfK73iSF9E8aSzuEMzHE45mzE+ByWfEqL1DMg7q
B2S1I62bh42whkNGx/uz+/0Jf0R9cunezmSNDUyZyaqfgTWgnuODJ74pM6Yg/xXp
USuDK6JGJx9odaLJzkjNOdqJcGWsFn+Ivbz7cxYcZ423McpnY+PKXgenLX6Gh2WN
UCUjfzfRKw/2Na542LnJ/r0hp1aNFfXqMk5lV9OnhSLg5xzQEgW08fbw7WNCdpG+
bfGphiB5TaD8QejbeYAWya30wa9i+qksZGkBFhnKEAYpAZhzN0G6pV1rTJOIw2pQ
nLEl12DL/AkLgaH+CrDh+Ol8gIHcGzmv8Q/4Nqt92nJ+g99IYwZ49Yg5skXCWhc3
kbv1e+OtoX0WXYdpq8ODD1LbXqPa/fsJb77XRqX0pmpWb2JFkQ+CdKZ/cPedasdA
qiuRZQBz5q1N2B7np6FAf+C7ZMP8UUXamjQxZr4lBxWtRQukcqadA+XrP3GXFWtW
pXY34wg7n3iR0zRLx77izBCOak87d3TYxr8XsNiqg9IbXg79Ls3TjbXOWMZAtMtQ
xINcLf4hBHC9mFTMRO2kKVB3ruMpjxLRkvCuaeU/atIgbE/FX60UwjfhQ6oYMnUi
j+UnojKLTCv/UDvKj0GMCEs/wAiAAwetOUVKFuXhxL+J9BPL0s4705HYaG6E4Ooq
xEOt0WyC/E5shLHDcSC8QepZU++F+q8zCLlV3v54rfAOfYuEVkf8EIeMKjKOSbp1
tTYih/NgtPH/GwHkeAkiKvz4Krn0fGnE64HwteAVxIM4hVqelCYfYPMmuz1xJ7d3
eZJ+qKbpq9PVGFZqgpaGqCa+nMoeiKmLCUEkW4P0cLfLB/UMfvxlnRByUfdNDnHF
Xiy/aYW8G91jlFX86JedNqBSXbwYYtv/EJKoVuL2BN78E8K5ELgiSZNFcK26i19a
q4pbms7qwJVjoU9DKaFAmh++QrGx64/NoCV+O3LZGlyjdTk11akL1PcTYDhmZA5G
/vJ8WBn5tKv6CyFWa4KOB/7V0eV67dVGXyfNE+Qq7xmFZS/y1WJ1FTZb6ZLydt2o
nkV4qBH/pfHW+BqUBEkptHXo+10xCeUXwQ+rH76O6kNM4Xd+E6ew4ZAWq1W4OpGE
n1waNex0omR7lwDsj8Wm6211pSm7ybxpgAAi88jnC4PJoT0pP1kgFTp5SuBbOWON
d39ENDr7Th4Wj5BsZ6TNmUqWqtpv7COv53X+4fH7V2SRHpwFITdRcuOgVum10vri
7rkLZdxsKgSn3ujqIs9NoDeDLk8EqcvHAtYbsM/MTQnUCBTQjKZ+geOPu7kEjoE8
s8+3Uuo1dLgqtN83zBfQuSCRqvgpPW+pu1uXhWrNJ+KJ6+LduvAJeDc0ZoUXD6Vb
tLCBEfBn2jXKfbWwVX9hNbA+BV6j7/UMwUDB6lk2qr8HNsX1zbM68vBByzWyDsfS
9J3+zQPh1mCJhIgoH9S8+61NPlj3hvsgokSrDO0aaZ7lGAcE0cI+9CBRG6bOgncl
DuByLKtLCgKBq80uBhUPVSfcHFTVlOVLjUkckr4SJF88VudTWCt3y31six1MnSKr
zdEtR11P+BCCtNj2Beq5xsFQ3NWzINARz0aXYFN6afOsWcjvzzlU3OfeG4xcjIUq
LizSlhWm10T3jmm5SKjmD/3pyHORas6rCgIoRWOyiM+ofFNg7SpukBoIroq5Jvnz
FUpVFmkyVSSvWu4pfiX2s2Eo3+dMPlQk+3QxUQMjoJiZ8Gd6QfAWnYmkCDN04xij
eHcEGjHIBMlQsYPJ2JCD2kvwjcy9V/zqXHJakPMlCrFDjNYGfF3G1+VvnOi/5prV
g8I2PxShpHxR0fY896yLGT9B29OS4tV6ypUPOT90Lt6JpECZyOdtBN1jlV9EoFRS
kgbrqNZ4DWprweG3Hgi5ZhRew2f6uXoCGm0axazsHsR76xbrPK4VZmWo6Mqll2NL
Iz2YnSN+R0cwupSE4jkI98vXMlmInDcycRJLEmHEMGq/BQvfG9K+bFUURVZ1Ql1k
6z5lt14zug6y4xqxQWTRFxePWopD9L68be848YYhsZVPXzaU50gU4KGSy/LUD9OP
KHtzW1PDhlh+EV5oKGs7ujYtA8mogmhiBNZn2Jqyt4h71KqKwesctIawZPTFxXCU
vBAYA6AA/s74inVdxi7LXqIEQMmHvCYqsBtFep5uq7/g8lt53tM3OtWa0wntUw6K
4fOHvHV532O/fxGUSEovv7v5WEmsQuL9E2MKCgF8lF+mRK5dpudwRlkHYoH4W3I2
Del4iGipbMymA+Lfhaki5p/DzEnPyurhARHfNJVhKJdX7HhCnk/6zf+xjZvQz0Y4
ie0FLXHlbUG8VXzGS8d0yaFtE4T08MUWMykuaPZJV36UeoCYQbee/50qwUWVQVuE
qUDi28MpUgrcvTRSVIdT57DG3UI9RPEIKBUlY+WWoLD8gsOfmlYQw9vcM2yxd4ya
St3YUkF60n6lPXkFs14M75nVSQ5fjO4sP1E9R+elt98hqoECelWlDm3IW2pskeKP
8ee4TAoAMlAhCBp2pmptlq5jlSyNX+LrseO7AK2/i8Ma/yWC7tkgUkancJVV/0qH
JK5BRUqI60o914Lac3TKeSxN8XmT0fvx7NoHBkQ4DMfqBWcooHlPPkIOuG+3ks+d
oiTGv1asXGdmstOC01J1SfmB7jF8Xja1JD8Z17/l+f1QZlVA6KzwKG383bBT/B8N
Y4MKtJEvzi9/V86WqLoJ2UmqnFL4FPyjsGLj02+2ntvcPMpwgWMPzerlGxoDLnBB
FI43fQ+eSX2/CqQwfEBWKYp+TB4WawtbAMlW9u4haHNfr+TVkAqkfkWxAVuDiKk0
K4Je1/KP0IFIjf1cTD4kOVSK27dbxxEdH/h74SOoRwe8MiAo4BReDWWXVQU9T4Q/
PIsYFearWp1+zS00hTQHMSrn3qlI2fGbcpPl7aDrM4KeQaciMUlEUYYIx1t+Vcmo
2KEAzqp4ph7ObUYeWrqbUvbTFhYwhFch5jytf7hWP+aZtMM/YBesC7bGMU90mUpE
7LwcZihkVqkhdJhZOZiVf44Zvnz4oRU/VO6u8HfREK4Xshk69aX+CdZJAO5n6v6g
vre7XLHsBC9FLMSPCvHRt8jqDsrfsgCCtVGqbHjIVFiWvzc9Xyyzj9490ItyXF1T
hYvOEXuX8c2AJtFpokkgxpvIk6YwyRQbY6OpWa4aDrhGw6eMm7ZvdpxFltaL5+DD
m1/T0XIXkQwgoSrmeIbVzfR3cSf1x2dbyq9RAhRtaxpJyoaz4/buD/NjWXIkh681
9dPigSJRWOvLllXCFcW9rOcO182YgLXoqQ7KgWdsg7zEtQpFg9zOepVhVY7iQs5j
G4zH0NC3gjlWYmBgA/LPh+6I0SZOhKLPVsXXNL2xUkAi6HOPk51KMVIZOKfDo095
HQXgOsfBkgZDH8KvQ4hxFhTtstcH/DtUp+J8o+9pwyCD6Joyd2jFSNT/1OkjdcE0
wcygsAF2obHvXp5m2l+pRpddrtehXWmuqAFLNpR6YawSR/tvXwg66j7qiwCtskYT
ecsw4W59lYizVZlahPxpc5gCqiul8/Z4K2jtCR4iKV0wHfpKJIUF2zLMf6BaLWcl
zl2fyTV0lx4s+ww8lpYDMDbV04chYaBt1OFXusebG9Q3i2ot3kIWANf6N4IyOQs5
1GaP9ICsE7678b4hb3L7YrggaWae/zdRcM6kCh3keMqufNKRpyhtURdLpB4iR/PM
71Cy3l071idJd974ocRFUdU7qT6hE28AomfVb54181e2ZISi8wYhifPpuAOLR6IJ
sVrdYeBI+U1QVTAzdbbztuVpXySmuFCoK5iItjqQOgIxGX57l0NyIl5dvhae1QSa
O/7dq/zxykTkAOouUcG/hQk1ounSQXKLpuDTi5C7xnUTlmTxP4NhTbeIL+sSGEJg
riZCPMATXAmeWmeXqXvFreBqYx0JYC8HuzcZt56BwnlA1T/9UcZq3+HMx1FCYpxS
q7vGgcWhaGFvnw2lVzCly16CEy2ROrikudiQGqcEgEEq35UMHWo0JF4ssZ+sD2SN
XvCUWR+qMa1qG4h3j9K8rqaD6sQ6hlijpVu12Rs9NSwHv11NyrK1vpqPIve8YcT2
U0iDU8q/VZXVYzRMGyU1j0RwFEbsiZYucA3Mck9trc8wCWUBRjKt/nM62q8JItNw
3GjWwUiUqDyXC5j6MYIjzUIiBhyWxYbXcbX49w9kzIqkXV8D1TPJhZS75jclcdO2
LJUjyKLRN5hei7fTttOq++BccDGRgjHwEO8tddTVVRP7EmOE1v+SdTIPI9phavAq
+enkNxaI8EiMAXIiseZWvMEo+7iyxvvUuTVIfFCL/RxRepP1rNNWI06L8M/5zt5E
fXjAk2m7hVRgcGMxkfD61QgPupmYXAH/MvdvWIN4fwHio6QO1SWBoED6Gb4ampeo
rxEfMZxGj/S6h5n7pdAUIabCT8fcRo+kTcELRb4UBMzJo1xfhngOKr2d3I4gF+TT
4sxbvhkkLHgQjXQUPkDBZMQ8WZ48ODZbQapI1nc5OUpEsTWW0g9prn3Gc+JfYcn8
p/F5khzV+EM/sbNvexw4jND0tI3TGetFQTf+k1RppOIXQ2F+4+spTXgY/g4ZfoIc
yr+gchM32jqFGcqWI8AVkjQo9mWw0rm7WVVUgjWVAaSIcj35BTzHFdmw2NII/1Mq
5o3O4p/qD6+5CrjzUTRxfC0FUEzK7XQxNzt/khMCIzA8bVIs7/+1EPCHZYLfxCEY
3DmYYPVPU3RPCWl6PIkMmpqb7fQ4RQ3JCiCHzMUDOulQXEKlx6muXzRgVdixRrTa
4W9bmixrnIn3T9x+D01smr/qWWJoQo94tDfjAnptn54LvIIbG3dmau9P7I41Sq5r
ilHMuPmFIJpxDMPGxGgcSHyi9Pus8NMb1mtT+4GzvnS6nRQRT9gIKvPBBinkLsAJ
T3XtQA7koJfn/2oK4oTSE2Mi9tP7oSRTKeYcF6swFuSsYPA4OO7YMvjDzRzs1LGT
8Zk3jETPZ/xp4ign60ihies7FnzoacyzIGs4K6vEGUB77ZykWRz+WsmQ5FNdyhPO
Cys6EeD/ZqMVw+Br8qSMctJeGw2U6kkPmsDi1cj3cxQnW7ntMHGOylZbKKKrJaio
70aLL/BvAbhcbwE+7zTuvcEphxiaDR7RClZf49oBBD5V5F/vu742jLqp7S/pFC4X
aLirvMZNqhTtBzQlKcfIq1hi56uJBpft743KHOVu0FfoFfr9Eiqvv/pUdJbWxkQH
BrWlmopKLDgx/C+JkQpeGKEOpwc20Qj4La9SzoECijA2Of6WWImAiwieUkFSibbN
kqK/KJ+FqE+BOpUKc5O50xlyJK17V78+dMyl85AkvY+j4ijKBXQA/N3s1yMysrlp
7GIVgbIFAv+YX3fGiyQV/sjE/DfKFppcn8OEnx9rgHeDdgrYfUZi+3Svo+6+XKM5
1K1PdiRBZp+lMgjrc0Pg426RQ2iugfZtFmZnPKO2YEByXWaLNNqO59WbeRGnpmWj
Rg374LBgzBzqrPF9McvncrSmbBdYG6zSIMGdfhtVBgh7osqONvTiOOjNLvGWr2fS
gfm7LMFZL8HOrMiKVe18CKBdCx8rKO5h7vyaYgF/LuJsBTR9RrYyaOdzMN06xJTp
Uz3JZUruO2E5Y5YqJ/nERkjbgM7NOzxBd1TOGzFbbcqOleWt0vTxVLpaD9BxudWv
JtOXCuG9iRjJM4q6DZRwz5Lbvwws/pr2qyMVXxH66LWcgydmRTH/kzkKpriW6Ldt
WCa7gyLQELEjlijXj4GMT0k7duD1zFxaU/rpKV82SLaD01m76J1aDx+unoGZJ+8o
GXIhbIY8fHQXqgTdnuq1diBjy32CHAjyeYbski333UpAmHa/M7DCKKSDhvU7EWft
uS/S+aTjuyQBhpXCgy7YlMgkQAgaQn9rG5WCeWf6XwZ4uFZkiMRR1oAbRzNX5Z7m
jldbrJDxSXL67Mbj7RCjD4v5BcXQ9Sujc95R9LI+d4ni/gFAIkXag8tG2kF5vudH
/YrH7G+BIyEYpj7Kq3M5p1JC6LYBGBzZYBU9mo3bxs7nzJ1l5iyJivGotWe9X7Vm
cJeBtl+1AnJAg5NjVikDRrfcYQfVTSJFVC5Pvs+BKWvOYXuCLLU5k9/EcYQ6/dND
ni7hxCigyrw/8UA6ifhbg2nlTKhRNf8hNuyJ1Oo3hKc9G/2bXhfQgRN6MOivRJWb
SuxpHGPRmLiJooCqi34JQbDXi5xHFXtDHCo+OfUoqea2KYsKPz4k6Minskl//F+k
k/nH8SkxCTdl910YEe8x+AbvFVSUTZtBZEqmB54zMgj/Ejby/9FqnOJbv/BdoSdI
bAikmUmKUH8xPwXhaRfMvY6/oaR6IRm+cx51I4SkWYu1sC4gGkEySgfR9kqnFx9x
mx/AwZFCtNhSwfu3+1UdLJEFjJlA/MfH0UiVfhqiD2ecL8iof1Nby7cafx5Q2UB4
082KzrkRxcWgl9wn5MW8qteKMRH72Ory47m0PZhXfWqx+OhNw76tsxJtr7IQ/83Y
nVSdUA6u16q2zPTuPzooX3dpVrwzaPNQeLqqI9aAQLkd/d1HnHKjF4fko4/GiXgt
y56J0vPCDeBMp8kpeEYbVqLFrjbGYF9p0Z/0QNFWobYc0tdaVhMvm3IxteDU8SK6
FWCyaZHdkuOy3OJU4RBMMdQVox1edk4fXv+LKvhqTJXlumR7Sn56XSgP8VYgXwSj
JZKD0tD4b22Gl6epDTdkzg==
`pragma protect end_protected
