// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:36:52 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Bbt73Zljz+Z943f8lFFGWRRdkGZ54tXmY4/XHM9nxAjYP79WWg4zeNKycUCGrM7J
k78P9/uPz1h1pJ2dTG8Hx7rV7oxT7fFbYEsAJSUwJMy5C1gT3PQIjOE9Ge13OS7A
XLaVD77XW2ggaP0GXA5Pa1siA6ethtDTVQzhk3cI6Kc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7568)
MbWMfvIyE3YPVdu8scwryFpAeLTmFhgMp1Ew5avEG3dhJGprOyjYcEBHKXk1RTW4
hMAOcxLO2+YRkczXP//v9x/3KQa5tivcyZvSljVDNRjxGfkmVUBJy72aFuT0ag/7
l5SJNOskjsw5UAzwG0+7JsFs/mStycFOH4hgc1ZWbaATX9qwGraAAmLyGHwROTGG
d6WhrXByIqiu6gIPQkQ4LCaCfpTEmOEZyOywdhddaopwQU+G2kU9sV7xKhGZr+R7
wKeGvDhc3XXaDQVSjYyc7XW3NPbUizgcHgGZjpVdY05gtPZVsYNXgCO4J56XUVWL
f6IT2G47dbSsIlWPWjHHmXCMhAa06Lxuja7YVwrjP1vdrxI4jM10XQnsmWoG9qzj
P5K9jYjDFmPO4nxbXbm3P6aWqniNEKudJj3L78sKCeaLbOY7GGDUt98dkQutEiJ1
nU5a1QroAV0WgeA1iijd4lWeCl6XPxdUJpZ/2GHPQfCbcx277/qGxhnNMCddpV3G
nwntVws9r53YBRIcjjxci7kq/rGa8TVDXmKy8zEFJ1pG1evEafh38HbiBvMVeYGu
9Nr91XUHLEJu9xPbpBoChnwfwLvprr/iTDk+UxtAp19n53zUkW+cE9ND3c4EUlcH
814Oo1Res+1qjtyxcMczfgwSn8WCKJ8Ru6ryF3U3aiLVgwgr0pE5CGyrGhnjEfmu
RBJSZjVZslj8BNlRYTvINdtiRFPIgT22VNgF0kyG7U99ySDJ72xRWmpZfcrOUo7t
NZfIFdHfPSKE1v6uz6J8TOxqMN26w+1A2XJUebt1S4Qlef2wVnuh6NorOptE0TQ0
92kOvr/Z3tMRVoxYbdofBygPsnuAT79zh/aZTIhNd3trcynoLaOHszWa5Ofk6V8d
kW6F9XVeJg5XTlkQXbS/uQ7P8+PxBL5d9TO/7gwD3A9RMSQdQfG4nLKRqhGNzHjy
G0ykNVI7l2my3K4/6k/j8tCes/DUVqVcvbE+qQtJLs0SsWbfQTFHka3eqCGmnDnl
dSL420qIg5Gp4GR7p4Zg88fajRxMYl8823EwDgwL4026oKNZvIrKhpe37JD790ti
dA3ys5m0BkcEdngdAhmKS8lV2KzpO5RLx+Lr4Bl+WXgrBWUDb2Wq5dyu3oHhLHDv
YUjHtyeUNxSoBTKCXTYGmzzP6GjcB8xh2B9F5nyEvCGolvDASR5qGfPq0CiAC6MP
cQajBliXXf9B6mB+kIPLf18bAmwVQDkkxBKJNKuDwBViRHxgADyt4gH0g1hdJ9n1
5eDbiltcL9+MF/YgeISOzsbJC1DAFqyEa5V2dmwb+0FV1/lI1T/RqV1QQ4FNLj1m
/nR/te5zNy3jkfCpCmhCMoJupih3yo4sJ1JWsV+Ql44/PwGycAd7vQusp9L+A33O
gqhI8tGIfkZooK22shblK8og1gfBBx57FQg/6BtB8toIlVGS7ZGWNdDgIwHWOGrg
Hz9pG5TRuWQ0AKDYbBzEahTPFkJY/w8QMfFcOkbENgvQl1ILAnL6ZX2AVnCmOMny
S4rf7mewQg5cTz2DwbiH18IT03C4QoJJAY95bxQHrV/8eqtOv1nj7wLcFNwsoKOz
11bIbxCtC26L/V0hJTaAuBN6VcROWU2bYZr02D+ZGEyQv2sNkiXVI2+A+Ue85CN4
xyIs6Zly/tBno06zq0mOS3pKq5sSbWr4M+y/LJWjmsyiAVmErv5y/H8qhZ1u+IvT
Cz09YkcUwc3SStq0UXq/QNWmVBat0qOOMM36K17EplcnEsPmW34/WWLFXOQR/b4n
GP/HPKMp9hjqeyKMvdN2vxs9hjDyiQewBLl12pJm7jtKQHXFOScHiyRq1OtrTlSE
yDWE5rDioChAcljnuPVoQFEwvGKehahjVHqshE+fuWbTuD0dnQfw1/kVIl3hhqGa
HIHoZPjfjovAK/AdERqLD27hphZ3xCDXZl5owbqh3fJNt7jV0L5m4ZgRGbs+xzJY
C3T/thTilids2MkJIG9aO9Lh7LZ4g3D3+u0WW8vrAXQarD0xMjEwnzyPhhxv+1UZ
R75I+2Ph7QR5oaDnYPtoe9siwcgSPtm8AvxeYuA0kObg15Wcuc/qBILGuuhd48wO
f+RA1gOS+GHqCDzkDGV6y3FhEIbY2vdwGysSkvKpWJ/5Lp5lYUqCOB6nIY1yNoAJ
+QhKRmwngBH1AoKYKjwRCPlQFTJESG6Vgc9jekLvda7uR6jFN69b/onlHJdCPgGN
6vz0pvNdAx7vR9O/KxAq6nvRFyfcO+ukyJ953uYrpMFyEm/lmPbbQBqVJKZBCld/
KvlhTJB96il3d+0bzyIVBSNC9Tn54oRQG8emeU9dXuJ9Cy2zJI4lxUB8HBsFevnN
8L1ImxLChNRC/XNoBsZwQHWaHKfBopPoRWoPQUNXkuO+JN6ZJZcaEtzv6koDM3rR
N0pDelq3Z7PCCJ0vpiIUpSAhDMUUNx+hGQm7ympCOyjDb4IXM1dM3FVF1QKchHGH
1Ft7ng07/BK9hikojUMZYENrFa3nr2LhAxn7DO8yaXLIAfMCFhNlQa4e65zJ6KIJ
bbRlXwy/lNHYcFo1OXYe4G2fBAZ5Ej4ESzwfCeSvCDHrwLOoVgS+uJY8gbOoNMy1
9fVDrOkDPkFGDxu9QnVhZcV8aw1Hi/ysfe5Ks19F2h9sRiF3wgIiL403JVYLgwkW
lPgCMU4URCdoAZWNNmlCJpHqkkY7YUZ0VCq4UIogo5NNWcajkmYxPn1FSkgtOZvW
e8XkV9bMWS6fhCZ1FQ0f1Ea4VaVDfEoyGqdDSpIicCmiNokIrrO+zAhQo1SR2RoN
ChDZzYweTIEbbMnFv4TAaIyoArqoGex7P8uPvlVkTcef9RHkXgPDU8TwvK4Bruhy
w1lryYE2da7UiK4Kf20b414IsmzJS5F8K6GbKKTGP/2VTDugcbeA63r74RKv8N0n
qJIXCO0MZM9jwpFkkXGLc/M7onDk/a0KGbmlfjqKIFe9gvNPaAPtZFowN8ux2Ro3
7iIgjzlZsunHujKwBiedcl0p7rJf5YXwctZqBtScODResNvNP/EvfLNGeNLum5NC
wyNK5s0iUDdavNhsozAF67Mq4jKypIQUz6Pr9/DqiaLeBk/fa8RdVRmeQGUECIke
Vixo2yoH1PGhvK6DOW3PX76y1uDxBOugDfg2qKY6KPaFyRWARhQY7h35ni3mHSQt
mvbDlnGXM+PKjCtttWP5jaKv8Y0JjoIn4O8xik8PI3V0rnRcJ1dfaICLfiyaP4vC
toY9gf+cxyo9xk7NWYe+KE4eMWmffAgF1wW2j1TZdLalwXNrLNq6wGMl3nDGVA8P
3ZuGUPjCCgRnJ9M4eB2jESS/eT1pVhlgtLcpwwYtFAoZcOQOcmOCd7oN2lyZDx9L
ZAVUNS6VA3KyHqYg8heYcQSYnxjo8GoHnwxT0q4joRG1PWtysKWplSi0c25xvr8G
mET7dq6PGXsLaRMT25ZFOEJv/rtxRjkucGEx0xBqNQ5FeAVw53rbdd2Xdqw3jgnF
yAPmt9R0fGZUddVuuwY9XmLVGLVHptFWyzmMGL9oo4suqHgeVsZ55lpwzkZSwI5Z
ojTZjfXuYBsYgkn+342cO2KL6Tx5V4khr4BES6V3L2b76/kj3TTn/ByiGq/gye9/
I46hiKDdH540i1SaeLpDyC6mVCAf4Z9sft+he4Ag2CSMSflJY70vUJ1Vah9yXmkP
LG0s5gALH1Nvkh3lrOLLG1QiaSPLPtvUD+c4dkyD8Ok+UGkVgaOSXj4M5u/AxwUq
ZmLXWQBTzReo2Mdi+hE+es5xVbk7vmEIcEEddXvfhPPx4vZIQSN6AA2ZLnSnp8Ct
qEvR4y4gxulA4TNpr5P3NMe0CZW0zZBX7Vk6FFAdzAK0mJdBOud58FnmG6YsMW4/
PbJZoCDHFixPuUfnoA71PhAHOuT/xHFABuFwNjvAMEs4ZW6Ymn2rkmrg1He+U+s5
qWGSBOxjpTk9Z1uVN8w2jbztboKHlod4mcGU+I3XE2H2MOBMa5VxbmjnyaYeOCpB
BOm2RibGIaPykdsUJKKM44L3bABGcjL+DwkpFl6UZn4Ew8B0oAEkqz/Ii46AfHMe
n+m7RMuXWnhGpnXMg7JVRP0rzIew8W0p5eKizCcAQe95RxkK8kfUlUVlFEMsGOfg
uZ/1kEuuRy5DFXMQNysR6ee97T5guIpXpGIyCYcb9ImhFWPtLECQpzUG54SG23zI
7PjQDEdJ44EQ/lI4pfjL3UYW6+Gui35O2uLkheX5tJXqRjr1kHF922kcqGppvrIV
6qiB18nYmdxbmDIF/k7UYSeT2BTqvjkEyHci1tS5z+qWJIMYgWshhEQqUYL+u8Z0
qA77hfI+3nsIr2RWl1TCDyIdeYmmPy1Vm0dhPfVbYrWMnG1sB1z/E3iBIxr0ucTR
oOzoq4l1goSXirfaDDt8+cnlMj8CTmTVGbvcXX/89v7ceJWTn2N1zmNq8AvFRCSJ
3KbtsCTcGSIXh5DmfqHVMnjxWB7ORLVNsKCdI3uuz54VpsgwNRMTPlCTqxMePu26
ZSQOmgh4ou7j9C5yRSxQRMDIQGJVZsaEhISO/Fo0hGOaYdCm651LVeqerLrGR7HP
JR8bP4dpoXk9C9Ly6porXMChN5M0Yff8dzAbBw4A5XG65uHFwUSJviHpY3mzD8Ri
/UOx5iipmadhW6RmChMYJfZLHWpPDhkqRlpLTK1V0EUxpMHou3rlLHyv4vYOEFG7
KAxkrEBLgE/Sq73VwtAFVaYJJC32G+fSAZeWnjXgqxqUyfQtaYFrw6otKoJjDjzx
7uinBasFFE/81xl74ewYYmf1fHVD9qDZdJ8z4pPaNxGUnNJ7AzByuP5PTajE9/Qa
uo5sLNv3R0Z/829UUAMChUzrF7SvV786c9jJPrRj6/AkexYiY8IttH08JZZIFRy1
YaBeLY6GSiuUS8XhMtYcNSTfhTlDYqNOeNPcnmKpZF5Gmdht6AK2elE0c4LSybWA
/b7HO13ADYtAgSe1uQbgl/QyFruiBR4DelHA5FztYYv1iusTbEmt6ZFG74RUSOf8
kfptgT8j/NMhP/qy3Gq4Mm5zju1gXXggvYn0UJo5ubp0UmBjrJ5rMGMlYD7Dzchb
EwhwjcVlrIcgwv1hpUPMNVZkG7YAt6fdDtbkXwb4pVg3J7F3+0/Bcl+spszr1BfC
JIgYXnrB+XcFsSNPG7Bw1DoPMvHrjJ/wwznlLYQsNtauTxbsrYJUxfBrUC5VWZyc
ts/mW1lWuQG8Y5pz8Ttiy08Sj+717gxbnR9h5t7ul4bFbhxK0Ahyppdpb9JzdADh
aA5oxUOcEjim82woxIayABsR7tNo36yqjSABXEpAhb0l0xFUCJ7Z+N5Nb5LVgGgG
wMYVsPY0e0aCy4jgFr/CVJowvVYkMgfLfXEJxQYmhLepHAsuI2VtlsG3Sxtc6tuF
MKOdrrN6xMwMJDUKnsnh7PfSLYZXloGlszhGYfN5DV4i4Zn6KsvFT38sgztxo5E2
EntdWQBGkoLdgMwReXcT/y9D3O6cDalfxLtSm5FPuilD5etbMyAZBhH7Vr7enfg2
moXljUk0GDttgqhsy63pkdX36Spnh9nLZDuZx2Nv5Ri6p3dFGVK4uJ+/wVxMgfbE
oqEKsSmPwEKm1RkPjRgnEj2fAkJ4Lt4mUawTaiwiEmi5lOZ5jx5EJm4i4qsvIgX9
q682YCydloTZi/cObbEj6bSCXu2mrqZ5uJaoOyOJZZUECk92u+3+b1DJNs7UmP5o
c4gf3K0VobOIMwEPo0jX5z09VwEYYv9jBVkgCWCIEkorCAS4Ro5R1vAlujLBO3H2
BI586hWza1WL+w4lOtPZ8Hlo5YfDv9InCvrC7iz+HU1gXEZWnTWlyciHE5D1Reeg
BZhzBFUegFyXqeYRl58KRnba+CjcQdJkXUzID3sgRNkgGP3Rn3S+k3FkIiVRQsC/
6fGEUxnCLQ26lxt0swZXvQ7W6NePY61ssN/JwqXGsRrsDeXX3Jk0ea0X48lfM6YI
3uT42Qu0vhOj6lovl2yAHFTtRFgl2WMbQ1jwNIoB/VW+VQPfVpvDLb1p2J1fHg4x
9x4Yb0X+eHEPQBcwcG5IWCGktvcZNC6Thy5zDUmsaMboYleUvHb3oswapnby7VBi
I2wXtBRoc9Gk7sOXitSp5+NjF11FHtzRAXCDqxffA58YD98PK8KHha+6E6N2GPxQ
NlEMlwFo+2NouRkyvzZZ5kwoEX3fwFupTvO+05B/GjKwN52DaWKoo/EVACC9jxws
fl2r6Z1h2153EHt5x/M7d4pb8+WOskrqevhmOj3qsmEa+30PUmMZC0NuIazaHCUG
+bHaxV+45cz9Zv82TZWTp8PS74xw1skG0A6hB3QSRtAQFU9mwUXzwrxZpSngCiaT
As8Wd/oCSMm/Ws2EQE4yAsKDWZpD5p5e2AcGrMgMRDvcoCuTPjujGN+CgBkOK0P0
q37nOIvxUJCZlcgWjUCZ2kcp6/vphqV0t1mX64eQRXlwS783o0auJQPiWl3UK7MW
qu2dCBowjp+O/FEYbDKWnVOm4dznKvgxKs/Gtox+mnmmjCfQXCsYsaeC8V4b+ibH
zFhfNz7IWf6h3vI9a+PVbePjf8HeIucX+Ek9wKQFtlfokG3kfuWQFVA963XAPpfE
3Vjby4g5V6hq4m18Px/67s47poSdszmIGOxBfeBoIFYCDGw2mYRjA41QXgSWSvhC
70TisXh2LiLFrxIoFV3tYE47QQ0TPy/gKOSwny2DQ2Up0ZGGsvwQGgszJVXXZkke
aHqxM2Q2/UumDYVbJktd0SPNYBolTkxjiKo1djK9c3iHroj/yAbJK1M6xBgywWJM
E3EcztlLEGkxIaPmbaNlUeYzaXWy4o2/xgPi+VEMeBjZNEwrpUEDsr1BagPVsR3r
f83tL6txg01FGOWKnpCfQUVLNJeTooUodBlznaKAgWjuBO5SPlRPIM50XbploF3W
98m1Rdlum+/n9mLKkngDl6tUK1HCwRqt5te60HpmdQ6vBmhXP7V3tFOS0gCJvOlI
PyOymC3EKoucs9vlWPqy0L0nvaYUewz60VdEYndi9Weg8FmsebcNHXtaDoKpP8kT
u3mgxjjd4k1wk1EY0sgOfSSNQDRItDWKjIAU0HMSyCNvw2dwm4vsPOHc53CdjNOU
UAt8vwlLL8eCjMjuNUNN0GKzC3huGWJFEKM1wTyk90v0h/vbiyVYcxcFA6YnNF9j
3EMVQGKxb0fcZvF3O7rUjQegmrPtCdugoOvquj3zKLn9lRFnOzo+hVJjaHHs8uV+
Q8se9H7l6GlSwzBy4Nlm2x8pvA6CPRJvczxM3YU6Fe/iX75+z5Y+qT7oTf1w3z/S
a+POQ1RD1fT7NC3jBeQRtQan3r/43jnYS9XIu6jIiKknR3t7DISa2cyh1X1Ct5L0
iqJVpUKFIfMnFr03sNivBlh0HbJfPdS4vDK4fQuxVcLb4dNusS6kwXHnTbKkx+h+
LWDDGjH9wtm/XAnMsA+ciAxayaNnwm2ZvSzWLLMCANpbF7u+ny+DFWTpA0nV0aZI
PrZoJ7jZ2uxDc0iP6Fw86ZZBThFiyv7UCSU2EtamlywkacxoavxOqbj/yPihHHDx
9fJsQKmR0+jaua0mMZoZaYVqIN2LjKIPYtfdbZmXljKfKS9ag4hdKnfYWqQdC3DR
MWYNRwu5L7OYwPLAQDhzaMF7pVgOo9MTnrIlK1sFLzG1g+IwR2pyy2YDkck53ehj
OhkOrD5fNw091fsrXx2AprvXpNrUWLTjGPBMrpaJf+D5sXnsPDypaLOTFTXTl9NU
dj+EwAjR4XUI2OY1kp7U6Ish4iOoOz3M2rox8On+f1heVDmRN3W1RX0kjb6suitC
/WEveKbAGXokf9ENj2DW1k4mosUpHK1iYlnvvtCqVvoVzTLuML9KqMreqDkgq5GQ
2nCHbOoRR6RIOw9Etz+J9veipok5val5pWBiaQB49Zj/CJFulK90/9Ps125SD3eR
6rJW11TpueVw20HylJ1weVh/kyd7uvaxCtEaqpYX8qvArTehcinLj3QgXF57NkAq
9tWzW9UlOyNJdek0pvbyPbpfL1CuqcDyQUXRwyB4dCsx643CxS2ozjHupA1Ejh3E
OAruMb/JZwYOJuDn8kajfb1tDBK3fgW+bBK4Y7OOX0xINYiXjCZGlN36uoZhQRr4
7kOaR+iOKHeFsEabCXBZl1msf2FQA81NMYGg6iMomt/4zyW6Gc3bPcsRTDW8pPFH
GEZaaPb+1iesFvVIEMLZr/HhQq6rNjCSqwGCjniRBJk+zqZfCIxs2CCnM3sM/KNU
yYWI1vudZHXQaBYprQ4bFfUVaEWwO39G2iIPzPSzy0MmRi+LWEKEKcLupp7hBq9O
+HT930k+rN6lEGGErnRhHbnzHAumxBByPgiDpiinQ/wu+m17lsX6NZtB7g2zmZfo
jqlxXqk5rQsW0lOB9q6RSiB9fs+vO6EdqxyonSgO8PP7knxZuocpOOWvt6lZMzZZ
iv1j3kde8d8vlvKVsTP+UljNj2xMsi7oHwVfDtcjhmj9vLWwnC5A8GnGeHoD4yQS
XIkGrSid8rSH5b1H0aBx0qjg+f7iRAnyqz5/cx2eCpG/Ky/iEv0Z/YQChjz1jS3I
A9XlYaA4N2K2X0o9VS72/bj+zwDdg2RMIoZcJvVGUAftu/wciZ65PeU2zlSk9mBG
VZPgzP4BdA/W3cTY0k9sKtIfNveaAualS7DzX3hjz4jiQpKQwBruYiYlNJIjjXg4
M2kanB5Rg0t1hrsG/k/cGd30VVZP+ij+PJQ8Dve8cXQ8bENjkte4+0gK+ceLPxvx
PNlWkAhLvZIlO9FpLL3q+Ukq/nd4X7QOhDi7xHkTvW01vS6iByxZ27RbM0hl49XK
RXSicpJ6ep99sOMCpTmszit8/rptT0eD7+5F1f5bCGzZ0reOf5dCA0hiEsBRpO/3
yNPHdbPU5WJTTAvbTLj6hVqZzKjDYcHcFcH8tEYOMNlPyFrmdBH9yY2QdFIyb8r3
hmVdp0vLv8XCS9JoaGp/RXCsde/1A4lehGoaXekvB7eOEGHTerTgnSflFrkW1n1A
66zbbWHhE03EO5j+87zewJndcRQGNmpNrdSAdHTANi4sVU6OD9Ux/zK9sPdQMnXI
CA8XOanB5F/pW4drLxgRcPMwKfolJF2MljxPuOlXXRqx+prsekEvxOQ1nPEwtFUk
zqNV3zzB7a+N/OXTkFB/6JrpNfbrcs5KdrLoNyRHIRpXhR+VpjH6dArs5WfWEhqd
VpioFMVzuHd/cbp852KHfrs5Sfpgbauw4xHCzAmPur8vJ5Onsp7Y5hAmryR2HxwA
G2t7EqyZscbj6QQRxeZE6PqUV1zyJNl6XvRhgRj+VZdBtkK3zQeZd1K4rGcHD/T8
cdQLemMQ2K9opSCGqnXQyyvHAsAz+5hs4gQ6/Yfm5jPFJ0KD0MuL3FZceMIulwDZ
TN78vV4aK1hI52PmH9mgBLFPKb4Jv6aHzW2d1A1raLIBE5kn7/ZonsVCXmr4z2Q8
0SvJst5Y33sN0KR4jXpA8e8ljQF7vxic/DsEYBdXdicz2bBpN1rZC8z9KyEcHERz
FXyfWmc+i006MyHT+I/qv/37nc1mRDzyjWb32kMh5LAVt7tUD1Rq3m5toUBZOq6G
9Qzgb4OZEu/1RvJh0KiZPtgrT6o+nieBX1TUD5tzB7w5pR2LMbUiHer7JwgEZwYX
SV8vYTObzEE7cQ0zZFlDNet76hOYr+zAni2tpRKjwA2iGQbuPbFvf3w1nZ93QN1H
i3KYQcgYUnKv6qFIq4E/EsNW6GjgVsBY6yhhKvfMrPGNgPrULB48uUQ+YV6R1SHy
LazE0gm9/Rljai401MW1ImltRKmmjC6dthGf7g3A2MothbwHss1u+qpaaR5OSK98
ya6ikP6jgXZnh39XL+3m1KCl6kU9d5AwB/l5Z1jOUpGd9rN/qs7HXDnEnqqr5Gaj
vJJdtODBYpAsurAm+4JL4e+rOX/brsybCXFDqsDiUqy7e9LQLdBehLQrHaJjbDpU
z0l7za5shvmnuUlLGhrBxKYYlWY+9oO/lorjNXyOHXM=
`pragma protect end_protected
