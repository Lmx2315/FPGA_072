// (C) 2001-2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
vgjZHPBfncaBTNr7hbZsCAa/6/p0DbHY/Chg9AZ+Sq3PlnqinJnyBs/DjD6bnNctn5T58V3xdoU4
HzJrHiXSUTQwhqIralU/r2equso/sn04iDTLrEEFVmi8R8uBlM5AdvKo6hYJKGOb5l6PsRkDZBk0
PiKhygdSXk4PTLu1bHfVApUULnTzqjl7PtCwrLEpEMqKuXtS4+UYo3dH5zGjrC1m5uFqfFvW24DM
0g5UMagQBx9FfDJpM5kWxRqwta0qysEyd5FVfpCxvnjuwXpXaot+SGA6YzVwTwVOSJ7DB4Vn30Bo
dOTVxzTT+ieqwgkoXo6dJW4CyJi5EgmF1lvb2w==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 9440)
9EXTonc/ToqpBaKOVjF7VmPHnIvIhxVI1yMDpbSUBcau415RZHGn/0N12PAULD2rMUUpVCI8gGoa
uXSATseAIiN8zFbAqQlGgomcdztCpivObNkG54dJDNu6RI47wSUHsnMcasJ6ltfzVvd4QObM98hN
clMbdJXu18cGjs2bjJKKURCxqemF/y+Zh200dILTSRFqZfCI79twcG3ph3f+vEcOC2KGm4ImyqQ5
BXEjtGFNGVmPs1urC89i7qtJ8jKO5h1ExDXZIGLVusJfxuBFcy63W33YogzRBKMiyI5PgSJGBAkf
9TYpr0nU9t+TbX4AnWv7RF7yy1/FJn4jmv8p1amfjuOkSUB5fKH2v+KAmcHpXaBjLinGdx65c7fL
SlK89BisGfiDYruzmxIh2iZvCSs+oUfbQZBw66KkQ2SGgwcqDnHn13IPE86BL+e1EOIp/en26Gsx
M5B3J7jEAFCKO7WR/6BdEXQpvVYjX6AMus3w5NtsYCEEii3R5m+8bkW3Y7uQA3VNuy9XOHBoFkTd
lzHROYaVk3SCNpSQsQ5aO42BIe9yxtTGa8WEUWO+mw8OvEwItPqRxjq2lf3jIK7aXac/ZuD8N4+S
0VJc+ULvQiqhfv4dX899EN+l9M4Cz+1JXnxxvuuO4h6fXkpM0v5QWprQWEHGiHBN5QVIoQj3fhKV
zFm4x4wnMr9QpwYHKJkRC2bItqIrHxmBh65RnUqVapkgaTnpObBC+91mweH9GKVSUNFDDDEJGYwQ
DXo+ifTisbTKy+nBSG4doKRT5615lOrwK+AE4/hfEiAzlIEgBUZ2e1ITfoHFRUttfrTahivlJRV9
miJWhEd12btWJCWFd5Da5jFoGbzARVRWAD+a7OGNVH88Ask/ZXSG6ydfr2REwfivAHBPEsNPEc8Q
zkbBW3DaFMYRf53rAsQQx5TcKbHVMbvb0xNcNPnyDAk8Uz0XQf240AmFavduyd1tqxhw19vdcV4S
+spWzpANZTsQNWCx5dlyH2/nKmXHTwJAaBXzG9LsDEbV98eFmq4iyJf/gEDdw3LFNHuXOQZWaE9C
BWcyz6R0FcaQEx8++OK5AW8VTXvUZLHl7RWsVTbTrsqdjWpYFdkRZIemYLzSVU5fVhoHlIJfYhNT
GXEwcYnT5CeGQY6j6Bf78N28l6kyxi1eW9R1lZyaogbUepQXQyQVw19uEalNMK727EEPTkC6ttn/
CcaRBfkBjFHaH8TBNEEW0VhDmGjKdsS3WFtZ6yk/3WuOagv/YeVVumHsVC/v7K0BC/1pYICwbBS/
qYjPJK++ZeOb3ht9aHICUeoAJsrNclQHup6+XdCxtmdTYG9DAFoQB+oT6XiX2e+FCyU8HeV2Efc6
CX0G2UgcATyJ/x3ypeA4MJkjtT6I7OkdUeasqHP18o2M5a/9PNVq/ZCPSTjzfIQSn/3fIg8WVrkw
Xk65QYr6PU7gyVG/RjwH3/2oPkW0nkVM8KjDX3DrMxUFaLmWC34hsgjt36D9uv2UWohYjh1fJavX
HC1zgqoqQ1B8Z65H7txVo3731BzmqgjGH9Hvlkt6+5HAZDj1m8tnR+spC5s4cWzGA9GdCTIxNqUW
EpxIYQg/DN22mraRVkc0ABQDrUKl/fkeevo5JlGjGQgLGdEtaPLTSzQ6cjqQeGJMkKOORXu3EYEk
1XMvYy4qVSRztM1p1VYw6Vo2LPsm+tUB2NyUg3nD6uzlzJ57d2gWytyLlyrLEzRLoPjLGbAD2LER
L2Fy3O7V7K/RJLx6mIzF9JQ3tu4UZ1XjiqoLkE0aXJFAb4ypZhR04MRVtNajWERa5naSHduH34UB
tVeJLJIVG8sIbgwRFxckPnCd3iopqvhbJcfEyDtvNtasEHqu6MvF1wevPQ2WMW80l7FVsb11AUcr
vlbSsRxCFhjAaznummmlHMtzu7cAZ0LDQtsV5UePAQlU4Xj9loMe/CoYwAyzExghTUtwy2HfU+bu
qDMaGitUte/amc2fuX64Egx4L9D8aMcgfLxF7lorYIiHCwRGTe5Fj9OIf8N+M74wnnrcH2f8CHel
WzgG+gRIEe7iUxx6o69AbG1A4Nz0qMcqzfcL4djgG2pmb0KfVIRZ+UzAKWvuIcKMjXpA9Yb4FtlF
+DI15oLz9SXlpwPSyxzNFqoh/2Vp+L47PCBoUUYjpnCOQm6XqAiWzfDNDFBKfIZEVB7+0iMpXWFD
n/U3gKoPahyqZ0s7Z0MK4bAtde786wtCFL1tevDPQyN1DUv+8X85RUxBiUMpZMOzTenuITzJKn3D
eZr4wmrRzZcXV/5IYRuY39nAD2pcjiZMSwAG+U/vQq9sOw7KqZ6STB9+OoUAWTYDS5jJsuDKXFT+
mK0fosrvLdN9b0fDiLO3JN0TZQc2+3FO1trNTA6Srx7aFACGGwj8mwfE/Wzo5ZUBQmSO8DIyI045
jgXDiazMYOPkrbNkR8YGoOujQUXat+Ii5ejMUee+qmb3jjnsHB+o4wwVBNcbkcrvYaZjYKV1lfmS
cynnKjwMZKmhI6bNAW+CYOVNtwi6+V7b34zH/cRsa81uaIeW1RSFst7hMeQgdR+4Ypl7dMd+aqZB
YqjDWJDX7jmaQBsRnQqLp+TCMUwulS35s/2fz0zAVj7Rt4tuj6dfX/wJk6Biomj3EJnXIJqB1DFu
ebp7R6pfq33tbZ5pHvmkgc0+Lo+nuZ+5QSMRpDSWQfienHMeCrMnGa3v9E/3FsxGFeCZOFdGdR3u
iy3/uXpU1EwoSUn8K8rjxDF3fIyb3hXvodam3ojMsEWzFltvX1xfu949MYPRQTCtrJN70fPlwAGu
HBMfG7CiBIdijEbZ6uLdHXECd9DxiX9Ya6H7ubU1P3slJ8vQRKe/LigH/mPn5zBxjfM1A9PNJAdL
dJUUgVu7Eg2Nv22SIABHSDn/4YzpO7ehSWIXAvPrVVgHrZqOiKCktNJIaI1U8lYtN21rgPUa/GNA
8o5uswrsACs5+ebvXgZodueBKmpTm6GT81iXdSQiSpX/VaNFBTw+YiwIWkGGI2Yd08IgAyZPvI4g
3/19zPMBecd9HpY+rOwROYOaPH7AEPw/CY9VvW9SUM4Rk33/ejzX6hME/RozmCgehvq/OkPu3P0H
RFUvwmiUCkCfxtGwMaL2QkqU6mdE3XUxmJw8+J+0oovOeNQcWINwqNwZuZht7IWsw8navO0e2kQE
e01bBN1uEXQeSahmMBlOQlPgXj+6Tc33+iDm0aUDU/fgliHVbyDoYEAhsw8JByCNHpIJSZJpPvT1
v4bbH22KvaUjcfhuwq0e4UFqqXHOxwKrOQZOHCNGZ2fTtHzsuUkvPofNek54XN2fXlUIDOFdKkP0
B6xJhjLgArhlqOLrzuYuZez4irRGDi5iYQWeg7j1x3gmVElkRkhZsnqWS3gy0KAgRKfzb2uIKT5n
6zyLbtN47yoaf/bkr6rCBCJbhnTxjk0UIsOIgYqNFWYJnyqs+Bn6xbpCTh6Sb5ICQhs/Z+htuAWf
pLLIQhqsl7izPeWptxz9NtrFA2n9CPRrh+Uk5q35swHJ3uPr1UAx7OAW8T1gYhWq2Z72ZWANozu5
4ZcINCv1swHygUmaHfG9myFsF+/IHLcWjh4qlM8j3qu3KMpyBlm45ZQHxSb1G18BEnxpFXHgVx9w
/8DP1/WCDzjh75374h4dCXu9SiFlVC/KIGF/B9HPDEXKkwqJVwNETLpUbQgfcg7E9QxONtHSHLDc
ORpWvAx1GEc4UWDMsbdh2S0sAlT1y8Byvs59PR6eaM6S1LjBZxAzel161dY3P+aj/ibPa6VVRDZO
Ic7uvr0HdCLKhe1EJIoligtHb901wSHTvzt9pS4lKTqzwm1TObnqtvULvAd3LkUrWQS0a1/mGHmc
MUBd2sibhZdvTLM9TQgxJWhqUQ55qqM6Llcg0A+vstwc45jQqaJRSm+M65Rzye8PCBpzi1l5XPsi
UqONAyTtdu0gNc1N0q9LH8V+6ddVAVx9h+EnedgLKhkKr9MphzSBc62y+qdBr1BdF+ZP/BU2aabh
HygpQsKP7HaPbsjlKXv9alSAEtCID+AoDjivsh4UALy0pKFGH4BoGSbi2/BTiRqDKwtNnzkLSNme
V3MYYS1wqDKJ/XkQ8oIRE1dpbbSiJw6bWH6Tfv4cfDwlQuhL+NR7zbPly/APRyM2e/1wJ7B/OFjX
G8ZFxtbzc7epuSGS8zZjxTtW3yBdIz1I9XW9vPBYuakIrpQnctUd0aDHFnbHcApmvMdfvTj73kXW
5LkvqumpuEOigcamdnRIIemDx/XpnAOIwVK6SYaHY2BimeRB/qKTL7Wt0/nMJbL9v96GGbLpf1/1
m138yGDQFI/vzmwqJgyAPRggloimIZkx6k51IANbRKdoRI93Kl/iCavKr/EWBp8GGjTj0fbRAW2a
pm3ahbrrsmoJkZ4to55DH37zdsREdgQshhsBsV3Pu61ITCoIkEwWkedDodnlGwUcjPWKuxAgCZK9
vJ8Q8YUCOuTPwkpt4F9BstjDeQsG1s1cWDp2yXZZLsGGg8eY7Ej/ptY8SrjTzCaJp7h1Sp+izdT8
ppmUt0pePCwkanmu8Ehjwuetb/2QadCN6WSgK3j+pzJObgmjSc+kaWPNv2CQt9j6xtCraE7HGWHI
wd5qgn8aemcsPXQ+b4YNmfhhf6oKj+V28AJeZd37VHRt/tZh5VQbfF3EfrhITv8wuGrIvXWycEGh
y16rBN+XKzK3ToXsY1XXSOkon3rUBHJAtOT67YFc13Re51t1XpNvw5hFAvrgkGzk2I/fTyda5nT3
LmiaxDyLpnHrAK8z5rBdzPVGBo/uGgeHbg28VhrN9G0h10TshwiCZqisogBVVD2zfcPA+M+42VUU
b/6dzkrBTrQeqKmyxUv9hjhIklhu9lT8LsuSSLlftQZgEN5CqCjaYM0TzkKSbvu+kRxipjq12riY
3GLGNrLVq5ZUj+nIBq36SE7IfDiMCsFNlZZakVqoOLZ0utSJcqw2yPTTHipab97MHAe7o5Jk/Aqs
iXhWuwzEMDIIM2e3dkqjgCzOf2AWGYDP8JBW0yxUcfhh+OFCW45rgl55PfOB+bo2nyvpD18wUrwm
Ht//O1FEfUG5BdZZI6oeaxxpAnNs0zXpbEdUXZp63sp3wwzMB1oxAKLxoTQ7UgKMpV7f2ek6AcCD
i9v60uGk+ELTikxXJIXH6RAoJoOLIYHH4mufftv2SmwnynbeSQmonC4wGorkpREu/iDaEVsi5J+e
xLTeVS/hpdbYVxrx+ywpoHYSES8ILx6c9C5LDPMxBz2etBVbrb3vo4oeIvybIuh3cFzkVNVxtdBd
7J+k1QWCsAIe0R/Xd0BFXYRjS1U0ISnksmk8yh/9ztZ9ivI6ZqElwASG2Ih2Wj8qfkWJXk/CHLwf
CK/z/LYpXD6JrFLDVZ4H8+YYeW7JMaPbEo0DOUcNQ1ql45OpQ+eq3VEjAVox98piQIsCFifGWa0A
Zs4n4TBsX5S4g3bV+kc7tuvXXbdM4Rn8AuAF0+iDpy4hiMKdcFR9/3gugTY+tB31eze4KLF3bode
OyW8MRxZTLgKwLjmpXkdUiOW9tbBoNJOnG6nzkPhV0lACQc/xru9JMqx4xPbfW0vYe83LA0kSo/s
la5VUL2rqdGAA7bwoDdmSVTFISMXwu7DFPDs9OM5bE8CQP/knFTmPps/mIFTQlH/uWNSnv/osSXQ
CWLANplV8p7q/O/2XdJNfmgCL+v/mtkMm8PCmM8XU/7zNh7mxsrfLPjvq5sL0an0jEJZLwms/MtX
eauDo3228OPZNC5nXjpyZ812ZSisrF7ddfCMkgunwYyjahs7bt5UmquDmpV+BJGbddTxKUIGz7m5
1I8hKo3NXTjT35JC131zxJsvfzyyhhnijNKfeDC5eWcFVHfpQO30QsH2LwMnUGf/fBoaVtx0Mbl/
09gg9+hS33gpJgRzOVhCHeZXqc1VjrzzE6FGKRE/lLrlvlIsQKgRVR8cwCF/rQBPrZCJlMU8Tf76
+Or1mebooCFoPLba408O+VrJ4qGfRYxnvETCjQTPYsHqtiUcFJP6PTEsDOREQtGEtBAVPbu0SHWo
vmbzNm6UCEzdNlYn9G0JLRYCwnaEXEvJKjAD1wUgE84MEJBMsFey5MrgwOmY0AaeNIKqwfB/edee
JQd7AQz3J4mZqza0QzaOez5ezlReYNpkW21m2mNgKo9qg/6YEEpF4teTNmc7a6jJ7UlUiKvJr/dT
QsZuRMWAuBV1X+c7A6rOaQQiHT39/HuIGsCcpuODpoKtJdFc4yXfU0QM7edLXayHJIh4bXEJWIZN
xlCdsOlaeUwnbT7XS/IdmeQnNP8o7N8m9/fXrAXqrH83aPRf7vc5xAiiBzgUMvhaSCSbCiJwhUHD
9RAL+YV1zO/EMKXydAJVL3ur7ChgyN20QhviB8l/ON/KI9AcAnhDdXqG+kd249ULV7vnuPxxUpBH
XsPU9SLlG+JZsEPliTAjO1UnM7vxH1ElH3V0FyJfhxhMHaMRbTRiSn9xTQ4PBpniMXl/xCEbwqzg
4eXpYRvP09Q5YQkdbumw0h9yVGkIBjvTBCdpMnI1xC5yiW6niEzT5pkdH0nutivqo25AAcGjU6EG
Gfp1qzUcUm2XMnZj1/yTZ9lcrk3MXZkr62dFRC0jLAzXZkGEDvAFH5nSjA/2lFSEsG3ngrtWJCa9
+op9xmxYyDKQfA6QwYKj0P7evAHAeg+rakPdOUhrmLHQ2toh8f9c8H1YK1NLF2GHRf8eiLSqBXWm
6I4PyZ9vv54rh4aBWv2atC6sKZKiCAPjWYC7ArY5dkn9pCo82K5C7L1gatOVBiX6XTCiuq0NI8P0
e0aWrSA8PYLYKihQTwQ0Zjt08oIqCmQRlOOvD2SY7IZAF9TT/MZaDfR92bXl8dza40A0Hj4x4SIC
VKBPxqFgk4Pj/YlxNuB6SNgZJIQmL4Z3+EC7xSuGlv3k6ub0pkDdFhhOqGWTLibn11Rgvv+PBEeT
SRXNWU5p86483XjZ+UwPnjhKzO88/1OhFI4soxjhn4BLUbLohSmVY1fRPC0iLWcSv976csPJW+Qp
4HSW+kVLHLjErkgkQeXsD5+XkWmct9MVYcNHWIIO4Wovj19kmdHD0WAKBHG5o5cHi9lc2Bu2smhN
qdOnKDluXWB64gbbfA02JE0hj94HCa2HGaKhxzBCsw+9pbsoxYTbC8dXROUKyJa43Wwte5f6ip6K
iX2iTlS1gaZiMau0bjVyvJcEpLABCJQFVE36jeX1QKsGv291EhkjM2Pf7qe+T1mKRdRkNwa1nj6M
qgQumttXK3fpf/E2P7vX6IU0S10V4JzOlRgIyJAmCzHqvgB8S5fHRxpNB65xnYVXR0NPhBcZ7I9p
CdwmWRo1bTtZxLA6ZbOQk1z2wcma4G5ided6d5vHF5bAeYTI0yYJ8AbH9AfIkMkpRvRtWCbo9pll
elpNfWalh8lNTRZtVcGNBf3LuVfwwoMUdhaYcoRow+kcoNk8kPvQbnkZ2aw3G3gFVfgpu2Dhs7Hh
MyDfa/IJYTeVFlEwXX0v9OiC9GUf+DjJyTQreD/SB2K5XWCmqcfhX2qdlVpr/vZ6Va1SJ+cx6jfZ
+IEnJtbZXLtQUlMdBMEiL2VRfXiHtJEvd7f5iB+97iRgluOi6yNzORcYrJhlxsfKxgcEvklEKI49
7bS3HzGPw/7tZNdjysMKgmVy1UB5y56raguvOYw7ZyiGGePyxqJg1++j7BJxbU9dYjZuexOltkms
qRSNF6uOLkVoOtWOMxoQPvApRgo6RtUDMFd2P1sPMBv5le4IWHTAIyW1AFCAFwDzFsypfvzPBtXA
EAvvFBgbewFgyQ4D1hz5EhPrTBLwUvfl658ZCvNzmzmocOvsk5tiAjxmK42jV1AzpQ1WCbPBdx7+
vjjnP42TZDb+58MaM8C1DhfeGCV+jcwzHgJ4EApKUvpBpKZTNkEJhQ2Xbn0cM0kFsvEqa9AwPfWL
nNn2j1yTEB+VlzZlJW4Kc5/aSongKlrYEeT21/mVVw16d/p3xJxxo0+wU2NDIZj05gzWI9BiiBKx
XE76q349JHmsfCx7DBXsAJ7mDYWT8T/SpbAXOigIfItFLSCs6+FwJ89K9dgHUVN7Oxnh5RGsPanv
1Pv24cq10UKUCFXhU9S1QgFZDj/N4W/nmbFRFBN3iqgggfsr1yAABe7ftisSDijN2imZA3rRldSP
KhK7IFsTvZFsBYc9l05Fqyn6UXnxChVW7N36GHMhtRkMB+gqlzPqS4F9xJNNqffJ+xOwA7ympEW7
9CXCx3/yGDCgti+3LQ7KIoeAwFUDmDt/NIU9z8j/3WdOxxptTrWRw+Zzojx92XrVUCFms6JZc1Wv
SKl2aGTuRSt8rg+pHIyouhdtRgOXzLsorODXeHjem+y6cOIB50pY9rinH1DXMVbu3CQXoFacAwH2
+fQ0gIEhYuJV/lPDuizS3ETaZw8n9wrDV+erJdF0SBR+vWkMLv4fLeyoG/q8w4mu6xXBQwII87JR
0FV4fLDfB2GkvwBfPcvYgTuK/n1H/nlcUr3hM8UC2j9ZBNWwSJOJVd6bR+W3AOujNHcbrE55X7+N
PS3mXcvJusP7WKVx0d1ZVwLXVEP9tHUlpyf+BxNsRl38a3NCJtIijUrMkIzoSP2UW5OOyu87dmBb
Hn4Ev8fAOVOggcuJEu+zdjIpDTf0qdOwOeYhsAv2z6QnBX1TIUcM0jzuaswkpFsxrhHo10vpgak0
VnTrlYiOQ5mnCyPAL7bu60JeAC89oTL3hVLvgUtZ0isdL1mHjRsrJlD/Fe1QBLbDXdgoSo7r3G6f
yBUvVIontaqWk2JOoOyld3UZx9TmGNNWh/HE3omoWsDuFsUoG6cl6urw/HPijikqOlapwjyhvJAS
N3ICH5r03l6Kh14K2SLg8c1sZAP/fjCmk56APNmVxYlJ3oUJiuXiUTgsVxInLZXZHZnyuJjpLUDl
GigDMZiFxIioRmxTNRxvi4lYmDCvhz04WT06mTCPlJK4d0kj/YPqOQeTkObQzOXyEM63MP3Zbyqa
WEgiBwE5LlOFXTj6zpZcycm9EBWah/FP69G5P/u7utBDXOkeCwaclwcjFaq4OJUph/KtYyhnFP5a
BBmSEMELb5toTF51rS4bg8c4Z8INPvVdQyvGXba/pFgt20xp116SzmHBfPnqeSnprigmATP/XBH5
LHfClqUZVUnUp+trjl5xzGVJkT9WKitZrpeDQmxD/krYpbM2M/6TaFQ/G3/rpnWx5IJWkkSz0Eo1
ofwzpMF/D+IUiQ4Sy5v6ffVF9qNHZ6wM12mAokw6rGkWwedktbmINQONhZwnAzs1D7seOP91WqZY
CbY5qoawJTbj5y/khRtyuwSwyOIx3lpjtBVoewZMpj4wXDcR//wewAcoJhjAT7AS3EJcimX9p/zL
kovH/kXsP4QI4OvydH6Xq6mLBE1Yp9jh6Ohzc5yhNxaNKOGx1iucq7/0uBSPztGzSheO30J0W8qI
ZqiTEoGiUvwhD0sZ5gOgy8Rx/7pIGwpHAVzuXu9DBHphiuFGfl4A9e+BwrPjZxv2AJql5yUuPwlk
Zvy0TrzXuQJTlFq5g1S2mVkAVWkNu6X++YWUDiCB0VHBj01z5JQyL95DYXqrk1tGZs9kI+t1X4wP
u3bLbzrml27aNaw7+S25935hbsb2OmJkPQkmJEv/TjgSNEWnY4ikfRsdZxS/sS0QskFYyMt39HeM
GjhaS+4PjAPkOq2fBiIHuv83ha7tVrjXk5c8XlFarwKO1V8oQ5U9dVWPdtSp0+oJ48BNV3xxc0wk
ZFeaU7m53RD+ZxV9OmwvAxOFxzCFErNj7pctisDFHdYMzx4eRDwc53cEpOiWW80q3BckHt4TSM6u
gwTMYBl9CHMyur4FV5GU8ZBQnMEWYo3BkOAVO5eBAk1/f+QT/MBwfwc4udA/SwD80M1kapAtfswp
kPanQgsKZuNuafkOdBtoa6t3tBRU17gQ8j2zOf2bPkQdeoRSmZyGd3UMyuYy2MKlyGWuea3wRSVz
3OGdD9iByYmDs22NcM9wgM59v/4O0UyIUM5eHKRTxoAcJGe5zXun95N5XjVTt1GUqx0Z8IBcceWJ
ShgEdPVCWl0m+9HbWTluBVIzt4h43rdtQaFSHXKtkc2VbPg/6cvBC6TVo83qNDHdOeVg7ARf3BQ5
htWNDVWmKdUUfG2rqihfqsNOCENu23supyPbIHY5AA5N8NRCfkDHlZpY53AgUF7UYdfh03K8FdO1
Y66pH4lhDDmF5l+7hNL0tzXgS7/XY619hKJqhzUjpt9eF1c6/QXMziTaMUPZ0GpmoA2ycv95Kb+1
vr9V9COe90D7PYixxlmSOF9m7T1bPl/CUQ0/SGMHR1Qk8OBpMq5PTPK4HFOzQNAdEqubjXJXc/lI
v9To6aNr1KerI52Nnbzo33kC559dX+BrnzGApnMz3STv/R7jUg0eHK9nrt9ToywPu3zcSzpd4zC9
Rt51S2q+WIXSbjwHu/rsN3ueZ6YuQJQjieYnLXyfSBrBqzsKfduSc1f/iqOAdHVeoVCj9oBzsaLx
JWEGAFcC7bPbuMzjrfHjU7IuEtjPfDOCby/kpupPO601j3p4mvLFQ9wUs7McgMdm4nV62FgKmf3A
V6UIYZd/TIhMdj7eWQsls2TfDzbpuoKl8t5BQoqOJ26STsOeK7IObmV2jxH7u7nkWNCUjzgTeYsJ
yqlj6wiFF8lB/LligiNOSorwCzpBKrUeWviUIfibnDaplDZUlIo2Zz0QiArRGpsW5p09evxNqg8+
mXFgVJXAg+T6vhmTPm/khn9lnpn86ugHy2+6xFaena6ck62Pni2acZJ0RfdX3ShweDRicdKvjg41
gK029NlHYKbiUGXJrIeI6wLNBucR/cspJVY77FpsHn3BfRB2hFKPGo9bTza8kYHlQwc6zz61OeXD
+doIg3GZoSvqGiPIS572cJWGIIG9k5tAQnJVa29Ll3k7GtL87SM5iU+JKnz0zBxgQdx32NFiVg/z
/D55pm64844zNZEyyepQ2JzzMGanByvzpzld+WRrZzJ5+ShLVJ0d5jjGQOcmD0UJhld1vFEuR3PP
idTKqEZMKWms1v8jTj6sG9WwRTYBsCSehTwvD9z/GvxsZYC7iW+/E4Ou2JXkEIOzf3t/rbRtdRM7
33p0RlljFFmFdmoj9m1Ymdtjpp5QZiBewHxyzPMsJsvvmo76ljl6/3Pogh9xETey5u62F7xZa/rm
sHvbfv6g4LKqZFUA3e8WeM9OsRpbUVYyw7i+a6X244QPToNOnhJJAphT0Mg0HipftEXBu8uDxO5p
VHV9zm6/MFvwNGDYwoIJCH04FchhavkqTBVAV0qi49MN3DRyieuU0EBOe+tSZL2m6QVrmpjpImV2
pOhECq/kGp+tgWKPOmLcx3qdSV+6OsyqVGNfM6ua3vAewNbCwNeaS1bCOsp1rmBJEYf/WglHd6u4
jnSsCNDb2+k8zNP46AWohzUETZdEzRKv+1bRu/tzqlPk8dLEwORygosGw4mnQhhXrM+z7mibOWQ/
5pm5AnC4sfp0t+DMWz3nznZxeB5QMDL7fjfBTixnoeVtVtk4aS4FGFY7mvuR60gYGv5n4456LiJW
zQmS3oNsVX4civfwWN8nhwRfcbuLICu0/XBDFe7SIR3Q5/+owOXmZCY1t37WAnwzPfvedhIKTnp/
tx005fAHg8LsKlTtcSAJ//JBRBKgwAx8B3B+X2mWShpcYXjDD43J0zymSFMN+pSlDpRa7C8ihxNj
ArDGulF6atsECsv4moxytsr6tZeNclAdO8hq+7wJ7KshtzRHjU+6FMqlvJze0IoUeDYIzMphME67
jWVc35Ociel/cVnaUPQw7TXDwEbtZ1aBmT5QPmljeD3V9REcqS2wHJeeKoiw3IQEf3mPtS/vSEVQ
Fya0+fMYmZCLsdMoEjhT5dZRNxYLLuJxgVvTbdzAg1AOCNbcUs7wBYye0L0ObRlQ/TgyjeZFwrw3
+GnuyFq5snz11pmzSa6yiYY0kGfXrPxyV60MAg50foPBMlJ/rdjkeNMcbHJwVVb/LxOGtSWI2ge0
jnkhv2bZGUM10neG9qXwlCOaqCrpHRO95EDEZvpgodtT6uNwbAM6w0XneLfqPN+zYmGF/5gJDuif
S8w6B1uz08mx3fPuz9T3dJk3CtANGpBJShkJ9lYYtsF5YWIkRvpueah07bUjnU5wZIz4yWjo4jVu
fZxtFcoqel2IXfVCxuEFVBirACe9mgD0zUbR/nQoXpkFAph8urQe3zIZmLemcE4qdLYNezfY+6Rz
k5tZ+ZbVRn9m+aeXe5XakVgDfzdGMUYjrbWfHeKHjp6tbAoW51NOvE58fsjTCxNGD8nGb8NRdsPE
102Ef1fjbUuncDVi+vU1Ecs4dLQ0wzci+ME0BCdJshuz15qJwtjE86Mhl2d4FblxS6LfqsGAiHsS
rGRnCroK0oTsFYfAvHF42nCxxKArvpNz2diZKeAlIeq+aCrzeMNXLZK3+/r1AFyLLaZsDk+PpU8M
6PjYCggAlOzsw5qP7QfKnUW+z7wiHPJoD3HmEtU6+o0pSh4=
`pragma protect end_protected
