// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:32:37 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
DGH9od1W51ZDnhvQ1C67UeRRiS4xwZH16ocyD7tDN/9uieaLDPjE0n0zA/JQy20Z
6scmujV7gBmuyBEqmAOVsF0vHx+NVPtND/BiRSNUkiZ8Xi9g9n+ShTDVt/qd/MFY
1ygYkp31SMW2TH+qEHG2YPD/VbRCMeYeO9DIkT/UgnI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 18368)
tVtamNVnCwqhOdFVA+inh5jEUiLLP3EMVboyAS3W78nQYwvzSWaPsqvEKuhsmSp0
LSJeLjpTRdkOFp1gQq8f4/ErhjJ1sipVRW8H0wRtqYXiTmV3vEeh0ugRZ3w1ZvH4
AANSkskSk/kXD3tAxsOZnP03uAtsd/4CWj8yKt3TQumLphyT9NIyPh0ISrCKVBmB
tQa33G5I+bFSnoDZQx1ijQoFfscQnZnp0fW7vEkqJJyfpSkpb59pyl2yPl9YXeZ2
T+ODf4W6fMFFp5L7SPMb4pXjC8bslht4E4diZgISUlVkfm5423yLEJDJDpwHif1B
31zSv5K68Qv/oLi4qtCRTcAlFZq/htvNdtyEOh27xSxm1UBFBF4wUq/cwctFLCyY
5mZTLtdY+FjX4cVzaXWR7SWxnbxEKKwC+r7IDKprfNuhHtlaMDaGlD+kQs1rhvXZ
iYpcD4L9PDojZvk6046cQQaVw9XbwviwVaKSLFf1G1jDQQMfn2iIR1fY7guhJqiu
lhcO65nPgYQLF/741yiBGt7ngErxLmP83QPybZjhiOZ0mMhoKiyH4XungnTTH2ZK
ZLEM64wG321iC7isZtNMd5o7yDZkNgxzJaJ3roCN/uktcxHwUrVHlwvJjCjDd+B0
JbA0tljqQZXqsYiLCPJRsZPEIasLgpJanqT3dZZ6xBmCJ4la/P5j+n0a0ZuymLSL
saEFCNTu92pUjhyadHtJrmF0Bkeu0AT0xTDu9v4uWv+EfQcpbOClFY+NMlotHARx
l+NFJNPxTD9rsAHeOl9/NbJyU3Idv486+Sc8CjtaKVqqicJbAaRlip2Czrr6pMfj
S4XDmGPBv69+/ExPOEZtYuEcMzybAFPR9ChCybaCnrkN6e6pQ19vyokjG0Ux5dZE
mEEsLUpf81VwX5xwl7D7nl+c9Z/5wy0cX5VII9QqWD5g0DiZmEE9odyiKLOx/LVL
tEeoB5x2KaN2LeCHFCYVO1VS4O4mTHCzjk4jgRgC1XVjhxh8ktVduyUzjf7f6rMw
uyOkvMZ1cIArCsXneMKVOoJFaEOMSfNFtAPq0UWXHCCxpmIE3y3KTfHCh5QDtFAm
y9d4UkOuc6c4MrbImzx5Sfa+fsklEzCgX9R8ZmJsR4QQhQynHUDvCyLn9NKAFeS+
+HVXAvWONVw0eamlsy0eTcE+5G9V/DFYw4H5sNcZ9/SLiPTQV1XldlctzxlkE3At
9yccD0iDFhntQXhgoAWt4u5q4Af36BYUfc3xs3ETydiUgzjVUeA/Mz7C1FpJKBKy
WDT6jYsYNJKsFdesEzmaz1mzX/p3o3SaoaQCj7CntKdmhoY0mrP345lPIBP7fqil
mOq/5q6WqcqeLSoPqeiVBxrpc6gRiGdxIHyR4lE/MFyQbIk04SSZ/LuGLSe5g1HH
vxeD7cpVZOrCSg/cPsOwGJ0vXR9l1govpuS+DnB1N6u6VHaaIH83iMfmpZPmognr
VfI/F8R3Ip+z03JQ7ALmX3P7sgduLVKZcJ+1lzc6qxQEsg55ILgamIW/r+4eiS/1
ouG9AT78KMKOR5bZsH4P7BWuOQhh6LWkmQdSLZRS2TN5LNnFLJmwf7UervbAlpmP
1WX2hrakplZjtO8zV8J0JB+QCqA6Zmr0/c48Qj4aQdGmI0PwxdtTuTWe474fcSko
yEFnVLSNmmls4ZE3P8Mclolh4WhgFqiThci46aLgW9zmNJyfu9K8vjFBRxuLbO33
uEdcbMasb3vBWLQ1qBfHW6qZgi1NpkYpsIGu+np1q6nD0tzpmc3CfJMKmbn+N6Rg
JkZFeU3gXtljJPFy7UnLvjM/ajts63Bo20eCs2h4QZI6ZN07lp39A0R2BbQwuYFI
xawdBG62TI3C6TeHHjrxo7Ab5WpqALtyp44Jwh/6FG3ndxozlY6AiSavzc/Yksk1
FFScd5YDJ7xHXHMc+p7X2JHEZCuqGAlL767Rrgzniggt+BYjlmRZEq/WJEyZ1Lmu
6IPf40oRjgHqS0+6PtISf5M+QT0ydCYyYD7Na3uNvdTquabyVEstgtx6bEBo6VqN
kUnvKHEEHDb/tB0CCIV0CGWVBFdCIR+3GSL4C+yge1vHzo5cDiOKaGCsjbMPm+BN
2Deraz96gbTIOGvbKSho3AJSzyRLthA3W5BH7lRS/KpR/g6T8EF3FEp9QJxF1j8d
Bl+Hxwljkm/9Wqh4sU4iCAVR4HnXht2LKw4kHZk3i1r8npb+YST2OSAwVtwVaH74
x1MMLet52tKqe/DKBff6omEQAQbwKYdq6ELAug43yoih0MMnZA2znJSGfOm0eyK2
O6B81uwRNbldr+UaoShHYodlU/RDqoO5VMdgPtlMEhOnKG33ukLZxB3DmPtg6w89
qDKR7uEJZU3o7aX8G76ToOOeNlAB3ZRKEB+PdHZ0yfrnproPoL0u3InD90kTgyoP
CzFQxeJS4wht+P6Q9v9yJvFi89f0BauKMCk4IHw/tYzOkkwMzp1ART7H3B0lIt9P
RfNYm2lo/ONn0RSaT2IVQmEHB/NmAoVzKJkDMoOqsP9YiYpGheulSlvnPFfnDBY8
g02wpNaQm5X3DRx2nl3novKY3q+7mp4v/WOBScNM3YKNwtnmtxmavemMzIhVqVl7
LI0wGsdADE/3QFe/6rQxmH8+O42HcODEHA2AT5v7X8FUYuriYJwACkCJ/rQUuEQI
XyRdMJJqf0VRp4+78kxhTiPzmi1451TAH0UxIYgLLX+FFNShIGJGhYyKJc5+8oMm
dtTHnLxVY4BubpUjOWthFapTmwRX1oxyw74dtTxKw0NPkJQIr0Hqz7tIpf4eQaS/
dbcG4MYEPXyx1j7STrGzlYk8DPTnPXysdXNj1pQz4vwNdBkcX213TUty01bIs1hc
iD6PCq3w+pwmFlgir5+wGOXYLjcx5VUbKtMh8SjPo1kNNvUV/CNYtHAQRgubYs/u
dqgjzef2EEwOh2ZULdHE8WTJRHWXcJO38/EjLA4ClehdMTZZ/py9dZgiyxilf/74
V5GbIIVUjzkeAcDMKpGXp1y9Eh65UfPDexTEmDyGlBZtDE5l6Na40WsZlppwC/pQ
sjPDdXLKsXGUafgOxvnRG+kcB6TDgCrlfhhHnKlI/4ALMc72d0mdq7HbVHXpwHIM
vqPKaZpbCSCLP/BpJ2ZxuC2cfxCc50O0hK94O6KADmt0Uz2uvAHbitXt/qXkAm/A
ccEe3rB0HaHfjJF2Q8MSfZmiOdLQlyr09VPDlgdiDkTfjETFzziSJX4Cy1ioWGki
X/ieLCs2m8lOOyDc+yO1xPdIFBTzNmEGGtVuHjQHm7kj1/CBMfzU8gGMWbJI2NUF
PzWGF3adS4akq6/JpoX/bGoFbCPg65lIh0dYZ2ao8YA7JjDjx529sKUiaOR0H+l4
gOspfWfgtw+KKHElrNG/PHXaEpvXylnUR+eByYockFus2kELJHGtFnhLMHfGDM6G
oJV5hMfmnUolLjxIH5P3y/+Mr2HYm9F28vXG7Yq4pYiPtJ1L+I9ZC0ws2RQnyP2P
5RDc12E0ZamMx4Ed88Ec5SjJq3GD9xR03Qwj9yVlUHkb9dtVcqPM9fEICQRGXNXD
fpZt2QP1BcjuFWJjxSP6ugjoPXT+oLCRJh/BYLj1L+VMhZ7dCMhZ9RuyaUaptuqx
woh3P4uHL5o0VDiihnLzHzzl28C5Sk1ug2P7LUM8wTVUdg3OfCrtaPdY1aB8/BPY
WVOk+7G4nVc0ElD2nQkg7JfYSXjTLn0n6qF9gHTcKTMAjFGGZ3oacvHZ5tzE78BF
xc6mG2sJtK8QUvpGeQD5+jpCwhTvYj+eQdc+hDAuDYmBhyagSqw+asm50Mjlb3wq
UuK8defk0eflEaNYqpF+hrjixmzeESVjEuygAfTYI8MA8pc5Bfmi7RFLzk/r3Mjg
1fnkOmGapfSj60jLLf2bjyxKpeYCYZ5CGaN/pzQ3aJWP42nNGh61FEAOmHuPlppk
ytQ3SH/9iMuLFC6x5ZkX30/JoO29j9ScRn2whaP55VP36v2Y4MJB2aLH/a/bdMsY
2sbE3rIZkPWTUPxmx+Swy96sqZ3wbwcklgQyTjHAb+zjEY6shDEeyZodRPg7UQ06
E7rtSTIfnGVQ1cptKb+WOkEHflGjqg3sMbR7XW94FvkYj48uYpxeqV+s9SaTJd+l
WL2aJWiZ1cQGeRWtEFOgDnVtsYqWXmYiszcf/y6pscvUsr0RUNFlTSQuLoJzq2fn
Yg3FoUoEHT4Xq2O79WXLvWdOquz3+tL0xRqoFGJSbmVd0ow0sD5PI7Jale5FH09o
Aj+t73ZV9+5quJoCD3sm9SZiblin24QWDwRPoLOMuMR21DmpEIhNNbaMMQVY2twI
o6gsjxHVOMbFCPtIQ9zo1cfndYUu26c0jDYffg6KxSmVywFRXtMHJWB5YiHj3XOH
qXbEUn/fjTmHu2nFKVL1OU1mtc8OXhT2RPilaL6vULq8MZXs0QtnUUFNStDNZ+Qy
TrAsCmvMHQEJXhFqhQPaBD3kCDeuTMYcs7/B4nvd4/jZplNEoj850mgw77KLLn2f
F0yBqBaD2x0pi1STRugqHJ3381AyseHI6670CHDuls098VyVV5/SXDp3+ViWTWbq
fDhqsQEbnTdVYSg5Cd8zCTTcJxGOCSkJLX2kEfV16RqlmAoFoGismQ8dBNG7kJub
s5zn+vwzp/8y5TDyYm28tXMATube/EbgEy5omfNPduTVbT3wbR2vMOEgZIPNEdRr
/qrUDs6RtQH8gOO7iN4hQHSpsTJuxxOxOPJYFcUOw0/SE7J7DE7V4hDkAysc2jiY
hYej88IwVhC0bw9YUuI5uRrHgy92ir87Rn7FwXayFcsqAvotXYgQWbk4/bYN7r5p
H1GV47HdD0DuLblK2yjbhZ1WIGOuv3MQOM8X2nA6jOAG7/wT4BRe5XSHdABXLlTO
xYmtZ3IgpM8XoZ/8IueDnmTPl75UnLzb0Mz4yvc1Np5HqMrypdHSBRBBMHHonjAt
ItqAHMeeibnrKOCq+h7zB4yBkaLM4Lz3olsfxh4nRt4BfOIPkNXDEdEY1NjRMuNk
fI1yRM39sQYPrBw2hZPOvJH4k7QrZJanOMhMUvOGhLyy0fC1Md4I90jY7CnBQhlf
fYMbf1wi0kSD+ykrAxJTxzNiwEatxMKD1B79NdSfqkCQVxUJNTJfc0vSBCZG0kDB
eD+cqdz2YSvYVeFegC3AGmBhgNX1NwrAApW+SpAKMP/pJ/0uH5nDiuQoExeISTtp
SD2K8xkuCkFl68qnae7slq4fVGXBiZ7Xp/Jx9fJqcefeS1Ybs4S8NT9Hdctr0A81
bAgYP/Pr0kjldMlIHROHBV1PkxJXlWqZfmPFSCUh8cyDfgiZSre7VShXgQLeNxKo
lu7lxRV4MC2XjRbhgkv0S9fBJyAwNuPJHykjINavbekl2ffbVpM80XHViVPolhiu
XgdC5EPUlUaVZnChkFyHkKJ+qbQRB18uB0Y/6019hSXvoMD1bAul2D+iRc0FOpWC
GWvj40oJf02mVPaMtNwIeHOxrq5C8NhMarXlvYs3okQreP1y5RkWADqikY9QaUuj
/PN7SQnJq/9bK1D8ihkseCfPKIzYYuffpzXhJISNAodblPS1dV1RtNQH39my4VfS
41Q2ssi1zgUqT3Ca2+N7u7G8uYRrKWxpT0NOeSNEOW9dBQ+lNu+dw7yg3pFdfftZ
vEMFuBYazPQVg1VWPJJWH5Mz/CH5on+xGhaEOX7D6iUblebOTtAEQAKOJ31Jc6OT
CAutp+emnu9dfjguH6BKk01o5DqUs3zuFwjNQE7lC89y0emUhv0Lw4UHf2DWb4qD
f5Vi09zoLtVK/K+1uFNHHl54arExdyZXIQplxJS6X7JmT9IZlO2wrbi7UWLM9mBD
IamvfXpEFpa2qx8nEX5op6/z1bJ9m0/aDbdB5jl+a0jn7ruf7+4EmEYxerd2bgDi
ubymjg3ofAn0VdprNZzPkHathi72yme7/KLnPccBu+C4P7PxxuSzcDestUFJI/om
zd9ZUXFO3P+kaEOKwZ7P1cX6JlSC6RLtuc+0gZXyqoqLF+st2E5XqcXXquCO7lT3
FAFjd/Wm3TcpbBVinMisIyFqys6GsDebpLH0BCISAPMFuzqBDW+AJgbxurHLohgS
wk6RD/IkrxJjT2DrB1GeSjev40U2QCzpvgmZ5zfqyRpsAM9dOC5+LbS0vuNPncHk
TWpaMyRNv379RZ1DyAP/RMQD8oyZ1xppaZEIu0afcHkICMmD89jBvq7XkBDi43Xi
3igM4sn0ubP1qZe4useKHN7u5IxdwqJ77ie5k9vBnR2Fi1zCpuVBEaqo/jzEDBHM
zp088ZS2jPPJTmRnkTLQp0R/TRiYvRUyxk20MZB8kS+2gpTlICL6xHbBBFJOzCl+
XgXxggKkTynCWBmgEo3IUlbWvM0/yT25REIV/U3iFj6Weoe0q1EsL/LyANZy2YOc
WdRAVpPWHkIWbWXQs8rK/RAf7pDunuVIdp9wG9QyQVILkEYhSKpkPhMmZO97Ygjp
WKF1/5niBlSliQ4zH4M6RJOH84p7uq9D1zHTEBPCpxYcUu1C8Uvd4YGurDPmbApD
YmKJmFBp2ByS5a9KwWbG6B9RBYv7K7E8bYiwcxcY35xH6NBoYtxgl6CI25q8VLES
q6iH62l1DtBMblX7SOjRoFrH0yRmpotvsUnTWCDanKwQzjcpE99p5ybRKewTpKbW
UkM9Klb/J9tD8mmdW9U1RLa6QVH8d7HopEdkXcbX+uxPH3KEf76fuwOf2KPP2e15
q+qA8vsvnaZRneZUpE7S9jEdYtyh2dDp/GIaYPlhqdQ+HflqACyzkFW4QGdWoBcW
lHOHnJ56nN2FaDrj58LRR1xAIMxqrXGbZkUKwyuk5/n7JtBBuEHOfi0QepgNu2vF
8ssERItziCYHll/00fVrkMFljQfdaL4ajEueSXrWxF3sSjMlC9c+g+NkBEG7Nehv
1ARLAMYNlBCNlkZM22ATRQq6WSMdpYLvYASVq3P6murcFMhYbxyRc2PDaFNAzOyE
Go+0GBRqAeJeLLYb+d/S6Q5e2hSRlj4QGsXY98rk5RTzrrCGa8SJBkjjTjM4BK67
5l67WmV29MlYAg5kiKVaHNZXCTXwRHkdwW5QW2s6bsFCjxa1v2QupK/QQhsV1ov3
QqVbSyvZrzjXXOtvizE19fRd/wono4Dcmfpp7kbCnUUnBU+r/yKtAicaJGrvPXN6
q2OjaDcn1Qd+pnQMngFMANEnUcBfeqGDssfVfokntR+Fm6j3E/xgSn5b6lvt3461
PgjwEB5q8kFHI6cA1UI9juxRm17ibBC+MFxrs0cOMwtds8UN3M6sMT7o1ncUwm16
Ocsxj/L2Q6Q4yiKgq/9lElXtRWMDRPX3GOw2fq22WqGaCy3J38aJnsniRBLIaQD8
R32xIrMW9F/i3LkK64gfUXr5STeUIxvob1nXiKj0CFhbzLVUT/F6sI4hj9Xhpv2h
vZxmOOP4ZLY9UU4miNRwIQxtOAvzpHOLIz5e4jq80hz78RUs88AmSdDlUB+YvuxB
yEpRuzaofDB/4Wo39cgIxuuaSsG7LP5QYVwFxlyzg9L8l8MDuiJ7hkUFUTSycPCz
ghxGCygO4TB0yM9FDZ/jzVHk1dVk07Y9Hb1JmS78JO5e4Esf8rMRghKYdTZIAYJ6
fTDs4EDn03hlVF/UUrDiMoKq9qbfGV87rVn4Inln5d6niMlxDjqE4vlYvVVT1VRP
mK0VYTZVmRazgysmmVmj6dPJUyRVlIiYBQ+CO2hekp5/pEinClMTsM3G8vWijwmF
wyssL8gfK4jn0aJS2HyFm2auhIi4xmL1UN+E9kM8VZtestxTkXmImvaBqFWt4pas
cpAYyOH0zwOrgQnBdMkskE1ZgSMa1qv3HuVgI1UKiCWXoFoQ4kx/zTG6uBIv6xRK
/2+/iBMPyvYeMZhM+56SWzoLBNEecQgft0KQ9WxpSihCOPDkaHCkh7BT5mZ5rH2h
i6ET1xRIT32zvYYvToLVkiSVZxDP3DNB8Gb6m1IGKmpBQFToVOuxICr7xn1fCBJj
a5uFQsUb/pSea/fytGQGMinmdKNVm5a5lXJcgMw9MLcClVaFKm2S0rzKe4oqDx4r
SlKh5X7zvF26gg11OH/p4O2zlnj/frTdhdmFqgNPrHEb627mQZb9FyXrkbRrxMHJ
4abvS7YqGeQNjk5eEaloNUcfy/+mdguzGdC3U9/kZHkKa6kBOrSqkOywn+W4fen1
E7RSdVBMrKyb0VFMGZMdoGiUOS8Zh7swPynXGH8Ld+i74RxHeHMW5rVswZv+nnEX
OCAQeqL6lr0B+zQpWe2fOrzth59S/4+Kl+ScyiZ7DaBO6lXS9/V+zbLhh3fu5GeZ
D52625/XW9OswcsOyT4DlJBZDVSwyomQUjcGXaxX40qKrV9I5qwey6BtgOylM6Vd
C4qje6fyssxW8U27v6+Rn+dKFxqe4pGy6+UXCh5QYwWhvWt/IZtdrst9sA6vxC9X
r1F0XQsNhTvDh3IJ5f9o5EOiHv9+zNNqkAjOspyy136eZb7s8yS4EB5+D/cLUWS4
QxC3+nI42JXp4i3chESFTOU3t24hhVWi3iSUxBku8mPVmpOKotL6AVJfRug+u5G5
KtwtUQHrJ/aCbXCp1hUwh/bDoXYX4g7bvjx86cewxSNaxaDx5PL8ihUw8ZNC5s9l
PI0Gh1agBCWCdQr4VST296TZHUGSlMeoSdZ5BT+eX2oHIkFDWsGlQjxQ1j3YXGlw
chrMLDjuxaPH5WLfB6De51+nX8pScfGGbkGH8chO0cQX6VFRmA3+csluWUSDdW6O
Z/ltpYjP5W3LLUYtQhgWoZf3mdQAFhGC6EITJLPfxogRYXQiaRRZ3ZCYm8CzloAx
hAnMO2aOb84R3/0y1GP4tXVTnXWNs0FLN4+hgu/3WdFcZNOy84CK/wkfrjkznAQX
4X3uxEcKuEfTZ6ZGEg82/VCMk3PgYEOavaqBrxcweujaAyE27BUAEYVr9bPy35FI
RpXKyANSSwwoyMjEOdJJUL8NqyQqKixjugTaZbA6BEhMGFnjJrH8JqLCMCZUVkwS
FElyCLK1p5RgIVobg0MjWG/5V0Ycr25DnFkcjbRRwIzxSf/TuqG8cO0V0oTPjisa
LX3rdv4gN2N6vVysn3rrHNyf87NLYLOcB4i49CrTDR25NZ3Mf3tab72X2mA0SS8R
t57N7vUso3Vzklwe+AjW5Stm1OtVoq7EM+W2pvkUmTNUzz/QSV8XhxMVwJmwXDe6
Un1dpNMRhdQ6VK2XICRqFxxAuSZTZJJbb3k2vym1k/5PR22KiSovKRN5+3NwKtR8
IUqeCzmDDN9bir1gXfZvwVEV49EOZ8TfS521ZstX0CXODzK2Z/qFg8xpmkt+kudL
Pdd8krvap7mBca/bkxUnsX+tRuNQHoTtFFJLQ+msCjSZyZCfjBW6s4xZ/MB4dksD
9w/LahRlBAP+Wn3FENTd3OadYWWJ0WRs/goWyyDTn87ZNR3n8A+6lmXHUZ9D1O3D
YVYOWmcMsVBY8lfxGkP9T8rudK1XDQX0XRjltoZl/j/plDKLl3qoMuubWA9uFxK2
VT52uFP+pNmYf0DqvIUa5xv3ms2ZWKTEW9jIQpaBNDmDr5hheP2O7fD8RjxCT7Qt
J1GvoBxBHgVgKHzuokEP36f/XZt/ko+3Id+hF75fZ8eZEcfUbcF/f7mk4pEy3zj4
HgWvE2I8BlqDuzBsXNpYR6vl3QZD8DP64NX3U/iPKlo4Vna8dr+JA8kzNDJPPNvm
EM8DZVpzqeogJHRvL5q3XGS/AnaFgZxHJ7t2tyX/WDNRnHGv9/HleVqmbgaxdXD/
Q/W+M7DtS47Jd60QtqWa819AnDmamVRPLjrDwJqjNH0v3gNzu1jtS0orGFeFXOxv
X/pifXDrjUOrOzkiMdtNYXZmSIRCBHPILQQMPoB5HmNW5oVMmX77a1+UE0Qp/PQd
EBccgyYQQ6kQTnGbjXyH4yj2X3NN+lqgHF9qyFHAHz2S2uKYTYBuRLUzOkG/mvOc
KUEMMBqFiJJCxgLQTgUIA/RZN/+7cK/A0ghYxManA6VFSXyVQAFzc1odcI2rvPla
d2mUDwuTsL9rFMzyYZyLEzLLbbjGU/KelkRsG3GPYQem+zRDo5OXI0FQT/FdG8HN
Nv+FBWO3P8v3zWWdJIHsGbKGVTB3U5t9x7dpVJ1P75JH32oWHiK7xav+duaNcRN5
5wFRHomUdoAIYMudTzbPawR2CtoMmz+Gpqi45n3fOxWdlFuup3TcXI1NyEIQhFHK
m+86CbCJDMiGmsy2BoroH+dJb/r8T0EJuSAAVxCJHKo8dJFBnody3BYqyywTViCZ
dOvvUjFvhdkZFefggqJ68tA4a6XsQzzHqDlE9iJ3r/pLxkzAzWzK/nJujge3CPRa
JBGqWp9P1N01z0KdUV/3WF3bLHvlH8U9G+fxR6GLdBRSBzSKXX60OZMJeiD5uNWM
KmQpvwQwbiugELURGkLtFr/Su+Gt3YEBsZry+HYo8E6Kjip8nCyrCB/qO9RJycPG
vYjGQsdlQaqrdTNx0P/dkeJBNXvVY5307sJDLPKF4L3W42q+NsZ1N6tH25c/6uh9
1ix+fwLOuYWlUbIJPxu55w8iJrCYkgvP9aLZBTr5jNal8QrXFnPr/zcLcSZsKevX
gKi9D9ZTq2hYwiX84yG5vpbOoa+kI1JycWmlbd/HO0dJxEcCMMWNvCT59/CmApjh
x/RknGuUPI/QHwGJP8ZKrOZzWCkDF3M9CaAWcXaulZFa00aI7IO2Vsoa9VGRSZom
lg/AatnL39kTgs66oXwuFudfVqU0dgUstSlfYn4fx+G8uq5QBlbMS6lRAwGlAlzy
+eQTnYacEdVoWRC+8J1RQOPDyL+ei0qTh9nbhHuVtXCoqI4ER2DwkBx/+KjqBFG5
62rvpMp2lztRiVsJi4mvsvo7D5DXlBNfP6vSmEZP8hik049SGruPhTWoJjCD+hEV
n2BIEefh1QS1QmAF8tyQO47sV5ryRxl3TPSaKzYrLWFQKdpZZCdcy9f+WPlZJg2c
BoZcddItPucekkIR/Bc1sgRKRaYTtiYxnnUZDH/tcDzOkdaMslCZh2kofZG4g8dD
0PF16Ww/9KJPMGOPJghQnT/VBdbJZgRReM0atWA+6uSErKiPk1gH7O/hUWkA94yA
Qf4Gew2W/Vi6pHv46uyfDvxDwECx8UmJKT31wfy9r0EdiQnXqbAqd7fXp4qzmJem
OiMCTwa00e12Fwsv/KGger+Mw517nI+dMUy8tuKl4k+vL4sogD3zfv0dq9VEFq0g
11wD7FURwmXan82zCKL8jV4wR6ukWh4fXT69gn1BV5BXt9+6ocweaikhwqnxCs2H
QpJoxrveEFOPjYi4k4Ncartg9SpNRodAtMC3+uMUTOCue7k5HygB6SSNuLpFq5mK
80o/pbhsXpNdmRg3AzPwtIV9QPEQXzoF2TkCtgFv1YMxrneh8fmGcR4SdYllKFnJ
eASIqqM6ypkLmmY0c0+N3/F5r1NBLbiJRY3rKhphLou74axVErrXcLho8VWkcQmV
ftV0HKVW662GCFqjbXGk7wtp/GzsBAbVF1KmAICvbVraH3Jvs4Sqs9Ng52181Dt0
cmACIn8CR+nzpbrGhmEE7pgGPFruItSggIMabDtYEbPiu3UbqsFiYAUKg0lWkx7Q
JBtSyGrJKK+w5Qh4j54b9W0fttNhFUALEZpMj1yhbXM6tywjE0xrpFlcKshvuRc/
sqBGumeLw2STGbDgRh/IJ/mMul9Ayiepm/dv+CqVMTXZibj4KOxEzxNg5mBbAxLj
YkbumF8T3+6DS7ChfGxyiq3PIOLxbcEQ/h3FTS2lSiREjCMYZaTXQCvs7v/7Cf5B
yQYMSURlB2iEpGjFpRVRCdNZHiuWHaitvNube6zTVgaygNd2K5n5UJJ4y5Xmbvrx
5tfjG1ouJhIMMGztypy07bGXylxNUmooi/WMLdqwOnUYSnpoBk8iUf/GEVT39UxU
AfSFZLpIRd0xzMKXqLcG6a6whqfUZl/4/Nyixybmf7iHdgYVLGkwEHgItfCkEE87
qyVIYwY3ZgO0SALqd2TID42QZq4+OryLsBVx1YwQI1wu4AOZiY4wLCRGOQpJ80W+
wk+R558Y9y9EH9VwSfs150f0O55L3cjKgmcRtzrtzEvwSYD2sY12ggJPDfWhd+X9
rAPBmdEMrzCC+IfB3SngIFLU+Ioz/M2Gk360DJSLW2DB7ZXyDRgx3Wj16mhomrLO
vt/87gtCxDEL+bfZqp/TmOCs9Hj7HfQRozam0oh+pYJ738AKqJpgE+cIYvv0JFm5
95Tpx03Oe6f8ktWzhWbSwXHaJaGv+BrM1hsxxkUY9n74D3Iy/Jt8rJCL/H+g6gxw
zv4F3UJQINSDOvyLJjZTLVCiJuJ2TcB9FCgab10QQJw6tMPzi3VZ8fTYVV5ikyr4
4ojYDVNpiSaM0EGKmrolqchdi5aMZVm50FtYeV/QXgJhkI2QCgdtb5dlOGB3R1HR
3d32giA6jcVlWddMXuIQkA8H5+hqgdTZluSasHjKVywe6E/vOf9mDITQ1zx/LDIX
BiSdNXuC4N/cKWqy1IJoO3X9yo6vT6QRjV8LrETJRWnWUbA/bpyjP3rM1f+vednF
CJt+99JjmfoCAK39wiobEgi1b3zFWwCm52Xh6Uf+p+Y29F+ud91LQBqgNA2VynD6
/nWAGsAMKuda0f6vrovlize+qepZiWqy0Xp5v006XY5vYWPiO234go/iEKA7EnpP
n/3/+POTdkmXzJNpjju20k0SjEGR0LCeGaQoFuD7KdxkP2SfL0DTkMcgZNOU3CNX
uFl5yx7SNzONKD3/PVx7KfqFwnlnum4V9ojbLpt5iWCE6WjiFB/iMq7m69O3xI1G
LWGjsYxjIFtUd+YEObusJybt4N0U3BHEQZblDwoB5rtCmQZJP8qwzDQq3ORuc2zM
OoWeUCh/OCSyQU0wTII//TZ0KM2A4M7ciZLOCr1w0QOAHXBfBzNxNOOjOG0kCBWS
DzXt829bZ6ynJHTa+TekbZ999GywB7Mq8CIc5tYDhUQ64Haca/o1ah/77hzYONYe
WuaXsRqUxCjM7xpGUnfXglvII9jyjzshKrRJN7ZHbsIi37N6V6++D4u0/+EjKQGA
z9q8od8QIDTcZXKcRrjSO8THHEH6rbN08c+jSCMxbvWZSfD2mwcR9CgrK1gXgG/Z
a9UGmn3l+HI87QwaSKEEM+kEgPWW/sukePEOTeG5pOChqDdKLYSp19uB9oRwCayI
IhnLg5kkV41koCA1DHOcD0elgvlwFVw0RKimjvrP43SgIvaZb4BV5RGuccMjwjEc
7MqUa079HbAy3T4rdKYIXbG5xgPpGFMdFOQsi+lDshOmAmIBbOAhUGZFydmWXJ7l
MBuUWAdiugPdFK9OKE1T0ATfYDZNLAQVclFV/xCXxMjnfeBRkg0o7XHB0bUwmoNo
FTBfNDGS1j+xkAySQkvXhL6SUOcmzEvmEYhP1LzM6ml7Zsb2OR1fRl89aPWC5fIV
97MVuWV4kIaU6nY2zN/qhsbF4ouRGOn8zgE6JVOIonm6xkNRMmZ+FdAFlxfvj1tV
mFOViW2dXvMtu8rqBD0+kr0XgNWvOfagwRvLTSHfAFE2/xBP1iWT9+Ie93QVp2cv
rgI899hHvj2GymFKOkEZjk2885Ut47NQ+IthB7OC5LaAtD4cEXMyPhef/CbJ0NEn
r6dc10lds9MZv35xvVUEQUkGyj26aJOXYJ/U0JLDn7s2K2hHU6atQ1C3EFfXrKv5
Ms6RsNyLQwZfnYbd3nbV5uaw0r6seVRUM4lAvYyOI8LkyOX321o8p0fN22irztBg
CSuRZ0RXMNH2t8LDRoP80AmtSk+oMblp9bT33DKMLLOrfjO5Sx33rVklI0DCdXAB
bRR4eys2IDBUlsngSrN+yEe1ygm2NbEaoQ8uCXitroogMD9HxZEqjzAOtLQ74Ltp
plcv4uMFkY2SOjZOx5NC+rNCmO55iG1/+WfgwEwalwzpSzdKd4Prytc/58SunNv1
m/OW+qLvsOplYd2KcHCYWfYP+s7iTdFCvwgcPuM0xCKATzb820XMGFSy+DGMnkIP
aOHaAI7jiGd8/yFa9SvslQPQJBa+/j89/5qktLtTUURWp/tyMSCHSisZk2O4L4zC
xmJ4vm76yKajR4WEHuOD/Q0IF+WRr+H1vx/zYPZsBwBJLSb8mcD7GlJz21pmEYZq
kTr754DLK255pxtIJc3wMi5LpMl2GLx9cMmyCR7LAPmdbHoYronqzuNN39EgX8Sc
HdN0fkWaLnXlq/HGnp62edEFC3GiHJjlJZwmM/aIfH5dQ12/qJEB0WWYGk/+W164
OKd/xL4jY8upqcSBpiFliJf68wn2NUUSMyYQXdDMWLAT6JiJ2PVKLIhD0iRj9Gh2
79ogllnHYVpuXitRSdlwReW11uzVC8aeXI105Uvx/zZP5TrEYLx+Wmv/EmnkYick
hBAJ+gkKpjyClGEV+OJcMvy6kiEIV6qk7tyuG7yYqMI8RtFziAivQy/lVq0sjEWv
jTMFakMCU0/3WyIUbFqoTrkRaP8GsYe6t2ERhR8qOkzHzX+WPO+x84XKSEJmQwKg
Go5xH0LSzTLbZnrUpQrjHk/7cSGt6rojZ6YHi6wWedXq+wPyK2wY84yZdzt0mrTe
10xYf4QM195xx92BR+l9kWUL8VQPfb3oFadVZt3vAAMHboLQgsOVfgp9SDiNPVK8
XVBQdxYoRoBAmJK0n+8sZ+g39RASuFxrT7Q6OucOQxLLoioPdP3atlvMaydE2R8h
39QArRHUQphmkU/K80ANgU7vw0NhBr+2I0+uCFGpGUq5Xx8Q38xSgSeBqFUWWwKK
pOL1zz5PRy5BiG23txjjOiu9N8XJ/j60uJwiFKpzRyR+5+P/3sIu2pIP+Ym7iP9n
2G8bTsB8dcYOthQgJFpGIQtU3pX2s+dIyUNPsMiqAwwG33XPoJpjnJtQOw/S2cT5
mzzCGyZDi2SZr9EItVNhbOeCl+ZhvyX592QXWEil1kukcbkfaop/UG1jRy/z5LD0
jnk7v7lxekXjyIpB3+Vwqvc7OYWIqmCOqs0kuWL37QeMatPnI210Dag1x4nr3nfo
BmEfHGZagWi4EH67HHLgwUfnJGkJsJSJrk8cOm123pZcBlo8RzVDEO0lBJCCyU24
inVfKouHmoXxBnAnb+B5OxOU+IArX8fafyVclgxZ6iMRLyS/h7REbK7/8EowBVqT
qVsa0ZJG94unLeLvlUT0CZOVPjZUzDwE4bAH95iuUzGxzHTJlXrB4dmwpO96Cxs3
bpnlg6UTCk9Ps7uye+jjIkd40GnTmrHr02sA9drGQ1/xOw+758P92yHZSX8K8FBd
nJX7VMVnxeMktaqkeoq0ZFQ3c+oq0C5sZqPE3P7gTmDq1f1TBxLnDI5cIdQmvYl7
U/2enDhNqP7tG1PnM2UycZGuiYuWSWpKwh+0hgipHBTymTPRw3bYl8Tu93iVwD+X
LgVc01TBjLppe4pnedfOys/fRGsQQOxmmwRay4YoVzEo+cdS9VggAR59WVb2SZqY
mpchgCwHLtTI07dhVBRaKvLCupF07KNPENzdo9cTqDHuRfRWZ+nJUGJzSFF6zLSp
PVEcrH+slhKy0qewh0lOFogkHOtwo5J8UvTvKkSUEwjtt0i06ixqIq2dOcmIsB0r
byJYxbC15DlmAlpg36bEnQtFdGD/xIh/tETG10W3RRRuK5+SmI4RyHvYMIIz5Snh
7iovkKz7HnL2+ywuJdH6qL9mpXdJ5HIiOh5AoT2UexsHB3JvDroDkioBsw8kKNUD
0/DUrdRqVWxnFcp6eimgB276XYbu8o+I9nehYrpw0ea51OX89028nQR+VIrFlGYX
0Tfr6g08HM18vXd9/IQLhF5F6s63xhEOdELN0IMRkp/vYtnoJ8us0KoqlOXpHqrg
kfiZN3Z5V0fz54EUWuCRFbg1Xxzhz8L35KuedpyDvJrZtPxmm58DKTyyCMbPrS79
wIZZCuoKR5bG1CB6sk+WF3mdgxUFRYm6zMoxbgzPqKBJNRYMPdeCmbM4rMNP4dix
LCl/XGIZOqIomInkxK78VyYwswQUwEIAU+bDqDGC0kjePxGj9ailyZe4GJBz8jfp
NgXLzjBr2u2iKHVfy/uI6FYwVbF1L1PI2Q/YpUoMjPY9k7//eiNsc/h9z2V2QmNa
0QGoxx/aprM5wdT/JqPHwmvJlEGftiS3eTK7qdMMXmaoS4n3yVJsbPj9ZCyvjT2W
x3T4u8XkvN8Oory8e6LrzEwYqfom2RmLchHimfgUubAroMCA2S2ykcldo/FTa0aL
AFKhklBoZHUnRgwfwNvtXlLVe/+PV5FLxUTTZLOwQhJsK44k4VGXPEdI6E2LjFIu
0JcHkkkkaWU4vXh7PKRnz838tfTFsjNl0UCML2NS8eFWeeFR72HSf1SQuHQZEuP3
0RHOAggKBI+fGElT1t+Ay/CTGvtkySm3aB3CiuCjsyDli2URmbTpNmJdsL6NbHdQ
H/uBpjn4Lmy0fkCzD4cDDO4TfS5EG4ogE54sP68rqOlI9eeocJ7QJJGWcbH5yqAP
neSVGMlkkVxqle5GJYT8Y+Li22/0WXqVcHqJ26/HJYcgqsR8h/Pe3FOUx0SEQ116
dH54foxT57zbe+2ciYy7sctXsnYXxl+EEWJKGI++biYB0c/mfkzvQBsP5+cFoFQB
wAwrjYcIH9upqfZ3mK5LVNtyAZ058RfbAv5QvrqDSC8pD7DrKmm+S8tItfjyOG4w
r2DqQhAy5Zx3NxXE7jkdqwI9iWtTczxFr706Q+9xfCc2W7QmBDmFBulDI3M9qJBP
R3g6yH++drIFv168kdKoX53W2th1l5rz7u7xgXDoLuwsMBvgQm42sdbgxTyVP4P/
JnK3AmTW8kjDhSC0MnKZIGvtUepNq8SDV/bTp05gM84+ptezltEGVU2QpAZiPM4p
hPweg+i3d/qmwdhByLn9AAVisqHbgz6LrGbRMkatR5f0dodgLqeAaTeI7v9RktzX
K/OfIXixdeWNrmlwGnwPb3UjMAvmONFZ+5UMGsLRYQeB4h0dwJLs4rkGP5md4Kkj
0L1bk8apMWdfy8Nk/4oxUylobSc5xBfoaRF6S1n7lZEGtfhyTdxexu0PvbsHlmnW
qXCilSfG3SxS4v3lIwILsBNNt43JVgLCqqZCFBp1hRfZZkrwRVw6RqV3LAtBx1Gl
tfmpUcAxSZ6yKrprrwzgLfLkFFzsbDafKoXyguE+Rb8MQzW63G7c8lhX+6iyYzI2
XkQvbQvL5wSTR+AxoD2D8RQ7nAjyZPU0knGqXdI8g70bmCS+Tv4xvz6hfuqeFDBG
avwrGP8lKvy2LwR+XXzRW8yns9/vF02wfBl9+kMzG/Wu2ksc41z6T1qnh2kwiidg
kig6Em0AYDCBXIOBMqZHO0+vw1OK6ZQda+u+MyfH2CJO35H60iWRWoaI0XctyOWZ
5F8a1soWcLSlAHx457AbrNTvHuDRyS1Nv2or5i440sXslbvEwXJ7VebzNS0cdf5Q
nBlZGELbZki0qBms5uD8uks9yg2ihX5qo50CMkWhzDmvF329Sqq1CftBfIaPpqd0
rn732FuF6kIifOV+YtYQSVrRwb3r4/mlWWfcV7Ho8AkT0mes91DaCCzgyhMe8c+p
/4+7noRxTA4q5VfFpQSb4ydrFLRG+79A10zcm1DXEpYWB+LtW0PnqHqvbTYvBnPG
jxwcp4QDO5TyOeXcY2S8OlAxueHu8riFwSKBrrWhP3w2b5Byv38uV5OjU0kgMOuU
9TVn55otB9cx1k0C4NTo4BF2sedgHXPqv89ZcwLFjPkxH172I1w/5QiyhSmkd4oN
AQKQwjHsptS29uaeX7DghEE7yDXwNB5Nb5BKmjJ5hTH1OMbh1iT6lX0g1Am41Ozg
lypiLcSvVwWyadwL561cmwUdXW+6gdQkSasoJi2uazCDtMaCxo/q/Yd3knLYKTju
SvPXC7Qv+gQX6/XnALw7LuLsD3+X8vHbk+PnVWwrlMmM0duQ7jVNLJNShJof2e34
5JZIq1CsH52P2R6lLx2Lf3Tzly9Sdg7jkw7wiWRDU7cpgq/vD1YYjQBB/QonWbNc
HaYPRY+XFzyUiy+bh5INqdrFf9XtbjD8Ybj6Q9lZh1YblbUCAE93FgMF3wKtYp2C
JnCR8WSvpJgBoIBf3fv1WcKFJVnQTXiQszrWPLAWtA2zNLzlXV8tQPXPavDNmQNu
Z6udRPQT6UsoXJmBlR/YLcVT/HQPCe4AYle6t4eLYtFKXY1BbuKWQeg1zitD8F2t
un7EX3cap55p8kkYGl93uc1X9JI0Et+5QwGVJpQVgaicwUDpMmWeAx/X26qeCWIv
qnuStsLS6Hw4rkhC95VOAEHFjrx5L1Rgh+Tiw3071iCZ8GHrN17WLj3rEETXe3q3
Mdav0/nJ6TQqwq1HAw0LIDQk8T+t8yNa8mNKIjbSVECR8S8hJrkVkRmsrEj413a6
uOArcmZ2mJvC2sfxQaixmxNJqreXw+1IivbHR6hWx8lcQbwpqALVxMzd+uNyLT46
0X+53PM2WddR/bpKftw2i746o9AGOB08KnSGX9a0AfuZgDfQQzxCw68E8HfLhJl1
xA5dpcmmeL+mOJwIu2SOLa/+NVU4vQM9lTq6LmHrDcgJidss3hy4r4ImuDERWwR/
uYBx9TNM7um+SM11m51r4BWGsV5tVkTQOiehxIPHwirng0GrCFsmwW5UZzKn0Bge
hr+WLmbDPfgptdlykAZkt355SwIsrJz231JtW+tlu271zLZnWW8yOQWC7hPREX6R
dih4i3JIcjp0fk4JQkfvmnKhmguhfX4U8/k7Wb2t3rZwoRUvb3XS/lHQhvWW1Fqc
SdsnpnqLyYwSsW1CtSGLqFrjMe1xvRYtsWsjXd4gg6OkrCmeCskoCleKpwGR3bsR
be+H6g7x5LYA8+xa3beWSisIwRDT0G6ubQfrW8KioNJH4oac7bufnJON6BzOjwu7
8w3yr67BN5bxxgcYqZyyHVr3uzbme1aW/yABzR6AurpFTuttOteOt36SiKhb6q4i
FTQl+/Z51qKVc0KWwx6nlrwaen+rWJFU6OWEY95TPCFy5ws/uFOPpup86zIWkErR
BfKLZ/f6jJgSbnwAd2VVaGdr+CgOHQfiDhmytqvrByqao02MgPIta/A32/h8Jkld
IX2tBQJEZTsIAO6sShhhuBFgrXe9OM/2DbQyFULZbWcxg7AEmROAmi74Qey3RX72
6YEiA63fjyDxxm4s+Tp+pjjYn4REHOd0L8vPXwFescxKW1Tch5/03rggfAHZQAd0
52QV88slF6MJLJxoSnrLl6diHR3164sRTlJJdLMYQUljW0A5ae/fcilWOS5/8OxC
8rX2g5bsWjMpcWmZFmJynqxLO+rqcelKT7K9qkJOvi3D6rFkTyyjCwTmIUd92Fqn
yiyKq6uC118H9TLJBY+wgUSC6IC0D8mKDbczRb1kOO/5GzCUH490CHIOj2OZdfGg
OJf3VMxw7n2Rg/j2dm9W5aV/ZICJgdQDLVgjk/G0lENyoS20nhzL/Y/WVAuw7jSE
Yt5sWn+/TYI/rSkMA/b2sdUVxYM0iRYVmLn3Aw5MhVsbH0cSkhSaGnk7uPrQsFv8
ryJ7YlTKSOkYSm2HPEYdkLobeepauo/8sW6X+u3HK3Sp9MuOT7+vhD5wnTo9Xr8i
RLGsp+1i9T/sOCrouN4himXdazX/LFfnD8Jo5JIwVEhCKIDwjshmc9m7HeWbSFrY
Bbj/mkVyPkvM4EV2z2AZmE8NwW0zLTXHeHe4g77MNzRBlGTNagYKw8YeqcldIBe4
lR1U6b9k06HOt+BstExg0WJxJZjMvwI0dn4WqQECFNjyG99Yb8GJ2AYB6tfsnvFm
qpALx7d07dT6Z0+/y3Lyc8r/gETkPaAJM5dmD6GaR7Kw41HtUpocfr8GzAi/jZwS
WuSIi7aT8rGIpG2ZTEpHeFUys4EEvMdlx+tzfbOm2ge0IBfmfcYCf3fUvA+FB81C
ISPiJ49iMX67W1PsJRBTCuwWxIdKcs/1UFBXrOesyjAgqN/JSKhiizq/MSMCxQ7n
zBdIOaxZMe2Qpw9DeQcwunccbmbUJk0AQSyZzx3GrlzZDhZ8zOh53PQxr8GqAr6I
ZeEioFv33Wc6w1Ql94S+nyulSEQZWIlRKkdBNaIpla0NwQZhlcUpr7T5ZOxfsAYy
mKELnXVBUhhtmJ9CgSP+Iiy1uKM2gfQIJp43TmojdI1gfaf1vwM74h1tYMxLk2Bq
Sy7qGBDR6kHzbEXf1fUh5QSLRA5smM/N9qJvCTgUig/JHAeW1pnlFdrH7N7Zv+fV
8csa1kPwr5CWwnb8mW3jW7aSqu6D7BpwKW9fnOWQSpFnQ1VpvAQfCaXddt7B3rwg
+sxmZkK1lBdmGPTJn0s1Jo01QvFE6BDJna8ByTjNZpvjx6znPXeD4nbT0qOImIue
yp6SHGn3ubhwDW2eL1c/VQ+0YfRraARBwbH2QV+9aicp7wHPZY6uiICQ9+n50vmg
Zf/rHSavm0FhP2YgbA2FLmYq13m70fC0ndVY9CeUEuTKR1HdIwxOi6n+qcw8ftFO
t0q/b4ixZhAK5H0/4Dv0zX4xsZEhf4tFOVzfXaZJm3PNDcilzTpi/y9b4AZ4s4WK
VCvV98dclc+Zp/pA11h9sdr96zxSKg8GAUBcs21S4C1699X7WWTcrrxsDgGXvK3c
ft8cdPnx9MIu1iBt+HgqdkVqaBpmGUJ0uwhm2IQaXG8MfqxiFr+CNoIcEUX8hB55
KMN/jxjcBWD3ldDrs/fG7ZK+x4wE65Lei6AKIxT9Bfez9FFvbxVkxF8Qn3Mb+BTp
Zd7Ub40v2qqtOYP+jfGRsGYkiwvPn8Q+PMcmL3fvDzcU38iCoZG53XKs+OtlZvSm
XkS5/CkkpH/+CttVNPN/vFJIKndt9+XtPLskR2wiLafsq3QjKqDIeo8iz9HRiRHT
aK/wGUQWZWYY5rgfi3mK2HVfDQsyJU38iAxJ52EjfO4Rv5bwEGGb42z4FBWE5Tz6
fJuLrgGEExQsZ63/Lh1JnF1uSHaD7lGX+eHN0+LPc5sXWleAEt1KEypoWb7/551j
8PQaSmlF5JKYdoxB4LzZ0NTMret5gg2dwEurFqJwRNSw3kH4g5fMocn9alUKuQIt
oUitlWETSs4ieL5Z0LqTZLzso8cfWQytTY0OMB2hgAZn4FNQyVrgx9rIQ1/fLCOx
74462KWENYp77/We8gbCjW5wk8HJxEXcHZe2YfFEWxIijzr9NU9jZQJwKnAAVybM
mCu5D8lRtQR5HWs9NtjwHssNqnj2Qp476WTA3vKtCIi0PPfDwkH9kJ0ZlnBovCll
te0h85Y95nnPM26exymLbrMzxMclwR+ouTpcZl+81l6M2HJbPXpata9eRpTeYwuX
YHSo1P62whJ7rZtFhqg7aQOqbDze47bjbc4B4VDUmZ7vIOzr9jiDx4ClwXEHHBom
OE2R6J/dFAs8vs+HP/2K8ir2vI1R5cEe3PCad5YJjI7ul8kbXTDIyWRsmNazAI0h
NvCT4wgZW8Qcvyf+3dtYQ30RGE3QHVAEc+deGB0vQQlebBVTR83KBhoeUQ3liNQb
8rxnvpVeaDhh2/+4OHKJC+vKDsfiiyrBpWdtSmrinM26rmojVgwRbe6i/MRl1/6w
L8Q8bIioDlFMbttn7TVAhXFuSdeMjVmNOLtv5QPxLAaQRv4ztv4QF4K/FVh80/0A
a2lIl/mdeTKh72ipOF+H/HciWH96acMCwntZsg1mi9JB/P5zf3KaZFfo6snYcdMk
H5KkVMv82r4BJo+bTWTDFHL21l4Sva0fdMscan6WGjNjTptl+Ogw3wuitk4183lq
Q6DouAK+0xEsnpeK56EI3xxcW2AB3Wu6B0u5St2qusJUGK3OKMauTkufsSqrDBej
048dJcb4E0+gXL1se1/U+Z4+cK38j8r7+SpQkj6nBEzFjZ0meHj8nZRnFamkNphL
xFjW0UbVL6zGH6GhMkElpUibK2g/6h9f6snv4je9K9nmLV0cs9FCt+lUwSCfMP9z
6kjpvectg2EzH24DTfCV8PHVQTqNFsVpwhNJzkSX/7AYog2GrS2MLOAltq8NIlxQ
75vUtJSDOzFt5DGTL+04CGRForRnvBVhyjuI+AdHztyf7UvtA0sKXnCGe0O0okRO
bRITm4y9BruASKy9Qh10WMCYOwQ04T4NnFyBP55Wt4h+ST2h9UcZXqnRVwZ3AV2R
DH4frC6oN3IOzFyvlb6TGnaGOlYG+vga3tp3JeYG6hYgUhXdkNDTKERW/TfRf+mj
7beX5e3XhCsKlWTLMBjcalVa/zH5Q3ZPUKTQez83C60eoK4ZSzRplJNUEMM6F/zI
TcGimrb3qPGiY6u0bH7bMgovmkYbuZpMLgb6vKsvnehzGIQAq+phfvhD1h1r9je2
tecRJ89G7C8ooeURK8HV06ppPlLOuogURsaNAPGwPcEidXEIn8+6rjUvwImHhblD
2McKWDEhrtaUHues2NaXJk8ejDlFOaAndXHzTNk4F4spxz7CFe83wKmkV2WXtfXQ
Y9VT3FRUvBcs0yuT52bC1cFcNw1rYC3sjMjPAXpX/Foi6U/L9rgXH7ewakdK2dyS
xYApq/cssiWvTY2BbOW1zMqu1EDQKipYAd9hVCIqCFmXdSo1JJbfGpUUgPjJ4SHa
/Oga8HCV0o/0wug/aYb3JFzqR3y2SfYx9dKgvdf56PEDf1An0F1IIm2sLGSCf5E7
rG3IkTSUev09pYXY3Q4NyhZ7vVki+59hDwOa4sCtjNF38cdrveHIuVeT3oLribWU
oxLPYeZFlIUsQyGbKqhfhFKaojMvzoXIYiEUHjNsIt+BY1EAcma459Aqs9bCkrrX
FBIRX0cqVsf6fYE60RRt5EBBA3qkBPubfYm+psq9AL2Ga5aZKYUSOdyV+gP8/HRs
Hs03edQJpCi4mygSzSpHvXGz+XtQ6Lz+89fMQtsBUNqPekrJIB+f2eRHsrkykXDB
uFL9NUvX/g4cEjKpifazq/FsQPFRdkMJkR8A/HcPwC9UPZpcQwOWAuUmtmj1NsE4
8Qx1MIkA92Gh/RXUIcBlijg80zfIEmiPmzsMmVUbgSLwvrJtwVHH6HddrHx5FO0/
qSE1+Tcpayx44S6J6GXt0R4up61yXhlO6a7BKDu1pe8PaK7wQ1NAo1Qnvabp1YFA
682obinbXJTiuUjWLIE2YjkOoci8/gr7Zt5M6dpyDNh+6qGx4LJjM2L9m90PGIld
aWzROdCsKuRosSZOjINj4ytPII7qJV5xY+daybdAzmIoEuqj+8s29LPwZ9Prhhx/
BuzWf/Et/3s77Ljg47delSeUWC0MVpcc11IQjCLI+eqHB2uUxi2Q58UmfihTQmwi
yOMDAloFlVS1PqADRg7YZoCB0tydUum+Lxt3wxzzBi1hGic5OGx4U4QUHj4Jt2Oz
EL5uX3POdv93rABrwUo5ujw4kUEtfyfBnBeO+nNpidZA3msftfyTaMLqP/ET0B6j
cApDUvmJ0EsYDaZRCdSxt86owfum/5szoAPUqGYkyh5DHZv8bGg6lBwPDcALPMam
E95uDyVF+arrPRG1/q+c7zFWfvokmRNDHdXhbeTws+6gM2udfbzh1jgX4GqpQydd
H/RlKSfG8NBJr0c1X9QJ2E5jDyKtFXSj36wsia9Z1qCKxggCx8Z8Q2PKdbfy/4K3
UIUDm0OJTzc5ee/JZkAJR7vNgP84Uz4k7EI9yKqNBDHlugK/bZZBm0bgLYmhcE1E
GdQasacaYc7GXBtMrPtuY51wRLBvKP529k5WLSDmflyhILSIPpIBBKNXgVwRCbGb
+NAOWIElVaWpeXJnbYWkjEnxIIrPYq50CZkpz6RHkfIqHjhtLmccrckHBbaTea5X
anAgQRo7XNG/DW2nrrHXyrVhDrrqBk/Z6ohYnJe56iaOPaplI1ri8LnjCoQkQls7
QvpeNQgVs1h6DfExt9GfSfXyBErwwWfsAVtm+kEp4PY9HlaXMDpQQUj3SIMOnbtP
jWO/jFtggnjJ7gmlThZNTRPWefD2GaPfV3Xe8KT6rGg4r8c4Ghvf1WyC4CwQ2dXv
lUjKQkXe4800j9Yf5ByRoghzxL6pab+5dAWNRjmqC4bzvq1tgbsn673hq713NhZL
w1EgsPVYB5IibUYv1zruDJtuj+Gw9f+kWsqrbmJUnNBGOZP4KAX6IdvtymyFuKk/
nuXZfx3ViiI4de7iSklVieQm1AXkZmB43BAZO65stxMD+cx/qxcR5uC7towa8A9E
DChaDe/rs9ecKOkG8yJBwyG9K8fib2go8TB62JMqB83+JD1qMUEK4m2A37lVFPl1
vgA9FLJa5rnTn9arNwpcGRcoa9NK63fmAhxAj36+kyc=
`pragma protect end_protected
