// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:36:49 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
TeOhNwNBHsLC96QIqGf/LN7A0vJLqzS6BPuiN7lB99Qz6BJtpbtP/x+ZrzCzgYsQ
FqFOxfs7mqRB0RGGwZtPczpVNgbO4wKXNWZ0sFKXcutqsy6zCmh5DCSOhYB0qgtk
JPWn/h4WY++r6iGWIU/5V7l+GJWGC3BpXU1P+UG8W6w=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3312)
A5aQB3U84zcAyzaWk6JS9d+9a1pbKe5Ps4dK4FBcbRPeaZWkoGD++7/M9ZmVcLt9
3WcUQ5y0nlZt5yLgmmq449XpnmQYldozqJ+aQqB0pi1+lv1UJBa8yitVbW4fiaAk
BowDGsVIJDn3jBjgV5IuuBKaSpoQ8XS1dJYldi+sATPt2jb03aX/KXu6K6Xn6BYt
FsLYAohwOLUx7wry2q2Dbx8+4WL7OhgHGwXEZCW1PTp0kvfKwBKt2m933pagYnI/
gxKO1fKXngtr59nxGBNLppc3sVaIJb0ttnB+CBqultNALhkWfdoLv6A0ZoTBj4M8
JUSA4VC6mjxpnqz3PVF3Q7ehStX/TkCf2mWFoHJjQ0ZVSkS78WSQ4ockD0e53+0i
0Z+SSH9r37SIrot3Ghf56st4q9allBTxjYdkOmyNWqqQHupSPHvjsU7ctaQnF3EE
jxXHdjMTFfdhht3kAw1Bb3r4NxxQ9K2wkBCBvAXukgA8zn6POpOeqRH2O+7uN1Y6
cYPNY/f7u5UQzuFKrI9tQqxmeVfEWK5kZLcgm/rws1bzGosEpRi5XVAYuTRCTOaU
E8gknM0lWVU/tZ2GuQZrj1823oireePI+dN6PYPuUZgm6Mp+rpPrww0+HhHNXfwC
SfWZkei9yXaKnhYMI8M6n/EZw9xr+qahLlYXsr06I1MUj55djI4uVa6xzfRV5MhK
QAPwd1Y76E7elZvoQy8Qq0iNOwsZCXoDoBmVXKu+tXCaoAZF8UDvXVCa68gIqqyK
MGb+9jLADpohBCul8UytUB9/VIvyz7Ysrcvj/8Q3ZNfn4J+4D58ANhkKxIXRmnlx
Xc1Tvx/oclA9zN9EQOEBvcuE48B7JXMOnfGl1WzYuKRryyms4JE16tC+mx6OikZC
zbpSDiB5rjzjbR9HdAEp0GS2ZDHbzLPWdeNGxksz1jNwGRjoa4z27pCPgsJ52nV2
YTbQ5CBq+5ut/QWbfuMYkNlNsdzFBkD51Kg52BnPS8iD9hGv2NleZa5ApWjZF8f/
wuCgsBPRVOYllX2vkzWlxyAZQ83wG8nvC7cPpz0SW8UPhCy7DIrzSIh8rUgyXaE9
lfplnqxDCmztw68HvlXie0h6HGljEdEBjD+67P9Cpl8OdaV6f5fYksN0yKzoaSWe
Boghnr5pnMif6SdLRqWpIZZE6FmQAlDQ1O4y+sVgNFnEiq9N7D/+TgVfNdiZio8x
3ydjpuBPZnN4a874z8SvUHtY4j68aNl0MlKSl244TTb/DfYemCKdHF6rl67ti5jM
WXcNrG8p5030GMUEcoiK4deaj2gXxekHmhUTzIl/JKxP4r6bsUbtAi8GgT9YPKzu
j7R6GqqKLEfIU0YZookgzqnjCkv5L2uZBTGKUTPZE9DS35MWLAayWbmrsppjj9C7
f1yG0ZZIcwLf8/RMHUNlSS8/33S6gLQ39rbTI6Q8CD2efxngf3/4eZHbS/LxqIAA
NWsS17r4+ATlFYhLui2wqzfP+HLfHgTYYQMVbr0qkeB+AlRphoBcbvblLy72nSgE
YkJRPdUR2A7jcEafu3g87qdt9k6Vw4ivuAbgFAo4g3IaOYwrD9NhsRt5LwrbG5x4
ao/GDQqzNTCqCnCG7IGGVUaG2caJQ2ORXVzMW55n9c+LFaxOWaC89jgDoZ57J4ME
44Gu+Ga1OTidRh8NEjPu+OJrQAE8klhGkJy32+AVuNYKCq4X7ikcVx9J15N/kr/p
g4jfJt3LZbTNE2EClymqx7XHzlyORMNfqo71QSUrwoxEKm2ERO7IKqYkKAR2uCGV
iowhvZK4sVd2i8kyrbFsNNRZFSwN1uII+r785DpbGkyTQX7lgmrPd1FFzKnayIjn
LSIRYDYcGpQn8Pl+Db4Xc0FEOgsv2jbhM+XWu9fNBaHbGnLRdLCEGrvWMnX1yAEm
dFbzD8d802KcUCM6Nns5sI8xWJhvDF338fXX98WhOijvs7+aE08bAZM/FH/keGc+
Z6JI1Ad02Iuv2fQyYuj/3R/CTR025Rnn+IOxuUJ3MQmmYy2EW+dVy7XoGSiW97Pv
0WEn8pLhRNqkAIOPdXLSjH6chqpWur+EZROqsUBLmfhgUgCUtYkBKp7x35YZodKM
RK+oZye4XID7++LwRwYtN3LdIEnFN5pYFmWw6MPnXexM5NJK8yv5xsMmRB3DgF17
eTZCloBJXzRWWIp3JRKODS/qKph+s2y4/cv/WxIYLVDofmC4dMGLs60wSTbbQ1Ub
74gEl0dFvubA1OGKxuCFt6nmSP1knpStJZT/0rnhACSQ9QdlaoO//AsVI12R17h1
b11rtkxBLBh2psfcfiEFk3cbk9w4itlJu6OLVB++WXUwtWhSduKgtTpMNWCt7e1x
76/F7yttVYLMPTFiHjCfMzmYnNUuSGJExvpvgv2se1TUipCqW+y6hM9WEmtHsMfo
B0/TB5y2Govp9PfX1FaX14hu6LnMc1ipYyMEYMTXrdNyP2tvw1t7CgJia8nALFh0
KbylYR1pQVaustsZjq05RAs2MVvWfn99sfVl3ZYhE2sQJPyaK+2n9qUVFrCKPDjP
TEZYnrUOir9JhbF5oRZfGDhvempnAvNhl8Ff/mv9giYRY72ib4AhfHgmi6+Rr3yW
GFPEgPd0sQbAP1sY04DwZF4ujP3hSqow1zYCQUw8ivxMkos7PDMTRNYOUrYzf8dG
nr/AA8rU1PLmA4RXktaQQQboP3jBC/WJrOrOq6BedJXAxO2zKk05CtWMVJSYySV2
VkQZ2FuSz5W62AJG5FTI+TV1Af78RMSEhV9A38++ojz7FMPtCoE4vL0GEbuuoknx
l0YQfIIh186Yp5o7hU2wj/d09+zksih3TOygZsebiOwFLRaYiLzyc2NL6pi1jVfe
TiWHJlO0bd48aqHzOnuybPHVkTOMyI6C2TbDkHA0KGIClEIxBwhjl1W4SrlwRDxj
CJLgmMEmova51miF/XRnaiG/kihupd9gxprLb4+Tf+3osDtvpGtGn1B2q5NeN3bO
3n+NcEuIPOHwuVgfiDMaUfEwvlbZdrLF3SFIpbbi7wesXWv3AFSMaTSC52ZITBx0
TE8VKfB/8y25K+HmnJ4GVccyKZTtHMP396KuiyckkIUZ7cmeLmlIXA7fyhjb43Z8
98JkOydcYKjGVo97XwMM0HXFpPcTHIV5PU8mrOjs7MnYfQQF35j1sG6znjkI8CDE
S0NoskNUOoY3S2a3AFLVv8BE8lbd6Szpl2aeF5BkbNSs2WE4hH16b3xHFLUcT5Lv
n64CRPCHCguEwyZh5m52Q5/ynN/DHOppmYBwGjSSkmKxcx305c6vqhl4rMR4l8fL
yHFC78dNwoT5h0+/rrMu3rikstirgqtaKIkwC3sq812INuAW4yeAxKuOpjKkCcW/
xFiyhSvoY6Gr+CG2lRwck1BH/nauwjkqCTv9sPMpDYR7gcGwq15FloEosCkrj+WW
YhaCX0IscIEst/icDnUtuBZ9g85hWghOXN2mbTphlEFXRpsY8BwkULaBJOXRxHTZ
utqlM3d6nJjSgyAuAPfYftTLDu+M6iv1QfkuilQ5MvoI5yfBqLnxWObopxbekCgK
33UH4yFVl+sjGWdYEu0ov3Hp8O8UOMsQ83pAzj93vGJx73xpiw95jlYv/KcalKxu
TDMl92jN60FgkcldyRigqcLkCelGexZ0ye6N1dGqn+6wM2FYiUA7DNCCmNkDt/75
Z1jDH1tcON3jIBD+YgVkeJwCuBRPbvXOfeeIW3LiCWH77Toxj3vXh34vExxYxmhe
dU63NqnmQfxolRL5hPxMKgfIufNNpgoe/w2HBjhznP2UhQMehbwijkr879L3Pnx1
NSqQe4ueElmxyAYKVlKbuEWbgOIzjhFoZbdVsHSpymi7IB7UQVSWL3eqc++ZjBYg
YEGxcldj1EpuWuHu0BWmjFon1ZApXH1RpphRfOrfWDbdjGf+/ENGw9OauL6X+Syu
lQyVjoQnsODQt/8NlS5n97H3ZwhPjsNJnS0Gl0Q36nnSMdbwOdThmCHCfA4EhczG
BlO61+j1ZYu02pOqMjqwaZmQxV65G2LZI/p4BeF6sOvIl9/JnoWL+sJVSfCIEpf9
zc/8vldS2FFv9J6UnWAeVObTmB+Zi4E/GYIY1WeBW/mKTnHCqq+QiqkjvtCkOGJu
E9HsUImJXwUTmboMeibnkrS2pYT1JIe/RRQI1JImkPxJxG/iW0itjy03gosDw6Ki
vdR6no/dIvgpS/eX+XV6CibE53TmrkQJDKP8zDyxFzAHvVx3xsAVehvuxoIb2e3f
4oOfBSJtAfvFyQfyNJerVysJln3+Vao+ISLDPXFvvjFXTqvTpuM1mAUuRjh9bzM/
QD/lmVU510L+P330tvFbtA22q9MP0KuX0QeqDNjjPpXSVhGFBjKqNwA13dnKk6hy
`pragma protect end_protected
