// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:32:38 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
pWbxQIGLhbcjXYbahiKBtEmmsI8UZn+At9L7Hmstt3CUgraBASuYyZ8QcZ/Whi2M
M3RRdFB1phBu2XEi0Lnt26JopcRgHC2F41SLyQm7VGUkSxWKHhhitz0WUzsvPbed
nKmN+Ei7y+ITF5GCZUckpUS60p+0Rkle8bAKLI7WS6g=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 12336)
RZO47fp6Fl1nnHks5UW6gdxiDyNQFU0dwly1npjYrd08vFUr7WivDPo07DVImQT+
kC0SkBj3zfv3zXyxkObFDS5Zz9ZBxNiXrsCCm5wWUvN38EUxYQUxkB/zlyQC0Ry5
XlwNNYMuddt0D16hjbElwNOiEGPOdLu7Hqy277x1owSJk51G/euhyAzRJWEXjNj5
fswhDZRDdmVgCvV+9xJpErrE/XjfP5T9EUz2b4r64u5yqAIZ4b/mz/9NO3wVtbEE
gO9ZzNvoaAeMPLDnbXaKDU/bd+3PHK646MH8mY9NB+i3csA30FCoNMJEwtML7K3P
57vnWuoq51lghPIhn16Wmq60qFuiMEyFwfwSpxErLHrQRRgjWuSMHnSvUgzFyWJM
4wwnGi6cT9sSMMgkS009GP6356/rXaA2JqdkLcvJT+Cr+9A3PUb2zawDpC7KWTq+
kgFXvC5aht037k1YSvfPrl8ZLsRqSZojHnlysQsM112Kp7K39qt0d1/a2MegJVKN
7pe6MYc8KUp2eQEHe+FMCTKdJk0AAc6NqiCNcYsdyd8Gu2gW2cqKqNlP3NHJzRIn
xYCOqvF0QKRQb9h9J0uaLX2RX1PTvMZbWLvySiwiJukqA4Lh9TaDf4KyiUUfw8Fj
yJj/6gLxw99IazFswlwP8kDdlmTBCMKnO05C5tcYLxQ2FdcVmIvhg0B05kIiS1w4
k2T6DhKpW2pBdgECPY2vdh4mtQqAlcPesRBu5ZHPDN6J+LdiUk8598PNZbWwxjj0
5ntGXVLmmvji4z/QyIks/rmPSllvNIGIHost/3EdotGG/fwZgrY//8RtADcHcBjK
VeVfOFnsvmi9Y6G3ZC03oKC2rT0yp0jRnelhq27TuIq0iz4bdVzPlpZe4H3vVPHr
Z4jWhn9MXeXZA5357RmwJPapT+HRh1usGXRqCMLFexZ4GgN0Dkxu0HGfcFgC0mBU
fwFCQkU4deHreW+PppdiFkPpBxRWM4+WgAOJQzXCfS7P4MFV3FuiWxycvaPjWyEP
zh1zPPVvornZtKIjbE8POG7Y9hSof2fy7yE2dE4mWDf9eDv89noyBTvvaIXwEjoH
S7MuzHjpWhPM/8mLltAuvA7LOTCyyKwMUJ3xH7A0JtkJdLC32C54w4QS9Og103o1
foVqAZfEtUKFaOPbC1uy5tUIOTB8iTCpnIB8CpDAuEyqtJFRzofQgJuwVAXTkdtg
eDfr4L+YoaY6mV3pvrjDjYg8gTJvBEKfKUj7t8xAcMQG9riweu3twRPNN2jf5DiW
aeRcNgz5XuzICYxLqAhtxsmXKPpmvN0pDGKAmb96mTkjiqCbrsqVE3k8/+qgi/VC
DQB9POqEJBdMjP8PR5CV/OaeW7iLwa1XTCfmSAiiQmMut9suv1BaM3Jvh0+XpeCX
d4Fir5fPsIb5X0BtBXVnREl6EhYAYbAxDrWSGADSB6yhBudx1u0eZZ5UdUO+C5rt
uG5qeabCpr3Zx02YviM9pkZwHjI5SOiyc1Bm9NlYKLv13u5pccf2tZa08kk7he2O
S8by+MMyyw3afVIfaKVoQL/AMYrTDKFUEkt84KDFBQJNSim2LRvBpc0sw7bBpyi/
22gpiQ8Ebctwn4VM/T/1edIRT5i5+O/RafGhT4NcBOBjN2rAF8jZ9zRh8i5199WW
IwCO/T96WVCrO2nWLgpvWr46xgOj1dLJJ7zF79mupkjpt7YM56LxExV+3GVT6sax
4qIIfHp9WyhC0tWA8vKlyVN8HazbFnYcIguzpuoBbXVuE+eqv/m+hFRxqDzgs2hM
mNUs4daie9DfrajAZVHC9K8yC4tkpNbGHKwx7P4eM6LTrH3nHawZ7v62HYCObf8E
X/2GAmhzrCNLwRFxf3C9hGskOGnsHkKbBLzxeKKe/lpcUkGS04qafzQWXwlXff7L
3C543ztWbfnelXOFJ+IilsIv0QKxWPLEclB/bp/5u/vd5rJIwnmB01sOdtYxiy0O
Iv759mAGvCJPfcnQlb4Pq/cMjl88mQJ1/QHrE8XLw/i4lY9YEbH/j5WtIFzuFqFd
Nsh6TF2zqJ1LS7eM9ZV40ScPeyOaqNLTtufYTiBeXXybyfeLJBKbu+j8xVzo23yI
RpBOrRxeKWmHtlSGAqRgNoNtanu+24XSN3SLbrcJG3MCRmZR640nFL603Xc3q1is
rG+y1sRMAJ3oNkpNiHVn38Jr1Rey/R3jqait/cmonRUtgwPXliDOWjmzzuDZayoH
pJoyzKOLpe4fXl7nZ5Mjg/xmizeSTrJSE9/sKM7lK+TXEKVnO3cD8MNNHOu6tspp
oYz0DbjMXtlzCqrIMIyntCOQzfGevCwH86EDfO5/yCTPU8IH8+CY5p2wFAVofrfd
kSmxrnhupqOuYwoGqlep95dbno4qK2dzAUiut12gNPaDrcbbrMyuDKdZafBMAkc0
u0aDEU664VR1m6Y1onuz55n5f0zAL7cn5mazS6hTJu/wuogeCiMkZZpEGTlg2ukP
slNDeoY6IC5BWhPOU9X0qhx5PjgdjHs5/Wv5BmcByWZzQ8k8TVOvyoODP7sDJSWw
ncTUjgy1K5Z39Aipay9V+DpB9V00AqZIVhrn8YnX3/451aOBft6tdgG7XPIElVbK
f2K98MXc+KF9dppDOIVxqsIyR7urrQshbL4IQrpbL34gxIaCXER4N7oEEJ7yQ87c
mpnelLYurAxExnBSUB4+QwhXsYccLVsMXuxbSEm/iQGTegMAGLekPX+ie+xGLmxX
X1hOc/tOucHibc9QIqyAhbgDzNG5jkEABkNUO+Y7TeCKGBtvMVmI41lDGqVSI5jF
2QJ5vW2X8gEatuu7OzSEvhuf3yaZou8V1pkiJcHJr2wC8rU47apMlOSdqZkRF7nH
9HYqhqZrnH60jQ1f+3/Ug9B6oWxw2E9hP9JVWkYaKs4HRlxpWHasSLlKWtUdScp6
fl4dbr3iiaV6qPZRz7OU8JDjPseeev99RakBGm8XsriCbEiqq/ivwWHOjSHgOZov
fJjaTNxwsUVfpJbYQyd6HS42hLg05yQMhnoICO6RdeGyL2hSQHYgeul+zGe6tVXp
DVQOKLeEMGeBV22gbzzDt+q3OlijnarwD64/ZLPU+TK+JfSBo8/lTwirWUXbbv+c
xEWKdOQp2BX1Dne5ru726pyLVRKWmUYWxTAFJnX2TcYxBHXIo1jAM3LqtioqPXtM
Ka3HUTaLEEyCDXkR9q4hJi1QsFEZFOScUEp6ceG2z3JiAXXmxqdz9EJr2TcRubEU
O4ILg8S/3kaXF/Kos4e3lagRYJUxqJ4MAmcjLIno73oMccKaxbmY4UaR0X66qBtp
NDkKJCAbbU02cwusEo/7f1y6sjuUBmYn12cnNBq2odRktPnPUsI8TzOA9kR/zCfM
Ru44fEVJyaOwAzEZGnrtlKPUZPLVYPYfOTyUT5DNlWez4c3ih0Mqnngxh00PQ154
8LaYxqwza1mBz9fosQd1aDzY7zCSSdYIOrf65KgHJg6Q0qW4ifvrrS+VIrWl+NiL
RlRyNGQqseaJSN0g03fDq2vhQv0Z0JNFjENSeBeNnIbckM9BCW9S2OQtEVLLnC+h
qdB10O3nEGZl7U+IEQIlQ0HcO/bXC+zZw/5ePN8iypYrSegcOTS0ei5QwZOlDLXg
8KGN+QoFVnUTJWNBAf4Q1S7wm1GOAclMr67cMtHXdR2auEwubWqHOY702nMnQ11u
p+FSPpTiwxdGfXOb9wO+QNiZRWXDRFpumR/rIuYWY8J7qjuiE3NdbvuZqPh/qBNM
yJXc18sbhd7wTT/nWj3iEMCPO+i4DsIBuPdOWi5RuHLECSGhzpK3cVFqw2Bcebh2
+PjcHw7Vcr9lUkCvnj+OPa9fqySrHph9OYWv5QW+pYWZcY6HY9zsuY4XUjGoiBz8
2WuvO45W8gEeJ0GpvkS4Iy+QRvI8S5T2oQtrOmurDni9IlQ6wGK6fDaVLRjtQIYx
6FDq2GAAWAxWJbCUIT0qYeoq5OYxVHoIU5z2p7du2p0AmefXOMoj48KJLN2+e9Lm
ZTutyKMFV3lB4R3hq8TRxXVi6cgHW/SHtVyKEoLUzXuwwseXhvlLwYrszk5l92c3
L18F/EUdlZelUThIa7DQ94b47v+tsMshwMzT3eUTD5yx5wtZXg8/kQBKJ41z2DCr
MWuC3p0ZTYkMM+PDJ1B1hImL5f/vKkJyjovzcSmfEuMcvugq6qf7caQISkUMJhWF
A7lcOvkmR7Yi6wWyTunPMIb/XkuSnrNeUAd8QXZktKEGNNtyEk6r3yRBh8cSNLAQ
FhTpP2sEsGSqrViVns0fvzegX07x/9B5G6s+UJl2QeHiw1043okWqiebixJt1Ebz
Px2tYGUcgosqJ1/+8mHSC8GFbg1toQU67FEVAq6cpyq/LkALYGMPXOeZlvChRTq+
C8s5E6lv2t+ADsgUN1y5kDEjw2uS2nyxQIeqQOQaCSNz9lKbUPv9HN9iVE/JGmsi
qYi6cPrSnEyoLgtYw40Ou/pqftkaGeMNReW2yVfaktg3d5+zDBNhLa1y45I/0RDC
8QEWdyVcHxbdjoNQuRAo7OUdj335gogM9429+A7PS8v+bsIxW7NgKsGbk8XbPeuT
pzzUT4lOMBW0J1JW2wvG8IxVvNMJcqi8bolLBeLBn0RWOXlvYl0m1LRbaWPD9xiw
csyyrk4YqgxkioFfWJE6SoBMFXxIQPhMWA4q6rjLLTyWVpgrTcSklon3rkqZirm/
+G+hnp6FkHpyYGWeVYI2HzhIwCWEVHOIxMo8hJMU8NdAev8EGMo0UafitMmWnCAq
gXCBLlLwhbIY0f/jJUJdBCtb3xi655NVRP+aE/ir5sJ6mqZxZPtI0scttfdFvPLo
UQlx4jJQDi3PmaU5kBcsidKZoAbfRw4Zg9dD+0sfq0iZv57lv8GtEqiC+M5v4igi
ndaaVqgtALpefMCI6cNcujjaRRj6mFHz2pMnuLGXP9hqD6fDkn8IG+R+aN2oY4/I
akxaxWAuWXkqMrCD8JjENAl8WBo9Z+qZ1HgWvXCmk5vEhmct4D9utckx/O6SvvEg
xpckgfvPlLvaRHtEODmuwc4Eccd+lcF26WvA5MBu7DIk+cMNpe9wW7rNDxZLQ0lx
jxwB52uMAX1g73+bbsAhhQScmGQWZ3D0fAo58zbSN8f/t+cfSKRri9Hs4YIPw/0l
fgk1f/Ml8U4CcdOvZLcwTf1FtgJACvxYptlxW37nlVhY/RwhQ3LVtIqtQQ0pFD4g
ehqyLC9CTf+Y3f8zVMM75aOP3LxV/BCLAnlEwJ284hB9pbtx6feuGnz0JdPy0ZRl
Jpsew14qLq79AwtEJCMM3U2t4r4lRbE+1Vcgg0vKltoMdT2591Wc0LXFgXUZQ5AZ
CkQGKIgduPf8trhcuweiAYkPnJgAKFHNdsZi+V9PAKwKBgJVH2z/KuB5F4hK3iMF
gk4UNt30u1iJ075VJIaEZjiUKYAA7pyuX84tCGSqbIUtenX42ara8s9IjyBk+y8c
W6G2U4qQ7wQIvm0R46VKmwU4ZWfyl3wWq+YLf5MVSsqh4E5YtXde7P2mWijCRGn0
Y+bLLFTY+jpLuDN/MVlvtMud+tu9ls7RsG92Eged0PrLMylThcY5aaMbUeX384kB
c0qv2V3TxzF42Z/VSF3OTmOnFZmdMfKFlzU2dcyfzEYzkLhG2KOahc3RqMd8VD27
KPkJlcd3UZAw6TYRuoQVM3LwAY8VHVTY95cHjKdaV5Dt5xtah0oGyJR0D1ffdPZ6
SScxfKmkNqUQjXNmzg2Bi1ZWrPq0OKzn0n0FFFT6hI7ZDCfUvjr5mLi48BaqCH28
VV0htkLFBRpiMbtD7Ot48yORPumZtbtcefX1A4kC1d9+WPFZxZWyheoqDLaAbWkq
HlGtEGLyc5pFQ7M5TVkqHjlXXNUKesVf7+9USQjRMs/cl5gsY8iLDa38XVBi5GjJ
k4576YrnpuqBF2oXI1NWpxOJcn2oGaPikOOkMwFQiaLAoWR4R7dnHmqR/wk9BS++
F52gHHzu8uQnVNMGXuLHe4RNmVwJNf2qFEoE38ijXyTn2A+GKTirochYB+jAqSNs
6QwTHS4S1YgGZqLQHK9zu2gcqYmPidkC8nfDinf4nXgTdut2PvMLZCzK+dLLWjev
8CiQRA0KFBjyUhHJu8IVtP/9yLFHwJaQoPAHdO24hG0T2CuVtXqMril4bMM+MsNc
F9/Ni4tuGtr6JS8c2vrBUkHzo6qy9dPieIBrBqG9J1fLDuBBFMIwRe1PGz9/Ve3h
0vIIOk46ExVUZ2hrzlAbV0GYIGpppCJ22XMfAQsgGN1cXk6OGbwf3NOyqVKik7K4
JEMJ0yuNjhsYKHc5QJyyhoxDU6vVlog7A+LJ7O5dvxYHEro9W7p3Hz2waNVtkjfT
rdcR3PXpL8FqS1NQUhSUpjsfxF16GRTsV6yt9JQP+sDu+fIIkhDCBl0EQEr7+t3X
sU9shqe6pSV0YcERqja8AQ3uFm6o5FqDBVxBaxHIcNYA2IaTbEj8YOhNg4smJAF4
tpF9wu0DdJLl7padB2dAScYLO3CUzoQUZfcTHtPzOv33fN9F0EaoabdhmYmOrRNC
QDD9ikmBkPHGAOiA87BU5BP7tqjqTCuWFZ7x7LkbBH/MaQnx/KB4+zxkDVr6xntV
XLcE13wrkQ7//oVyoCJHgLQE7L/aQOgy3MYcSKPtaTUIww3Ith6kR3ZmMsuoYpsK
ZbUb5ghR2/vdbcnC/38BOM05aSu60lVMqHpnlX4bRocSecUzd/oMl1TgjqIbhz2g
vz9/OYyagz35YhrzbO1ZNd9WhhB1ZqcEqnz4jg8yWw2bk4M7GIaWoprdghJH8j/j
cQZv+EVlfx1TUheqEiv2ChDWulfETMJMtlJm3l8bw2USMknpBElOD24S6fKcNa62
xFgJU3vVJStdnIlaWwUr/fHPgbEFaJR4/Tj/l37NylT0KKulB6N4cHRu3F2e38pD
NKvx6sEBaaXaVIgUDMJIlMi+vJIce4scllAOkLteUlD2NGgch0LLYUjdbWSPgAAr
Tc8rzyjFCl+gkSWXbGq/ETjyiuCvyfpgmoWHWPmnrzH1nAuKCLl6Z0QOCPVy4qLy
U5HtarnilOD04oMO0iL/j4NxeSV8GAmkas8TqO9fftlaEZtSEVsQKWoOfkwR7kZA
uAB12CWF9BY9P+dNNLDNQ3OGIB2KYOtvnwT8DMz0EB/DBo1oYLXMMBz0k+S//qy4
ZepNvBM63zqhQxgEmsMaO+uGCYb8Q3FjU2Lb9wtiMp0o8iGzO/2gkMNsdg3/aCOp
3IFEzf9Sl/VcXYTAaAq09Im/mg/Kx+q89bdQhTLmbddCz6SwDPv6rbTx8D4ypNVE
LbTCih0L7bgK1iXugBTXhVX7+2mNqTSjGE7T6dSxK0Iinb5chfc6NcdGRmjB2r9n
S8rch/gwQTX2BCIXbRQoekbKETzEZ3ytaWMLgYtn2HzCT64RcR3hD2hly216rw16
bFHbw6KFaAjLhycIr8HHhA52N3+pMBVDPGuW4nOyIZs1M4hxDFpz7OyXRkyOtloR
3KL+PI9v0ifDlB4YDiwfCrVfTarJAH6le+Ba/wUFBZJhCiHgyaOQ/HllBsyhadsQ
1HK+hy0pLzcUpsezAm9gdioVnouRVSp1rF/NGMXsMbMbYxHkRCQ7Ll9nyMKL14HK
Rkm1X/OS+xFq6lglOQIIkilxwt7mDJuoLtz04DmmVnMlqQM26VgNaDy1fMG/7lBT
nepQrsKlH3VXdHXDAbrX88to7zeF47pVMWBFuuwdhbGDF9SnvhWk/2oBeS2sOWiH
cdbbJcX/CYRMCfXu1/62+DvHoDOS560pHkqhYbyq32gEDiaUYtSY29v26LhuFv9F
O4ov32TyFqsfcKdbokjegl0gx5DuWQbLRJMrem3UfWifaQNUZFz8X534uaTjza7A
W96YTuz/XBDvZscrxtupywUG1Yg7hx0SQVYqsae6EwTeGuOXoggHA7MihXzjMmJs
/2mLp3PvO+FHJ9Fu4IAaCfqaua4PhtP7+G1kIHMcoLIjBc2KqL+MkBIxW6giiuiv
J20SNpPlJW4LifQFHWsnq2FmHT7rT+b3e4w50+6gghVmW28tiPanT/9O8y+QqDhv
H+P4evd0FQIlGZOX37sSgEugTSG/qs6ahhhTqXc0R/VA7cIZ161IwA7ovhhbGBlq
d3ogvMJC5uFVWDK7EKpcH9PC7NSawzXLvA8z8OesecxsyuiEasHzFPqv2P5r42bD
EBmfz8DPVMfV263xEaXV0Xq/rNSjJWfHzjRSJbR4krZSQ0f5/tNi3i+EAoTNY1ql
1KQ9ENK6LoET4A4pxC/JqCeIHnlIKsHqvgOn976zcMxiaWLzaPNUqzkgSLGUY3uI
CZ7mQioIjkbt48rTZWR3DsCDoHlPU7o2oeer3gOWrvwbO85XxiKht3OhdqUsAohe
Z8QInMv5XHAwBgca27AMJs2FkXRSu7wCDd8su9VsfYBD6cEix6jhSBuKF8v9RQ63
t8vfe8j7xDOQ1ip5/z4wWns2NNEcMd4dCwSXTzQ1fW2s3z2obdG/Nu72QaT+D93K
NyE7h42AjkSHyjc71MnDomdfhqiDP77yhohVwYDdLTyVa5eBBGSFNVIl8Zndxft9
ojyaLzi94qoUv1GzuIdYAI9MxhfoxeNGB4P0QSl7Nb5+jgLhTvj5RLyoUuCgzMXm
aFY02rJ6mUjUW62LJn5px1BEnd1m3ubADXUKtx0/oSCsOq5PSZAgbO1MU57zX1Uc
4eljN1P+YazFWV2E6srprK8mJsvf3xUM7EgtJW9dyF1GQ0EJcLtGQ0bSxk4uTZd8
kCZHlRnsi8ZRT96vaDDtep4BR5qNFZMjWWi/cFU0e7ZghNST4AwNP1TdD5HrppSx
bwFswa1GnU5OVbmLPssdDaiqH5Ramcx3OqUVAxhiwGVx3ai7wZsFdfvpTiRWai6r
DhRRhnIW9oL6VYCkPrWXBct3H4AN/BvZAhIbYCZtuFai+Tq1EjfR2ExUa47QoM3e
ATlZRxQU4TaylWR++mlDgb5Tf/CCRmgBUAY6YatPorilTxKzWFsQZbYC4h+GM9vb
Q1igfEQUMHoq7QtPBMwNY2h5oIO9E6YMGoMpATSnKrJcvjpASNHV6ynypGHGIJC1
9tKakjD7wrs6lsu+B22M8x1cgPrE4m2S/pJHA+ZojKSXi8fMQytJpHNQqAlD6XO1
8yNtLKiABNURYDcsyUJiQN9dEJBv6iHuHtm6YQA3aFvygyFzDBDc+wOYm8y7/mp+
0YjvIBef5yJknHitpzS2KZDhA/4FqMIfpqODB6YI6bMrJK+9Lr0ScsiKnLClTDUO
2Fcz8uETAIUCo7DF19Cc/wuSgpZ2zzfHJ4jNUzsOVDwpsLZX2b4p+xVrJvfjD1mF
YDNsl7VNmyEc0drptJEeVJTaB4xs+ehf2Fp2KHQ1WgebgYdbMg27wd6NFDFK5zi1
kiIH4Qi1e9N5F5zy2BFBY6UeYEJbFjIgqMPiK4gfuJO55INuXpLdU9GCPV2H3/1P
sGr2j7fbtEFFtkuDRFFyVGdfRp6LiHfDTTaA7GS3RdKXUNC5CVt1q6zypwdIuEkB
SOSZxRJCNkB5U/OrdZmvqPNMudDBmylpwrZEVg23LfpUaOmXus33xgZcVMll4ku1
tlrFhIWzZiw451kQIrAhb3IUXIm+F4OKSSomTeKcdtxN1Okgjb3pHgutD326x8U4
vDYIbxy06nFA/aAIgNx5Yh+hLW3lTvbSu+i/KEYvfCudWwEJm7o7y/BBRSDY/cbr
owJhEfqmibsEONq23vvK9MJVck52w4ArX/EZ/s29YkTtyfBpDvhP7AyCz/CiVquG
tFBzCuS2SoYEur8HJD/mJ5PPy5IBUn2GVCR6aJrSXPhNWKTissKSIqTBRUPyT0WT
6cqzI67MNaQlOjy9JwEhfSdpxFo1rDlkHKKSsIoBLx2/Pn9pvX3TiJ0yubldqGMx
D2giX4K3HDtU+8tCDnvkv80nE7zUjpUfm9S3DjGJw5sob6648i0F9t5ZAfyJAWy5
Ud+aodAKfXJUOrb8JWYth4wBlkkvXcB5+/brS45ydPRbxCRvlrccFaJliuijr5Qo
59rSq8+oBPqBA7WftNLyJS0f8ulIcIsdSHjxfzhwekPoX+fB1zRXwzo5X3fV8E0P
U4PyTx8IFU4UH8mX8B4Nu4VP6BbC0l+R2sy9uNAdmK7+U/9ryp4ctcQVQxVH57Ko
8JfULcNyleTJX1hQU9nSisteKdvWyvAm7jov7daa8rjixerSX3RMpiP95XTEAxeB
HCj2v/+C1y2daie9bNgxM++CiH9qjUF0w4THDIvvPoDx05J1ejb8YSs6iLEmNN3g
lDZyhsuVl3/DwXapfP2/2sT1rZuUxgaurWVjMAQbP/CFoLZpNFBlTpomYhQnn0N9
iBQum9mvsK6OjXx+aaty7YK7JgTL9Jnpjy5IhovSDJtpUfPyadNdUaDmIDg/D5Eq
XoAyjCVnXnBYu8n3d6xGGol5J8Pc6A4jWEBxgWivwMSZeqn5/TeOFXtso/UbcTD0
KoLGRROKI4LOfwRGZfhW3o/JE5puOsgAFxcXpexlfk8Eo9Q6aCjLT+CPi04xkMMu
1aevz8M4NGukJ/ojwKBTyIUvrKOCvUhw8aCCPqRcTzaeKw1vgWHSaqkG/xFSNyzx
2+Nd6wFBq0y24HbPuJTGquiSV3NTMuUFXvDhEnuiI90SbjK0ba/MMsUiBhMq8Ssj
ZGgKlgAwO5Xzjuoic55Kr2FC699Jnk2reOpF4AhGtacu8poFvP5rLABd8ZBQoUCi
K0h2wj5ypre4HiEUJv2i05cj9YdtrqVbkTNoDiIVYgA2Modh4tHVYhSOViEvrK7b
jP5Cy14tqr8yrcFPDE0QGnbCuz9s0BEypj9jKpMHV06QBscqEM/2Yc1F/d6WCSnQ
Hh/FIvqfGeB9SyhYRZ0Q0qWYg3Xoeq/HN2gXxbBTbwsSbjXIM7HkEjyYykt5b9Mk
PL354ppygDcZrxw3BursWLE4U3iJlH7xI5nvzOT1WC94GnxuW0tIZ+yB3cauoe7A
XOqz40DCZvjQS/muFhJMUL2cdqNU+e+IUYh+3hH2BBXnJ5p69yykju+qhnZSxntY
yfuXGMuV17T9EdTzPLG0ys+GdURlxeMVFFrfW7GI+ZtONtJUjf3MCGsyAtKVloyN
pxYQj9boELDkVte1Cr9Hhwo9Wc0wuGqD9WA7FYmf5DD2v3DTDF8eTk41WPCyK+RF
C9uep2LytnQzPwJrj+/gR/k4UZb5uoHOu34zQ64xy4DGjJW9g4cRB8GfFum++GR/
USNIcbtZSGG0UZn8JDKkEEZcKzVK/gMYkXIHLS/+qVyAAhV7UPs/sec/kMxBv7j4
wYjsrpUWVK832/m8WVGcT/Rhrg+9Yv+9rbFDWiM1NzDqgztG3ulDd364qv+qSeAG
tBP2o9RfPMZWPf9eKBZRSDa4/wRxIO5okUxniNoCSaiOwxiZoVLbJTlvix5I2cub
ZxxFaTB7DZ2qWhkAO4IndYpA2wQykV6XzL0v5ow8KlTQ3YwY5khku9/+LM0umNNt
vFv51Ad9lpUxgRMuGjuuZ4OqSDEqHJFJh2MTGNEIctQltHf3YzQssFs5jcJa3TVl
si325GIKwrYQOXbthhp3BBpmDeUlHE0PjMtM6BTmSrrIASFyDOsQXPGEFhVg12JJ
WTt++AlS+ItKEeLESyyl1mlgo7pKH/2XeFX7aT4TnbcxqUImwwsBIKjMp2jLi80L
UvaX9346PyGx2DkYsCELvpIVvIKnIPK39OYrdaCAjrtaz1LRd2PK1iUend0k4hO0
PLRR4tgzznHbdSmwO2r0rxQNLVQgB+xj/Ov+1WaovYNg+2DwyBn2bOafC3ZkwfJF
udas6FkkrKC+q6xW0t5rkjO1HgDwKL6XfNamU7ED1BWshoXEQnrw2E3FRtFSLrI2
CVPbzspXCarvxQ8DDKphdG6+O6JoGCA364su4KImabJEU57p5lsPr/i5QRK0mEKU
80sKv1MLeedPceBNyLNPebCrt2v0wh3S0gy3tW1PFFBhVt2jMzG9rxbx9rmGkUqk
KfyA//1Q0AISEx1m81wNNTZ6ingEfp+oSkUyBhCv5hw85rD33pm7+qdNlp3iGZrY
x3sLI0ggS0MKo34xIV6/LTIzg6/IRwjAdZmetEVomZkbqqaU0c3bjDEHPqErZksj
5oKMmVK6go7EXjRXHTg66EFxxqxQXWHPLFQxxLhnDqwu4LMs2vGdkcLigW7QDuvt
pnMkIpHLZheUYb5sVW0z6SEdObEggMHN7KwCaLE5iOF7xJQH3kOyo2yc0FpI10eq
G0axoORfCKp5nEyWObcDeXnpgMKUZhlPCwYp2Nt5lHy/L0PUGWC09j+lJ/Wn0qxz
6oxVcKIxc4DXb6OQNZ2igv2qRy2wKSQOxzj1IcU7RPOzGGKCp4B5lmiucbSNyHPY
xhBSl2BEgixm6E3yH03xWKCI5BgVZkJ8K3tTBan49Qdc9l6+8HxkclvhGherzb2x
uoIY50Yg3RY7kApjxmJdrmHnpF5kJk2PGVB8MBEGGQwO4D5WgS2Rrrw55QqhNC36
E771l8Q+Aeg1zlpY/rDMwefY16JRSr3+oo1QtG0A9FWfTFG79PRlIA7UUrA/PF8i
MGetILwUep3GJFdKd1odxNt3HlI09W6kAs+eWM6eRHDp/UOPc3sSQ0xa0A/Qu/wD
d2lp4Zqg2TdOk+oWr2YnAxtJtHkHwVSL7Ii3R/6xg9ouzNDHyBlp5j/PaeV8zdKv
+eISaPWhreK4iq3frdaqthJrO7MffMB/sjfhdXHoUP+ZhdAocAtO+V2GPOvImVKN
ebRqFgYLmAaGHJ0W1eOBRqY8vVvcDIM9RBXRpTjLlUYTnMBXZNioRcaQV/cAVHb+
yY215rEBdIpcLZHV+KLzFDtSXY715XOWm4borMYv8Tsb0sc/h33Q5MIqRtoqzQiL
09X5JV0nAeqG79IFlmdv8+mBC0C4yru92++LhpUn+vXKoOydtoqNXV3tITDKc7dy
K5zfdIMokh+GrRJpKQejXYVSkRdGvbs0GWhnzXBqVrZH/B3zexIZa3hNy0CrTKKF
QkIHov9Ik1a/AeeCl/qoJedCcMUoAnMJ6RCoBWxPDEUiM8oCBjcnXED2mdoO4i6S
lGXwUMgxW1HeejNUtKl04ZAmvfaG7UbiX6ApzGckr6qmmvF9YeMmz1Oup67ybIn2
iDETvrdehIIEswo5SYHW51zTeU0A39Cfi/LnWvbl/HCul1hPKx0xxrg4g0BYDlMp
UP4/chqc4cg5Jh+6p9AVEdaEUGYw2QGX3HCUtBmrnOVK+s2pL3qu7tlg7dTDkEn/
pmqy+krdwhaLUiDIpM2ZNcbfE8P35sCc6k/SEk3bzfkdftWAZYvdKu4hAq9f/A2e
YkEnXtwkBCnSEE/ZRA4qG36qGW8tj7MH5vKi5dfAhmxOeBtLZciSYTVJ56ZkQRzY
WLeuNVgSnYb13l/NJ9Qt6JClQiF/Dk0wfyM2Lsi8keeL4n0MCSBlJ8Vfad8GhDkV
8qsPFENxF8QHKMBtFU4PBF+bCMdU6m8s6YqGwkDxK2vivK6MKctmwi7INk6vIW02
5i/lrFzoZA46r/ZiIISCZqDdSnw6XAlTu2eks1toWnx6CFClN7DBiR+GqbguQKzF
wuBFwST+KPCrOVnuNd0lP2C5m9IbjsTv9ZXe1mZnDBd4LsigqibEpWYi06N8hIUr
JE4jvvsOEt4U6sMuNRn4Qmi4EVpMxlmHNrngRwHnOAdBrWVHvxs2Kzll8Urr722o
eId/O+ZBJlc1tVeziB+U2/5FzK8+Z4Ko3HM+/FkKDfCN4vhxZu+E1TDpl6i/dr79
4oQUGxvn7duo3Ati9lvsF0heFI04CMc5KcDNSWqCLDbL7R1Yue2+U3irbMfHDZH+
8YsLxnNrzcfHaOOFmN8Nx5YcmHVRVi+maS+QJmK1/2eOggBXviDcaLqpSlZgDcpK
qVacO1/J+E5E6rdJeJ8b2tOf8+MBCfUomEIMpHVUAUQ9SGgR42MGZ+EASNZkjulm
oc2QlEzTU63h0c8Vn1Hj3KKUYKmNNNnVwgJ71cGZokNgqzv5BnOb4mcIQ+EXSSb8
aMu0jNmREKLbtDjbEEe8NvDj2jHDLucNSDy6VtLmE87QQ/WR7oPbBzVCLrKnY7X2
ZfkF3exxYKou7wPLABvU6GgaYtSfLcLFPDrwxmNH26vm8IAKF/m9b4eDdAK94RmV
0gscHeGf9ZIsnAZt1DQXgIcCHcwL7uWZGAwmdnDRfk74pNcPVBqX4EEZvtk/5SXY
mQuVcM4885ECEwokTWhwXw3DArFSoxfLkfyVdD52dyqn+sGR59bC+v4NuWSrUwr7
BPNFhNzPUAMj66gp9Ss4Aaq8cTFHwwkvm1LmaZLK5dsuW2Dc+Ix6KRut+4MEuNa2
DJHnV2xwpfMnMLDtNDwMmthqF/QvSJqJJPnGhK1qbSkZ+mPc8DauI0Gmffen8qFY
mN8yhv+ukDYIUkRJnyMY/kwjix6+PW3v0/jl2utUTyfe4TdNAzCmVG9Edr6SxA1A
WOUifzOnW4Vb3/dEb7LqB5Po/y2o5I5+X5h3uAwLYjAuldy3OFwAD9TdWGX4rtdn
/zFLL5xW9/FG31mraQweyByWvOY/14HNFOs3kxlb7K87k0iuves5yIGq9uA+43zz
9tDLSnTdKB4fyNR4APnXR+vWsg8l9geRht+xawLUWj/g76XlivlD2Un+kJHAOg+N
8FzKOP7xfdI5ZlPs1jbGO2rAU41HQpC6lFpvwstr+tVPEUXFXduvOorfjuFCui38
pTTxkBgkunlltGrf48KTg4xo+RLWrg92QNWtg9AoKl/JYLtDowrWjjZZopm1mWfC
VA/7lvPCUN/lvq4tIsojbYlx1/U4c2LPVFoEOe4tkRnF0Qys/biMeftU2w9LB1ps
j8CYT9bwOkVztB9wRMtyRAOQMDAf188Am/s3GKx9YN49CLVfhcTiLPgwrmzaIicu
mvPlooHx7QKeEkUQ2aSAHO/BQtrqvaKwhbRjbg+4aWMCUSSIjvlNFzCwPuvUQeLm
oHy8dczuFyCToEoPMcVuOrLhr75669cIHfG9u6XHRgnzRy6M5aLiIOKKKHg3OaGx
lusqrOxpmGzJC1OXNRCivHiThjbgxibzEhTZzGV4oLFXJmEixFkPlwqTxEii7NM7
8leKjyW1BUXGRs1AJTEVvTfKmu6yGD+/IxcU9q1d3Nw2aNjxxWA+PEZuvlVD7Uuw
QQLsevVQNX+7UzXu9KSY60O1wKGPKQtK+DVvfXqN3hhGCvaDhFNqo1eIxuTU7N/H
LHBbJZQonkaQnaqfpbg7vnRv1456BFMf0YvcZDlEr3zIPxn92k4w6newliO+K3CP
6GL1ZvoKF8Dhbxt6m1ZU2kZTAKgN/6H0Ge7I7Hc+gYikHMo9QrUAm/qfu4/QLf0h
j+fApfU/HFJ2y56DXiD5Bvro7MSr7Fm1pxqrtcKWfGYQQUv3pnojL7M4RoWy+V1p
V40v1e0MODsiyGQ8dXQ3kuixTa8jrzphmRV/l3UPBnaDMOnfLPJ4uKnZ4NnsgnX1
4o692Ym/TbkR42zLlLWBPBSO4lB160+G8xZL1YZM0Wk7nNgwfEZyMRf+Ez9fGocj
d7IGzHGH006gVznT8D4jE6LKcCxgpUskPvFxycbvDBrQ/Nh4svhFTOQWLaq3t6Tf
J8L8oTNbXaGX3rXCRDYMM2kOr4nPDH86mANP9kzHTnaPkuazRYZtl81qNbx4XO6u
HiuHmPV5ZXBkbAu/9HkVBy1mq9xRXA58wtrD8X5dW785P7Do/L3d7YkCt6mJPWcF
4pFr3DzNASq7wr2Zxo7QBy0vr/bpL3dIN1lF14D4c2V56J+o/0Zk16l4heiIQS/N
CyOczubnnz3BlI7st3LUMSn5+QnGnEXwqCiOUiOLalzfaKIdvljl4hiMrDHPPiUN
ak2VGb2OeqS27Lol7dCP3OKE6lAfQxeF7SGcEWQGe64dxwonpObAW8xBTkh2T0uo
o7OfCuIweyGrY9arsZzLBZDGzDWA9yphBfYZd5ZHA4ZdX+8h6O600Ta6LwCdWVgK
PXxfO517IRi6WZi/OkLJJa2Y5ulvpCcIKLYtBbcP5Skk2dlVzZ+nH8bxtGQ/c4qV
wnHT+erXJJtkU7oHt40De5Ji48caFnXDb3vsE0JgPEqbJGluu1jC1gGAKECDV+Pp
4ApdhkUnzah4yFxjdviLKXda8+tgi1fbZ7mhW/N18AnVo2/VWF65djYgx9Dn78Eg
/u6/gddnrtek1qzBjYUH1yGqixy93HV2Mw6ptpnMXZJ1TvRBUzXBsvMs3bytVbfQ
xONGls3X3pGyQM7cFn09SuZLrQ7haGOYR/QwUQ4lG+882/H5hNg4oQq/XzasonZb
`pragma protect end_protected
