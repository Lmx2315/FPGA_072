// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:36:58 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Em8Bgi09aLX/5wCSnAe8V2Chco0TFin+UCqvEVjjSkCGu6Mgb+elGtDDu/xuKgo2
hxRIZXlqoaU6QsrWi6uhTZ5MlEyAYkHybrx/DS+Pez8bz6+AHRqHdc3KkLOSPy5T
QFH8MF/yT9QEknMCXVAY8xvyOjGaQ16rrmFrkjwARO4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 16304)
rShINpok22xrm4TNBe1lod150ImsCXrt15f+0xVCHCzk4+F8iyR/SXj30n1hOLDz
DcqJbnW4DmXZGiOs8Fh5wYq2N9rWlqxZHtBzhtCu9SnNbKtx9WKw7119Ne1nhjs1
qyLvnriNCoOCGNcOojh5Bi766hoHgphh1zIvFMJM1nU+jz6O+B6kJgqj8niy9Q/Z
MRoM32SICjPyqzZHK8LqD9kHAKSw9P4IFhCvyW3oXjKvxXkCrOZxusZz0YlwwbUm
pb3JqzjQw5RR3ozxlKanqxRXVXd0EExgCakkPDCXpPdhg4hssFgABBZP7Cn/X/56
ehoPofHng5IYCamogKWiyV4M/ibjzyw9cxZwl+KrPBD2KNxMNESoVWPG5AEEavW1
ns5BvRkszyV31VAqVyuVNH3gUcI98TB2ySSh7+Uj5YryoVQMIBYhJwus+niDxThS
OvOY3Qt/kIOL65v2EcIz13fwFOigcZIKwHfHrSUumUxeugo9+9MlJ7I42vEYtpf8
1ULjY1Ako2WyfoKrL/HhBVydlURKGdVXFjQcqd7+tJebiZbxMpFBhyZk9fE1gcom
8YUxwRn6uW5PR4omrHv3XrGV2bSPeBiJtjYh5wVdYvSeJ5STEiwLbEOcgJlyNXR5
mIdvTT9Dodw+eD0ZI02C9AXYxSPPkzZEc2u/UZpAIg9p3yGgkhVUvaA9mbgx1nFu
dfO9Ztagm9O5eGTlitzj7P96obrWnZCk4lIbycsxYqOJP6BjIQlIRNE6fiJ2CT99
GHawelDGaeD1VRdZhKirZyPNm19jaq24I6CpmSuLf5zYdM9C36RSEKnxfTIEGV9+
LPKeALOjliSuQvT26Zfh1QCkfJJBywlIJKHARdQVw4uYu4hgMHdFIWuS6FuGGUka
TFDkF7Jmh68z54u3UB5YYDeHdKErp2YIu1JnChF0Ey9xBaQeGU+s7kJAgNuHsfo3
dM1aF3+MhNEBJCtsHg6B5iafKyXxE/zi6eeUkUrdLUUFcT4QEE/EpKFtiheljCub
Tpizf/Z9uuMpaRXliJuEFY4fMOMiLlM45qy7dYXn0SLNmaUBkkBKfzZNP9VYB/fC
xnybl7MFqYG68IqDU+Cb4A5+BE5UGIjhYyj8oIvyIKZSxJxPQmo4JODnbtqfp+GA
0LT3RW1aUDh0G0fju+TER/rg69zm4ejh4sYtEEHtOcr1HQupDhGABDa8yA9cgw+T
wazhnMZQzbvX0ddhdoBv8Y9FvmnBfgirHt1shFaPLpgBXm7j4XrONHqjG/7op8yv
eHO00jFeBdt4bAF0fK9ZVTpOMF0IRbJs7STFJwrg1w/rBmE0OXFYc0fMpKBSThG/
Da2TMd17djikj+uOAzZHNqypMFyWalZHciYCS98iI8XSBrtz1lrkBrOCea2/xNPo
6OJfqcuBq9ibO189EgIUm8ukZqNBKP8n+6cFMjH8vNn/0LHZsbwQlVXxQedDF7OB
yLlvFjfCWgrPdBjGwNI7lD0ftG3q3rryueKjFlbD96hV4kHxYUUN2CDIYsuuNMs/
urmFtDNC5NB3w/2O+ODGFnkd2iVKdqeYLMhMY+oRcUwE4qGy+kTmlD94pIpquDKc
dW44DrwrbLcWQdHOCt9dkKRzJJAGcrVOKkHkm96GGTdhJmAm6AXyM6FWYUyTKb+b
9IEvbCiF2jtQ6KwCJsU7Uga8rf1WaoTkOfH57ud+Cm4RcquP6ZzqQUu9sN55n4mY
QUsu1JtjiJXTUWUw5L1eZy2Dcun1vuWiBKmm3a5N8fEwiK0n7crJ87P00VBSFPSY
QN8IKdPuEC7Bk2QQS/AGo94XfbsUo0cWO1v++V54zY1z0/FLCpmzLBkZGwMysERY
NSR0aXc/DDURMboX7aPb73O5BqmADBDUWDDsvuPvPLi13q+OvS4NM0msK3GU2FjP
HKlsR10hHPrFohqXeZLgy6YOcE8fY9gRKzJnGwo8lCaGOjQoDFh6x7PxYKR6u0td
z4ycnumEY0kEhyZsWac0XB6FOl6h2ZmtDhTO2dzZk1he7UcTzZtlYUw4QZ3Gddi2
1o5HNnmbQEJa5CU2G8bojQzXmbxHZVlI/3hPkjwEkAK4y2yvTEXtnPiqTqUBBWla
vk7GgAsIE/+N740Jn92KwdncPW0Zlek28q+/IM2UMDPnjw/v5mlALDLnSGxfFkG1
nLrE+eZQXgceQGvrfNf5mekkonHdODd/UwSuV0zfF1M5nDRpRmzXTnL0bOzLtbM4
XXZb7gkNmpfncpz+X2GLNwes1E+ro8eU/xBFO446srzKaynFLgRlhus8OsEZyi7h
8+8Mj5HRMBkaJZ9ayQBTYIroGFh+BiZIaabJNkArKESO/sZmGH5Oa/S9QsK0CBzD
LrnptQhv3++zoeakm0Zz/f+g3o7lmVSk9Wx1nOSkxkMYZmBN97+uKyWMzehkEiUh
tqtSTPbj3te6IemiGRfAH6le8ztAIi1c1NpGU0nHi43/JcPcXljNBEHfD2ImvClj
8KRH9PTSOLRVp72l1ZD84/bjDGHp1Mb6gbg+LFoQalrYz7FDDMjsZlZexxWsNO/t
AKO+cr9P8qGaamM6dH8KvvgtQuHkzGurFnJpLQ83eNvXBfRRAEoHgDzM/v7U5+xi
+/QYXpQ4uqPdczM5LhA8z/X4jQTrfZMg7xPiCO6uj6BpatzmM+ufzRsDAXo4xMfQ
pszq49hUn9eVAicx0/79STyMMmN99oRonOw/vhSuY3/SU6vKOLvlv5phUcNa48wJ
ec+z4x84lRL9UXyisYI5hsMK30c7QyTUDMZo6xRzrDPpbI4/rXBEW3/AgGGyEzwN
Dch7J5Gcqu77FOdl8H8a/kOORnXnKA8jPRqv3n+b60ij5ife3DKu5BXdKPyXlYS7
S7kMtTqT/5R1Wb6TLn9JOjIFs8+lzbg1V43NvZo0eUY43PL2HDJM12rv0uuoSpik
1V9LgjsqYgbAiF6ju3/97Mh0MP69p2jvFiBI62HfRbXinKJRDoYBtOrtyfzQ3mpp
pZj4MkD3InV0f8NTBVEHfZ7ifjX3YcSGpgPmMmrHgUIk1NnEMYLUg67SK7vJal7R
ff7InA3eRkjNI8MxAWRGcutXJ346ubhR2z3T4508wxxfj4k+jfrQM6UD5wxqIh44
F7rrbKHH4gaO6h/XaVXTCKr/Xza4cw9MbrCJnQrI/IPV9nE8V2JOdJbvXZ2NLx/G
sz1K5dpR60R3ePs6PXzM0gAwMIFJhRKx4r/Q4iEUO0Pgq4AD1aBTfw8g74B7YVUZ
QYijCmmKnA8/bWFK27g/Lpx1nAub0+SJsiisbddlkYBvp4q3pKYV7dRDRUpCf6KL
2Q3i+2zonebCyS1++apWxiADyV6O4eMTLaTEOKlV/EH5TT3LsDFlViip32QR+j86
DvTOMXfF+L+0tO6MhP+Uqnh6FOtjvYEbTPZ79LPKlCa4zGMdliM3/jwGFb0aMMnb
wCnshhcr2P7tDzw1almXws7xURa0uR951wJkTP5ye5ZwL2yX82qgl1vWHOYl8D3V
fYZgmmDZfl3AYli2ZlbhNZoaVgvM7YvrtMcL5BrMGdPT66YZ4D/43fnZ010kSeJW
3DGeLsIXvF9V8pUv5pEA9+5LkZVINlcN9VuysT3MjZdRIuKaZLgmZm35xFBxZOjb
Bj1QX0pqXmyTtB70xBedHwA/BUfoEW50PKNeavk5woEogxSKqIKypDq6IrAZ9DWl
pHMful05RWLhGCcJu1ZfUb9TgVGVRz3E6C2UAa66U9UwOy5vr4bkqiEhnbnDQmz0
veg8nxtWOmzIloo6qigmPzrTZ0k7vvaQ5vsWZzawlHG8GebUaAcCfr/g0XJKyCfM
IA+Hrc2xoR6f3AWWUjP4mH/TqiCeLqicmz8ta99+nM5NzBUGy8DlV2uRYrQ7eLj9
5ahyzUKcqrhiT8CA1zGyRuJm3BgPwp+7RdcIj/eqPMqJ0fat2tai2oLcJYybDqRb
+u1gjk8NYLeqD9nkgI7j9zzGEDzSD1nVlS0HcLrSuwDV0Vjm2ogIC5xOm0gKINIv
B21zh/DXqARvl38Z22u55UwtuX2Tb83JBm2HC94JrTCSt2peI7We0gYdqLRwp+qS
o8daL0o9nAalFDCWBMPsPeksfS8xdVw3xFc9GyqKlG+vqeW1l0hGB5oN2WBf40Jb
GgRV+++UWK+ZC12B2zaQzhSo4W4qVFgVRJy/c3eTMyX7FLvLfgzfDNeGk4czjn/V
bDYeiK3VrLXbbBswPfNlZYUqTuH46nG/CyUsuge5wQj4IIVB6dHSZIV+L+4KRn0q
yp4e+iyKCYLHSuwG6t1szFmQifO38l651WmiegVkdMC+xbSRWqsJnNwDaoeJlkyk
yBbKilahGaMzoaFD+eTuQHRvnNIeQhnhUQZm89UGQGpO7Bdj/ZH6KmTXozHT2xak
tBFJBiNLg+I8MfAHesYf7BcYda7VQwyX66d+ZtZzoJgEFcfZxeA2G219C3zjJsJ+
Hyhi12wLxvPDwJgwt81ek12E648c1kQLSIYpt75OxpP//x3YjhJEUxMRII2VCFrs
6vB9wW4Uykl+0nOwLnwwCCavRwm2PepgBNgbyWy38huk724xKmCsQaBSZLYGAU/i
ejkF5pfvBtBKIW5FiQ15Poa6jIYiE2U/geR8fU/CqYs4pT4DRB7uxELEWD7IUYuX
CBED2E3Vw8eGoGX9KW7vxOTXAdhS3LakVolfzr+G+3nuzxsqk+Znugz0eiKMMF/e
9lloL+4QRIhUA5Bqg4/IUFw0tA5NH6w5lwkW89YKzNNCgMKGqjZg4x0rnZoc8qox
wmuaOShbuoRNR8MdY8R5QpYUxQu+/b3r/n0senqbl7c131x1VMuDl+FuucG/hLX7
se05fwhDjOFtNQ8XHvWFxQpQXI+HWcR8lxyEE7SzZtguKSE44OssSzJIx97/28Ty
WXwl+5uZ91t2p3O75Zx/5IgKUkfhqeSBc0ftlApzC/IhneN7UC79gQekdZdH2sET
5XG9j49lpV5a56OLz/SdbozWJrv+4avWpFQb7h89TO5RUPuxxke3iagDii9SZwrA
SgRmaFTNvwf/q84D6po4DArIm3s/NIBGoSXeK+MnJTKRts4MhOqlt1cqoigRYzJI
nYzcPeSU1USsqrERFrAeBOzeyuKT/vI7n/R/xpNzx7bquLLTFAIhqn0HpibAsgNx
jolQDtP49krULfDk6Et+2VxCOTTsmPCZXFJIQO2xQUdQqgwQA+2yLyveOQD/m0oh
AWk+5F9GPTi6noBU2mQFUhmDsXXrgTu90spacA4bSyRLUd8IVwPyDyvDc1KiqvRD
Y7M/o4v40FQoPgFvXqdUQOLOp70Y1426iUAlqglUL1qLtp/xxRIJwwfDKzsgck5W
Fwu5lr7nGnVnscxgme7c/WsckKTrXl0Zg6/hlYWAk3SMlPpMrRRnuDu5iQ0e+oON
iXmFNInutqtPX6uyr+8wMzPoLFVG+BVCUjWV5ig9ySCViNdxUhh2rjdFEj22z6rW
syaCrc9mD/emOfoaB2T216dyA8ohMprt4x7cOibcmG3TH7d7hPhlmYoOS1E7YEcV
LEwL1Brr2JE+WnUwI5t+NTMUTeHmPAS1vF8kARMvil6ozXyThYMvbhj5Bu8+7pO9
HAgRAUDIvHa//a1yOg57ykwsBfKOrXELZaJD0BZBuV3+vsNgk3Ad3oiPKEhSTaMV
I4ghqMS5fzCoBf9jIqtDv4xLFSlBhb4afsWleZTXogvK3XtYrd+JjEm9VjY1kQQO
6eZhdARwQhBeE/7Ks6qvo9mGyJ1O4RUcpYydCQu53FxrUTZPLKTFNniwHB2QXBTk
uxDwwTnNCxzNi8p0KiRlAo1MLcb+KWle4Eh6lU77Xo9lqCopNmzwRmgJtZoM2m51
NYfcApSxaEz5y6MSHoRemZtICI4p2qTzahUTkszXDMf6mGhQld1pqmiWX0J7VRVi
ihuckaDcrfYDxxzHB7oOKvevnkYJ8lqDtfJkcy27waIrhaPp2kGVZlMJfuxXRgHf
JK+BpPxanNlJz1/KWN7fHBSONVI50Jhk3ljcQu1s/r70MexgDyAw4rutM5L//FX4
k1Ps8k0jSdE+RGp7yMJ7rvHXYAxlatKI/3+sOvajOpAiw0EHeywsjiTCTnmlgki+
fh1deLdguoMJtYzK2nrFiXi3z/pqDu4ujvAu805yiY3ZdLkFk0DY67heS7vuZF84
R6q2mlNGIRbshg11bZe3rF6K3ehGmez9OxJAw+8CgScyt6welt4teKFPzrcpxrHd
AP+0C476m8GsaA3DvucDiK45khI6xVb2fWdXTX1ihFGb9T4fPzXIcrDrPsq1IdoE
NK3369mEaD+Fcw073LpizTm1M2PDWYjkagBRusouDEmeX5iM1OsSx21aLptlzXLb
eB7O/rkRa4M8ZoudVLmiqTDjNmPet5X9W1dJ9RqjuSeAhEwmX1XCnqHXgjDG+DkV
Yvrczy/cw2nKx4OoC3MyG9leHiSgTj3lAq6xwtHhnu4JGrvGYPhgUCTQuu/JGV0Q
feRybGhCJYKG/1hwYxkLBGYUHa3MH2sERO9yTiSlj6iRZ71jAxQGWJfnULrqwJ3O
93B/ArAv59ls72OEiBvz9oDlHpo2xWfsjtZWnhRrqSV60TG960YdfxeGwZ/5KOnj
1NyXLS1DGpgZsEkV7O+UdcqAaaT4COI3jUlONYsHCiWInEFOjyla47CeSHgJDfIo
JmXYllZyJYEGreYTqbY5LT1fK7vUrE13cVhPTVokoBlMHIGh8RH+jj62D2fccF3h
Q4iOIN1+gvr/pISHzce2kdziwu3bByMzMOn04XAlT95mfaf792FZs7Ba2wiMCcdW
eCFF9EmJfmO7IRmJyoopg3ywoEt2UIK8yFiEvEyIBn3i5WyMk9XBsXnrWEEfrTTh
yBUYe1UNA+rOE/CPhQykRHMVUKAgidAOzKcGs/TrGdfMW0er0O73GMiN281pKYrk
WgoJoNijfIALX3sW+nS/oltn7ZI4T+j1hcQhBxTNz+si0/eKz3ovJqq2waGpr7qy
8pgyICklcnVPESmHyD3zOxMFZOBon0/I770hxkS5ucbuGEDTamjJE2iUhuF1dmXF
CCve33XvkGHD4DU1iDwP0UyWW82olIUOQmdcDtYyHcX8x5+74YgZkFcZr3Q5Oale
NdDM4IZSFJSg1M8gi362NHZVXAflNpB/praNtZV2h6SgUYE8xg2vAIZl1CdkvIvq
dX8Xlri1O0tTJMP9jsyZCEVcgP5MhXYGf6+xTFFO3mgcrL5n1s9tSAqvxSES6lg5
G19VJT13C3MXn+ChvXnGDOVVPj39H4i82q53bUUgD9GPeZihZrt5xbti/oktVDaf
GiT22pggO3NTR6jVeU6x+62UNW1+UL9g4jDniol6hTitKAM06oItimOSmaACAHUG
TnwIG10vupXAPLwaSHn2Jokm8WybnDirqHCXLH++NZ1H83wuoG1VZD7OX2J/Z8zl
SLx6+H6oGxVGrRvG6vptYwz7reKoUhQP1p0AI9XQpi7ybt264YJGik83w08al93x
y2lJY4GlucA+FKl2hYlisBwROl0bZAnBwztmf0Ygj1Hj2EMEUkkJnWWivnO96a+W
Eexb/RzuqkDbyXhl7YcErgsLDeeQW0uPyeHbbc5Pwqdl3t5kbj6aNnU/lHPeLmMX
be5KXmrTnT8FnL1wVEdPaFRmTj/cExOf2lTczxzpiTWh1nLTFkijNWRrmvp+SIZb
Z7EiufucpVG7t+MdukAxbuQufTybydMOVWqZ+3NonXWOfv64OSpRmexS178VocbB
CH2TW1AlhloOGORm/PARrrY7l+Bh3vxYWIlpYYtU0iqBVdHfjRHcR4hmwkaYJQ1N
O7eYCJiPAfKL3EYxe+pjcCJtcz0z9u//wlnygRYgmpyjgpmQYgaHs0hAltKAPaak
I7MwGnXnfYQvqZw+LPHCbA6ByGWo8TUuYZ14P3/mxpR/A7iKN0Q/ewBG01XtUdb5
W4g5TzZE9c6hDk1iyuPFMcTU/1B9lgNV1oF5cjNI6+ggm9H/5SJ8KfYzIFQ1yEMw
3MvxmWsT84OfzaxhTAuxRjutEGHGzfzOXfgrok7CCB091C5KVA+RhY/f7CMM5adR
w5g2zNtFssK14BWwKKlEYCg7xIK2XykGAiuPX4H88baSVRT/hwOk3GY5HhBicf3N
fpQ/eW00Pe5dFG79GyCwbAGqkiaw0D50DHq5u4xYj2dJ9agzEyFux9NvLgAS/O6m
Fznxflg8Lv6WoMjy7G/vM+ZCMH+MDiEsyMLk1HowFUZNsy8zqA/vcerHvDUUiZEq
QwBWXXLxKUNECfKPvGyFsp4UG4ydMeG6HTIHFNllYScner/Prt8+gplaOrPe/30s
zu7Ul4gi7oQsu3GF7cJZ5VKc1AnTU480nffySwnxk2ohIkc6hxuidO1tEJU99aM8
C4hIoJPUeKXYMRM7O0k4Wj0nNsSFOX0pgR6AgE3DZjxQDgIzYPLHNnhZeeA11Ziq
f9sorupwIwGIvcrmT3vAZb8N8LArXBXztsre0/2DOZCijK6EhTpn0vhDQnuWwB5U
2WL5BJrjlCQNVJk+dzXpFMTp5BNx3CRoLeHE1SSFEk+cKvNI8ifBIeer6NnjnfsR
NRgo/x7JsgmPrS9ER2wRFZxzVyR54aXwmTT0pS43DeERT/p9c9koDl/dkKpnw4xL
qgNYfKKf7H+7Jyl68tA9794vGub0eDshPcd2zvTX4xJegS0ytaY85KIR+1ovj1rV
84xAmrqG5/wMveCUNzkrgZmUPl/Tq7rJloL0Hy2hXp84vJRagg8RNPLFdG3Slhr0
3dPPQZ1UaIxL1+YbNKZeNFAacoSd9dNE9EKKmKVtfPg72P1lbwJjG1xmJTLc5BA5
46EE2MXXaN/DOjRiB/lq4XPdQzvyWtQ3MWpjjm6sn9pw9FTo+TXC86aQqNWSL/Cq
yC6RBt+j3LecXVkI0hFQhqjXajApn2SKSen3eJexFbn7hX2mGcpRT3f1zg1Wv215
6U67F/p7/YJxEhQvsGepB8EeBTwK1ZI/VFoLJuKeW6qhGMy/lAd2rGsQpGVndQIN
3X0iprx/sOZAjCc3JS4ngEizEbwBIIliBKJBIH1EzwmuN3lEIsKrYwTi/7ayoQre
uQcxcUPLhRLib3c+eC2km0YMTIggtRv4WDVvmUq41c/O+3ca6R1v9GNfLNUNPjUA
n//UCCsTUR/90Oic36SMA8lnoZ+0mgDa0ePXp+7z6UYIgPbG7dg/wEtVdGIa/CKC
vCSvay+bnfK6rEOa6rfQwglyTFiirIjZ8mxUSjwhHBAh9u1xE1QKFRZSjbrUitBI
F+m0MBMVMTBli8IVa/kz5AH4UEZbdHk/5HdAKcdPnKqcKSkmwAvyCi+h8D/3B3bc
UX2FIipe4RRUQwidXWuHjCU3CZyA3o65LIxLchFCQUoa5S6sUcZSAGwZxrms7k19
uhIMJp0qZXeI2QsUduxtqw0LebdGMofMR+cYJaq/GHGZ5tRqpbnyTAwsV8QgTe5c
L+d2ozqYdRKPvx+LnUgeRG4vNTwClIRhkEhrq/dt/93QU7IEK0aWEVA5OJ7AU/b3
nlAHMXnFjU42LbYhXtgEP68oH+oKSfTDUnFzm7iHwmH2SQteow2mHKmzPRPEFpFI
Pbh7jenZeHymD4FAUogy69RWOSWUPOMgEm9NFdo/AfBdBIO0jXPXdgq74U5QToVh
Jx08jHrWjWL9QUBh6oj7Kl7RMy2hFiL/n8+VvvnVw6X0tNxGEP04lEeycRANrbOZ
VQ53VSlwfpLiLUKvBP34UoMCkxKkQT26FvOBqnWfLdZ6hqfolS9i7toK6fxzN/Qi
1L4Zb3EhDxLvyHCES7PY1U+2Fpq1aD2ST8st7n4e335BMficXYd+VTgiS5nKbo8g
YlCtAeVk21xnXecVpeSJM/AOEBYXpBnNFhI4ZQdAb9mMG/bGr+BlF/fzzK5dn7Ko
4qfEuNhwL49ATwr54zFAQSMjDHhlnAaFFtmcLfF6QWNgQWFBfodQjMBlmTuRyKZW
rP3LjIaljVxHCYHyk4oJW5fVEviVpjIwLsTalRilydqXcS5IlzQ2M6axg0YkdV3R
wKFIuG0hb9AioLLYsHcC6WV5n5AhDPPG5/6/BZO1snYYPTmVAhCgZh3Ftbtq3E+O
k263Zh+Eq0ea3PEw4Cu57Qy2IYp62n9Z1xlTh+Wmdc2s05C/T0VcYMbIu4r9f8uM
ei68anePyURQKWwysYudjrcSpbgjX+0U4qG8w6JjryhAy+nH1JRvZqq9lFvRKEfo
ggQp7FdPRvnMHZoR5BbrZmPilDt/e8Rn2FZT3PWEVia6ENMCgpGj1TgNgNfcwbvO
2QDvqjli5dKe1yhAtOsz3hdXGFIpATj2reTvKgikY3b/NGiE/8tAxNjt2cxmI9ko
7qIQFa6upEGbLY5aYUHA0kEUtGWRgqFmU4j8JBNa9gOtnbVKSD80Tkf6ssZZtBxc
Gi1lgAchxOTsAXeAMOMtCkyQ0lteWIpbekku2KBh0NOfVbFmOa2J0mWoarp/uYz6
QQI/X8asLWP6ntAJyfIvSx/MVweSXE1TijfYzj2GVCfL7xBhALjsLjRD/EHRZGms
t7pDxYE3CH3Fe3vLoECIcnxnfAb000i4htKBwbNdkXW5OTU4VNH9HkhUo0X5L/bv
qZEOp5mf34TZRsMp37B/H9wP7lYu4CCXU7z/GE+vZTQMkK3Es3V72XqWSJNp9qxt
3euR5+dEcFoyPPv1/Seujm51avwRhfhNnhqG/UAk2eP15VLlDoQ9yp3xsuKtSWBz
3H+WMRSwT6uqw2JLkU2xB5Vzi2GQnojIuBuX/k0v7y5iX3PEGgLKCEp1LexGhQas
r3uLIjYl4QI2V2zU2FwD0pJMy/5q3rmzdGdgXk21CGKpLtcHwkiqtaKu+BG1cn79
ZWnl2C0j1TJI0sgH1+0LG4YjhawD7LfC93LTlD/DWwtVqUWnFFDV4M9EVez8JGZ3
GrL4Q33Cn2SEttxrni3W1SjFlDl9BO8fMK2ox+xyk3B2Dq0ajHvycEbNGy2SYku7
Wj75kv/zTYWwA18+eUTU/11VRTJXEPGSRrGixbuz+bTiUhL6CWZWU8p/m0xHej0k
mDCGHDovA0m7iwgQGdBZ7AjC1nWfYFXMuhtP2B2irdhwuFHVbxcb2xNvPvGr3+mW
WMBTcFvVdYWnYsSGMh1K0Nh5F3icis9PEWDh3C/Rko2MrA9SLbpCHE73xeDKqgxG
oxJU5iBYkl+Wso9X1whdJ6dCxY7Bq/TUnL1SSnael4M82HvqIJ+o2+3fKhIFew8D
HqvSGiKvpf9UNXE/Pf082eGMHiUWjN0WqLhUNNgpX7Rae5tzbQJwp4CGZ2Vq53DS
qwMjBwqL6mLLSbTPWXxfp5jz7tZsdmkWhsxHB9fXTP+9KMCZ6i3uKc007Zm0Tg9X
asbxBkCA9b/S2wnY4JvI4KYinFjJAscCGbHyqAUqGN6yZabdDXj8dfnGi937ACZd
4fAvUfGziOV8kHu7XRuuf3aLbAfSvrEj2K1GHmImnxMGBUHVIRD0DZyCroxEMvos
hQuV6/mLv/OI3mlQNIQzj3gWcw2X2g3koSNz4rFrq3emrk9rnsb07g/VjQ/yxQRy
cB5pTFl44oQatmeFfVkI6Xy6epIkk7Axa1ytFL2Q3PEUEPPaNmWrv0GwnOACbD0T
n7+CNkMOTXwjqhk7UAkZhKXrZykOYzxEmZ+y+npNPHrGIitLO/bixSRphfzaTaB7
jEGK+a0wvNhVNdEQwTDZylUhVnFK/HccOf+Sag2b+GpkE4cBFIeVyKmEuepagY3V
pKhGSvuaL2CV6wCi+54H5KV7cjgb4ljE4En1gbUNAIUqWj0SsPaqG5ihl5RcYKkJ
B40LM5M5BOF2hsfranOkkGq/ksC1i0tGDlNLOtSdByo+TxQ/sjEOxmS7SKJW0JiH
JxtZip1JHlgikX7YwMeic2VRSFP4IFNrqnjKgD5ikU86q9E7/YH36MCPduezgcOM
aLRk3D5rKsE7a01kz9Yi5LNsk7VbP5OuVr8/C8Jp/B23qJLMaVzasdaXa0J0sf+O
b0Jms0NUSjDY1mvTt/Jw4K4f1+CswMIuIB5kPPDmSZCTqBH873x1DeAIZ8bPbQpk
EolXFdSpylE8KFF2tL9s4SJVK1cMp6Ai7nOACs849iwrNqhlo299tWnwFx38W62V
kYZZQ/zwOQ2Cp8ChvwbqeralPtIbcCIZd52pWT7crEDttSAktVHIluNycy8HIld0
KgbFTNzAoZmJ6INJalkJ8Lb9qOcJBEOzzpqOpN/xRSOy7HxfxlO5DiiUuRfHf88J
VQ5dWX/MhxJigtnthqus5mn734pcJl1JrwLn2USWLcYS9T1F7/Vt52ZAAh1SvY2U
Z3x80gpxFNnzcz4TIoD0bev8ZPyJTfQ9yYACC60Axhvd0FI0va53XTHkKkNJn8EW
wZE7Bk+TcDznSsnpsQfV2FXhIizqTLru4qsZt3Sz2ShAxAXXtLLuL98y8qq7U5r9
X5AhcsJRI5LIsDIJsTD6biVai28toc1OeeFLJZiiXL8fJkUvjaDN+2yBB1jZDk+i
3cByY1HEbANsN4/SgdDLXVi8f3cNwISpjUPdbZ/rMYeGcKKloyBYOjB7XO8Kuz9s
sXmj1U1cbKA8tNdf8fPK9MDUm1R1Ka7vX9p603ql1//ZBHfIdWnUVcxFufytrgX3
T3cqi223577tXmpPbxYmr9gROGN1frkJyhX/iJrrIIDtqNsxej1buSuI6G7bsO3/
nZD0ycSLVIw8HXhwJsyE3ge4radZrM3gxs14zTlPZtQ2Ppptnf322QsauFyirDhW
QEzcsgaplAGaSmxoQ2ZMPFeDRAfYp7TGfD1FxMgACBfNc/lyRKpZYfusAOE/RimS
BLrP5TINj/tpkkVEwufzNsJ2aoDV2kNs37V/Hcf/fkwvyVKynplqS6ro+RL99Etp
xD9UoKmGm9d7N+YfgYzD8ni+eaGsTg7S2aUs6M36a5lxF1XlZJ1iq5dfyPvTzLnY
GH1NIlgETWu7i5a5yN9NcPU1hlqTtDdx4kG0oKIzEEVoLD4kodFZ8c1lJPiDPtfl
KELefl7xZK5/dLYVxrU1MBX6WBFikdj76xPFWDjVxhAVV6JAqWF9I4jk2m2JVJ2j
NVmKY01sdbv9i1WnatwBQAlIuMNSwq2eZjNK+h3YnogiJAYs+vXuVhvY+h1amOWz
UqKU2gHbRMRiGuXR3I0+NyZRmafc6vhXF23l1iSpLA8q9Ph359ZW8yd5IQtMRFHH
hjc1xq3fOL0FvIX4HvRw2z4gujsv1QGngUbjlLd7MCfcUuIpXjGrii9ClldxUHH9
PTJ3otfB1G0aRi4CTQ5JA7+05L5+/ySkvD/EAuXw0/sS8ghZjVK2WlD34C6iHoBb
wZbVDWHfGuI9wiaRzXLN+SVZflKqdWB4GLy2R4iyGem0/knnyDEdIXRxe1N1SI31
B6WsqWqCyhSau5LNojovyAoRUxmh1T8BWjm+6VA28RwlUGYE2iPR3jfOz1shwm7D
aKHQ+EKdH/BV+TL/XUJybQKeXrWo4oTf6WugK/Uj5C6IlR00Jf0PUG8owK2hMg9h
W04mIPJUDLqX4A8w8U2LsjcoYH7+K0884+rDqul7bNjMLfrAa6/af8mbRe92r03f
ns2irnVwhi96FMvswx+xkioTdE2P3JNb+pwALrL0U22UkAMW9r3NIMEJ7nd/kwqs
FhxvEIAlonBrKZXz/VXHTXloAknynUpaZivwu+nJbzR9MHhgkr5rsijwPA55XuuG
lITqtDYBzoB1xyFSmyurOBPEmnWcEZPOtGDp+QrbcAnY3URJXEB59dQpeKrHgJ4l
BJbSdN1bICYionvFnVDIAU5qYUChBBNLkL/W0dFMs/SHPoJxM19kIfDZ5jIP8SVJ
eP8GbKJCJwqG2jnfJpW8YjkrHJL19mpFBX3Mxq9A5D82Onw/GbA9abPud1Exk2Ti
BVKIH1cNixU1vYgvwtnOe/diF1vPwCR8U6MOjYxen+CzeDR4QsSJPrLciUsn2XGU
zNqYhdbF+4X6VWqi3Fuq+z49mZVUfb3FcABCo/K9NzRxdCNrKWVS/yaA631WrNmu
g6n4ODV0xoIoTw7cJpt1lsQ+neDmlWIKf/iL1IkGRNMumGFP0RQpBcY4rrN1bh0d
8k5nCpkJ1rgg1FwQrDqrdeJr8qLtTIlQTvWxvS1rM8xW7FDfrl+kz9dbRsOjHUAK
VADIg5wSRzCIMTeX+K05sGcm/aj3j+GAKuVc3krcuFSeCUiLi9Yo59/xEzleAEED
iQkmNfs8+t3AN1RoaOrkOPJZ8hnNWxWoQrX3GjE4KuR5u9JmGypKUrcN8/3UsajU
s8Fp6tafs5qFgHN8c9kAupGHotM/K0uC4xOwCMXwDWdfh4P7bWIQM4i7mpF58mIw
2wsYBYUGzjUFZ18LY/8XFP7Cg3q3v2tEtJHGbJBpMX3YPx/uOJ8DO8nC1l9QLgpY
CWrtLQ7q/fNf5RM/PjaRNWu/o5MUAzX8XnBf6fd8GdFQIXvUFEauUX4H68+9P/3W
THroofzPlMhnU+UExBq93SdxwaEvt32TneQCPCIk36Ka95UiI5GNZfsuVhbRCYVl
wcaFOJJ94msIpuCDKObPkD6u25iTn4n7E6o4ELeuxNyQV92v9fL60IY1j8z/EQ9i
qPBNATaakTjsuwC+EQXxTKHOMEnoQCqAumhi9DOKQAT0k5pjemoKxhxMRU1oC+gS
aZQivOqnwQhIB46Na/8AqcMKDfZu05+Fj9vZMNXcPiS2tm7K90Xrkw0A2i7JZjSC
Nn7nHur5xzMGA+PdIdiySePnDb4X3f9g9Q/4MLfMyfn39q6xGoZiJrFt5aIMrt2T
cEXxXjYhjUQDuiCcSeSEu2PzgyFDLIOYewT0qz1LzPXe35Roph1KGKZsKiwrRNur
/L/wbpDBQa3e1Pqw6R0D0S2nijjsMyuU1Pfju6v/xagQLQScEjDZ8x/+Pc2shsiZ
+AYoUQZfwHJ6Dw66967lPbJDuH49xg1gBfFOnGNo0VlSM+zvNmvJJPkDI357z/S4
vt8No0NYnwfeR7222Kxz3B2TeOMQ3p/6NyTnnJ+qRJlIB/SabXm9ld9kAyobWX4i
eKboZNGKx9Q1NBK35Q2cSj8Lyh0y1DdLtjqC9+JYiy6/saja3zLdLIPeblq6yyIV
Il6bw6xLXDrb5Ap9hEfcmyBLzxeyjxOHmW8XiyAMi08C7PoIbqiZVMLoDjDvaWmi
DKe17S2wF/TBViFnIC3NjtcIHU6gKUII2lU4lQ5QwqqgHsrF84UqV0qqQD8jBvOC
RObOUZpdoQXX9s5LdfHFSYNbSD7yvM3rKXEyhzY8aKRFFprAAmpjvWcf5xaHPp5x
FGaqjiI9pNeqzJ7oDNBiR7PpTPBfbX0Wbl5FT4z29PobzcyIIy0aNcvu8lzZK/pk
e9KcCuTmKlPKmAIWrWiZroGK9A8B7DlVwVtN/W4VCCqOGt8Q5nplTrjVcaG5e+wU
ljQwudluouZfmqXDSi9MjDIOQUdNCmZuq329VIuxT0nDNm6mh/BNoyH2YaJpKdIh
rWd1uR6eyhWOIRNmt6ad2x7hqMH/E965A+Pw2uJ22Ci6AYZ08euI7PKJR32b+kZH
qr30v5KRvpmtVMnnSsyxAJNcm/WYhhiw2MX5/MG8z6VYcXXCxhGFw7vfH5fnuChv
Z1i6Zmtz7tNOypRiWxc7EeC9hSUATNfGZlMswYp+UvFNQF445bSe9MvgvEjmP3yF
LSZdw+yUP9CV3t+40Kal1iEu5pF77VGR2tcaYR+Y2UqQLueqGPrYxGa+BPr+00LK
67vB2lgBlcG0+jBL0cRiSjhf8RU4zQneR5f7U10G+d9dMg3fJJIPFJe07f7n6Sde
8Je/58gn17OabI3Fq6HVHxwCwvSc7m09SW3zwLAnmHE+caRvmfZvumjByFRJb2ji
pfNx+xAucaKisBOee7ERyV4DvZ5/TWMDChBG7ytbxPuMp3VNDJT+2MSrRwx3pQT9
7vqTY97kYIWvFVz54TknAevQ6o8Lsrva92qjcOEelyr7SSp/NRsYidVjpDVKJdcw
GG57nDvFuMgIVeLbaaGYydqzlYiLU+e+cRAwMqU1gvUPorzA/zabYR7YhcS1tKUs
X7TgwTh6JhFUaNH6FirF2uUZCugioWNJTtmUccgNlZlsEhGBS/VJjwEhPerd2TIY
C7RGGED5N7ub8K9HEnzLsIgSmnaAUoG0HpSNKHj+IT9veD6X9djftcFzW09QLMma
TOKGnhQdjBZweEnjRi4p/HnPSBjSCfpBodKjhoRCwo//d+dKXhBDjk9QiLorriHl
MwQT4xPgN/xPy3BS78ot/FIkoDBSm37VgthpZ0LLxXCg/Ast73SuZoULpNHOvxRn
Pt85a4YAaeT2GYuJmAYPV3b//uZDTPoEVR3u2tQzJeAgs/3fpyEsbhJbT8RReN8y
hrWT4lcpJsh80jaLTV3TrjwJdk3P2FG45HsQD0QOV7gizJDd94Tn1BndvcfV2DdL
xu+HeIAaTx2OeHKE7GH2idiCUzdFgpT9yY3aOE7TJoIrC0XtoXMBdv+pbLAFpq98
5gpwvfgpDS9LZ7JhQyw5x5yjbi68DdLm/Gww3Nqi1S47AOwd33dkP8xmn4bBZ70w
lQ+r41T+ovK1RMP31DF0VTEPVS0dIoCAIlrISXo+4oPYSd/g1E/OaHk9wGmyVLjV
F2ul1rezfDxbO3x7rCqacgPDao+wuhCM6ATy5CgtL7PI3JbaTWEIuL9TU9DUUhbZ
/mDN1LOwF0FRCpml2OOCZxgr5fBhDw5yFP9K5GwteGa/KuwrONtmpvq32q2KAevB
MN3OZqd+u05ku//T8WtCUHCHRyI42uab6yKadRzYTkkUBXbq/uDHqMM8XEb4m8lE
8FY1AwkwzgZpdTLhFx67sMIDEElVvvnwEpN1skSKVhznw6CoP4/dmhJrm9gSES+i
EScAw0wh2IZX9EuBpARh1PqK7uZI1RD/HdY1TDw9txu3JcwhiyJNh4OP72O4x8Y/
R0/DY6GYV0iHXK4zUfnllby2Q9LyMBuTxCJxRtNac3D98CMp6EmMXskWpzUbhSSv
r0O3zPPlSTLOlJRb6S18ONQSdh9VWy2HyaNC80IwXS8GH2F8uqDRLTmC7HsMgjql
my88xrYnjBzROqMX03iEok8gH2H1ZpoWKLONSM8mxK5od/iH8XUIq5BBCvtKsMl2
Y/I/Ra/oCvfxiw4oTvi7XXp10CphnjdoRQ+sCW3v/rOg+FMVe0C4yjc7yKQc+v5J
dRNl3GLNSJTXG/T3/buuTaww+9IXzyTSr3whC9qr8mqFwGwNaTcWpDrOf+1Dg0XE
5pANQidDnAhDX7PqHTdzNLYCDLFXnNdtoRhKyK1Cq8ijZ34pkyDLxw6gmUSEhMpY
Ib9YiTEBUnBcMF+Q+AoE9HdnEAkFFqS2IcZkH4LRhzIe5bbH5y5HhfDjZ8tD6nb1
ox/++F5guCz993xolEfTFD9xP7tNbcQnD/jpyc6W+Y+F1P2NsFqfajpGhuKil6wa
I2jECwXFcENZTMjoJYuC6nhMlP/Y3Ek9jUx5nKWgnzFhPO7S2UPrc8Z+xMk6uo5v
B8NADpd6Q4TNfxMC7Bl7gaeX9Xn6DVTDO0ZCNhvOEpw2LoihbR06Kj4Qqj7kERGx
BjevlRD67zJlPn3n+JjMTWLbK2zvqS55Fw3Z/Iyof3TjnahXzRIdrwfFQv1fePw7
eXk1ngHY0RjmI2v8lyhfTP26ldu0UV05X83owSxlwo+5yYdW4Xlm62nxLnGPcwse
tXt9Kxoj65KH0Amg680zvhZrsoFosb3SNyE7kFJX7krzJT5+LjdZh0G3Q6fkS9nc
ufGFEuK3OZ6wWnINyfU2cKxKgub9ZaEEj+MEUcbh05ify8vHJXdU4BjcOL1eE1d6
3xac6jixDkH6Cca4KcJ9CCpKrWrtASADTg7fx4ql4QusALgp0vX+0IvCm78pBlVB
wT5k2TlaiDKCc4iM2qYmq/ZSMwQpy8NR/M/3F14C7ah/UKQTr3SPLP+kxV3HmmRT
3b7aJFvsmOlriEGSId3eu/B2tG6VOPOjqg5T7Pykk6JVNb4BmwkVjo2eTv/T35C7
53tHtQpVYPpOBg3ReZKmhN8rF8b5VBK+IymTIdWft9niK0Wz9K3GukE87Nl1sxyO
LrdB2aC4dcV3wJpH4WVC6HJTxzALHooeUyWBTlJFBSeAyXk78ZsPVjUCYgN8G/Jt
7tXfu6sd1VV4LnQZ5Qeqbco2ttqjT1xtEROuJYEAYNpirXQts7olTAt2Lay8GckU
XFdXKDVuyWA8Rme38QrilkQr2GhuDEz9GTku9rYGOtmhiR2OG7fO69aCQXcAezPS
kUP45ZVfI6LIkswgksDQydURlM40Wrfh29Qq5YZcSadneW6X1KZUo04y6/W+J4wY
MH2ygYLbZazIfAMp+cR7p0MhaHnupQ3sdn5OZc+udhqsT6iSlt2+HUNcRQnjNIDh
tXak83I7cLiOBikORXO4a0osNY/TEzUZwopaAN212cbv5gmCgkAQFL8nsWoN94u3
SlsEvop6v7U2Wt1c97m9tVUoNIoqbBX7KGgNslZTUFzikZCoNwyCOniyGjAEmKGq
KbTPOzHN/f8is16iUu0aIeRQsD0cAKZBOIIwhl3pzk/Xl7Xflm6bINBw4tVJmxJL
MqfMOHp1F46bttV7+EJrCiWWs/mzAsPrDgIR85LIiZFb1u5eDTQorVDHvdH55QlL
3NuHGgdCxKqbZpK9a9c0ODW5rvo2XLHoOUzNU9Sq4cjDdjtIp0u7RcmVkuCfLFKJ
ANdbMGYU8CRZV5S4ptXJSldRVEMLu/q8WeEtQjojiCB7+DnreLeAFDo5N8QgYfLB
CX/EwuD5GvD9x1HYZsVXN+BZFuHcI+xU2igi5kiP9VOsRqMRw6m+Fw6d+fbaM5Wu
3VHz2tDKYGqDI+LQcfuplaksa6ukw7D7KHHyhUXnePP1xoYiqQL6FJB4kMRIy11N
5AYbSbJhzotzFpGSD/qtO2O/xH086BEbnkcJnMdGu3l084nzBf1dqPdBPnFfJ8sz
g0r7drzAW/WxaK7KckKL4YnGoBnF8L1oksI6rwUjCAbIm2aSBadbPI/cY5hldjIZ
illGxoGAYaCg6QrYLpx7wmNbfPP65NjnAAzIAs+m53XQkU5JZaOJQmR6dNLj2153
/ITOQbzTG5GKX8MSc6hnoJsrosIyCSqfeI7Z7ei2uXtsh62Rps61r2YePFjEufIA
IKRukgYLgYn4KTegEnS6sHOah9vHzBePt3R8bwqwKFbP0cXAZGfDvMarQUCMIjWX
P2L1AvXiXxE44NeNa7V+opZH5XG6Kv0cw1uDNrOdUGXK8TZ9ULViEe/3en+JQ2VN
ju4xRTN4reX+DTbsZt2Whe9j5glRfB+Ks1+nOdTj19X7JgJKTy7CdL+0zcOjtcaA
IohHNsDzT83OpGmMZZ1Z07BAHun1aIjcfBrVO59DlZprH3lwFv7YICBYth+GYMm5
Xph/BgVObn4NMlBM0PFzx90nWn0eTQSaVcDulXOQoEY2RStdRwlPrAjk7qM7TWrQ
EExbwUwG2F5eJHRDcu+hdenFzTC/HqnZDTX9i0HwasKqzqQAKZQK8LEQE8ahCdq6
RUSxmetwlwZ7PElxzf5DJDN9LvRMmLyQd/j7QzMLb96dZzfVzGWOE4DmZRGL/Qy9
jumegNepA1HnPQpSXvnJMF0O1OBMaoTBsJM2CjAx662GOThrsX6BPpJHZTKDiDZS
DlExy0UoijF33Kaj3Pz0m+TRl93lWt+lZsMQ0vIUOm4AcTgWVDwdpEEcxUnwzwal
NzSCu8gmN+GZQelnZ5C3n5z/xgpo2UibNUdM8Yajn/Iny9/pSniRUn79VeQt6cwe
Jjjkmfu49HLbCd/zdsDYI4TfgIFzsSXsqZKjbZgaFo4lDHdmQPwf4izmfhrA+1uX
uc1i4V4lQTY7ad4khsXYfnuNzaLij6QrMj3N3pZ6g8TjLaIrLyaBdqZTf2l/tJD6
q/gRpYOY7jN2MZ0Kj5wmJgJz0dVZtmOdH1KiNSGlFsxOFiAZxPd/0kb4S7MevYxG
N5KNDcHQdFlLoOyO/WalsZcIzAJwiRO98Fix2ZqX5umLqm7sg9mYSTKuyDkG4POo
dEObUBUl+ljWyqJsG479EoS9kmw3+kRFFvgyFbPSQOhNPsc4PcTKaksd45RYfvUO
l4Ajdx+yUUcSg8t8FJB1cvTN3VZxDTXf1HPdqv1JNsNgOk5OyGJBhz/SNOi9xHhZ
a0CiJddnjJXTf6/SnvUHCNswLAy0+oBAxm1ZFtuuwLoEx3+vzqiZILGk0Ci5INBG
nTpLAjCyErS23tYKm/csqvoBphcvEz4pX7KgOi3OaAORKAb7+gBxfEBoSwoQKJjy
PBUXOSszK52D6S8WI8O3Xx6996Z1VQ5IIEec798xXr61v+Jz9l9fzJXWYx4grpi7
Ya6c2pvT5NkB7aKgexpi8ccSoJMGqeZ9mByGM9hsB9/vA2azxJZu3H0M4+xGwSLm
Sar/Lj86bg6zetRijMohczu9Ao6mYwk4sIQb1pYbvDTzh1myxKT2+CC6e6slR7PG
2AaFlzDow7/CrFEMAtXlGmu78t93BpVjlCixg5xmZIqJexfm7SCIAf7wHZZBO2Yq
OSGXMHxsDC3hIcLMHONRZs7ThKxuUBQFIYJtmbuQRIYLXDX+eiY1Edo0GyZU9Ago
IdBF9anb4lljXw77MjBLBEWYQf1go4GkPoQQmIBDlcZjl5dxVClYG1VXAkmP9Ryw
+uAnvRXnznETFm7qKOdGOPBpqjgB1K+HbUJN1w5u2fbBmKeZeP+Tyx5GGKJXh8qf
STidLVFxiVVXJl7Azo+tM3H/ukUsKM18G/zvcrTF8VkHoBPH1gR26WbFSNaCw/b/
C7AX2avKwzEhnFFKx6mUxt5MiVc0MjxqZoIQ/5ZX70Ko4jKnwpd/s5KfzDFqYfkY
8H1y0JVkbf0CM6JLuofPzXMq47NMwSTasP1UlMDFxsgZyTC13j+DprtvtmfNpyfh
nq57iqz+GIjJdrOh9f7V4MxnrMFSEv/8dGChEioLrv9Jw22oVxJBL3CkYmdDL2hO
fGAcVgG+/mUQV+CoK4YppFJPpgLjwqzp8tWtWLanx3aOl8m32LwDqhavh0PXwlMi
jrJmsMFzBYHHokn5hHo9w0mmhwVs44Vp7S4GoZVdrt/suxXVrdOADZ/x2/cgpC8V
L5O92aRI8KZnWEiArVVhiAkpZ9opXyYrrTapSjbRYBdfJg2h8E5JjZ7vgeM6yC1j
CUKO1QLEHZzNBV9raU/ILlCTGo0BZ7gISd1dn9or1rgREaxef/lNw/00zbNuuEvu
mQ1FHNyHy/UGVk5vle6mnLTXyv5diI13EPIuA2Qo3o6qbwuCy+GdTOt7Vf2dHcER
Byd7zVqeGI+t3mNB0zi4uDMIOEpIYrKL2obbPrM1ADlb+M5wy/i4+IGRSBSBGxSU
tKjk81B/+drhtSo8BzgXDANEFCz0IjRz6oZlzORIDiLid+fgPE66CTx3FWiUoG8U
sOhJ4OBzoHX3xM9NVmUDf3SKw8ZapWBbedNugBGY15E7jSFWQtFWcI95+zQcBnFd
5d0VoUuMeYEM/gXHeBIZAPHP4wRA2RE+fp0fwRe2bnY=
`pragma protect end_protected
