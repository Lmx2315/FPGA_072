// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:37:06 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
C51Ev5uZYjGrZd+gehL/QgcpKQrkwJv9u+iF/7s4Hd/a/5mFRyCHvQVlOPEiV0kw
IKrBMFc/ch5g7GslaPobHR10hlXDDFg00r8GH+mqg/GwkDcCCogZkCV/a1wcWzwN
XhVTfb2uYIkmgaMmXeZ7Ylm/flnErlQP42ZUVfZOmj0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2064)
qYt+l6ZGyDKyqlV9SnQBbcdji1MTg+nm07FZvQ27sLBBKBEo/uUdXQaZvDd4ZnqN
k4+O0iA+jNov1HoxqrO8wBzVOzLWEqlTrBHyNx78+5zlUApEa3q8PfKgWHQ34Kff
X6UYv88gYQ8NPnx1/Bs/pbCIqlkAYL8h3PM+skdJIDMs2hjXCuogREsLeBgNQdOw
WNs6k0RTFa9vJzBA9N8z4EbiEOKubGhv21/3VbUnZmFStVeSdw8Oy/gRZfgJjua6
PTFL5ZikJT8T+wFymcurXQLzcO7Cw2aTiT/bmj6MnD4FfkuoOzPapTh79uq2bRTD
fi8dAwOAd+o2r7MsOJ5PqiyzsrfpOyDah5Dr9+ay9MIJfneIkdpEfUf6n8I+XxeZ
t/tmQVKkNZKlvLyD5eUpIUF+81tVvC2pA9sD+zg3raXbXYpkjlvXgV3Wh0I5JnUz
8gQvK7mmBmqWe5FNk0lAiTF069bmke0OJNMawM/gtF04BPQETQVJ4s+vu+JlQXY/
6pGEG3/YXbV+PJaolJY2wvz/nSVSNsjALnjnnUN6x7Ik2S4y09R4buK9LnAYH1ea
yTQ1h9sfOdQ7SlsK7MI5xIA3eq5xx0GRUNr84bodbyZb07/a6uaqLiKa3+lh1RYf
NY6I1AmBJirD1bVIb2RsHO7cBJPQcqvh6TBfR/GbLuudDnFpb2ldwn5UX2p1GxxF
xGxo/YHVtr+n91KKtB19R5/dV2LFEf8Eol+7goVQvv/VK1tbKRvAxUpk0XWqeNU1
ULdXmkNg6H69TvL3GkzgAkwd5WggzeLiWfxMArmT51SufQD8jnopHlHnG3TKx8SE
x/tDGQfSS9hSUYPKXiWe0RR9T1vKSfl7VvmvjxEF1LGNgC49fqBRb3fJXluYXYgn
tPw5vrBGdz30DVA3OuDxYOBHuXTcQ9R+7sFxQWnIF4s1L4FR4wIc5w8Lux6VJ4ye
sOOQm5cpVh2avigS5LrPIBor6JAMJHmH+s7dRlhZV8+lfS8MdjUUErLgrS/on1in
9XLFQICFCjtff3mJSrzAE1jrBtBcsPPAJSYs4lOx6SJXqbisnp8QySKw1YJsgYd8
lyJe7c3Atr9tIBc19SsqqJyz5Ub3+6vbTalVlZF4SG/0ndoYahq+heFg7mSPuCEt
9NiC9sBUobHp1s/f0q9FXb2Nr69hrL+NdGrC9nPKIHYUtyDi0a3dCntSfg32FdHy
rDn6SzSZXg7Hje9hNhPgYNvGOiOIGDFvIpNz3Adj6lptyIQfUdCvBM4fHP7yRKI3
sLis+U44FUlDnG8frwwznLDEdXAiHSdoAfxcMwqqM5uAlwu7b2wlJS5r3qVJan1s
Temfy15Dkx/KzZQSWwtKm9nP5sduEYYbrbPvjwCvG3k0Y0mHsXxeKkhsIfXEuhC5
qEbZ5/JwN/0o3JXVAHzgy4wOS2V1Ktxkkfe5RAinMjcZLcpCb7F0T3CBe+OkA+B9
aqkZdC+JHVobY9AWtt2+G+iQPlyRTaDGbwPjFMzUiWNEgO6UM6W5/HGkW+Y5LDAZ
Xk0J0kMWZyfv9O/+n0JHD9t53hpIgkKCX+vBlmbV+ySwvHBnMHTUtNKh/MlhKFqt
Ot8zdPrfO8aEOSArVQJ9y+gjrF9UkLs/K1+8Ehg6gsQNz/qpJEDxZNgJOrN2QkP+
DK/tyrTjRfKIUHJcpq8FNYhTi5EQyV9AavFza9tWo1Y8fxYIp6G7Z+wkZQgwF+jb
67G6WHKgax86nB4BVHPWCdUl14GDZBAzrAXnTz9DBZfstxFFTv7NTpuIw3MCQEwf
VeERi4tBu4bMSkFUfrL0bdHUYj8WSMRRJYO3WnfjMBz7wd1U7Q22lzoQPqgYAYr/
K3cCDfGPLBs+x77wo93vospdKnCAzAqP5gC7JyI48OKU8FS8rnnVi2rH7Vln0JSL
0C8v40NE5zS+teZGBd62x4Eu1SuZ4EgHS9HGNH3QwG5hmsF7INJjjqZiazzsyyXN
bf7J/g4qISihMQrG0DO3K4/dneeSxMsP8MkJ8wXknNl/NnYs6vp+31rGbA+rCPP4
lJDfYCtvOl5KC9wuDirxqRKKiCJ4JTqbMO4o/NzuJ+HVLQQvVD9ypgLPP95gRtHK
HP6uaRbVqT37YCSxSTHM++k6hH38tJ6u0ny24Eo9UeMZzP6URvLcaTPw/uvNhype
8wItMoHXBf9WviAoiM5nl5MferIFgEsjxuIiXhlbc2NIdHtptSxNZkUJzHAXXfpx
5DMVBKKNYWP+f5N5lZxCp9afPAyTtDXSDsqDuZ9gU7FwlON787MLxcS7M6hlbcFe
OOJiK/hm6i/2cJcnJRG56NLER9AqBDxzIibCY6i8XvKEL7N7Az77s58qyOk55vz9
UwO2To1jbb6A8y8h9DjbqvT53oGKJTTQHbng+0sGeKoxb/iLqWZPswL1ozL7VdhX
g5cr0LH5x5hgJ81Xuwpp8UxHGfTx/cdDSgKWmBPnK3mUw8cwP0p8UuGsrGfYnjds
8RmdGaoWi7f/7fTMzTxITuHZnn9J5NJtm0TzZiL3JPWAe7HbDhli5WswTF5FrrB4
PDjq+Gz25I4klm2+DiZfZ40YFc5t7Oa4PwfyGbOb/TCbvRQtjnKsKjqo3TBw6xlj
PhKVTtxdDAPeXyx5RxrTPiOsahNQRBlv177RAH7UBZpUgPqiqfx/r0AdBKkd7hdV
oUMIMXOXFFBjOTysafvTn/btqkSIy2yJmdNQo3M2mOlBr72GXSvIoG/dHKT0WEGf
`pragma protect end_protected
