// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.0std
// ALTERA_TIMESTAMP:Wed Apr 26 13:33:38 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
dZO4zHjptmnQPibK91d9hIoUDW4RN8nm2JxOZ/2b6p691XJ+pOYdETZK4KQXW+TQ
2jMimdIERs/mwqg4l9AqMo5WHCY3urxF52pPQV0Oi9lFZg6h96WOJZ/+Ql/n6u2V
GXkCiM+MbLdMY6i4ipsOD8H0/veSqGtLaLAWzYr7aac=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 33696)
QggqPhVCWRFX90IAnXyUmi1/ae8M+vdqVu4W94hfTPWD8sbIVt3h/gmlrFCqfm50
sXPFcSFQQaTds6Xe+4jI/m7SLFIbKsvuZej4yQXdhVR/NSAtilrYmMZ9E/6WePsK
tDXo6WB3BM7GH3hSjmj0Wk4HujbCnng0ThAKdxQH58X/KvOJOizSfZTkReW/W/B7
gr5K8Sule3premvHwTq8GZ69VpAsaaUeegH2ZZnacLRKxjzK6K0qhAlOZHbSGHZW
jv6KW6HylbMkm4v/fN82NhLOpiYCF2YbehBORle4El4MQyY7xosBwbmYdoHD/3XJ
K6z7QSl3e2B7R10Q64eeXVhNQri1dHmzEYEogv4K3QjKpcO5WAyC2J462whU1uqK
0SrhXzDzA3EEwh1hWaUdO+mKzpJ1WGGSVav6hKQzuef5kptFOg35pDZzWMwLahUJ
nGI5q03b0K3I0yjeHpOIqzJKrCUg7oH8IoG3bKNZzyNIIBgS0GHI0aEdimG1w+gy
xIJRdL3XTW2FOY5Usj9bn6XvEjpIxm4EaJmVmAXMSRH7m2RyR8tfZ/Fc7Xeyei72
zRTwJ9xPlCgO/09c+41brGwV84z4ngpdACBCIYAw5ZJTXAOIi6k+MFejubdL1XPh
DmI6SgHxW0Yp8abTo5fe6V1ZcMx88lbEmFXgNk+hHbXZfpIEwrPAb9Zw84/ATXQK
0D24dASwfmfUc19IDkizV0cORNJzUn8hPOhEcH02dVZTMMTFk7NnTairiGGArkut
EHnU9Xd9/R4HK74uERKFSPogGZEjrmAFIepqiYYPSc+l74XAzg2zKiKhePxExWkU
2dW7pm4sOkcQBM+6YUA8m8NJZ0n1013JQwJLq0/EE0aYi2F6qk8uoH053+ckJNWn
3gw2NXSNEuJc0xtdKaAZk5at8CvqekBngGrvxN4swCqbJwYrt26V2HcXGXVWvl6e
p17v92ZtY/nsNjQsGIyMs4rzqNplmtgIREz1i0mZwSGbPCiUrxZxb9PmsjOnpBnx
Cus40x2cGsbu7d1X1TXhT2Hx9R+m0200osIkY+kXhSjKGa+hc2wCi0bRZ7rF70rB
/MIrI93iGYQNGVnYnHEIuZyTG3v0OOlAmfbjVLIdbNqyDYMq+bL15946Po4AlvYl
UB7opOAyufD8q7NTcL2aqxlig+EeA4jJHiRLgw9VD6QQKoM/6QJwevpH2sVw7LSZ
DEJpDYIsGEqmEqQkgi9d1WL1nHKdvcJwIsLwT/h1o44CqUC+G43T5ehIUKhpkDRo
FTqdmXdR7SISpQGC6jooslpeHjgrVhVaRitjJyMmTnifQuFhOUXM+8bq7j1EoJb5
DI7n957urfeE9wYHwJaMUw49JtkcbwtOCwzxA6GcmkZhh5xfosNf82L/cE9Z12DJ
iwpHkaVC/xajXlJDQA87ga/RQdZyUmOaKOKnn0/2MzfC4CQEPS2aRVw1HsFJZYYZ
pNXR3rwnsy9lVxPKifqYKhY6smNO+fNg9itoAIsLl3Ut3qcAwYns+CtFhAUj200e
VndtdT/Z2v3zQQEBUSHP60qPdvYHd54M1zvPgNUdy4lkU7OGGxBw/mLdKRGVUFuM
SwaOFJvsvIq9K4WGN3mpNwwxLriJ3vYgxVld0DoS9THO1BT+1HNIQ05XWFMFyf0l
4GiW2rknMScChIpXTqRbuZ/frw+JoqCybubfx/fY1ZpzRXGfllpYDozxPqG5x7iP
n1QsoECzraT1yevvUCC54rohQrgdssDBbm3O8uMj8pxM9e13UZslFc7VQ+7gfJz+
v8Odf2fIsiO9ieAPYEum9YCmrxZ0v07d6/U8Q/dlo81pfm7z6V4MkHaRPIwwo4al
AFlOoBHP9k+6bFU0ws+3zSVFY5MPoGhjOngRoLuk4kDLdfF6tRLWZt8bIgXxCvXX
vZqKdlBSHw7N/xwsLWQP8eVAyu+jM8D0msHSV4SKdJPWcJCwQQKuDlRdazlA0mwq
QK6KQNtCpF5gw+ufKSOzv6ew3kl3dqFKmbAZ+pxDVl10pV8SFAxvsoO50TpMD/56
2BJk/Sc/O5DvjJf+ABl3z75F+wxrYgH21WVFyzdZmJLVG665lx8pHapHQ15HytZo
s1nDZFrgMgHoT4HWohwewXbjGSdwVLq6Fi2/6/lBsyM4+LmHid+46YZgrzil+xaj
FSFW729R1e958sFDT9cwq8LLRjnQI6DsWkeNk7rgCMLYw4xQ+rdYn4JzPpknklzo
CWPovDyn3/a6PmsgFVmLLwWPpgiKaUPitkvcaA0VwArQg14KEmLxcdTarZdYkl/C
fQc9fUTO9BsZVE5g6wC3HEdHH+9z9AeT3AllsvBUd0HRrmjMxXOmqC0CjAsMpI0V
1vhy7k7LkVTZ2xivFXfcZlYjDo8IFyDbIdqq6NSzcFJrK/tLfoRCJDuLzociWHkI
EbFQN5T0oaI3TuHUGk03heCzZaq0hVD89OvjbTD2NkK5Cn7eibIpl032QjQFUG7o
8sGxHEDycHTios9ZkeZdr2eWNjpHix3FE4fEaHgUmi7ekPNSrbi2/DXSQ7Pw67qd
3jpCpFJUc4BeaYt3mE45Yf7dQIa5Uw8vl9kk9NFbInGDo6ezFgUKDq4OWcXf9/Zl
mheugrhnPYtNXd5HkgWLvspX8gZ4vIJtzVKXMnV1Sy2HTFLmJINBY8RMzrOE7kXG
gA0Bl9ZyCJiy0s0ca8YMC1EeOZi2NQdxefwBh5Pkt8nn/Vtbw/8ussqrKWflRNuz
0I2EikWKRhx0KQIeBCzeZh6N3cU7b9xE+D1EXSeDixJ62Gg21IEMIa2MtvE8fWKO
tITZpKrN+MBhz2DRo2WaQJ/B154rDBCI9iXF9fncHMQw5qwHuLGWxtxhXt36NkTP
a/B9+syif7Ya0tpciwz8AjHV4a4q893eDcW4GDRmPiM2t8TMmsZkr4ErIQHe1pUS
R3CCwPnLUiEYYd3CNzcwxM/zu0o/rdI8L2HIYgf7sduwYpKZIDhWFc8xkqgpO8nO
b35lWZy4v84yo5A/4OVyZ3DqLGGDlqhKEvRi3pY/GhbeOZZ+SkbQnn3N9K1x6nay
o2xySrS+Pv8CxuB/Sa9M8FqHcJFI8LsgMgvZJBpyAZfzFrGifbUHs5v/qiQyyuy+
xfIPSQRbSP/8jOmVfjyDBAIV3A/XNzPShofrKYJizpwypR9iPfk4/TcSi7bh6d6x
an2GGVIcb0ppr9QlO1v5CsVYDpl7APm2A/5WsSbQ80gJl5FIB2Pl1zL8Y2Qhmt3y
dvqIuzBVlsIVidgE2UZ3EYIdX6wZJhPvuNpHWxP9keby2Dxii1FgLiRwjjS9fEn7
OucoIY6Z2hRWj4tq0c372PcaEhUCBpGQQfZM+Imz3lhfZj5jPTKdk+5qU+Cq/mFP
M7qDXFeyHmbvvXmfF2BamV0/tAVan9MT+AHN0iwmBcZnldapnRCtaLaoq33DYdqL
DQabKSiSrypR08R0UOFhVmlcGDxBvH+01DMpXDG9SSV727bSCKT/9QdMAkGweVny
L6tUpnDyLz3iAB12T42XYg/PWg8t0rvcOHSV9uF1Lh5+cRfnnwLYj9yeWLIVgmaV
Z1DKjlU9ZjrFOfyYeZ7HFQv1Q/XrOsPaCOiei4st6Z35UgmHj7MC7zJgCLKOv9Ug
1y6yijKNwTc6y6fHdon4LbqTB62GW+KoKnwjV3kOTpcAtx/aKri4evmmuNxacatl
lM7vbHPzFjZiMMJxFZphahkUJnZPdxZa+1NC6X/XqkPhsvZn+7UYpz1O87DBcQ2k
h79cCDX/zISpwE3Qq9eSdwtLk3Ith0XU2jO+jZVFCoMMcV5rsGr3nDXtiTYiXwBt
Lm2hZuzzvjyjvyYZMvnilcCB9EOdtL7EQyjz6O3SIHRluTlsqia3ufrddxbIHU/C
0fdLMi1RXRpByNoG1XHZFfb4byQksTSb5KkAvfmK2BtjmqmyWNrqn1/iz05YbnWH
GNfebRHZ1GDR3dgNjf5kOPhktscEk+mzYac1OIQ2l+R8ok7J5JfzPcoVI0ccahea
+GIrdOOrrdeN7jlwKkI0UsqYzD0k7cP3voO1gwHUBWjqdO5k3+U1tvhJqnu8UUZk
p/9x2MP/yyY/QaxLsQJ2Wbfx5iN6punPGpA/FNJI27owLcQJp7JCWmWevwdIMCHL
qRknkVF3I2nMMdx6W5yuC/O6oQruhrD65z8+98B7EuereM550/snlAbBUz9xghoF
/GGf/IbcTIY97LBK5lxR/+1x4FIcgRLeK+F/bpJgxcyZNc35QmvjQb+yqTjoee/L
hr0bfScYHjvxBFCwVqVpMk1NE0oDJiQaHNUDWJxQEQ27y5oGHHidCJNm2E6+Fpoe
lqfd7oBQFrbpilomok6IXqMl6T5raU57Gvaf+44nE6leI+C9g+L8pWbgNj47YgLJ
XaEFl9mMqQOI6jzFJx/CYQTWcmvskI/FIbiiyhY0IYMTJtzsAIP4EmZCayDUToG0
2OhxSLVDnFkGcivEzj2w2D6BOHZQqGuH0lG9aABH2dgovcwkS1At96x2XXbAoyjG
/HIX7n4HPZnYbnQd7PBeXImfkJ6i9EUvJ6AeX0dBGyT6AtiKKRgXX1swVsou6p+/
y7vj5Mk8Gozz+2cGcVULq9YsbQXwVRwarz14nbivcZOH6VvoS5llf5wlX2lIfMJo
SglpAyxPsC73KX3VWExr4LYmg/uZ8ZHvWkELJb1JTrGvOevSGHqjMZbg+piOG2uy
MD7jPP420NPxUIyTqPcWcpA31q44sVDe8wN5j4R9Mztge95Xn4SQkDjb8GVauo68
m3/Tq0bbQIaRm0Nv6vvp+ONGTLPqftLk1iHyvSp1dQH6WAW26F4RIimsS8VSiGKo
bfpPQ1KsvtUXyg5kKItxIff+NvVcMVhtmL7dl/keXufh4UuVFeYMMmCk+mfjwKAV
4Q8oxcHQpRf1v0ESC4bB5O8JLeT/a52NmdoqtiYT05sX7mMQGDtPA/8N45guronw
YP+howAAjfdCCWGyqXl528sxIkD0QsCwmUPBieU7WNaDbaRYYQqqlhDPuTimJ6mQ
2trEblIYCoIXrLU02Ptbnfszy0ST8zJ59qP20BWWb751nNBvryO8EjHUsXZdpQ/q
ZiuxZLwKOfQYn+w8TfCX0hBDZACILew2lamFSmGjTvKI++pvdAy2Fw6lA59COq1p
vm5IVdvhD7jMIgzigic052J1RYP0UOVzMkTo5MRH6HElSyVr9bob+nLS5d2PO9bU
rWGmlTXOA+MZ0lRxkT8MdOs4KLEQyln9wgLqmaL87vyISeErP7VPkOB6g4T6lcFK
mqh1fkfuvxAUGjxYfDScBP19f2REAs1aCoGRXkYWWu6atewB8f6CaTaio0HCqs/K
4hxQTFDQHKhJOG1i7GMPMPplB7L/FFmlEV5DgUQOLB3w1IuHvBF5eSHV2fLJPMap
c3sDdT3E/l2JL1RlFehNkfx36uJ6dkpkdFAojeMzOYYzEBcy2WubAxaBMy/dDU+2
FKmSvz6YyVUeFHOlnBYe52ejTS+lU75DFZ96R8XA6QcgLRMJ517V54dcoGMg3V1e
yNYmzLCYphNetIUG7yqP/LMWfJIpZBbAseEgCqzZQ9ICxshKp0WurakIv0f22yWL
l5LYvPdgjKZ3YtIH/Wu9MDCOLbB2Q/Z1HaQ2QRZknxtp/CqgKyDjIOQQcqwm3lFE
YESLWBBKlQY0Y086rt7mW6zVqmllg1xgdXrYkcmq+37am8wusrd0OUQXEk7IcQ76
Un2XPXZeTBTUyc8v7lfLg6oK44AZFzR55C3WiDc4Uefq31bYn/d0vd89xvsomq+6
QFc+D9ii4iLrF9w848Pr9dlDqh2THS7/PhHc0Pk11UzYPlS2yAval05X9frtagcW
z9tjYRlseh9QjcXhiX4sShx7UTaD8trvHG7Wp9cb+RpojD6tTDGr/4d4KBUfBDmi
K8GQk2d4Szik6T5lYMSw+0c/71FtFEZg9V+OjzK5DAN6F5tQyB2W7F4EN4DOSSeF
5jB8JiMU4SCtCShktpxXp0dhaCH5WvKAWHzn5iyGQCnmeRjLb+F3K7shM52Uqrf9
MVmi2qU7OuBFR4VL18rp5g5jYX3SZl+CmnGzmDZxfrj5qG6208tLdOIQNd6BeywF
M1sJgEFrOU8dQMC6Ftm58wWBGsYG0HdFx1HTActfbC1pXnOtuiqJjpdtNG/n1H9X
Vy2xNqxRnCBVYWQO71U5MLbDeDfws80ntI+nhxbmZ5LtM/JsGm1kmJm1k6ep7Mqn
scmzgJwBZ7972Ei8lEyl1y+jnaRmGNZ+YGkw5Fs2ZbFdeTdgJryc5FecurCxh45k
090nXuGPFKpAa/Eu2wa/C6mHO1MHN/HiH6IjYiZYKGBfRd+iLdJzEOWKoklEqkva
n9NeeQOH0wmK3dd1WgCHCXF6hNBKBckqh7wlvG5aoojgS/1uJo2woTDXPcMPYc1G
qEIcGNPvpfMg/METVrTASx1VFIZ9FLVwlJOSCg4fsNPa7Nl3IMX82dV4yePA5MEC
LfjHUWaNlM5ohoLIA3lyTak3cBxDtoNlAv4ZezsJg9cd0u9FdtsLd6R5fkqLqAYq
ibnTfOSPpA9JtshiZqxkyeQu2AlNd8o9R7pQaPUtnyXHaW3H2WAXil8wZ8QKeuwp
OjjSCCeMWgMBS2nbUiq2V0f51S2Wc8/Tq17CyLzrvDJCyLpOXh5jE/NmG1TRw93i
W/vCQsP+ku0MyvjKNKoMYhrfpmDmunaZWFgqB0598JHz3o5DI9jtW64bXcDu7tqr
yY6RCIKLObtuG/PAdS/vqDC5ggx6f4Ts4mihTJ/8PVCF0roOZvWk7TF2m0HOzdDV
KlYqOItsj31ybJRj8E/KUTDyxL+DeEAYtGBFwTZQ5U+8wDArnhOP3wJhhVJHHCYI
ZEBseTHpdrvNNaV+x3fUQfXLLLWC06Fu0AnxXyZjPq+lVpUWRIWqN1S0XUEayeIO
J51BSxil4kdtHFA+OIbnvs6bxw0GffLfd8AX9pGYO+0JR9sf5iZ9pYaqtN7DadgD
dNl91nkhB9gaITD+1AV34UBbR3DweD8d3PclmsrODI83qaucxpOGFC98KmFLQ8qK
LdsTrMGC5t9eQ34aqI1HpMnJf21cqQchpaxkuY3jBGEqt5ZfG9dolXbshadlZRwN
LLqQytYAn0shjtkeG56bd/x6F/xk/5a7tbtdP5llrubM1b94jws7xAk7WHx9lPT+
gledY3zC8K0Uc577MtfGWNvo+Oh9E2Hd45KiMJ4bfrHqE8ZPYjGHBn6Q2IHiej7z
+vQJCbUdSnzcOEMyF0EcHLwZ85Ef9OgCSBSvbNTf3+wOAv7gpD747uRAKNT5iXf6
b6RMLiFO0aKcPPGgF8oAnPoHgw9tL+ORkVNq27YcX4PV1TpyrrNd3u0eXohLxrFj
XTgtAlN8juCUCCGfwpSQMzV90JioRmO58CKmwiE2EGG9WA614jnM1OAO0N+uCiY4
PNMu3kBixf+u84ICjHyDG58Pm/u3KzchWblUOgP11PQZ9ydWBRzKeW+JeQRYxmBn
OpA5qQIli2HmaPEyP8Lp2+MLe89trnH6n3fkku9/ZEw1brBIanNFej9DPBszI6uA
l85VUxYJxBSZ4hoG4DbNJQgHd47yB3BrU+jpPz0WOiUlI0LKz+7hvXkYJD7ST7mm
ViDTzUxkfHnzzxp6ChKyAs/DjRM2Otj01GgusMQUa+UTtX2a+wijAW6G+MkbR2Pb
uTOQFT6G5y1PUqn84CAlP7mfV+6dkvECCCw9aChrSKfepX+JBx+qSvpqni9NK1Uu
J+767pE2GCpm/24VXtslD0NJ3q/CdeT8VM8vIKMz54t6GFQoJhWkTLtds6dbzTHm
hErNBiMcaYhn7JUdEbR05itsCEArhTCb1jsH8DQBfM18pJ+AqbrzqvMrxG57XwPU
BK5kDyUM9F75Jffc/yXtMpvIXxUiZhC+FEwzCnhcUPTJ8IueM9fp84/KyFcUuSVW
HUbZyR9LIqVXtCJZ+Ai+Mav/fO2gV8gZIK/bNAAHcBKzQrsP9do1Yvf6YXP+oNCz
Q4Uh2QyIgcobZX+WsGshfKXZuNi2Y05OCs5m0awXTavDzsbs+/zfDDnOzNYC9Nzz
LjsiQdl8vt2WMPQJT5uCdLEthbpkuP9B/hu+l6EFJMdckQjb368fMz9CMcIr922W
O0dNut3849Y+YEnpCfTrlxfWdYZH2NTGUeQB7Qhuu+96F4BNEmbNp5PkV0/VQL+j
Ej0mvTfIMk25m7VJuKKG1PfUMDyv28CXa2MmDfJ48+0ggBFAAc4l/m7SfIdjDlhf
P1G2R+bbQ2d4DbggXGYe8D1Gt1rB1po/gWE9MJxNt5PEtHtoD7yu5LhB7LgCr/gd
3bki52tTwcHlSsNNpkEJefbX7jEoZohTVWTgfMiebUmpmhvYI4l+qXL+XKPrtUfi
o9wwYqzxBQnRDMVz2Ng0Sq3bG4U5IS/CoRLWR5vM8XX1NkQdiLZ8bav6ALhdRA5E
7cIPtkam0BfM549NRv6Wb+TfWgG7s8v1mijiPvKYnY1vPQfOmpjD5egzrvBWSjRt
vEsS6DdliD60svLhd4yjCE0lhLrXwyj2ULM2rBq2T7PzFlPuZe84kWwhKrq4cmRo
eDbu6cmNSBYn9400fR0JEYACoYJFQ1Pz17Ovjbr+DDM0JCJpPQcWvilncYWeyoqz
Lspe+uokmnKOPO7Oc2mMC71MLNwnBNQG/2TBdWkeIU8yaFR/xo8hrhm3wZDcU+Tk
U5m35ScirN19CWPStIg2UJrJbOtnLSr7DX50RkmaGmZRXygFslue8h1q6KW+QOBm
YnU+w68v9oWSLXfelNmuaNM6KTZhQVeDNH0COPPEkK9oknSMNIwCjz5KoTH4eDvf
kOD2mpTfvZiZbKDhtdLYe8xYpbQto9UUR25+HcTvNK/P40O5/EPd96zFAgJ7XOdV
RqshUDyz2tAKxH7CAnjEvDKfC2NjX9lBmu23xDW6qeGlAPAbi8OTky1TNkHcQEEK
J/1ngC6LnnJ8/pjdKYgGg2AuWzr/C3UpfTZUbPoFeVSzR94O2l5xlLmRB81f3VH3
6eJJ/WTYg/4v4+h0Sja9y/PrrObEhL7gH7weE+p3R9tA8AZLB8vjU8a9CMtY5KIe
dSkCvSOHKOc628/Dmk70gkMx37s0w5fj0o+/GFvWoSfp2/CTgAnMkA8TChKmkdku
+QUFguKUEJ+bnfft04m0/KoQwtdOJ679GYqDPZLodj6nVVhzP1AD6ybOFA344mTQ
gq4Mab1QF8D0p+AEamuF8Q03NVYmhooYSMZmp8LPwbXIVujumSwB6SXeFLk/2JS7
9n/Emc/1m8pyfSfcIutvKTka8HyPPfuQxOz7PjkL/xq1aQcvO+DGMnJxXRo0a+AN
aDaDib86Qhal1w6N99chGfydlJxdkrJJV7YkRoZEtMkpFiDDhp9sU4zSQB1Z/T0M
Igb5h+FdIWbOABQvk5VfdR7IOzUKqXobUrt+aqgf/phXoqmFe1v+j6ghmUWH4F18
AXvL8BOqZ1+TAXIJ259HtctCzhyxadPCFNQqTFsUDGZR7nw6XVKRX7SOPltsTy7C
Mw9mfNkVerAEaQxYcZBQB1IFa5SZDV6kcyml//zbDv8Npey4+kWk6J96vvfywVn9
9yWHKygWKibAomA49sQ7zdiX3jRxcWcTroahh8swAOIlNLsR/R6YayeCHT6N0cPN
RV6Efse/2uzJh13/y/GLpBgbL2+iCaR7eQaDvcAnOGOe/sIzdhGbd4PrhjEsic1t
4JituxPut8I/k3mmG/DstF6VcEdbF9Cyv/26O5RVgrfSbsO3VZxoAbDO1Hqc5hRH
i4DrvJp94EUUmDpHp+4iBoySqNJwH1JzcvgIJlsGYk+IDzou0dpXj48iUn9nW9ZQ
6781R4dEskJiP/fIOH+9Zn9NAOEMEVSa0uiSb0S/DwMNeqiJs6SJPugby/FdRuGP
hCSO7GW7hgcGZw4+2Uw1ObwegLHDrbuRkIJF1KRyjc9XWUFKjniJrUXf/x96ko41
on5RJa8tO6Epz145VKQVxLhwQnRFZ5iDLam/I7qubmQSf/uAMKKodNkqLLC66Sol
qalJFn1+XIuTaUNjmSNL1A7Hmi0P7B10e51RF9PjhEHSP/loGlCm8j6ZV0fJH17c
KeP8avGDPynwY+mqQzA0ybP49NzJOGflUuEBUEPRCHhKlo0AnhGeAo6vUuG5pjS8
cpADj04z9KyO3xSnlzd/FQzKcDEiGp+/Tv918Dws0S/ii5Kt+pYeyVVtSby4Q8mi
SonchgivfGa1b+MxNGUui2nuMTUaKy977Z2ZvjJKl1dOBrcuF5d26hbGu7QsM8Zq
5OsGjdYMYOgD6GPVrIxyhgkEH6HQo3IsENwMaA7KgbrKRpYuai9evXHMTYjIyJPl
dAFjSZyP8sPqXyJzO5li1vSZ5g+jwKg6GLDj6PXfUKiPiJFPgoJhDhrXoSnDh9nc
9xAkEGoSqRYkcRBmDfUEPcRxNhvLNazCZPbqZth3dnHPibrzfM8nGPJq47k0n93Z
IxyGsi5Qz6DOJgVROBlruUu+OuNXawAwBjVn3eNt0YZn7ZFYTwaR4ysKwj8gxqfx
HvhSJgqh12VyXT8XITT6tzjOQhmQkgHm/f0WCdEmiMRt2635PphwsaV0N1YAt0NT
Kt2QCcIANXZCipKE/ObIPYB7oOssyBUXVcvCbesckm/EuWmQ3UlJqxYeBgaWiNUg
AMZ9kDQT+uHL0TNqBln2TlaFRtkvQ8Dnpes9xg4+py7V/S5kB9seKz469cEQ7HeG
/AX0W3qOaEJtcOKz547jLDfBVCYwGGxfK9ZxitMaUG3ZYqfgtU7cbwra52wXvl25
vl7GzqBbZp3c6CrzlYjSC230hyDRtboRiy/SoEwC2ZKWcPSUoOjrYdbMVLvlZVeQ
cqWkl5xFdkXU3mENlPApSufy/PlEe5jKHavWSsp5d+TlIxNh+Dv5fJ2eH8Phfh8T
dI3xJz540vfVaEFnQxC9iviFcP1kOrsbxKpntlBKMlJui2phdpVmzrqWvK4pcCQd
JVUe6dSR+7+p0gg0J2qYRRhNoQurBaGw6tE5fCB6Pgd6r5fEOBdkxSBvtHf+6DOB
/W3mA/OCZni4iKgrXiF6+geQlGHo5zPY87Iz0DQ86wjfJGHpE++902JkvlFXwwlP
87qEOatAO7qw7DjC8FvsgQk2nPg2tSnUhOD1dHrqtyECkcpVwXY5eyTTAp/iMXCY
tXU3oCMf7jMPIhlYS4ptNebZn2B+rFuyUFSPDjCLQhuT4AH0zsjk6oPi56FHGzx9
h2KAt0LpG4m14QQW8EMGHsS1+rhSOJ/EKf7aKCkhoVh3YcGTyF+90MqkWjsci+nP
wL1K4RdtAkwIoMjOUkA9U+R3asRIRQH7TA7xI7gqSMXjL+KzkSdOmPH+jhunXWGe
bkaoFgpCfh2XDKCfkkhkZt25EJJkJ57GRS4NwtGck6DcNnix+y1ZWf1kUW/f9gX9
wT4Hd+RFzp18M8t//0hiJepX9Rjjb++lpq9OsBB+pqIlZUpR/+yjSX52/swib2k8
nflqxUh7AZsQsrn7bk9hSIfp0hl6K1xPnWwTGRQguhKNbzcpQ+nqDEcwuJmOqXeM
MtPpZu6ZICQ76WokJ/LM88R+HiV6Y6U5zEonQOUUYY0/B3vubuqG5hTqZLK26nQC
P9l6cwZMEAlZqpHMwXTafdb25Zrdsi/sdQf5vA3hcTX5+I7OztUd5XWTRgRyYWZR
SsvzuTtylH+o8ZwZS7+ZSxThKt9dqGc4xJPV8j81h8W75vjYpUZn42AntQYGOY9Y
tSZBKMyNogYY8F1ZarWQ+bHHrUo8HNm32TkuIO6r1uPox1xhh9KxADk9XVVkTIVh
NcnfEihKNiVIa+1AauymC+iYStTf7EWK4FNwdGKZrlXT/rFwTqCudp8F7xOmUxh6
Yh+DdpdUWidFDFupWmGmL+Hkwu4maY9RI1sFZTLBZK0+6Gxat8dnocXTsKo+kAlh
0tpOYOz/Mt8kYYAhU6VHXydWnIgTFa1VV3oemXaR+59tE5jioXuPRCixKo+AqBey
B2r2lFTddM6scFonVm7LEA8jIsWtXE4CvozQ//TDKSdv8uJmQmtiQRaZqkHDEht5
wgSTnzD76180BbYZv1aoAFn9VkoJQXTu/4ebODpvfu9gtX4LoV4aCqF2/fxVNZEY
Pne2ibnvWzmKBlMIIDOsU+vc9dd5MJr3AW1bwtZzada98TMwidLCirMW3gRstcTh
Ad3d5qfaVoBKCMSYEwmLXZGZfYxphcpjtUTrAc/II9mYK8V/fGzBUQ7mlpOLtZdh
IwesAt9RbaHRQdxfn+zt4ptBxpVo0uOzNkv3osXS3bayiT7u8+GVhVUuRnsa0qzu
57xcJURa1l9K1frfWNurAARGrsLIR5cShCCFBHZHu9NzLN816uFd0ctTrUDrvboG
9qjK/sSK7pqeN2hSFxZ3hj1pyp5ASHp2gByAVAl5aE4eDipcyukjQWudS9Vv2SVu
VSMORzK6JObbj/f5CIUm5m2M/JJZy7UmjDA78cCxxffLyrj2Fclylue/hg0bfMpn
SEqnRYY4242khLEzb5quEm49H+XZCSvyGqHDSdKqhNozKEe2OuFsNVy0UbW8+tLc
6thQ+cSVEpokhBN8Yx5qN+x9B+PzUOAbF1FLmCVIwu8+jpm20NsL/nlNcoIlsav/
x+QIxsryVuhu0X2O6QYHv1Te1jy0rrbVG38l3n70gYq3e9i6WPswdb1WmwlqeWJs
CPjCp3m65WoidujC1HfcPWTcZY2hA1WSGMVrIq1G/MBp0LEgI5t7ql4eeaQQjW4V
WGe0XC5SNOWROQAayCEKfdsuDFejxoiz5kaT2f8oaXY1beqYnydFSz8qKoQ8QHML
YFzglN76iiYfQNbbAPRuSAlLXRt/k1IAOV8IVpkDjj07IbZr/ly3tA+9VepN128v
vo09B8i5LSJYds7KT6zY5vys9mc/j4A1pHeMEc6gVtwO+G44h9o4zVg2hVGVEilY
YajP3XwXq98WzZdVTN25ZRHM9XZ5uTtchTxh3XtRNAzvvzFj5fK+GI+5c+dnXzOl
5tLUBizZvOh9D+Ar6YPcoq2myTOejxQk2Eg166YMrWqptRoNW7Fwx26rBwoyNXYC
2xgEsdBdRzcTkEHbFCXsDRyrPokuzDSpJ5jZ0wCYI66ao86P+Z++h9vitoJANwiT
GCJQ9qzTpe0tD8DxlPvOh6dHM9e1CDyRg/H8PAtitZCK9FLsm0huG33AmIlujXj7
RNReNXLzv+2EsSlPepKXrpbvMYJc5tfhfn9et/oIUAVhMpgkV5uqHtmTmp5hjixS
79S41lcvNhxY2dH/CpuWlDWzetrOYryqtLlqF6eqfKaOqEvYD76WWr3Dz4pWvsLh
x2rk4+EwRDXCBLLWY5dIlybUKcSMBmuXRDYXg8zsatrHEUwz3dxp91orCda7P9XQ
0qjW9G98SfjynxlcxGnZrcXNj7f74DRfH6Jyt7TwwruXOSyDFd0h81JdEqpdYDUu
w3VuYr9sp7YsuTMijFhNAdgJWTcWLOpmRY+JGipu3nU/jP4s62YGvN/4U4kyp5D7
rCB7Nq2lpYGPqdt9GTzwVXxfQYCg4XxgWKicSY1L8EnaK/Z88HyOe4DSANc8Xd2W
1zxRpZ3OPlXB1cpJchBlR5fwYhAv/3vZYxp1kDH4pMxZadS+72rlOFveZUNcSPEx
d9A0NiGhEeooCh6oFxGLvVPTvTQm9C7vKVEhK2KKEqH1mZ+zmUZCIy+yuDli7poX
/Z7QPIp8yBt9wRzypkBN0HvqTNMrT4tput+wvN2G40ni1cBay88zNxrYQHlFgyzM
rxQDeWj9qtJ/W6LZHlQIsdFhrmBy77enPQWAT1iRxq1/wNjqgBx9Mx6dxFkZTOzE
gdtNVuzZo8bToEx8yQofpJcCJQx3sk3X2dQWxdCON48IwjXSQUy+CdGqBumPjhUp
CF95t9N5Yr5JZIgvGQlli1wdYCOWRBPTOCKeglQSw9hboQzLVI6ZPnFyQmLEkJck
8U9n+IYWBaiQfbWg7ODXQRGL6TzoJcCEUiztUZP4hlgudA2gPPppO1aid3eWb8LM
JPgrs6Nuh5YGl4lTtwG1hLYp53V52avwL7NfTsMEpaLPha1y9WmThU1ByBM7Sh/s
eALYLfbXifJQ45xLMREUdbhvmIR9vqiRyKqPto6HQ0Rwte+ioduVtwDPS5m+HXBs
Ev5uFMAHgmSUn8gjiNPNicUfVw69Gi6hLtdfool+81RCkIdRkiCbtLRyrKJZ0sI+
0ZgpOFBm7xeXb18Kwld8n2N8uWV/fWTFgA8K/xajYK0o5yNVfkTib4qDON+haMVo
CNy9WuCtY1BbFIQx9VC2bdqk18hvjzMwYdqnhtVSoRIF4pkOeDkAoPyI0YBVwTOc
iqflS0HtYWET0/ZiD1n2G2mOu+/hCieoQdxizZIfdXXgu8ZP3sbF8tLD/m6VW2aA
dvTqHP0J1cihKnvNYifunGif5iqzRRwGSBYWN25GZun4F9WOj0hAFNViMfBcgrVP
sqA5s91yJGB+RD7IvtrjulUg/wHOo76Xez8HpyA8DmszSoOgDhbuqC6kQ8u6v8dM
A1lg47g4/uV76vOkxx1jPUQswDqkh/gCy22XHbo8lf1MiRSS5uk8z39bfzUu317j
VUakS8zB3y6BiehstJvSqD7yj+RwME6uF2vkteJA1BngBiXLKIiZWcOI8g1jLnLq
JhCe/lkOCc6ENodknlpMeN+iUCNfA5TPvqbsRBbhx6cIvD/pp66VLIehusk7nd+v
oUbxHs/Rrwp28+OpvHrgVHhV6BhPZ7B9zHB3nl/3iuKFb79HjhrC4GRyky3HHg5p
i72U7UQ0INx1TppslOQTKzJwlRr1pWxRpKniqXcPm4O5lI8RNmeIbM1cI8VnRbwm
4y3yvCZqwv8Ea3qBFi5iGUde3xSCPZT3XjHj7FFjJv5Xni9nruU11AgBGXmGBIJP
cds+tmaEgsYU+tTSWuoGGpq0ii+ZehsUhOA8WP9RJWqedHftHILR69aVjV+bqs/4
ee56I/Txklssa9Quw8bX2aFw42lnhy9MqIkaGFrobGLYQ3WvvBFn4D67uTRCYA1f
MFkJrKlecn4lor+gKSa/D7nyS64tiQMfkFnFiztJajY+sLNAFd42J7528A4Mbdid
eQu+PISu2pye3HdfoL73L+sVh2hP3URtPZLQtgztRxA4eSJ4Tj7wF1c/89Diyulb
6ZfiDH5nNc+YDoOYOS+FNMcyC7aYslSpGe/6fFGcAHfDGbG8QHtWxOLZ75y3RbIx
lPBJu10/V264pAM2cLXzOrBbtL3EoHtI/T9LYeLbiMmLCLc/MT9BSCEHTtt/uEDU
b18s3/dL7X+mxPBtu2bdppPMUYVIOUwwR+Fuywh2DSOxB8leX1DBpaT57n44WehZ
8xGZrrXaBbmnk2AaTVVEeZE9qAOpxIAoWFvv+wI/gJIpHNUcWg7HTseEgmauRz2n
YVoJvLahij3cR8G1YXeJUgP+VPhbkdKF3Znx6iGxXddVS7MjL5xpAVGcz09vYTzG
6i/b73NLIX1dlTwrHL3U5kif0UtVhZULUIW+a+BKnRbjRgO0kspoMdk9SnptG1GU
h58DbTuHeo1E+W1motoHvDkoq/Wzq5kRwxL2sbqg6NnDmN4QA0vNtjuhGny+Fx0P
uqDmumcJm0r3+VotcCYvh8yhZTJomZF+OKmuqP+BmXOnlQ/+oaPi2ybiI92BCwjv
FtL1y1b1mbvXwkggP9pcQKiAaEracCS1rjovPA0zj0JyavtuW7SoS8+Lv+9IAkps
6m6fVctnD77I2rxeQEuK83fcuzo8yL20NDXTkauD9fh9DQpWEbfOiG8T9j7PlBn7
BZRP26E+vfJab0DafMpp7JzaQd47JtMRtF9zmf1ORGytJ1hgrko6bBNz6u8VwdV5
HJyzgFNUoCeH+BWwWqfEibv1ln5L4rn7RUugtqzEMUWs0vEtJjGpBIYXrnzTvIXL
nKjhlfJoZ2ZOD9zz5ekgEL8LJUPuvhSNVF92Cw6A1c8WRJzh2SwF0ZdbiL9YRPA1
E8lRJwPgRRNsAqnuggmoBRTnS9U0ciSqeWOvKWQ/x66iB/ahL+ZenrKMyKYjGjtD
A+uu6e/hHdkbFrkQLgFu81c6OkVhLN3MHHj3tjM0pQ7zWPi5Pl9lNwNvwXEsrUdh
pIpc9vFTRxpM/THexH4W2O6REtGHxpocV1IUGHeCz4YhRHQ5JA1ST58ioOPczH+I
ZN84SJR3LjXW/ZDhlf0zFeZU8RCRW0eF9rRoxINIIKgXJ97fDfMQlqqnsgBxhs70
rfVD5/5LKMalpxYaRfjtMD5vkWxjij7c54MArlnR9GnfjDVkUzt5yFvsJufSt3yh
IShVuVXolUU0kOHlt7cv6DMpS4WRT7uQhMRoxLAGb701++DMIvweW5zZ9uDL/lwz
XsaZn5rHLzJaifHy5EE0rjI0zgK3oyY4Y5MtlRKyWDZjQaxNYn1Fq4vThsHZ9I6j
aZV6vzWaEJHdjnylsnqphzCK4o1T3vzcJ7/YclmbBPODAGSQ+SuhQbokdAMdVqxK
uAJFYZVQCxg1zRtCPJczHCksM1upZqWIcKQYYq05R0SLmU3iluUarr9mSROTtikz
vU2RLbvZP2kcrBr2MX0kjRlJO53csarMcFs3tHybVAbF/fXu8BJLBVQ4VbZMO8IX
gEg3mKbMMMiEpgRpSYUYZDyjjjgkX4A8KIiNr5n5eOjLfPNX0+uzTEuB/8aLW4J1
KWoB5BH6WSsvpNoIwtcqwGnC7ChRV+PPUE2JKxOVFnc1AVCitG/K4iPM0Ee6Cf4L
SHDHGSE5ygooMv/kTrGC8hUuszdHe0DkT1qVq0FWszDNKxFv6EGE1LeYTpcU+PA4
JsmduGaA06+0hbH9Ew3Ky1jYJFEQLXIVNFVj9uqOEz7AVAWO4iaFx0k7hwgENNMW
UeUk9lRFHE+yjS4yXVF2gvPHfriugUJbulNoLL0Oy3r04c8HdSCKxqDt2gGXHTvX
eem3pu0fB0isRYQUj0DfFmZuEklVmu8IP3bhjrkoWYFGV19Cyv1mQ3xWgDyN8A7R
WxH29t/Ut4kunaW3jOiAKY57YNYYInZmaFRzV0nbGUTlWIlYPmyBwuXaRoYcmxSb
mxQmj4jHmm9N+LYXtv62XO0tX8oK6Xc8mcBWlWktYx8UliGUwLI22aFmFs+yW9PE
Ue91HwPjO/BEYifd4zWiG2axflT7fJoqn33sOPpkhmb3rjCszE/0G64o2Hi89yxK
ilAQ5Z3al2igdo2nlINpoylekQ4hoaprYkMB4PcaBtoOn2DQ5cAyYeqq9TBfGmy0
J9stBGTSNXkwnHOansliZR/9r8eeV3Tbu8r7ahFasdNtoeDn/YCf0jnVArrS3JeF
rDTSsOyYd1UZTChXuuksP7GPZamNIIQ1iC1GnKGqxLQmAN6pdkVP1bdG+eVU52uC
1lrV51IVvqU7VZboZOZqanKCVEE2mA3PoKL0Tl9WEG1nrrOxrvfZoFYn3it7U1+s
HmzZDSbER/mmq5QMaZGiwxGIXJoWqDWAkwYReMUKwvrkPtIm7ps0zCIbNsVoi9n6
v4yM9qYpUMwUiESrteWpvjd+98yGyX6qos9BAhMztbcMy85Wp1jzzOgIenuiZpdD
yNqfoCzuLTuugpAYu8AbWquOTkI4JpWuRd/O6/QzriTj2DOZ5pUST5zGGczyC86c
FFzgab7YNTH7DzbZbD0wt08RTtjgBtXg0T9lPHVlkpmH9MAwLu+0NQ8sDHgJT/sB
XTdWNfmfoMyXnp3SfNYOVKUm9q6VuiLwDlvYvwYWYPm7+bAVRRn1JKol94NezlHS
CA7eR4Tn2yRAsDVLEqlKZc+i0cxST1OmfLMLaTf4KPiSyIsFo3U2AUHQi2Wt86oK
4Acb12OJzAtXHEuLjDzr58bUJoNuhiWLDQy/c2BBfpYU/R+tTRHLzPyudJZZDnAR
SuhY0wwd8TeOE/35ErfQ9FDf7Yo9TFafASNiQN3rK6D1HYf+enarl3ktzb98VKtK
46HbjaOUEPkiXcW9FPqZcU4QHdLr/pkoPQFiIBp6oH/5bUXyMJl4zw1l166p58es
MUhnCBP7TW5Jh/TUU4IoSjtpupvGbzJdpuyr9Kq1MdoOQl29ngcB5KOSwdypLm5y
XjVntAJW8kPktx8aAsO1++vrcFqZYywOfuhounED2CUvrGui/bxBGonVXOu3tUWB
qJ2oLeUVhqqm6BV4XZ2hh/qJNViOnOy6yhUeQT5Q46VvlAXrNNVyxB4R/OKzsUEs
YVnwqR2tXKCEvyvAwLmkCcCTcBcOzWIfyCIGl6LI/o3GnPJSs1wtRFeWd9dWdOMn
EQEtxo+pYjyiwvQTxt7cJHsaBijEIrW+7Klf7G+VtruxtKqN6fGHMf6L9WhYZw+D
Yr/CumDpBlLAjRM7Wyuciz41g4AZCiTxrnrOzYG29jBASLQsbzzeUA8cu4thuVyx
9oAZT9RCYT4M/U1A+K8daNXGmQDvyt83PbYMHdiBfUyUyU6rqp3AdrnZWsdOXr/n
UbPbXbFRQ4GA1ZDq3KnmOO1xhgyCaa+RjNKMKEhvfpisfy6rNg54diu2NFXR4BB3
EllGzZfixHG7b7+lRggvNGU4JxuLBHETtnnL4SjKpSoK0wAMTrsIQshXknoDUaCQ
suIE4Ubh+KpkWhuvO6zjmQeJ8cjXOJgTbpAkMh9D0mwji2xHxRjtrBHjpEjmMzIQ
JpZdtsjO63LhA1IOdQ34Eid8wPyPA0IFXEavqnTbov1L/ivFxgVI/CB/6AVTbtia
ez7M+wd13YNanS3oPLfO+C+xLCb4QMi1ZxcLdci2pUZl9uYR2MmJP2S91SD9H4Eo
ogmqAz0rOYLK3ZQeXCa60wy5M6PNBrZbqk97gqcSZxHXEHVntCdlbZDqXi/gUIBj
QGNpk73tvB8jg3Z49yJOXpMHFJMl3xiFK3ZeGzf9BivAhmk4xp2BdV2FqkguRFcl
rXRjuE+zOPT/87sWqk5vfSKBIN/O8ufWgUm+4LKoQkD0zjtX8iB5SdJHSWgSBmp8
BJ/0dKK+x6L65T7We7SLJrDSF6Z0MzqMV39WCzsoSLYR4cEHw9AwCAwYhNWzftKW
ZqqWmTrDynRPVxWUUtyVzJ1u4QJTzjxtkMilIfoME0GZxGXAah3244T6OdIwpJLX
Pi10Ywl54rtSk1NVekfXknQweMfSUSChTV0CHjWoqCevahYM3GcgJUWTC+XzKU28
ziQ8j0wAwv+c95dWhmW8HwMQs0Xw52hg4R/76gAfpCKtaORWAX+pPO0YaNg5GHey
ENsZyAkFcbPKehqgJ4waIqmWrv6kVcxaJwOLQYo1E2WYWI0p0kehuAdh7moNj+2E
C+jyPVRilsGeNPfOAmF0KDpHWu4T0kJBX8Crx733GoYcSb3Xqu0dWLclvE9Jl0si
3dyrNR381nteceNBW/6riSiUGR7Dt3pBrF2kG+7H5pcAZg3n+GBpQ1cUOo673p5k
dkCVJgI/tNY42t+/Ad9nOEp2MnpjIiwmcE1Z316rdsCfO8PWE9Sa4KPQBQgxYveh
0Csk8n4NlVTNtJLr6IeGDZ0OSs6pIOkrDTKo852EzCtKP9C5eAA//i+FYLPlD6Jj
TMkvRb6KbOdHPrQDUREB9r2RqxNX1kpm8yV7uj3AkigSH+tNlQgO3lkJ0iSQ05u8
RSIHnu2WXmfHZ4dTuqsk+LMOGZkZ+UuBXl28gLIreAa/6uAhcUMLxtdzYQQe3prn
02e/hSInqNi28rCLRHr+CnnlyAM8oR7AYAqpQMbSLOzbixazlQHX6+N6guOBbXnp
MZmLgcv0UHAfCjRVqTXjFS65aG6HVe36vvL05qnPRjc/EPj8mwfYM6AYlxQLG+Qj
s+9ncXSAXLP2Ms9ai4DmRKYrSGlSv6StuK+LS/HmzET5pImya0DdEjpuhvHks6vm
/eDTVo9e1bKulyM8IjM5ttdjKWJZfgcMhOCpo81l7TMR3bOxeRkUddk+3rMu3xA8
RryYm2A7KFfnImR3Gnu+LHgWJnHGzFdS2CSVM+foj3+MIpyQ40dg8B1XjYr7NZC3
1S2cGBG5L1K4U4MHUf+zmNQ+9Wq1KN8VBcaTE2J72FEdVuFtMtrpJFTpxm5/QEMI
04rgQctf1pKrhntolOOAT8+UNgsfic60IkusQBG8uM3patc31Rzs3dJFp3mJdRZD
al1nrcAytTsbthw55qzwT3aqJt2fDP/Zssm42oi2RAEDqWu17AagDtTswm+CTZkj
01SiZovNNea1XbyyhwVEXwgUwggsJOgAQx4+YAUUyDRm0NKRNPdhej9DVHdNMKZj
B0fQERdZjQmkHJJ5bZv5Eoyeyt3YeK6D8f5XlmBJLcqJ8KAD8OYaf90sTJJ7eT0z
QsgeD6HXGKHmKPUThgeAuHpL5kNJ+5pJpPrbrAocJsoXqAD4B24NzUADP+KXg6Ao
MQK6drVAJEDCBY/MHvhtiJWbXjPDm3K3WgbnH6bzI0QAApOKL1jDRlEG+wNCFIhk
ANlHbHoQ3XyQD9V1kE3X3j0adrhWxREuOozWZniWlhuAAxieMuciegJSZOK7y68v
aTLfgevJv75gd/4arEIOn4sFFjDAiEAxstsyPJSJkdndWLv1HYATHnfMF2ePARqd
L5eJhj0eQj+IM64aa0vxrsW1xnYp62Ts+YfDKN2VnbFYpbWD3+88Z/4mUmkl1KNf
PzCZMQrh9rEY1SEs+8A093djs7RCRoehvP80wUTWnxwhElhfvcbsbqhBE3boVvhm
1SJaBif75AyDDKAOYzq/s3adOki5Li3WCJg2JWh7A0x4Kqzp7adf2KXCKN4doAhv
51b2w1fgBQW9d7CK2Kwoyy8gFH/x8XG+t6ayvW3qXqmuKRL32BkuzqiBkR3sNrXl
jXzqNq3dG5m+FwJYHuWLNuAyzPWerRnvyAEKhG8fahlGwzcoZpdXmjKqBpYUXBLP
KJUdhLvgh8cME36Wsut/yClvKQvWSs7ScGDgJqG1FH8hQ4vPtL3d373u3Q0WLjhO
YcehFKaLfuax8JcwBAFojkVjyXXmS60KFCSzP4g+Scb+7GGtnLzpdNUqunK57sOZ
+J1DZVdhZkgWDRlbGDf0PRb8kiohyfWNYHqb+IWrNIKYAWqJ+JtkrF2Xf23klJtP
vxVunQQ/VTOhLLdukUOXdAw6vj/Y4ND0yiEJf/KmTcVhYRR/A8+zGMjWeRIPkx8U
ZbiEvh7MMcEUW9OFhbPkQyCBH33HJwC72Q+Eq52/CFF8v6e+fJRnTxTYn/dz9g1j
FAnd7VfR2WjagUhKcAEqbXSNJP+fwTydUmsJYIAyp3btw+aIEkXOR3SarHC1iYfJ
c1zbsadTeN2X6UEuXiljWs0k50WOXnpR0/cH35Z7K5fuDNulwQ4k3sjfsXwiQX+1
W+hbZIZqRkbigNFVdAE24wXLmVbAQuSfOtljeO/jSmyfBvxGYKkZ7sOaAD5FqeTi
q+sFSGUEaI3zKJZGnUK1zmBI0HVNG9RKlo4+IapkDBYZcN3qWeSHB8yAqJFU5mzy
vmXPlrf+9So9dRfs26sxc4ktyt5TKhwv3W/hHinL/GiKxDXwgw0SEscH3C8QXa4N
eeobZl54YV/mks/2AcL804tph23Pr3/JtH3wQ9THoNzv3+h57c8Ph1Dy71SeNitZ
pUwjuTbGG1hs0SpBtOmbeJylN3r2R7k6PcLfHvUAekurAIZelzv8Y2YJZjnE2D9w
92E5+KgjEabIXlhagJ6BZmZ6CqEoHHHrpZ8WmFICnL9NKEjJXWVkWnDA9+elglMd
3A9cGifY6lueDffXXT74mPINWthq7I23v8E4kR2L2rfYz5oXHtpTkHLxPd0XoBCW
ybeVJlxpuK01cCNJSwq3I++tOU/e6BMxWhkgIFKoFAvIA06M1WUaXv8pUKKhIaTz
bUifgOodACxDaQRoKW5WinAeZi5J9pmo9nUG994Xrep2TkPFaYu/VK73xUaC02e7
6TXvZnxx6mA0v2tz8LzFvn3aHDR6OfikS5AwLPEIQaPXQWo0OufNh9V+tAroTgro
16h0W5SUM+BzFggJ9TFJ/5T+/SXO1RGTQ27bR2S34lPlM1ba/9KRPdD6Iav/yCkZ
AGvT46etkTRMA8Ihf80to+Dj9AHwtb9ByAhNNodABwZfqescibbehZRZeAEC7/Jr
i2vGZslx+X3JvxqI7mIp56rC3TtAah9DhocLJDbQOX8nCj8SxsX6bM3pG9uW42AJ
WVoyQUfjqyp4Z7fmtq3TYnYNejYHk4fCRvHVES+M9SY+lY6Qe9PzxCPIXojgBys3
++ABlcb6+G1aQumCRcPmBL3/wSQcxQcvV5w3Pq3lmVMGCENyABeQbCY0ojJIZgW+
kFdl8bWJ+MR/U8jSdz17MS0E6os9QxezqvbCi7e4o7d29hedceX53VEd7PJpwpAe
G6pDegFDD/ISl1pQJ4kmLVprOfIHg7C94ucjJEgUhn0IElZ+CTvp4/pJbkyjpTyc
StF25XKRH2c8PgxOS5+G+G5ZzGMvLGtDiMWbZ5T+0gyEVc1Zr5AtwcmXzrtydlVB
8ykyRfc156aaji7vSb6A+RUWEVbpe6mGnAdNwFHNXB+3yp4UH7OKh4USs/Lv7qAk
tV0hX5SHz35hwi1DiiKUp9R8Fh3FKfGKPyDSgvdkJ6xqiPpx3XGOIXNDISASnTZ0
UhTJODN8xXmElh4HxU12qpMCYCjnhiCo9+unQyV7rrLU01vMmLPWx+NGuyCHGbT8
1fn34snCm0ltIPAVZmU5xuj/RiMVtBx27uuHo4SNF61UuHBy6oGnq0d8CK8xtIxZ
QnHYE/osniOiosZFHOFae0WcnvTjlCnzhlQ4NIBsH+kthIj1WF4kr85QL0Edcykn
PCRgX+aSZpD1JpUs+IWlCrVKPB+vJ1wHZUeGoT36bnzqZkr3QHTupKVG41lf9XEF
yDYKDItOk9ZaGP+XphhOPudZlrJBGHTcLXs1Oik4xGaLI9Pfmohb0/na9KK03y6x
WUUGXTts2chX8nR8E+AqBqi2Ep/FzuxL+8DYspjebAqIOeeDYIQFRkbna1Vj6NhF
Fjyw+ffykWshK/cFlBeb2EpKCjbJ6v4vuNxgY36SPbAIrF7OKrIccqSTnc1kMHw6
KbrtFJGBTYz2Jj5OmQNMPaDSd80Tz1dN7ZXKNwiW8SmEVUJHtDuHrFTuoSyRP9Ih
Zqlc6DJwJBBPaZhTtQqSKcqiLxiLFeSNWfgCBk4wXwhi8hN/3a9yjqeuIycxCyl3
W9D9pqU/PIJlnPM9NriZjwfjddFMd/O3zXKwNxFDQ9yT5ckJL+7ccbb23FBp4Bov
3iuphyMFqhWEc6WDnrurO5nyLwt1bOGL/+zsKwba4/nZHdpG5TGMD6D8H2wNhTCJ
EmzeKm2pOrcrh8XshWB5nt1slcVEMDB5sabbM3MCg3irASNo2d02wsREcHndwUqv
4CviiKiv+0wLv619u/P1nkLUvByAS7J/d4KIqToLEl5QMl4ePamkNRF8yNPwDNBg
a4pkolaTH4ykoWvvu+FffiNpIcW95Za0vPmUgTnUEgahPDQv99nBlQImp6nOGSRm
Rg/Fyp0tO1n317Rj8sPwDJ+lYCDJXuZEU0h1ZTKZMhKy875UcpXsgDdKtanrLI3P
9g4Bj+BbSGBJA5nJ6eHYBX33HKRK0t/Gqvc+lxruwnjHAcuXNo6A5BAvnVzo3LK9
1i82TJtLiMOQbFrIWQkJH3UrmPu1WOGdp6Tn+clKL+WPIpfG8mBmIHL1XqEJCoed
5RbGya07c4KkIrVRU3aWiesM5gvd9448FlG+wdG/X/lQeO2R3tfGovIXZ+Rz3dus
dUiu5WO3dhVEb8E9URLcnT4wpcEEOJQsVH0PlVVRYKQcxsos/YRtwbbBypViXPn8
Lmt7t3XfclLcvA/+0RSL6ora8EMdDfZV2w6kkHnWd3o3kMTPP0Yj1yGmN9FL5/7w
LQJM99G1nKtU4mc0OlOAIb4szNX+vYU1wvm/q8Ju/MqjDb7mlXNY4X5KnrKaZQVU
dJ0icTWE+P4rBFYg44V3xw3Jn9KIPkxGb0zbUljx2/h+YqNBwBSqfRSzLiGdf3d+
pK6sczXIbURCv2td5gzk3wd97HKVL1DXVDGWlKPelFmMrt+YTrquP0utvFaAXilR
h/Y1rRn9ZgJokZXuxQkrJNIpjQi+ey1QhPpK6a4vbncCdXCoQRid/53TiR/HKAS3
4hdY8aMruNyDQKdiL9PRiI5+jhomaCRQjaK+4mxxg321UoSLwIQfTEzhPMS9Ah5K
tMRkb4lZMYiKqrlpx3DRbfNhvvN6mN8ioaKGR2Lxf8H4pM7qmpmWRl+0sNd4dttR
NYH/KvbNr8DtjUXCBOdvqyK/epRMa5fxXyF1F3jSHKIacNvGhGrU0CTrM93wQsnK
3ssq1ldPNcnoe6UVKTp2Bz8QenkHKQXON/JTbEbQ5Mq6FQGGfyG4sG9kF7NUuV6a
ftxjf3iKoqbITZat3Jdlwz3z3lK2e2dVhUkvGMz20CKxp5knzouD/4UZilXnaRfO
QUMrHW6ryyLb9KnhYtYaabeEDLfIGT0k6Cx6U8IJo2x8L2exuBU0zesCKpQtYiKm
Hr0y6rp/M+iQ+M9ygDy6kZuf6CnGoCFu53Bt7Hhj53H4iWigxGRNhm01HgWvsPij
WVcio9NAES7vH5/2ok9scfqURtH+Ork5XxRExdeH09KdK0wuUZwuc+/eRPEvYISO
8Uqt26cpWl6m8XfQt0rtvNtctWtUTIpGlwPr50YYubmH5X98Zy8ofrEAhyjmGoXz
Byn0CJaq471eixgSw84z2tqhZewfSaw5t+YarPFrliXcFyY3H/e1Thqiv6Rw31Y+
voSfCyuT5sAvnTwGvls1ZS1nPKotFtUR7qIba6eRXijWj7F5/R5CM6v1dk1WzTfa
Oz6ffpUWOOpqdn5cL6bsOwalTP5Ag4AIzTSH2jmqmPrB3lvK+5le8Z5IrLNTUrvl
5htbGfo7YfLcpXDY2AUhXiy+Grz0jqpyK2Wa2u/vql8KkOkB1bIo6AzeZc7DE6Oi
IPXg5yEEk3McJ0yfo0BET8EvB7DIhceg1BjSsMqTM4PgOTQYjnmgyQ1plxUJv3Pf
qIMxOZP4x692hCrKZMgaDLfVtgR8xTzNmIDczcq7BV7zXc+j3UB3HCqh4KhuQzcE
OaYoocN7QOPhunutbAOEsa/90WRrR0YNmbeMGDpWyX/Y/9B6WMwy7IwKmRC3hZqa
SfBchTwFwwyhZMHk+7hSDEk1eN2toX0p3QJ9LwKEKlshrO8ujgNE1ajxz38/S9u1
uV8suDaETPLzecZyNDxxl60Pi4Li6yVKw43Jg6cr8zleDE/XaXZFkLcmj/R+jHkj
v45K6rAEsGGoiCudwNA8zotVeEffyDR5XplYw2p33wgP1DnoKzmyRMJxY8lCv5hg
4UsMA+zm1eLiYl5EPRATstvGNguCDsCSK1lRXT8n/Bfqs6WuzK4sBFyqiEgmg3Ji
xDWWbmdToa199wEbxyWr4UcDJnwHt+wsaSn5oTpmLzDIcwsU24jlEh+BO0BeTYZN
wn22UEqEBJvSESwjWEmPsbfCbKON9onWxCFbmcLSDMxgjWt9wNYeanKPRSCjw/p9
DofvZ7/ML0gstQcHUxrP71nGPGLzz3wN8phPf0TiBQpzwlbNJxzGC87OlBdKTp65
Zvm7EGcdOyMGwYgq85fUac4+2rNHcLSgGnBGPH+pHTZdwU9hruMbaJ8j/j2msdQY
mswmiHlsaUkWf/zJ2sh5gCy3rQNf1YRUPY7aA6e2wAy77oe5c+3+jHel8PnjcjLd
8APkRj/LM83Sk0X1aq4a+AtW1J4rdSjlMQQx/imuoU13H8ohKJMl04V74C8zg4ib
ycKtaAGV8iApStPTOwP2+JM5lCht5RoZrDrKFbKMGDWy/2qCJppbmGUAuYMNnYs5
zyKlv35Vjm5w9wJKjDGXyjMIT8xBlT5mqO+d4CE2x3AGeqiFIxpnqzPH1kNk8rjd
gG6VcF4gOpELv8CSVEvbM+GiPY/2Y1/1UYFT6eBRUdsOsUGTtd0145Pv3ycsxSWF
ZitDc3F7+P7ln+RY2cBgiIZ7aDiRrUY1XYuoDZeHYqULbuykgo3QOinMnJopPuGd
xWE605ZIUZUXLra+MjMwk7X+zD2S18w8472GGyslUDkx/thRkGiRL9ic5ipdm/Ij
f8XPp42uCuAaS++j9kLGcCdyfbAdYy2LZV3U8716fS5F2xjCuvGIcDqq3+E1jIk/
YHsS4O2AG/6tXGBHGfpTLqMiI2MNkwkXh30SpIaC94xfthtATwk/CSraZNBHvo+S
AsS2i37wZTGqXqYktoaVsh3CnL2Kp2FpWWaUopIisDX3Vjsi+iY3aQvHgg6WIw7f
vbBO9+HeHDRmB7AUtlc89EoAnNUlqa4T25ybUYWr7L93H3+b6VHCsGqJMKkMXlwI
sJGw/x0A5ttEltFeXrXGHjKnn2Hj/OBxZyO+mapHXQegscS+zce99f4GOVBCDbTL
mocVO4hcRrsNQCu7Y+Mm31ynawUI0hTjQ5XaQ//RYaUc94rvwKBH4HReu897ZKgh
quhgj2VYv0vEf55TY2Au9iO0rFzQ64gKTooVLnZ/esCA1k39KQvq3mUDa/k+9YnD
sqUmi9DdxWHsqcYZPw5KUn5JQngwYPIfT0wficWWCgN4KKz3tuu0Ff2JzIaSJRUM
TOqAWDOBO2IUhE0lg03Pxk3UaQcsUiu8rdCzRnAb97m057aK7skth75EOMGgoJET
oLy42tp3J8hteNW2KX3aI/q2X+reKLpGJSMVtzT0ehHGPKxweKZwGl1pcIwTgv3o
twN51/0wSS4nFqmle7D/ZqO8nR2bUjZZriirLWT9EA5AwbAW8obKuejjKeFAwt43
8wqGL+2DHfteTnqEHaMQ9VSnMjGoAF4bhOMJH0xwWSyTvWwzrIcAYZpJcHb1p9E5
kCorJh8KZisN9XeALHVd4fFJ1ybRjA7lkGPdd5jLxdyCVSLUGNqFypc892tuKzQ0
R3ycTpGovM+RhQjXXd9gnP9XDxA7ljVYbCdGibPG9bYqWo15TA04nt+6L5iHXbB/
0IqX76/vyL/OX+FbyU2CPKXdh9wQi2D2o/8Dneoj3QEU4+V89aPOcf0ogwgAtc9q
0eEzmzdlPNDRjCKyAJ02rg00QGko8di5XQZiooNBUZRbzXjpwu3MwU4imx1XAmX/
kL4NZwUKzcFXbThUPxSfbv8vqdJzOnzbCpvQWMHAHAqfKSAUv8sZ+sRiYLP774xe
gE9J5fp3BJf6uAwNpjWgBJJHn90OEsp9IAGFSQvXOsuyCqLjLrCRoKFINcoV9hCY
hniJj2kK7JkEZPDDefihZ0WeLjQHnCHs7x7cI8qHxiPdqZusuYB2PRQQ3ewGeCaU
PhIygoSunubgZWv14pqH8BNiWGYxbLaWKKh6mVkBY0osZX/Cmv6WJS4XFu6nHcFk
bmJx/5tdlCLOOia/kvHR0NNIoCBERZLQQxOYRzwwvpn8IVyVHeipj9N8EcPK4fmH
zs9A9Bh5ArpQo6Mllf1Z9EgfXl4Bgzww73jaLyAv/r2rg+nqB4tpSt7tyEpX+XDx
+VEvZmeae01fSevkrjFxDBTSmhIx9JP9z70emEULHMrIkCoUZWlXD6T6S3WEuCFK
GNWLT7+kbOsvhpuBOQMUJK+k4X3Tv1w2tpLd0mWJv8OKftuxTjhxYrw6htAORPNT
1AOKQzV58qPgkS4uNRaj/HjY3wuFwVbsS1tna69AmD67Jx/rArCZ5h+J1nqHCI1R
9PU8jY0xxjbnG6BObXjrKyLqkguYopPI+nz2Xo/dTFepFZLeOGL4qXLL+KsZtNKy
t/p4AqDtZrYwmyzTHPVeZTtCYX+HMSkbM0rlHUScoPs6hN+IeCyjAjpYMEB2Xv+b
VFQLTeViBRjnJtRmr0Exl1bAclL9zUAHdlmJarZm5Z2pqOPUMlWgHITi6b2h6Q+E
wMJxJYBxR3YbB7TtMu4dqNcTE5AwRWaX3U7pPpSKvHz27GI1czhlGAOiXEYBPiNN
1aC/b0mVuyThQlhNWP2e3VI1xY/gHjUgOtcIEre7ozMK9Izs4JnU/wh1SsiKfBcc
Kehy0G/c+g1FtkVdMEMKvmeJiiKcazzmWuxiQqnqCBjcMI/CL14QmMCPGizXHwjT
IjYF3CrXk9eNgMGF0Z8vKpBgWyysRHmw9JXGp5jyZLjg8tnm143dNQbL/3LFaU1S
63B8G3vIxBcevOUpSRxUuujLLwmX73DdjuFE8bZPhhnyX8SskdmBcFZL+EnEi3Bs
UwwJ/nhQ+CwxGFSmZim+KsLd79gVEt35NNNwz1on7rAeaZ4zl3FYR8l+3EPLTA2t
5o5B9uh31vKSOb2+beR8sshFvw+gYLVW01KiCzV/wCy1CgJ8E56JUkoxMKVJNBC7
teKaTpWr8UxrWHsXboeHXOXtYrL0CXzj9h7WYKKO37hpjP8LzqtMtXQF/nfTJ/yC
hqXGqLBGZ9IH8Xa8YGoEfgbn1QCj3eAg6JoU96OB8IQl+Plu1o80k24AxStIxpFH
QNTCACarZXG5V75SoqDz7g9uMJ+ovx0a8zmrH4eva5XQ3uoYj57bpLhtrpbk8/zT
EzT8P/ZPFXZ2aMDAHtXdyWESfzDf/YSdJXhI4I3nR3SATCJjW7YXgjbY5EzQXpWo
pSFTkjesqB1q72DrKetp6ZSNNEdi7/Ezpb7EFzTQyNxhoyd+dDZzf1q534ujXgy0
Av1SGNaLD7eDTQDKM52iGuycvzmbD1CJ1AbEb6BjzT3u65KT0q26RArlFJK6KJlD
p7b3HZuVgep1Etaq1I7dh8IGzx8PFdrzsWDDD8n6W8vePZrs66FA+shMDyTIj2cA
xegkLfdjwOM6gGQ0pYXnY3I8ORQYu0Jrw/KCG0i12AQJZYi1+xjraNmtRC7B9Gd2
TNfjbYR0C2msIjNHo7nqcqX5iIQF4srMJ2nbV4VeRS95RYpj8EDxO6Y2WjinHvxb
rHOE5jQWNZ0ldOJk/p1k1/QTYiwqyfGN79RKRcvOicJp88erWC4komF+38hCvppo
OTQZqVLQ3SBrn3NLc0423ne/Qe/TwvZBg+E5f1YOvkVOLajHWiZglFzfxF4YKNyK
8GAIg/rax0zjvW8mohAIDf4dHY43J3UFLuWOfzrd/y5U+wimKPjlAYWHeh6MjFd5
s1dt4Dgj06WMzhPgHG1+e3LSegiusL/cdIlF2IsURf6iV47osa1j4aTXEfBh0cos
WENBnHt9FLe4EdaFNNqXw1ccVrn2DO1IDnfQEp2z4f9rVk0Snxg/MRMF2YcfO7PQ
J0TaplUMh3GJew93GkGNj3mTzUmC5TjbIwaVWUnknLiYNPHp6uBRAqbniqEo6gY1
e9ohO9jkxfa8mnQA4RdshetHWu0+m+rVLl2kyMRWnjPeLIYRC45q0yLnIAVpxDMP
sriQRtAMGpBWuQUKa4ZLaAWupKJ+SKByoor3zgLczMcnA+8QpnybtgB93qxzrfMF
fwtsQ9qDhnCJTYzO5bJJAPDFCjc22T9q1ucrOoLL98j3aiMPu0TA8cn2E91KX15H
fwG9WXUb7x37uQj7vuDa1ojtY3r5vz6aWyMDDZ/JBwHVCh+fh4RIVIZNfFsTJnVE
o8hXIT6IXtL0DnXztntFdOgIeMqg1tepHwI1zs7/GUmt00PY8HvtqVTmBNdJueGi
MUljKatWGnr5I7kYfElXWy9nL6AgQnkRpDNaVwtv9Z6wlzyCX4USDIf6R2G0hLBe
W55wee0PY6fX0gZ2FLXRxQv1TDuWYMvEj4LHZX1JuMAKdV5YCpkQC4E6ftpmYZad
ZX2nW1NCIyzMzqYP7Btb+wUL0wg4aReyjDyxgBpb8bXiC/eDj8pNef7BD3ogagex
M5FUsI8QLfzgNr+QkT17zx9ymzgMqSkfNQnQLxfj+ma+ca1ql3i5U9g3cyN4dGT/
XpkBXqGXjyglBWMNO2k7FJKu/BC0NGdDsccesPUq+wMP3RwlhsvihyBrx0roHeLA
0fJKPgmjWbyvUNHfK/QF98BjqUDh60yR/cVtrv7aO/6kIRnTv7KPP8KQhPKDQhmz
VoBmX17EcFpv3rHtkC74cUoeCOMmpevepFeKIMSAkoPxlhT2mbLTBUyIcqJMwN6F
LNIdo0vC86TacvYRA/O+OJy5qpCFH50mr7zqf34j18ibGoiaXjBqasfVguLPIkmg
WUO1V6A+3rhX4EEY8enXQ5qa9zQK0QJaLNXzpsKSPSFmWWtei+UiNXaE8UB1Y/IN
gIdouGvEgd4Dc5ue3sYZefVzKWQzLUwqGMI5bKfaG1UhuO5nEIQgg09S+ND6j2r8
jc4Whj1Ai6DrMK+/LxiaZoQaagOugwLxVa+xlMUt+fSBEHjmFxccZJxpIDUY7dQg
xt6cRv3VjUi1DUoT7OXj2eP5K3jx8C67Y+o53DUBugXp+5BkvJftnkNzwa3Mv6iB
piAMeh7LaJAB2vkhvpwkwx+kPuqVyKBGCCF+0YsOB6gk/gAStY1Zdw67uoO3hB+d
o/JcaK+4Bbido/qy/mwVomudR9HhrL3innKoxwPaNTa+DBHAfGKAwdhtKk2j2emc
i0vSlExVcLSWzxnOvC/khLMiflW9n4OVFcfXHQoC7hXPFUZxaNq3lQs7xI6+5cr4
ntyLkIgdhEc/F8scdAEfdIi5c5SGxC/TKOCr5Kna7kGNLT4mrbbzQs8TElhLxE5y
9B7N9sx9HVZk8NcOw7wjaPVu+kY+r8WT0iJafAZ3PCQJ2xZ/tPm9EzC2qi+otkUO
UOT76byEzBitk6ZVY00ZURsDjQUlc/G9HhYM4opkB8D1VsnL/6fHnKnky0qnCXeW
lySFp1zfSLK8BM4+fJk6VzFtOzlsEbTzHpnwksTJGX+3qRO4jwPVFxWWfBni0ojT
LYK4JWM/XGm7l26lITG0oJTvp/f0a9I4Wjdn6zx5/QcP1E9rpEg9LjTz3Sz/FkE/
VR4UlqhRG1e9H9OYGNANYD6AdRZF4/D0brzbKXtS3FXapQh8fW6WrH+C8zD3pxGW
dORSgpDr+aPjXNN6t3uk+ep1LrdaFCACjPTSz8AoRreG0ThUXavLcnS86ITt9CN/
HdvQGHURiWQJbNkdHJSd6wk7y9kcOIB5ieJnhesKwh2IL6YkOx1CNClXFdZaSXQ0
/37i6deMoHxAW5XRwb+M1+IVmAutWoaN1g/NTZbQhtjdIGSZ15Y2/XKojMPJTYcq
W+ODkRM5tsdofTV8CQxycb39chp1D340uuymxab3dCEyAtYOcNF5KWRLfrPI5MMw
k55vxMSZhnWjQON3kLp2CAPI2GxrRJxtA+HXUhTsxh+cS62qDxJZijdVWdTQZHEi
Z7wvV86urLqP4Pf/ZrUSil8FPnlGAM7O396lP653Tk1vdvRFzoiT4YxXkzgtLCZM
yWUnGqbww/KDFsEzobU3l2KiwDtFc1z9sqGjLO9Nz429l5yqx2YIdNaC6K5mEigH
yq+w2y5o8JqsgM0F5tk2qmDKwRVUVsJWsD67xaZW8f+CbVKAN252ojmqiHu2DDSY
0WBaGUNBUwew62k5trluDGVSHfM8GiTh0e49EI9aDnxlGw4s4il1+3ytJzTon6qq
F/T+PlKu6i0g0mcCAykjF7JRPeFnMzvSvmOfV28ZNmj0joWc7GT6nYhS2Ur9l9Tn
lgI5I/7eSYM52hGxCcPyycXaVzJdzuxnwWk7f/m5sZ1J3uGKUiZToJTJGpFYUGeq
8o/7KfYtp1+1GGiy788UTPc8Z9kDz0vKdSV5a/vqMK8dK4SogqnhrUNPhw/QxJ5T
5XrG/36Go18epw+c+8bmHQb2zvqgvnkYif+7ZedfF/7Ek70vhExnJf2BFVJ9RFlt
jiiids44Rd3F9IaQapv9PXmb0TJrjRlLqlAn1ZeTcAA1jTiWoZ8YjKEZAHGtO09/
T6Uei6KAaKi3UhtFHe3Azg2ik9UGKdNlP5evM8RG2d7+pbOk6Z44JFBK35YNUCdv
71Sy7FCJDm3UjKcK6B/ImFilEchYiiKt+Fyn4pG2mipmfQSgbFo2CdedjcrmBfUn
gGvGL8mh7FVM+J6sP8NQuvgOYE3ILnARnMPrrgo+Z5a/yRi/bH6QdpFweMkAcp5b
IpbsvcrNlx3egG/2EWhOGwThB46QpgQbCcoRJJ2w6xoP4wVAXLqLvFpY5CWfBH7h
cwHIflpls7bZGwm2AMjicOk0rAlxkNfRUH5q9TJMgw2n2Fabw1Tug2wrn9a5axJ2
V2cjBsgAkjiTKeKLp0+w+hesn3IZFdHwM0e9amqrS6WOgshMHr/XIMRCOjaAXnH4
XNUKzJpuRQDhbv2NvSeW5sBfUnzUgSJpGKuT8KVsiSw36LBDK7nIbGEziAHPIJRp
xrvw1+CB5l1Dl01PKxPOj2DUPRb4PxcpoXuxB7tkVOdQiZ6jY9b26mHlTjzSeE6K
YigYbcfEZf3NjwMZI/zTsIEFf1fQ1nPQfaX+8Sxc4lfvrj2pwRKVHbTsTspStDeS
ps4D1+rnGAihVaPPY9YAJhyDD6zlmErxbrJO4zQUWqjML66YMh+mkyIC/CbrrQBZ
7J2cFwoTo25PXNjMiQnZ82JxJLKT617MF9JoQqSSe2VJlJ9FPhmAGLz7pTUy8nmo
Mf0CdbA3XRBLt9Z4/MF8y7AkvJT5OyN+BEHgPNASdl3XMcMrjyxeUMKVkgL84WfE
XOOWevNM8ZdCvR95+rYR5PJL3pC2nR6p0TQYq5fxUhmPxRV5MuiWi0wR5t1GnTAB
28IpkwFnlGm5/wMhATsbFkGxNDpOz6Ym3Hgvc4unR2E9suYHf/G5irsQpY0aJ3Nc
TB4HTVwRu/+sPq6wOmjCG42J3qGtQF4t1TrOhK45eF+JakV3qqemoIrF/TZpuOWW
ozlaFBd94yf0+WkbIFcHTTXz+ysPpGNOM/03vCtgHMI2W9afE8UfuQ0sgCxuoCDw
2jguaZP9vbqJjeOtTDxNI8APB5jXVaxFea1OjS6x37cS8EtldhAhT+q41uLl9E4/
B9pndnD1L2yeETH2VhdMd4ESAcg0KgWJrqe5Dxmsx4xfA1gvvVO8Y7I7/fJo7pI4
NZxVNKW7JGDtr8ToiYvXwZ7xu6EPD+Ti8oLqRlCz7GDWQjiA9Ty44NvAIMuJtDNj
pFDeoDGxb5UQOD2Z+XpAv9GTqDeAnb4hEaK8qdWZaITDms/1IIbI0MEzdMU4y3WT
14XV+dtj00YLcDdkzhlhgTc4C0ZCwxOGiE5v39+E23/370OSvq+47qKt4apgK3sS
DznOpcl9Kbgy/bbFsgBvNdLtrG2gqoWB0iX+WbIR16Eu2gk6RxtjQuV97Kzu+CnM
QrNmj5bCQKUSO4L7w0hY+8h0t8qkbTzc8bRCQt3G8lvirG3o8JG/nqEi9wUmg0GA
j2sAUhi67kN/uDy56P5jEaL+N4ib9s52uJ5uUpGfvxvZ8ttIdd1W9P461Qka7N/U
+63GW5OxZvMyhNHUtIcunTXForw5e9E4SpyIe5v+lhQnlpG04NZUh7xFIsJ/cInO
2vNFlo7vigRK9684Mj7TDC1sKoHeg7T2HhcB6GjDhIsnV2c7G98+N4walCRiIXVW
VUwXETIsXpA8nLQ439DY3EsEOdZfCQaB6OLdpApNJItbxIMWolw30HW4d444e833
EJlC4i6MxWM/3dU2Elx13J4zAxPOcbQl6KvYPv1Ufe+uuFzQH+Ui79RGN9d5U4/C
dyUM6n2PbQOAnOMA+wZI2IYz1+OUbY936596UAsKrvuGZSoVdm2GFEKbpkhm0tCh
2akbeDv3I7qHqsEvx8MFq2zzVulFS2fS+ZALlUcujJ+Ia764IAz0XNzrqdopOXTd
GgqO6UsvRHZ1SWe1ARbeCrLN9eWBfQAaUv8wEMUyipULeWST3rDSvVBFDiQIYz12
plPf2DQHKsyZvfkQaSQArUb4vj1CdshhJahXgVKRdP/6k6ec0iil/GzuGmf5/0tN
61ZdspLuOqGbAk6l9R9jYRLnGjUUfqJAf0GS7NQoOkw8hdEn+2A9imCUAugq8PzF
JvFj+a0TD70Z9YzfC70msX0MZlYPxHOrRsDSY3lo10hJCAddpLtmiod3qL9mmtrB
IKYnpZ2uEuWGvT1bkxca+XgDY5z1UT5wmtNHVJUP2qVgzVu4wrs2P9DeGCZpUGa/
7wM/qAzXwFhDkdJe1CkmKwIVuyDlm0pqT/4Qp6Rz966AbbDFIPHD+Skw2cQDe8wd
0K+HpqD8Mk8Nks7LkpKDTz92c0BB0chhTpYaml/yJs3qRjU+AQcDrULofrq9AkZT
rpjuZ97+MGNVdXv1feQSh3A85QxxMTeaj2cZ+q8h+zRRtGII41X/bCJEgozEPeww
p8UfewNg+HC7GeCXqKDoQc256m+binqzaCgVxgJ6b1wNK6rTcEjPHDPc4KGiPZC7
W7qmN3DECb+/0z9MiAPr7tvtnT8JiCgysZWxDSlus482qKkHuKkhjYDb/rcQEXPA
z4xK5uLmUjMFX2NiyW5NTDx7ZuijUIANGgRVsze8ct1oR4fBRsHs5W695YmNODwD
F07aqAdKkgqwaMjxQJg1BsGiaH/oF2vJsRCS17i8BGSWcU+eqK5rOLGKktHKMdkF
0jsKvU3GOhSXCqIBg+IRwQsoH8Mlz0TkC2SQB0QhLGFSesUikSB+G2K8litXAtwe
7IFIiN/Mr3b2CeejRxCPSb/MP1/1Ba9lt2en/x3k2luLtVoPk2kZM9DuiSUoMMGa
ZrmDoXtyj5OvPVG0jLwbxe3Ieia9jftX9mPY/taO879qJX8KHAL7wRUsXc5BYYKz
ALuOS9zcIe2eQUvhIAlCr5jEtzUI93TtOF+CED6ukKpIl9EgcDChABhe4kuw/qeO
uLCiRSD9o+RXupqVAW0cj0KhS5W+Cr/J+NwEgAbk652wlm0Ha/YHX+sOv0UQw2PI
nyvx5OgpaodLfzkrIAW+CC5I72ghNmvjKCGfrKCuGs6iPSxQmW3tDJJQGRCreOet
JvxGZTG+FxDu9rSHxlVDc+I2oD87MFK4z2FkARnHwknuWHs3nOZrXfdDZB3hSlCB
UH49Sv6ADIlYrEZ0QW/4BzRk5Bhm0twHBzJGnOnYxwd7KflTKIAau4tZ4WsEicN+
m0gTDvT4K9qqSm7UWBHD9NY39D3txmh6m8hVkuk/LmFkIMNqJGV1zivXI2VYfJN2
OItC84Viz/E0Ahnj3N6ZVbL2dMA5knyyq3roapFrfpWWg0KZf1ehZyx0xoDQbb1F
A9CH9pTJvhdisxUvdSZ3PuwfIFq4gqOXHH4k2qTr75X5LV+7tcn5FXhOF4NHOCA4
MIygYJFF0HEncDoVu3BdMhp6PNeHJvoCW+W+ouov6qUujU6WB8/Zm850o/OLRoZm
L3ogtWT6GMOFekXBQ7eC/kdPtOBW2xD7LeB7UUyMCHihPjBsuVumvLxyIIOGseTC
vvHtsZMw5xv0P6jjpS0xVkSMQMjxMLYNd5hTD/3fGHemoJ7xH/d/QhoiOgld1fR4
zMDlvawGy8esQZ3dELnaK70iwob+E0jXRJdpd/GDYrxJFpeSjf65XmhNBIVKr5KX
Qb9ECkBG5uTHL0q94HGXwQPTfPLUWM31z1jNSNi4r7p1hgZzKgBu2CATjTT/9QfD
Po0TnBnoLrDRT4I+H9hIIbxh5XEDANVgfkVepydqgHED973X+jPBoFywJxyERda+
Lz8oVKdeK2ddKpTRtDHmq03O+qGbG8V7W0s90pTXbsPQh2w0bEJHoiMoaH9FENHx
bqgc+wT9LfwjXIoKjIBCtR2On6V1XuN/KvLdXNMSop+uMaUqg7HtpQDy+5rPGiYI
8/FcGLYdrwHX9jpbYIIE98u0C5zBs35jrxO54WovsN0Dl+Ke/685h0uGzqbeNY0T
u7edHyx7q1E7PX3Dok2OtqLyxVGxj9o83H1m0TmaOhU453n1uoAOxp1xPUks6e6A
9IcOoko973Qfff8V7adakZa7FuU4lHx2TAWgBaksGXePtHDNqX9Pkl5hgeyX8UkZ
WCLQyVwJ3aRyFNaha0Whk/MQAihXBPoGLRFkzI7R1wBT0vnpElvZoD18MrmYMRRG
VCxmCH3NBgLC+bVdDRZW43fCxPmELF1Qc9Gq/3cNF0a4W/vFaamDJMaNkMUDGbe3
20eBxkjNE8oeto0nFMDzng7SZq0ap/GWQSkyeSrXAx9PpbFVZ8b3qoHewfBCvCix
kCvKg7xjMxh3z6989y37yWqrh7yAIdkvXg/cioEFGpt7/2CiIvMvU0T4oCEkiQtx
7DTrU2+eC9EVkztnpYOtRpS9sBlWzFGpxg6EWb/rNk4oJhJmed/sN37pO8wXwNTD
jt7cECx0vKGignvPUjWBYVeTHF3BR32CVDwpQDIedOTJTPdBiaVAEwH/kJVIt6c9
yFlkQC3L9aHWNx53zkU3MMJL4paywDaRy7kS9qYobNxUbZPu4WaxqjYZjb7oLuzo
hatA3TKNDuJU0gVizyjceTaT+9H54o0oeltV6mDwTJp1rn8PgYZjYkdQ1u3QkBcE
NDtgQOkd/WqRrvNGrzhoS1YFakx0wgrKcHmpPGpqTG/5w/VUBUTlnmaoudWsth7K
0ajZ5lq3bEd4SnpL1yZJ/j8XVTvlSK3H4YvdcqaHjHbw0DphUQP6dg6iE/+nD+OY
6nWtGEKv8UJ9zNvCCgxTLA92/wrhion793rWimYhHAFXGpWjUs44v5WZPoihI4wP
Zoc1he35hHLVuwL1yUpL+7k6I5mxLrOBfTqsQBH68fY6gLKtdasU+l8Z/gS5v6F6
XPm+ktFpifFcw5yB55ypcg+fV5tMF0oHLHaLi1nBk5jFhGbi/Zk30mFcX7SErCTP
Atgv6j7rE/vHtK+00kdh8W0sppMSJkoIW+jAFOI9799LyF8DwLfWiDgavw5D5h3L
U5sUU+sq9j2MtrkHbI9fw/Xf6nToH0HWH9nfBZYlVBAkpW9T6hUh13kFYijGDTVX
BdV+LeoFN7IxGTj/AXzb5Y/TU9BWiMAYzGt/bOj8pGEcR+etzdu0EJaSLHpTy30l
Wdrxoh7WVY4C1zXjgGLG+bquMtGoix7qM3KYHsEQP9FAWZHYd5SmMqE98UuoBTvs
jrvM7V4cAuflRqEk/C/t/F5drcHS2i3mWrXyIr+SoMnXtzYOgMgQzy2f0LwfSPl7
kMdaWa4lVCg/ztFbmGR4R8XGg5ZeauB4sQsSCBJQZn0A+2Zmbv7m4O1QXucuaBBH
DgVNBOa+t1rMHjyjMuui038U2eDh5CwLgT1alAL3OVGAKhwlH638h89mvBgEiqlU
K150Kgxy9xDeqD5ocuh91WO6Uesc+cRWraQlHQXMCV1GAuhgFWcooJxQd6TGY/Od
yuWKX9lCtGg9gY9soMZ7AaxgMklbmMGjRtcsnCcwpsFJx1s1fOUTj+RSnehZFE3X
fZzHzi7yhwI+7idYX/b9q8dKcK4GMbVxZSlQAGCnOuxge1qDDGjGNJ9VnHd2pewa
iwOgcQXi6tyVSpsV+o1IM3CSbAJCMU17Rq667q/UzcXo6f2GFJGcTqeDsMQmSCtz
tKvHLjZZXC/JomDICYmgsQK9ZWQ9nNBaK7if1pKN6/HCo2IGWmNQMwUf3iG5fCaC
521zm2iJgvc+dJg2yMaE1uRa20VUAuHuFf+Q+uKtaeti9rlDmbdPFycHvghvZzNu
CCLPCuhwhR1oM0kGZm4jo2K5Nnhwr8HK6Uj6XIm8mhbv6RvUg3fdpRS3PfpX6aDT
K5UauJwwlOADYB3aFdg/E+tAOR+BoCeZkIjPXvIQTY0AoHPCrK0QJr9ADFtgZHpO
PdEjvUzGa9Q/4mH9UKkbTthYUmYFMf2iDHOKrKp00TuDJdD4xu6MOt7m8v658cl5
+Vk0S5iRUxWL+YjxarEXmPYc/ylaUn0o6A/DD3MP5UhiMj401JMSYt42VnRVWH4p
zMYB/sghGetWEfNAstoWSjZzl+UFgqyPjjTVxeLK4zk9Q5QEF4qOH1LJO+l6LW0F
uLjD7xMHeXz+k++AUyxfgEYVByQ9Ct7J1I4jzaDfeItHw0Hi9rrKL8iUphcosjn6
dovZ2k9sBpC5Vt2VYbf+4I/Q+DCMhJUNFSrEJrXTE+wXyWmkpa79nuwjbn20OcDV
qkfHJo8LjL/ZOJ1by1rI6SdH/lRnbc1ALtL957Otc73QJLx0lIJjUymVylcsdiNe
7Zw2LRvz7G3rwBwubjvfoCh+zEgUZ2yozoQ2XyvA2g0qEo4rR3GDeeWjVmgI0YLC
TkF93T8ZOo5XZS1Tf4XreVvPPeCWlJy7uyTjxFMY07lQa+YyBNeMG6IaOzQttA6P
j0hOGWeBVtESjzR8K+LtBFgmgLknQh8dwi+Vgdi7ivFvBlF2dNPMbNLBtc2/aaMT
RxpAaLxg+ST1ZkQEEY5Ll/YZhB2u5oSxTID4JpxhUeEYI6nGwGKs2vxevN9IeTTH
QipH0h8UAzkKa+yhTu7e288g1yStRID9L4xbRhBfPOFDkHAtBulcgPHSbCBOlcU6
xKH+IdDHyazoYIWlD4/uh/Z6PEMmEkrvf2/JBMnDLl1uJttECaREaPWTASXzElVo
WksnTtDkrAU/riNw9TyHuBrYPtuFXzivt1Gh/UJlzm6AkneVscJbWHPS5q6VxrSh
jV5lSwHGRpJUw2Ir+xSd7VStC6dxU5UBSmefU//pRTaypIEuHxxKvwnSvTwr815b
5qacK+g/W935Po5OtuFPukDfbPoepIsxGZ+oGg3zWpXrvZiAwBuveCDtf8Fl8ZzV
4WO0Uc/Z0Wk018nY+KnAcAGgecFjKj6ymXH5WSmCJhJAO9A72fmJbV8sh2yNVkDx
xBpdHXrJfNnshwq6GKp/JI7eGJkRO3RONlMKzUZNGLIlkokkUg+t2qc61P3tLTqs
hiavMt//YdycWs2aG5a4kmLJJwukl2Sv+4XPxp6AS3OvkJAtR+ORXEvn1RWJyReU
tay2v4xPIAlsseKuJgSLr6N3f9PV+qrThH2wCHDhGsr+DIN/DFqW8mAW2Uhsm4lx
ID/u+Cck4I9A4jZ+HfHgKCOxKYP73yOzRZEGvMEZiSylYs2eE0TFt8bKYHQ/d4nb
n3Do4L10I6hKLOaylW8D3u8W+9EWSl3IwH8yOdhoK2n4niyQnasMJhT9stTe+d7a
QIayt+B031cM7CxpA4gN1yJb9o7ZhmBg7dOVYXBLjbjz8xdo8kZsQUhnpYisuHvC
CCRXQ6SQJyVtRQv+C3HuTuT8fgT446bvQ/0s02DBoeJ/HTAlv1maljdYchvltY23
S0y5rZDnNySMWeNEIEdKB5dPS9I5cTFtdDTmFkfxeNK3sXSo6Qg7Bqsto1Pod2Oj
QoHumcpIh4fnr78aVppw7vvi/uiHJvtyu/ip9WZVLIO9tsWFPa91rzbPfkdneav9
74TxVgwsplGrlKpYenxN4xgKKsqYKSd5io2QGv22f8kE4nPKtNTZw7XxWcqnIvBh
5qKEh/KWzq2s6YtneiYL6jQmAf9+62pibkmuNYliouQ+yI8AZ7OT988K5FzbmjrZ
nA2GYL3TyYBcEgONMO2Gub2nYK5qBHumzzvAwWfRn2fdjH9Jnja9ihv0f6CldQLp
eNw9KsJjOZweAkTZGpaoiWBDxC/FEA0ICq6AU63oY+fcbM/8Knq48pwlVkCtbja5
32G7jYt2Os99Wr2bM7YcG++0ISbMzEDGg62FQ843R7CGD27FAno0A2sjcMFkm5OH
5GZtFQdmHNcSTidofKzPaJzQ//uBo8MhUuP4XxoaljSTCKALMqRvW61lp9ixjfGs
FP7o6J+2UD+s7nvFXzQCvEAKLO0r0SUWfbKuCsM6aDmgzK0d298SiglEb8k9bOhS
YL0p9v176vM0rWbn05IOWTj55fbHngV41MZ6/AZeIjMg+5fDOlsRIWhBlAO3xcd5
V0HpLGTFUHjiY/lzvdOvoyrNu+oXHbp6siR+rA+vPzBHMezF//dIJRw9HCWeSf0T
i8qqCeRth/TAMntCb2dzaWJVhHUIEzSj0+HbMzl4fXgAOn1EYKlgS65p39nUoPhd
5I6GPHDNkgL1TbKIYTiM4fo+SUvl24J5ZICgXw5ng4TTAaP/xLYc5w5jMUTahPkd
5lSCk0p0MJIdDqCZmg/nqlkv+N0GfqWJNZzeKXjNfU69SCWIbx9CqTx1tnX+4sPK
9OFqjY4E67zvO35Z+nuSwbo8RSkVZe3K29X5hZ2aEatkIazW02LWrlWd0GEMtE5k
1gRaHxGPOzsUPHau7siA3bl14tdlzfOJTacpNWDorjAoxR7IuWFfdRrhpdcqR49U
f+kZYzEBRjiQg+s8LTuPTNON/WdwwB3sU9jfGjepWDNhohaQVr2fQNwycOMjQod/
45q73PGb8BHjfuTu893GUvpDM+BEoLAS+JeT8jZhQCKp2kaB6mdMNf3Abkk2RXw1
EX8snWArqHjfX+VzwoJTv0fcN3LMwolM9jblPqzQU5N4dA7QC3wwXWGwMPvyE049
jYIqNr31sma6IuoAlLu7I/7S2Eo573xbZx+4DwC0+axEpMdbUJU4dY0PgLoaUTKt
C0ld6cbNSa47YjC79OBVbS2xsb/hZxQeIJ2totEqR8JSyNkng+We6rCWbCiDS73n
25rLIGpnOjcD9Hh6UDjC1RdHQtyagBuGPz9JcMZnORTK/UpgYmAhjH14YgVeP6CL
u/8oCAyNVmXW2TVpJMoPuJ8RKLQJnTfNxqzd3VFvIpp0kaXqKpA581jr4+VBzsBc
rP4lhVzXxPHdP2iwrlYF30JoFtTRrNo3bVdOlNVa/VuDXVuWI01vomkLJ7kiQLCe
wKPMvH+FlWEJnDW/2NRopCFmGWyRb0XUx87/4dxhMiRIJ6Ixud8P/H1C/szf9989
8dWIupTzwqZQuLveH74nduQ3cZmKWkJC1LvCzxuTPJehKdMkLA+PHaW7xAWgy/LC
mwkmMZJ1b0ve05e6+jFHtmSk0kDIV6OAdDhRNh3CojY3qPub12IdEfTVNFjA8cs6
XZ8A8gBceo3Zf8n/1gYNFefeChJ9pcEG2/tFdT5MCz4hcunbwmsdNyvDfM8k0vfB
Sfp5wQ+gXd2LADgP0l0PVIWRyrNBNtk5LZijjTVjiSMZLrTzNPjxUTeTfG6R42SK
O3SX2ha4kGLu6Zf7w9N+qCvtWLs2Uc2WCt/VZV6Bj6tayQi55i5mFBEado9ZCYi7
6JOM8/o25ZH6qKIBRWf1cou2JpNqu5N7gVAd013l5pidoy3E9V//YByCr/ZVgFo+
AO2iaunvOT4JF3AQOMuhFn/S/ig9auRHngn4IengYLvJX69Z5YKg5C4jE4jvChVK
D5Rq78g6XnsTbOjyHjlcSqnGtij2odisvsFTcvJ6GjdKcqbB9CBObJ4/rFNlPn5T
lfxs0EaOzn8/1GM8RKfAgeWCpr5nG5UP9vVkmMvPQmZz8aCQh6byWUQbB65SKUJ2
jmIUGasKSDUtKo+t/pRBB7ERg2C3QoF6XX27gOwMROLPi1PIxDYn2D6IEnRdkleT
QteJ0UyHVlp5DMjoOpSrSOtETUK07mpMPEpOFvp0ejCDLOrbI34uWxFA7B0wmq3l
aojzgS4O0SVd2novr9Tgp2QjVjdhuW+l3UXOl/DxRTf0XhScyecytIiIxlH4HD4I
NaVQRw5GcQFSAd1/fR2iwumHs6Y5+9q5Q7/5wCISaM11Y0Zghsx+4x3y7uUrP7Dp
tIZ5tRkHl2kH127LUs9wW4E46MwlDwwu+ZTWRNFhI5GZnhykGwp+cEvwYHBQnn0J
/Nqqs0odO4e9uXsf9MBIEP1KfcjQWfSeD+HmocQd+n4Fpm8jtzTMKh8WlZ9DccPN
Zj7snkIKBWb4apvLwj8URqsiYxhDmtnvmBuJ3LUwXtok0fIw8iolnwjQUNvdv4sS
zwozOj/SQjC5KUbwVF4fj5K/d1RWP5TFymdkp8eUAScTZS7WOZ/87mwi8uZqdWhW
0pGCgfuMOMilitmEywD8Ukt9hS3SMwiEaEiwLsn10rjP51xVkSMpFhGcDBV/aBHi
x//88QLwP5acWD3o+3+U5840fd5cvRhxakqyn9bcVg5++1uHAHrreVy3JyeLJLUW
1b6gEsFBzO7gp/LYOhQVujJrQR696PXUOZO1Pr8K3E/ZTcSBhkz+ub/57ZXO/kcj
nOf6+bb7vhi8kDSXdAjdRqy+Ruvs65HdzTjSMuxcCNlhyj3e2RMPlsa6D6XE18OH
6L0VxsqXvmzuLHODNlE+SeBPBi1l/NwLV93bodo1tX3120IOtWvF+OsJF7rYA7vW
d56ePA7ZqUrYXfEjOqDWrQatIYj+74KZZ0jkN78/yW/BqRiQTk4Q4vHNSP1eVJmH
qF88wCga3hcAAkN+Z3bf/wAyX6UPniNBh0LtqFniRAPISv7t4m7J0Wb4tD+kTqmU
iIRElSBp8gr8nF0Ex6N/KeJVtP6QPWvMT1exapVEMy0d4kMo00czlOXdniO3/1SY
YwjPB1e18AwDHleAxPSD7ziJEy0N2m34C3al7u10PrYqPF15s7jFY+zNFh6Qtz1t
XPQpApZEVV6n1n33Pvbie/DlGDxGinzznQ4H+7oduz9eG6fjJ39JkjDJwx55XPGl
KkrD+kpQyKy+JzknmkBjgiPMgR/JNy4bkpyleq9JE3wmrYL5wz8KiDRJn1ujunTK
IzA+6rL34Enzp07K7gNpYX1ZY6MbXc1K+RqHIKN9u2u38KoAged4ps0u+Pp8Rlfu
D+mfTNjHIMd/BGe6COQoTHydUZ7NTlRkpSZX8YbQBw7CTv7uVu1LxPQplt6WRHOI
aYdAt4yGwf8i7plpG3rZnQOJ5scB4I/8ogIbSE9eCJIeBZlLCipJuwcppxjxtUuR
X/hMvWoSnmue63NaxKvDu9i4RQtz6FbFCT2pFjDwkkxm1oVD+nmK3QibFNb05LuI
7xQH205TCrifRjJLU6oA8s1B9xMCd/LpHbCiu4knOr0PFGYgZTfbRkYRph0o9ky7
NJlrBkfcbADk6uQN5UEkhbf2h2TBZSJQ22VCfEJxxO5NnNIxkbAZyEJn8VRjn3C1
dE64WL1r9kSVd+36DzJliea+coUUHS31xI7SVVi+5Th6IVJ1orUXBcbXMebm0MoX
FhFzLYg9GdHlRbzIt/jf9+vTzJF6TUAhV/99qoWE1gJfORa3vvK1Q0Y6TDTvD/UE
fDL66ZLxOp9T5YRQmFKOW8NU5TDv8m79WwZ7cYOiHSdInIIyIQliRSw1SvtD8b7H
Q7/ARFHszUf25aL7m5Qp1+4YPz5PQQjBcHwPlMGc7TKEziutlmDXWqe0cdkX2Ha9
+HpBRolXRN/NyFEOUO2C3Ie+ncijdXXqiGNUXYpVL5W2ixxfMC4zjM/cIgDr5APz
+iLlfkfvJ7Y4tjMyp9iIFeSecjUX0WtFt+YdzpeI776lDRLdczG/MrDkBER0NZUr
YT1wmylK7r13dm4OWOvoVB7StQxaMoTMRAkCATPxvO4GsuK2sbp9Ozgs1VF4T2LL
s43F5ejhJnwLtzEy6U0vlokt4tcKXRKvBpNxp2L5r6YdME2/fzXt4v8pqYMMg5yz
bOVWCrA8LCROnVkajPz1pPiEvZ7aFBiMJ6d0RY8qE57V7wv7iF6REohtm7xRGR4a
E1obpebyDTTVTQp2mCzeOjyy20UrlygXRFupIdSBPESeV2ZTQoqrNqytqCY6bvVo
8VrQSaFWMp+57iiyuIDIFNfjVkMFk+SAwqCiddKKIuPZJvwHxHG+bDsAS1Q75GiA
T/VFcX/+ozAozxxe7Zkq78ynkLag5MXCZICGKXtHPUTJPry+QYnG0KWl7Eo1L7ct
gV5G37KcVh8qVZR5/iv6iJ6ugwnmIKNxlpC6tZVyEFs4LpD8MypWt3GGq38VF90C
qFGi9PJc8aBa39yFfWRSg5cO9snVC0esJ7oFBDkrUgiuio1L1AsHky58JQ6MGKkk
irhNOpPUCg7jiFECYuR/XtPqfZuJ66PUyhxCDq8M1qzj2TCvjeTvPAS1/k4uhTuz
7AvXPxr2UdQi9KNqUXNyO9qX+NayJ4IIsIL+i0O3HmfmGzyBcX9kbr51zimhsxg5
D0Q7NvW3nqQfjqwGOScxu1i5MVPKjLuIa4Zd6cVf7DHCtEqlYiOeFO+Yyj/gl3zQ
5uozOSK0YSwdxnzUFmYNB+iZJ1r4QSfA8b3+/mHqSzx3WugweGitJa/7JT/X8zZb
SwLs4mGJhLWBWVFwFN0V0NGiNsnIp+aUWprJaCOdW1AcPldk3n4EG7Cubm1tLc2H
Lz5ksJwnYYYItWPrnVXpR0n/YHlbCfpvFg6Ltn0AVAuLl6FHfadmyZGHrbXXeTQr
zCrUQFtOfAgxbnWWaelLuLWsI2b84zDd3rc/Sx2SoyfYQBTqo1xj0g24bLG+69G5
MSy4i3IsdNWS7jHDeWA6rcdYfNGKk6sFo+C+y/noMjZndsT3XOhLb/5YCpbL/QIn
quKfeDVUU8JaAwbqwXBL64q0t1GDF2w4iwykYrQy2Fvkw+vFhHfkp/wzij7nftsH
Iz6anAJ8rmsrq1gqwvoGPlMBuT9z9EunIwW5uu7ME+b6FhukLgHHEntAWqfqhHC9
E5x+aRZsflCpuY2pvJ6yX70A7KZdoSniv6MhQuph3Yge4Mp4ilsxTkjmBlqN9eVZ
+B2lOZdZavDr2sn9KQTkXWxMj8M+HIUfggcCLcUJIFTUXKBj7RzexWhQml5SnZYn
OqpPjR6Oupza8LJEgk5/+T+IsqGUIzyxmFj6J9ofGchRQayShpX8At4e1CxpKKpw
`pragma protect end_protected
