// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:32:37 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
nh4aWa5WIEV5HROZrfJd9F+Ezady30G7Y2A+hkZnwt4/PnU2vqAecEoW4w9i7x4D
Rzf0zs9fuXdX82BF9+2gLcAVECSqzM8ok6a+JdKuw6NKd2MUFP/S9q6r0rR0X+TP
XYNIxiR0fmr+PAn0i+dxKdqX02omh6BvQcVdDOPXj4Y=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 176768)
kLQI/ZMi8DFqH0Y5MLKe4RI/EtGUNDhx3f+UYzjzb1IyijbqfZByt/d6XPo1LdSt
MolscYmirPIWma6ataQvgDKSEq9qx+2PJUWjtW2UHOLj4jhJuCG7cyGjj+/l5bqK
+mumS0YKVsMsBBfkuLhhpWcPzN8JmqjEIYJHS4iTUQwgRd8gJvgG6fXJkIWwKsC9
FPcF4PotKjK1/DjW3rxon00cMRwJnWLxsX2UWqxpj00lqQY2Xl1pLYaXrt7/hzh+
sLT9xrA/u/D3Gs3jseNa5t/mNeuRaslfiXlm5HU2S9joSrJBd75VUgVfQVf0Oq+7
k4dzd8dA2wSUCnXshG5kiXLAdo7TgHqjFlqVSgv9P9QLww4FsMbIPv6rlcXaQjP8
e5M2XU03oxPhyZzWZmmY1SYkUQNgTSYUFm0TU65FqQi1+Y+2tDnHHBgm5e8JZtQY
b4rzTEv2R6oOunVZj5rX+E5+75QbQzJCBDtHs6TUBfo6AFLG5SE7bJoFghYJqA6e
mxVaf34l8uiAKzy1Ij8OBUt5sbTVx0atG4q7HSz1URUHjg/2ukvDsu6OaVYqDOv3
xgI0cHrMq0Iqpj4KG2fqqx/KWXLfV9KUZfAZUZJHvm6llk3Z/ZWDECh4FzK9Ripo
+TKdxzCBJibb1q7WiA8439NAx2vpzlx9altWg/sMeLxD5B487VOSXb7f2DXiOxrL
EIjZj43Qvs2GvkFEJeSLpZ2X7PZ4ugWKTlswjmlyIkIMLkqaCre2pTgTqjdJFlpp
OhWa97xss2emsx7mnmX+PIOuOKig492Th0uo2fEwBqbb/vVr71HfpAius9o9essj
2LLyJeJWaoTSYZk3NqvFTd1z6oRkJTab56pGKWxfjkczcjmZdOwaJSkeAz1KdyNJ
U65aB9HSysOuxj6mq4XSTS+Yt3LG8X4Aqhc2LC987OQZEvLm/ROpCxAYHA4wgBvy
9UwryHlsg0ANoJa0Vw5JkosbOzENo8pFjfkcxMx8fwnXbzp/FqdHCKPCy7MFbZyi
NfejPq7cZxZf1NjOjyrflRiSFW2dlcPSL2ve9fcfKYZZOg3LWvNwv0SfjAidlGV/
wXDPv4KOReCAUJJu8oRBXt5GRu2aV8EqqMSIqOLOePk7Maw1+SLRqVvLAymAmy1q
FdtjxPyiTr1gxDFBvESQzG5v5BKezzVl7DWnc4MiNGHIb68Kwoz7kjJihnCBrF0V
rgAhSEXiRKYp2FdDqzfQizbr/xmbCDNsM7g/FJUnMy8n1I2vj0X8x8bBBPDK4ns2
dTcJJxRQnYTrS07QfI/8Yd8T9i3t5ZXhWw7xob/4LtWhQimqyzj6dfsQy7Y4b5in
iYcfCKyJkD6tsorwjGkY6vfEVsVSEbrl8x6+k5J+/PN9Z0L4rZ5FuTcNyV6pF2CV
TrGKIKA0TULe/nBOgrl2VNgzTlDbrbeyTAs+8QvDNmhOJ+b/LnWArdnLZ+kbohT0
TpCueG4tXNR2toYkc1kpPETIkKLtSNn5VVrhqsVVAXd4QiTdcQ/Z/0QzJ/dRgma0
sjtkMJwT42P4+ddcQK329OBE83uD2EgxniwV4G0j/gTiJJej9LOC5UhMviT7PHP3
cwecpz4GtRQuYBPPmVuYHcf6ThezdGxV1BHw92X4a6GAmEB3MzmXaDOXCKf5VVzv
33WeGEZ0I5qeS0uqHYghUZZnIHio2gDt5DBbZnvtrHeqJBQikgtqMi701DNHOtzQ
7RB64b65KvMKHkoF0yn0yW67TSdVsAaC3qdhFsa5Qds0D1XYZ3m9j8fVSCkvvNZU
pocfUUUwsFvfhigK5rwPxjzUxb4eJ3hIIU4FSHGHGKDSNWYYWzXRvWHc2Ex+XPjq
6+KFnqwEDGIl0jCXtWIKUXGZs11WN06FQkROZgVn2LLNo3d8n3AY8RFP9ryspumt
K8RyZXc7B2z7lZu1fzMVWudahX1NRYX/b3lXslrL1XpEtp4eirMyM2mYqyda6yqi
3KuZzmvXZQJ3QUSfWM4tL4J6iQCyGI1C4MzzHj5uSxLEpvlxwyIv+FCAlXExEQil
QbPEwq/J//Ao74fMJBkeRd49WRGNnt1EifKzgNqgMrlXqJ9fSAUMJ30EZa8xq83m
o2tDv4juxywdE4TQDWyBmIZz3qz1/Dnoab0g0h9p3a1EUzHHWWaYfRZaEsAbba6v
ZiFBRvxt8rLA2ikXRO+kd4NgDla3ka7vo7F6CKkxWr/ZqLE0HPFUMkDaB8DCNHnP
YPtWhlVQF6oO7tNFLs2NP3I/CNMWhTFBJTRLrmACQoma8kEPYNTyHXezmJ8QNtK8
vMiw+rGGEKi9agoUa6ErCpeinOqe5OIZolA/Pybx4Wsqfs5RFrrlc4BzN3qrsJHT
vGGFbvz+YGiYxNyfjViGdRHQUs7Df+6NaFeMQKcU5YAZc4K6qvz8TJDdjmWJ2PcI
8jDNo7sVyYL+UpnobUFpGnzO3eG+cBs+SPtIeC84tUFS55IU8TWX5uVDbq+GApVI
XkTtUrYDqLflAhnj8znl3Tqc+s9xeoPOw1IqhF+UpX5Z5yuUVjgQ+BWppmH67BCM
iSbHSZrRifX5XNnNN3vCp/GfZaYN9Xc+8x8lzp6krRj8l4ZKVsFQmPk5+wI1bZdT
iAp9TxwF4Virk9Cr+kNbzTDH6IEFVwe4PgWKEq5jQpcyjS4OyTqz+o27FHs8Cj9c
YDCLSPgjM/WczBNtRra56zGJ8KjshNRYiqlj4Z3uIHkr/BQXbpo16mVC8AQ4lg+o
szTHUZS8iB3H++kEXO5MMHPIzqAg804Tbw/q6qrLqmDmDgLflRSSaMpgZTTfL/AC
E4EdwARIQpMCNr5JLddjlQEIvL/83I3sB1AE3CzlHk0yHpsUc9yF3/cM+iEJ7Cz2
3IsnzZxS4xgnYGjFhm1leaKd3VwJOBaK46tk7f0vM6aYSc5HL2Oo6Er6AsXFuyQW
OaxZe6v0NA3ryzPfoc9e/Dr1wpxsEyj8dbzmZ1Eh8gwtJyn+RuLe3qrfKzknsKpj
K7pSSYev8ayvf+UamP+lBaPeWTYBRHOrYjUFxkWB5GzS8CRpMc/j6ltWZCMfi94O
sqAmrkU3moEAqXCNDiZY0nT0sVsRKGf/bldExb+e+HazWoMELU9LF2wKk0dp+4t7
vsYVRmMYnYmbNifJN9Ye0WA5Z7w7Zd6Yihy7KSVHLPRHQx6jrxCnC3Zx/lGFw6qk
dY9l7G6LrTcI1GyHyGa7FM7bEsUJik+hGs5H+8rKDGSr4QJ6NVq02zpSaevblWzb
t1DpMMyq+A8x1qZTZXv9aNWL6sbDEgFfvXCws1q0PVqFL64edT2xQvNzc7cxBqn0
rJa38CIny1IgDiG9LABMtx1/USyBcaABwT4f5aF2FcvmurzPTX5mbw1A1jDtWhtg
Lim0O5Gg/Qc45My9n9tXIFXk9RXM8GEvqwMU0+8h5l6lGe+piInq50uZlHgwXmbo
B/5e33FTy560n1v1OEJFEmgMhR7HGby4qg+eKdAGYY72F+kH8ZDDRniTO9JDjRND
OxbR6mFx39CUBnlA86/inUr2wK4cCEmiStSKynkmxQrCW5q56cFrz8Kue516/WZ3
wx0UnUlLlPikawL5ytNQbEmcY6JfG22VI72ZBROFQQ/QmyKXgipzUUqvc8IpI1hY
QAbx28GooEQGhxaTUM3vSDP59xDc64kLUybZUmKSLyzK3IumvYvPjMmYjf4nNulH
KtdwrzmF+A0/lTCJUfR+u69FrgkOjtaL91a8lWnVHSq1C7OC3GxWJDb0GhpO1/4V
6DlI+HAg0CXfmMlhfOOVyprSaCTSrlpfbVctpW0WGJ8e24LYu6u5oXtM1HKdiRF9
aOF48T5NnGH4M1IOXdXsUui/CcvKwQ0vBjr8ceUGBb94U7eFWxLzsr9ugfCgAHRF
ygHsg6qmkVRdKRoTjEwMAbO5KnFO+ZoT49xub/F5AFTfA0V96q18Lp4Ha4aiT+pf
7R0brjz+NfH6XT5qb5IPhzm4zMEYe6CuQ6x7ht8t48jzFvrCaAOWjZ3wZarX+M8e
IGvq8TtJSpwjfz2w98+OZqLlD3DEBVfkG3Hnn/W4yaMIt+3IjuhzRk0yr0iMUKmU
T0K83S1FlRS3i6AaGGCvi/6fvZ6MVFy2YTejNuBfaxV150JZH/TdklZidu09ptHb
pnXiSZ9RLljV5mjUCTvjT1J0ZSsrOaIThT3Fq0YeSnBkABXplg2nBk2PWfrIgT8P
ysAlDhI6B3AB3Q29dJc+OdAsTSV5RE1LJOg+cVDY4wfL6IQlWnJZMgRv9i5NQmmO
vqIolvAGojpnFL78KZxYw6vEyVorcO2bgVDMDDiqgIXmGblkrCvLGECXKKoIG2NM
FJLs0Q2bdcT8GjLaiNLmR/ps9XMMBwrAMNzchUkepo31iLCx9d13oQdJNhztQ49l
Kt1Hg+5rKB/AFnYS/zdAtqqVjNCKjx+tpnojBHYWZQy1jEQMNrcd8jVQ8UkP+9sF
7M4xprq+YSA3y4T1GCPHfhe8zZghsvorxPkLVL/ixcxZWo5r3LKbB3L/DWiiZwt6
EGFF5RVIrpix1ok/Mm5TTKKmxmbuPx0IqYajrjx8Zlp1xcYhB8te+4p8c1oCZFSc
Fms59HkBtneaHGejUnfg26DVWC97pi6AyRc1YdKMygkcZteMuqGqt8KF+a0q70gb
ynmWq40ixOKYWsT9dSRHxkX1+eLMyXX15nGmE5wZQ/HRlhvIQpdlFby7EJ9QNXiW
q+M8EcTsf11yxd2v6dZoSHk0wxGjU+SqWc7fwp7vqiO52Sa3eGKutlZMoAFwRdZ7
5JS21XlynvRBfm6AmqlMS9EnixHCYoPR0VhLTp4TFyiVUvqOS8wgDz3JgqWdy3sh
PX9HiQIei+pcLyL6/55jT9krdVMJbR25cnZbJBaPu4fFVW3EiFVaOiHDYRsq5xel
vPFe8OTmL1t8lSKVmgMfEoFL3iYEuKWvzuW5xuUcOqmvmZ0adV8XQUB0Ad2OPw1X
rar56UuoAlhdGkhrXkEWRmkjhveB+v1oewQcu19+67LSjmOXriJ9xA0/yxgUsMav
qVun0iMNYpGbpzED5AjyabMi6BLoe8D2k1i1VGluvqacn7G2wEtWwJmOQ55CrUcz
u1DwuhG+l9C6l2aqUlibvAiKRNaqFit4jU21/NT2WslVDoK8XJ3gC9gwNsNRFpP2
/g0U/KilwNIazzIXCvqYd/86MWmzWQ+VARKJLI0+ordcnmpBad6WwVpjVOid/n0x
GMkNR5NLWK/FTToS+W4cxG4SHuKeLbnLhquQJOJRVMjfsZTTitNh+hHYsiixNBPJ
5tIOjuQNjQ9ccxQbf8qfFZv8eQdm2VA60gvCYvjSQr2WxYVuFt65T9wMU0uw2ETJ
xslrSYRy4vUj4ZshNPumZ8ygpqHsLgd9F1g83nA7VyF/7RGjcJTw6l/Zgs+xdPFr
V1XS4foF5vawKYEBhE3U8yStJoKkKLzUml8qGdAuVhLf1Ls4eGugMA6S1wVzY2FA
+QYr3LZKkQ5sh4Yk819W7xefoat3QruEwWHs9fqMdRkKSmhhhcvkr61h8+MO0G6q
wQ1KPOXSz/KGYwxXFWR1ISpRp2BCDWttHGAZHPOpzdqsX59j/nj9Ob5sMMuV+Dj/
+raJ1jAG2fhC9WZJme0bEyJMyPGGRUd8b431nIP0LfjfF7g6pBm+f957STCWghGC
s0oWK/OKtfltRSIxhm1TpZqFytLzIG/8J//oSSNrDnRC0rzTi9yY99UGjtTCgtoo
vRiVwHGkCurAU4m9cvwP517BjFEq6Wf8UO6Ma9ESSBl6gvOh9Qplp0wrMY49WQ/3
ArM5Fpn0SRtg/8iDs7SD3WpeEJxhrgi1BMyMYBITz0FBtwr3lyML9afYiRpnBuAK
9Cp8rJCBiQKiWFP6LlHh8EE2VIedOVVbWCGkiLaNwIjZnjUZZ/zRWzNDyRxqsaQe
s5UwLVa3VdE9MDV1yoZ4cyaj6Rt3MRWjXAxD8orwqpOkkPrEjZB0ydKdEeuasibe
JZahmbItzDTF5ehowsTq0dzQlgvTmQH1uYpegtSTkBlYyvCptRgbNsE6jEgvqGn6
O21rB3jW4GsEz68t+pZtYCE3uf/HCi10nVH7I6s/u+cYHnnvhu0Mon4tRMnyVTpg
u5Bxo3ooko4NN5IYNa9EO07JmNBHjCJpv/wxJlXo4UGV1AVOS1Lbeda8hoCW5Ni6
+I76+/RkGXWQ9u9+UpZE1rhxUVeSVDAO2Q+0fTpi/C97EeT0dNyypDd7lyC7bAOi
pxO7vgbX7DpU/1lD+CryUTe1prg1iFBwOuzYSYnIe+2mBqvYcZtdrRqOxaQ0Nxub
59oT1zbPGajXR6fEB/jMEo8WVhcg1eW3VEE0lb6xz538o4wF6CN3s3I9wi+WK8ae
oov55pJRgFTtVQNRbnoYHr+TNo/YK77G6Q5wxKiaWqkbu4vw3YzeBoL1YXjlC1Of
uMoKtRJ2SiRsC2sCbtA97Hu1+Xmiee7Lk8vG3/mE/qkcSLsE++Z9InbTug9CihbZ
zCKMJRo1cTXmPPfdlDWoQVo5qrujAhNtxzpitQcKjLzqswUKmZXTDgBzkB7X6hA1
+ZylktAp6/fBKbKX6JSRwDnDI5E6K/W7sqLI49sefBtsPb3lqct/8Wpj83sa7Ppj
jvzuUrnw6DE3+g+bXEMFaK50tXS8DiK9VbdD8lSISXb9AYKkUEYvMcr1yUukv02j
kRgZTAJjDql7J+TJ/saN/0pSdYzCbKeS693A30QXtH9fvy7iQFRPso9Gf2hem2j3
iqPtzS8KBoHraRpF1nOKILcpjfMbu+9Z939Wng1DWNZ81F0BfMVqKuAh9nLrjEOm
8/NMfb+yLJq2FDyBUWytb/2u6ybv1lAvUB56lCER6y+zufaHv/MpbP2khNF4R4DF
AkB6+qunFhNgpVA3QH5zw+Mg1D9iYUm2mFFxsQO2cGEwyDNtpS1YZZ2Mcn7dcHCe
XKEfiebUTcdCB+hTfZx7/bll0VQ6Tk2bcxab9T3nOM/5c1o5AaWJEEQ48OfaFzDn
EFv6b1hbTfk0B4YU5bnwuZCLZ4XHE2qnY6RfCYDA6qyxJlhCg0klpzVZF3VTZR/A
Y4Zn41bqfMJctVHsc6Si4aOFokyhLIFJi/k9Zd6E2U/pGZMsxp6MlMUmxv1665jf
ATOdm6JFplD/nG+d9tAY3XgJ7VbHzAnt9sJNCw99lLfu3PnYEJJcP/FYYA8S3az3
t56T/fkDEuL7TjaWf9cgCWCUzDNx3+oBYWimP8FW7Yo91Eb4+WLkDZFOpeS+qlAt
Q8yIrAnnqwmWaTU8LMnSu98AjDdqzR/vMFtlOjVgSZxIkVUrDxnnaL372WdJE/hW
s4jlr9iDKK1L/wVKwS20hTJfZd7vodpYajC6nnji6dOn7KDuQdHd9sWlPiNU1HHi
KXNF5kI8u2kjZUb/IqRywLy+hi+J103kHAa7tfrPawlwV1lnQyL8tPWoJ7ASaNkE
uxvYBCWgdP66+l6AXL2I74cSVbb3fd64CxOg1LgZJBiMXg3XkuFWsQiXrbwN1l/f
aPAxNtS0gWBDlapFshXru2kbg2H7TvckC0a2TE+gcE8WLEMhhbbMTMOAS71YNN7C
GJydL9w12AF5b1IhOW9J1wC4rhcM15KaLkOHy7NbFYt5h2f7iaj95OuCBdrg+tB+
JLFVy2gY5/f35G7ZlPAFW6uvmSYBjocuwB2ZPxQ+Ny8pCYv6LgID4rVah/nhMn7l
IZ5yNt+nbHTgTKFW7p0FzlVWrANWyPxdY4KcFtimkRB0fYgoUfiOtsrgJBac3B09
hialau81oNelH2fuimb+/7FOZlUI9EwjuFhjNjUfhXtgNRx/6Aka1wqJD+r1r4Z7
qtQxt9rBGqfvZ+SsMW1pWIITw/bF1IktaHImsb9KPmoRoJ2EpndnQUNhDO4vZRmc
3VrIe/H/05ZQsslj1VUG9exZiWXXl+Lh+yCQVfmOJGOxTNdJL6uZCALlyZW3rTyM
b3aZ0DQkgW/2qL2tqdjvEKMoDj8K1N26elaEpF8yoHuyZ0Dsh0jT8nVofOOG5Epi
jemh9TrpoZ2dZ/DGO23Myn+6+oF+pHsY5DIybZS8t+PJESAGtkgkjdxP8cLVF6wD
cPDqyphzoM2q6tANLxHjMdk2SNrwg2PrRLsUpCpak9KU2K850/AdIishbWGnFM7B
giAPEdjtGiYYq6m3ftGMofJ064y0sk0/EH1BhUKq3jiIm680nHsWE+fSiL5zH0jm
ZzFSqshlMlAf8i41PGrSfDglEG05IkdPm4lDWdsmvwUxFnTcJKrhQ1AE+ytjbHOk
bhFtWdeTOCFEJIupG3r2rYAbrQihEUDVsfCWPwEirEzp4opmgtmveeI1MLABloRu
GCCZYoIFTAuQcLWLQKVkoms+NHxvBn3GQofoouUiWAYEpWY2/wuz690VLNY0rrEB
itWe5M3O4JHE1fRuOLPA3J4LqFVs3n0Cs8/Y1M7Ap7looiGkiI3FkD7YhtzcwJW2
aN5oIVoP8KQG+7sf689AjSma3wxGgE7ElXitDTM31hdYInqFPCz8QMP6KLshOcC0
46TzrPlOgpSgoIMC3EyC+iBaATAkpJ7Mj1/2deZFlXbNnlqn0sdEp4KR1RIS8WAY
ZUu+03AWsWIrw3O3A0tWTe3iQDi5fi97SH+d5/EK7vFAIrHTd4uDZ5fqLdN+88po
udKrICpIbyJDtgDKh/tKwkL8/xvGhx4F7VhzjnC3bJXvhBABo9kjMekQFaXdQLCG
bGLmxyZXHFfhHMqKmY6JiGVGAb/kyE5KUhiMcaUaR6P0c34bdP9q+WvVdZu7TgbA
lds2Bi+eou+yp15wdmmtl9yISsGJokyPGBxUEiyfRyFsOJAHnAFgNiwDXaJHxI/6
9eWAW+h7blOmHM/FMPdt8oO7rLcm3oQCyQIqgHzw9Z0buKFDHC0ufaIArddzmJqn
z3lRe7okSBnO9ivHPGFxscrSCoosHz2WVOS6rEFKNHUMfBZuteGsjScbnWhpodyn
GyB0HKnGTTJ+9zgqvexybgUwlim2/txjwbFxdKObO9KuSZ4teDDr6ot83wNTbyCX
ywjv4IWxNb3+wzrcLrhJ6Kzwo3Q/6q5rgUviopEaLDivfw5p/qpanrQNeEBEoL2J
d7yVJH6/tIt8UJmmkFjTdpGMiSB4iSIL2/S4JYTFfPc0twAaPuiCTGlEU9kRKGA7
3uAbAUR7xd1j2RuBTWFynh3Hhjgtpyu3jpnoUwmb3gVQEZ/E3k9wwqaeJwS8TGmH
AlTOgzlMpE0OcAX0XmPunnGlupZHpAyO3nGId2HchivvAfwTocAotAqtxkbo1nfT
NX2B6WEJoMOztF/Cb/MFcQvFd506Vq+fJjGNE7zqWE3oXXHFSEtJ8rkxPJ0u8k/c
6uHOvU5+PiWH+yHlvuWM4Iv7ICD3L6yc2QB8xDTu8ojpA9kfkYirp2FlaK21w2kL
ujUXEY3Wmo1DctEMSyNlHsAuy7RKRetnNtbZLfTbQaE3sNJpXpJGEfjZMcb2HGvp
sIogdILVA7/cgU24tZyrA76NTjltlmyvOqS6E8q6/t1pIXzDxKOa7NztEwAcB8At
CiLE87m3s1pGxetdBmQH5uqEAs19BjL/0SftTnSh9I7z/Zl4cwO0n2qxk8qUVqpO
8Uh3TzJS0R/WsB9TNY9orK09Ax18CZmzrFagS54PkbQsP1sxruoFZ0//WyGSVuYw
HFCgBHdd/zeAA+jEfv+G7o/+6Dhq/oRVufTYr0woB2yEZsrBciT7WeJegOgVhdFi
NH67sBBtId4vDSKIa8P3ys+e0VUcsRT6e/TYL98Pk+96R/uGxbZ3R2+Tj7vvm/Ng
HCuhK9UcZQi7SQ4t33/5nAeeG63nKA9NXOMDF3zpxCw218sU/3BKKxMjA2BJspvQ
sygoVJ14Q3EkBw7YVufHDxIpgnyu3cJXEBGsZES4YfbgxsL2c80ilef8HA007jaO
nC+Zm83MMtEQnF4L75IvK3VSAkrWeC3jyHUfZaFkgDiLwmjX67y607tPPc7weFGS
mOeAt3CWa2IUdr1VVIq9Br06IX3ZjdoiJK0XZ70ZcmSYZfeaxFTuIwz2rZhM7b0M
SsRXuYbk7U1JcBEtobVXY9A2NsYUEJJIginrw0VzVq6QMkYIUuxZtmM5hKOLuHzQ
EAO+ZGKKVqm6/iUPGi/9ULSng+TDUbjCFayYDInQBHdNEVyalFVTf77GzhBfc1qM
wEfVhlF3lHeg6a0EZo3/iu9hmRWzmoTImN3B3e6vM+t/G5DXyao3cvKANaWnaz8j
bSFmtvJRVxrXOoHArRWoCEp8gxAqXudnE/e4Z2cTl48lY2ix+rFNWiMZKRaUdR0I
WunthrFnZFhzufyzFVxWF5kNc1mUZnPi+H68z4/yqiLTbEaTXX64zjx2YNzLWqAN
KRnJMAca1UFza+XIdsyhZst7Pyr3eXfd0NYN/bY++SMlb9O1N+ochlZvfWGH8Eu0
VIaroccM4EwzFqRi5IzYH96Dyz65GbPBOBZOmZTdsSMuA/8VVsyXiZLNKFxse7h1
gW1q+XYA7g73p2W77RoDeEvzmg5MuNiwns8LDsV3sMpPQpdRxnIbKqPnyO0HyAkk
eRRQYSPDxRiaubtFG4/liNcLLQ/UNY8MjuG+82IUA56GJkn+NA40Txm5CLSxE96X
/gcUp2ojGEjAVtsTmqnSznCX0IsFUeHDzvRp7LN7YXAYp70mcHNha3EiaGNscEWZ
vR3Wcd0yJg4D+3aOLzunBzPPO2W/eYWqrIoANe2Kbzd2EtcRMZ8XITh2/62/1DDA
yVi88ZdjqXZYdYa3dOLgGcLN7A+1FDBKyXDl+c3qO5iHGCgGL9JtZyhjx7ZrINOb
jBoCdq+ZO5jkeWjlMKJlHp2AcxrRp3phgTVO8wxmEy2Ij/Jig4LhAWvRcdxMflln
TJcPISp2DKcKJjLKVEwsYjavurJvETqoHJz5nUnN36DNPIypMfp2M72IXS6juPK1
hMMyu0fkt58Hs1iozAoPBt16D9ApCrdsCOombqV3PBJAyV1EBCcKP76FXPFnsAsg
UylVu9p+RYh2LU1D/S3TK5IEysCyF+RzlkmvGxv6z+X6sq1CP4ro3yV9NMwJW5mu
XUk3wpXLz4nnAu/ZsHzZ/I0ZGdDaKJhOu03NQZub5MyAMCmrvjq6w1Kmy3XvYLgf
1V0I6inbVR43m0i/FmRoAXpWFROY93kOT6pTW6/AeTljyI9xn9CmQcB/y5nfJ13u
HiZKZ/mN1I6qSatLResN6VvvCUrbSaB97iHevSVYSGF8A+qM1OxCS0L9SuqBEkWE
JQAgiR65bpjLlrF2L3wN7TUzd/AHPw2kPnu8Ho4jzZ03jl0Q8jZ1lNA1YgZQZ5yF
JK3UmY6VderKRIx1QvVAp38WUW7ojUwiR4YJ3U1Mshl8nwXrn+UpxfSnE3uCa3Iu
8lU0CxW3QbIMXB+RGrC+feIajJEk7TymabUbVTZdsscvC7N8/PV/d6VN+0Lfmr5w
F3Z1AkOl+VH2VmJ8Z9EG2R8fbKGbzTZo3pSjkHnBKLwiCgVoIDcmAvgcWDa3vmE6
rgtDkaHz8FS+Tb8WrO7lzP3j5zXMbDuPsf9SlmHBe8K0C4ODkxey2+jVXGdIJ7vx
eajbGpryyywy+IfJ95p50swUp2TXb0mmXF/9CQqnTfiSoERqTmKxAcP8OlDBOFem
YptCnnq6OkLVto8EjHk4UxAgZhwbVtaPiSEYRxkKcsr9Xf9zj66SQVVNXreVOEcm
MvCk87m42nTdGIrbuIHz/FIJFXLOO5YsheOdSKtzZ0Q/rUlgHsnTg/C+3zoy3mk6
Nj0bjoxQqL6eA34SixApRcQxnyDVNq1aBEDAwtLQ7KKTeMcIZ887JZN5ZiqBVRE3
Pc41YqUIprZWkxfTykdsXEt4dJbFEgDM88YBBIycgy3Fj3zc9/LOMG7TlOtIc8Ao
u5wyA4KFlGMR3+wF4KDvy39SSdi/IAFaSBuIeB0xTJr/80VkiHWJKyBdwihE84kD
cxB+NcHSi54jhOP3U1tkI+LAinuzeQ+a/SmTqppFKWcvnv0/0qvendgOKnI3QkFG
FJhyoc0vDOfXVzuyv+A5OpxKcBXfJ+H8tCnPOX4dJMyeYnKdm2mbfFZIjKLt2xM6
EmvNko6vo5R7OzKJCZ81iUVlw2C5tCLr1GQmWwR/yzflmmtjhD6Fp70J4jOMJbgS
2chpaN+Zb2HzD4e00vt7/gubd+xaEL99vWYpsJPQ+J6t7dJ3ZR2/Ee6407pdevAi
nIfgJa2LWQuvL5Y9BCVRFeSqS29g6ZS7AZL9o4WzEIbmyXRrDXnaGsP+0CIdDdKF
hctXJu58d70Pdm7k/Gc22EPQ1ruwQRC7atd3X37USWV/c5fSQBY1Ie+BXgMi9XyY
zW1dRu9LupuAKOCoL96Tg05yq0YNRYD/vgYK99rrzibckBvnxJaeEPcejyph+RLP
MG80Ck7gdQbqqQ1PIK7HN4cOZH6KUyjNbKEig/LEYnWiGS8xZzQoUNzciUVVXD1f
hXPwVy9G1rid5av74C2FT+bArJFtKTeqjfTZ+AUGjjhaPj2WNQ6mh5aVFrsDnNGn
buTEXv/LpCZ0dIUqe1FeN5ws4KeTpW7L7F7Bsi4+OprPA0O8613LL8hpJiZaCB7J
SzNxOqVnon+tO7Nrxwox4ENapGcHYJQfchO+cSCgq/2HNl7W7BNWADD2jS4GIQg7
7VoDz0BSQMqppAPNjrxOsviJrcCOLLGbT4EFAZ+fWhLNm8jmwnFFB/jKU9jEyiDy
99cKf2xSFjwnuwhL0qpfBh9Q0vIX7Ld2KLKzd4CgcEzBIscx5RUXYYw0fbqMMajD
4tXfDWYelSzYR2dSGg48zK7VFHH3AwBoPzfraNbFOn8adVvmAtEOLx4ThlqQ7Wgw
Lu9dxbi/HjRo5wvv7zbImX8N3MHtqg+UlwU9+K3ZZxlCUg3KYYbT0500UJ+4UaNI
zToAtkwR2DQVbTZIG4fEYVBZMVsHdu0XuKHpL33P7gladallBDWlQGjDlIP7oPrI
z7wkY+B1nZ6cTYgmje6AEopGOskhzv7g0xsKBflnsB9B9TxUDl1SqADa1DmLFsah
6JVHVBk+BNKgl0qdjOUPH0q7DXnBLSaEFgVt3RFlzIojSsWi/63cRT54NF1PS9fk
9NXBzyylsrRe5gQXyDVM6xc2N/I1CmL0tmRqPdKPZNr+6VPEQ92mgORb/iNHwoxJ
JTp6gWpbSIZ05kCemkxkT9fpR0C0X/SxTkdrHkgIBICkhi6yUaxRahXi4hPz1EQI
4W4AZHJErkadHys5D9iYXMZtLLZHHvct69LN2GeJt2FFga+AXoUAX+plmHEh42np
hU39ifn17kR8zQbfGG/Jb0E0i6WKZeYxqHERwT8ImDtq4WrvIAuJDFj7PtYXlbr9
I8shdbUyaxyvT24tJbjseXy827Awez0ZCz1kzWk0QKlvDGdCio8JTQc5u+fwkiIr
wNDrIbrUvBkzqn1TTiAV4saWcVY0yQU1Dh3C4ty3xBx6QXBCkHTkhVhtD+0zsu8M
bTyemLKWCemGynpBjszKZeHWCEFpnQCOadZYFV+jv3O7NXcgdlFmKALOAwW26KsQ
lb6aLoVd8LDgDyuDuaeKKYPboo+MdQSQ6dFo/cKlrz/BrwF7cZdZYoT1A9uhJerF
z5J02OM8VjZUTUXYHkdf+uGM7+G4O9IHlWVbugihNZ6ncsv2hWFBxLO75K+2JK8x
dcnbuy53/vyr5zPVcq2pTQsJu0lDdoj0UeBWlp84xICCDLlH7/42lbi/twvGhIG6
7IoAks3FMBKT/1MIyj9rBh4YnlyQ7nXmrc3vTH1HUM1gCbdbx4PvvjCowSI6VSvT
BHId9lZ2XpOXAIfXozXehJdIAIexc17NoJqaVzhLf8Z4D4Zez/gCEjjmDVAFY3YL
CR8aTzTYXp5UKkYSAs2Azy1xMal67qBEj7vkhFk76mWYRawl71zXO6Vxx+vmoaJF
qDsIQ0FiGHdQrdOoUVfJx2sKEOR4WiEqXxg1TYr2Me8Aar+W77D2y9nhSFf7D77Y
bKLI4IK6EF4ThtbVIBph+5GidjewMXFoD2sSR9C9XW+gmhl8JYjgPjGi0O/pVIAp
E1M8Z6UiGegWUzyOGmuwxiI5lAyvy6dY3eNo39KhnRhFJkUFZ848nILXlbT2J0Eb
P+NKhzD2eJeafOaNIrES073HB3gxqjXwOtpBU4Ol4rZzUdfy4+9R53rs0bAGu87v
vhMvZ5JUM6iZYtpCx45yeFG6t650VnIzVDIzTlZDKs54qUTVecTQfQ7vnmZ5Kn74
POQcOWLKjd+X4z0QPTuMT4jfOAmqaNr7KLI37/E34k3BL7NyepD0M1hKSd9xpyhS
4N6ecKW2KD6udvk1BuhE1wsGf/wXX9KJJsQo8k+B/51p9ePoBDTtP/5luywlP6Mm
7d8q9vLkvY19HjSC4fNj0yS+n3ynXn+uSrtfO7ZhJGIUgR3deqnHJ8ioS1hY2fxu
T+jw5ejp9z1vC1T9oYsY5tr13V0ZsEBFEFe7xR3sIPNgOrDC2FpjpwvH4FyC9mER
YXHy6SrfVGr9xnnhn3n0bMrhXyQW6KrKm0aVcrL8xhqUUhtmdje1mxfCzqBOLjIQ
2mPONo65W3GdhfnbDEwfr3coa/ZS3NdLghBrvB2s9Lmihwe4BkGBzpzXyAtMgN+t
iXDOrAlA912jwRJp31Kh2DBHdv+1U03nVDw5/7UwTnPLIwfEMYYtB+zzKX34jFjS
ern5GEr5NgB/Y0Wwof/mCjnaRLCRTEBp1NspokJM6RrEanWIllWpi/Chskk9WzqL
evqX2pe4Lpsfaxn3WXyIFbyNqrrt8js4neN4CDrvwCnb4tgbLSYEzBDebqdUyAca
AxYQj/y8/umdu9vROr3UBOXvfIP42pZJIm+sjve8vavIxwPHuuTaAdp3aDWTNj7d
PBkJtbTKiCYPgW6lZPrgJqWYj5HNfHrrogUdPsNVNhDS/zu8qIPWzm7QxYQ+jh/3
6qUlxL4fqJznb4K2fS4ghHSuKjCZQSEizXOe++J2D/zIHKA6MNr6/cQHhk7wAkHj
pp8dZnOIHC/SwYKKIv984JPbxwC+Znqx8t/XJVaRwxKPznlcPy4Y4Ka71Zx/n7sA
saontMbCXrXNVzIrLXhxSY/CGFHki0HfOmT+0o1zOGKzJKpsDFKvbhVlDcbgeHUq
6QbXwSuIchA/YVbybr9Ny+w+y/rw5dadohChZRklsNc/IE4GNZnvmq+CdhCIFKwZ
db+fQfHCFiEzQIJbgDUgJaEyX+CXzqASQFNO+fyTkBYHwmtN3WF5FPoJjgv3WeC4
wib1HFbHL0tf9RKkSDCXbN2FzBTy8nIVreXWscw8Y83gjo1cPqAinwsxxM6ZL81X
AGZSAu9v0pw2QY8wU6kHT+3AK4OtuLQp2m1sMAp/INethUxfD6ju1zrvd3vgp6dD
2sBRpCpj1Yo7HC/iozeibaXHztPFby+3MD6d1vE65zB1Y+CVCAFTNvzYQ+facplV
OJDmZB3Lo1O2XFu2z7hJMF7T8o/YhF3f4sAh2GTwSNAyYxQz3Zl7yEIQzKbQHen8
kZa1+bu2tY2Ek4Hc9UYKalXaqRq3voLNIpFlpSaDBu4jyTTYwNZmRNGiNr9p8H0N
LK8qiDSXqkYSankdbKu9EbJFaX72P+My++rUGS9PrydCgRVA4uZVak4GXU5MhTTA
5fYqb2f8V98GMXmj6Jmj5CJCiJlV6jBIZvk1ABN55K2bRYKTd5rYyGqiA9lbq9Ln
pvIahDOBnRpjNsqm6M8iX9C7GpBi9GO+fM1qERYzOyihJBX37WL1ZwqYRVG5Wp8c
XRh6WI8zzFUJqLc+RVXjC1aAn2QG9jWy5rOMsrWcBXf/wwJEvbXbNp85ZU8KdmL6
IlACR1SnwqsMMaaWZ8akGndofScK75hARdZo+gK23zq7WOMWYh6bqXxvyrZaGMy9
BGVkJVCFWtHAVbgeR4XVn1x03F/uBiipXS6ndsU01olDIqSsienyh/DV81Ncr23q
kNzDMdght3BilzM3UbwDUOoPNWTx7Q92uWjhJHnHZbmKDS9J1CbpCNiOfMgWMszg
BkbaIF3PbPs8XK/p1DgW1cYfS/q8317yRR74LxXQENlznq8wxk2Y1GTbfIGCPWz4
/VdnNmBWydAJBnUXZwbvFoCGOpERyS1timsmFnPpz6Z9MUlyJKPw7Ie7CiKUqU88
tehthVFfwMXXXHlLfi+DZoXxpR/N1WdPHfBvprgT32diPnhsE+M3cma/gqFTRTNs
clZFQ0+BMK0TZ5v5z2dYb8jONxUP818BFEEpvSD4xVx1hlyyxVytlWVvhoOImYB8
+TsxxfhV5vUo+11ZWierBHuw6seqPq0boOJ5ZcmnVcOu9LfpktUCPDraOfTspLnx
9GDB1Weo7Qhw+KiSM41eWE6V6CnBN3Eyw55U3rztfU5SWR4hkpjO7pN8+uqIQ/8C
c1nHozaJfHk6E2mHhP8spYJAu+bIuf6m6Q98ry+Atsrqi2mVDFHLryzf+miak76n
ZaXKCgwB1TWZ0XlVAO6rXoikmqS33PaBmKvWk/gZwBVVtVoxO1UyAfuJgs+5Au4E
FgXD89kZmsXOCS3UsP37hBBA5SKakEolD34QWUm9TYUa24qc2Gjbb0WcSrW+0u4M
3U6HDkpUoxUFSMNnGcrApLhcVNLxffAogB7NNbYIWJK+Ptfazo+mYWN9YgsK4jPT
+jHOl3KqQ4xHiPqbftj/L7WBR9qBAwwSrbifBKJx4PgBbUCFbEDiCOlJmxpiG+1G
ZhN3gaF38YzWQEXazXJFi0kSCK05TnLRD092Sk0KGtZ5z+GdEJbG0P+4EgYUfEzp
KunOkoOQbnC2s3Mq+pLL6rPfMxo3ZrGBE3K2LjjMpdGWiGt6StV1qmuofQkpPuvQ
eIbq8Vh26TKoyaN3l0j+tluECQHyUxjdliJb0khmWr6+aLBDGxvRTK+Wus4jcZlr
t57RbY34upBxZUXD3zr+l0H2XlUX83xLuhDuEw9WNoEozUQlyXGOyMG/n13IsIqP
SOfVCG6RKvPmZWzJ3CIhwPgVJPY2wPoNQpvEC5xDJateYwTxREfn1TNtUC82ZxNz
xlJuAa6ysesMD+L+PgvBxBc8IX5RN5aIwr+FgB/rjU1CCIG/zAMK8uHMd/MR/fMA
lcuVO+/bDIaJgMo2Y/ILiwKAW/SZIcdgE4tLhj9/g6L1OIa0orHPJWX4XjL+bjg0
TC3AcDMBYnlgqpWWHhK5i3hCBbM8OUVhG5R2S6kCBJfp1PEKOPQ/vsJAVqJ/sXAh
JYU3KwMMcr6xJ7eHADuCzxORkFimAV6qQJbVl04URZce6tZzG5ejlVwm1eFCnMa5
dMmN3Mgo+PTS5DngWhGFzt2jWDyu2X7pIpjI6adKG17+jmoLfDYgpwrVdVdtNv5c
PE+LS0EKB5FXEvodnshlFSHv9DqVjJzbtNDee4Dh5WsioIzCFn4FBHa27uCuN7lf
nftz6xZPe5ih2WDxBJX0ntbx6wtkS5JA9RooEKzO8jousURNzoq+mm6/2BZ/esmZ
ykHdTX/BOwneGvqkwliDHgVYU8bt5DerySKowPAJ3sDA0D1unhumcmSQeNf02MlO
Z4+P4Avgu5en6b7alblY7i9kiMR1qq9Bhg17tx1jmlvkeJRUs+JadluL1FhJPcFe
rGsJUU0v6epr4hWg+YBQp3r5J2tuLoC5ql4icf2O+xEI0Khyli3DAVKGjAHnpTtv
IkW3hEnidjNf7+VJidKhubme1ItQFNfqllbylyZOiAUAsUk/epnEh4zIp7tykRkf
Im/jnvgeQ95kNhpJjyrkZ2JdG0Io7ybNM1FUAM76U0lyY5t0qo9HyZPMG90L2Y+s
Q+K2Ge0mVuOfy7uTIdp+SbncGfmnsOKtNDUclqfUURBANsoD/FZSLZoZNhwXvWS5
SzrlDWI2MyYuDigPqU0apkQeNA+yGewSQAZPcQK9gWm3Tp77/EUaXZfCASMymdsr
6vxvqC/vLYzWCNQrnjHDuKCsPog4AbRgtKoQocoLgR+PEb60+dxlD16hY4tTpov0
rYzvwBCDRdc3NsVPOlhBgPAaWdgCsoTuxi3298I84LtMQHHsWwV+iiW9JuII1I2i
bfe4ukIoewJJAdxiKjF5pvXXHxvxAy2D7I7u16uQ34GAch4+86b998Oya/6yKHcx
y8oTCdwxEW8DbO6ymwRfJaDLRY8C8s7kTlSLbwPp2oa/30DxPij+GcN0gTw2b+YZ
TijHgFnrfwpt76UItPUaOLrOJ6szSw+AEtqdrEqxeSmJ69DIMfG9D7h9AmKlDuQQ
7IAIyLrW3JYSN55328DDcaH4FQvG78ohcBptM+oA4lQlRh1qtQ7608vrNCHYc2KF
7rq5WOrz9BRE48WgFLnB+154K0O3QolYlTf+OdmUM4qM5mpr20wei+K8CEvDD9qE
uTo+R6fuRYEx8FBaNgWD4E5OWkbGAKg2SXlRQR4FZpvBG/erD7DWfCSKHMfF2MCu
I5Z8wriZ/M8sH8e9NUOpKN4ZmL/by7ZbF7/CHlsBFJrlEBQPQ5EzRGevlE/jpSFS
gJksFdSfp0gZBy0W4S4fgPkEs1jDpzn/3F3hatXwqReHcvJpmlHzeze2BUV80d6j
j1KzCb9t5oz33l+yJ9l9I1Ok8R3OpasbcaPmHBih4IrbYXp38TnKb02z0pbzYlC2
SXce0mibDoF5Fau2sZNfdVqTOlDQ1ONSmGTu974JxR+7B5ivhxdqeyggFE3VHAvE
RQOu4w0BazOZ79Qzz3jzHE5WxdVYnGEUQFyJ5KbEYv/YGWhFAjv+lkFp0yECwWLr
3E++YcGgYCCGBI7rJB+udE4iX6RH1QenrPMTtcUXW+E7IMqjaPprWmqS+QTv+oY0
mE81SJr+/DADKdMZHpegSTwQZLLw+cothfMac9Nx9JDxy1e2CyUSqa9BgKTgWEtJ
ugzJ2TytSm4xXhZlqbpiHgSDJj739iYkf0VcKmEyJmtwSBKGpxhS+VNOTiBTh6pK
gM10S2qWp1IgxtlE4pNyU+AE8bNoXe7dx0X0MWfWL7LZGUdrN6IevuVwAE85z27c
VvBUPYm7Qdgds0yKoNV58KHb2jnkBN0m1ZWAdWTtyRdwqwKxr3iw4owmDo2yhDko
c/Hpi9jjU74Dd1RavViZEL03cC79uCMsIaKz0IYS3JaeZCny26NDCqUYka2lc16I
8NttjdwU2j5miuAw3b0x/qmYk943gKcjJ8Aq1aIZTTG/Ynp3yGMdW3eSM14Uh7bL
avA0PEmRQ4ajdZB76OYFfUxZKYzUwAhju2XC6NC3Em7tm5mGcyTGnwwuj+zVEwqy
ReFlPGm5Xm5yOT/xLtSM+DqPgMjrEhnIsbQd2FX6LOlLaE2GsAdc3nkkUF7IyZWG
y3EYu9aEY1HvwrDMpLrVJyJHSy17oYz0RWLzm7wk/1+9RZWfXq/32maxP2rNfl4B
B9oQdS7pGlk3uF+ZxNbCuG4wjsF/NP+oPN/YiQiuuyBo7KmiR9QO7jiHneNDHo9T
+7GuCbNeeJ+Evoem3Q2bwIvPJb6wUkA5kpNEVQ2kJC+nqkD4P87u3whQqCt5MdTy
+GtlqIeu8+40vlTMh2+G/owmqk0mAOzGC4g09sGae4OWQVQeUaPfmvUHA7LHFKpu
Iavdc+f6iWy3bHlaihQdQGY2RyvCiRwObh2skKHoWp/YIpMpOpmJguYf1RyLjxfU
Ik4SjzdnrLS3MwIU3hL76wH5s/P931D1TfYGtB295cAwhwm6pMjLPOQXBd3W31WW
WQDo/vJ6VCpvk9rGBeztzwpGKP57qhDUKKy75rBk4Psaf8u0Vxihz9ikf1N1Yvxe
O7cEZ6HVUB/c4oqorlNAIpfz7ihb8KEU/kXqDZAuejdsWlnKAHlbW9EgOw/M4lR2
rdbMnUG6OofuLYGgc562AEqQoia27NaO8KwMOnwr0wLmYomMtJVIkFkjaNnEAm/v
uqTo4Qa1vRcj5c6tfVJ1301HbuP4glOL9HVurHSDSnFmzfSo1EqA1iMhIbyTOQS4
WXnzDmed9D2jP54Y1mAEd3DuuAFYaO54TQrH7embs9v2fPjsR91b+in7M0Z9xg03
Ug4DxMwhhJ8IIrda9P24qgKw5aE95xhF9f669108Jgab6xdk5aDrzt8o5p+VBvgS
TYGESxtFvRZVI2+kbp3h536tE4tWFc95BWx5FsBagoKSZnIvKCQ+Sc6rfRd4u5Q3
XdYPsWMPOYkjaKA3HDruHcPqQsgY/JAcfEpQUCz0hCQ3hastAX7exgFLebGYYtll
FIqsoqOk9lhNqBMmWYpk/HLnZd8nBTQEETfFek+ACL/H7BVa0xK7pKXpQRDoPFkj
5xXUV6VH6XcEmaZuTea4A1WBPb+V/JCp2fDgDnQpqxUI76/rYmoyyHzRJGwkZsEz
ZopYA4idHEgeCzoIkY95PuXvOqb8Zq0khhWLz5k+91FyqIUuaY1urCF2w+t2yrEk
7MzlXELSOTi9yS/5XbF7QKDt3xeXbjG9x1Cc2pq3yd4a/PIVQRJR7s2BkfGT3OV/
hZCf6I9k02GZB0xQNx5YTcbbVYjm89HSsWbEWUqy6HCCQrC3fo6iHv9tf4E1avEN
Fb98deLJtYgJFw5zZX+yw5P8fPeqtw+OiNfbBynbXfbM794d9e7eVNTT0VAhlB66
CVLyGxPAhagsU7O8lo5K3DeQ0XvXSRFiXkNJ0EQy8IuaR2jUWMYrMXa6dPANy4Ye
+bbfX4L/8n0Ma4FI2zrErb4Hm+AxSxe3S5anm+4OPzU/JgMhRUHy5AOqubmnzPii
LRRWAJCj+uG4tUlwmYNQsBJO5v8DvZDGEzioJDZSwmZrIhrIFsXSn8R83WX335Kv
uPFlBtd1LD7fCokmH179YHXozvHC8Vso930nT3f2GFOi8NN6wDMoQjEhXUNdOosX
VNQ3m0+Bp/1U/rmzOTV+6iZAb+3XLqASmw7QJ+qPSgStDMys8zWI9WeoxwH6bac7
3FMcuY338UqTnqgjFymFr0AhknsV6N6cEIcrkZA2yNsm/M8d5gfV6m0jHAkzrSDd
jAOll26wNUk/rNJJ68Gsm3LYPCxAAN62SRDJSQE/SOAzuwr/i4X1TYSfkZmuITyf
26a/SG+jGx2dVSwSKUx0DQOfZ0Anq0n/fc0RDwXjn/K2QJr41QMll+N5VEUaY5b0
CkcUHGwFNoKeYYQzKfJicaUQPJlkENnH1QA+iExk7lrdWdxKTWWPIaUHeRLCk67E
VZIvV0+Ocky7iMdqijcRiANwgOdKnZ3loDWmhhi9Au95j6C6iIH66AWPQ2mv9CBX
xUmNks6kL8Av7jPhVqdNUkSPN5IcXEKPxByda6PN0KjTEeXGtxlPIO8UqiR8Oq5x
e0R4sIpMGnvHNj/cL/1ZI2FoIeT+gCtCYcf45G/ljED3SWr1d7ulvRL1LW/Xv8oK
NGWfEOZOAIyusunHbCV/GbDO6BoT5x9YroWz9YcS36uFqw0mTPnydGn7EYa7VYFe
Y8xTEYOqpa+SpsZ+Ab+PsYZRto3LAarvLQ+EhkmQwbkwOwko4/TJLxRgQGACqWX6
SgDNeaGJ6rlTFu+4naxXMIvOK6/wD5YlDfj42o7nrLHprpYn0PV7DMfNLxHhz8ZO
B/Cn331duQyA6CByw2Wluej/ov89EtjwsnCZv0erLN17bqlHGZh6t2SwLnkKV+ZE
bB5sfR6lU9xUdMh1wskpiJutdxLUNsGWN735NUMMuiyuc7BzFx4ZIKF/voAhNpOA
QIFXAnDLNTsA8AZO4TcJcbgF2e/3J5jRTBLqNu9eEyUneIXAFpuecZ383zouacah
/Za5Xx5/CldThUVt6zIe+tMQKQF8ZzxLPovh+W/3i2EdjdSSGNwPdvECVCXP/2QI
GkiE+ih80xJeAYS23b/z1JKItJYlzPE7vwj1iaOVhnux9SxSR6Bs5i3Qt/sedIXy
0d+Iojq2BsK8jpD63VolMKUtkIiuKiXG0zB2VY7qgs8LaD+PNP5U6YlUTpO4jAlc
AOnlniyOPpb9u+G1E7vPwXqjo8DLNtogpIdaxkkdIKLELcLW8ZzPuDM6+O2FZVxD
JC+erz4Avc3vKQetS6+LKqGdNDNjPv7KbZ8/4NBzoGEcDBDl+HdIMRrFE06yK36b
EC8avYUZCOyvfRyhuvwLQq++hEFcxerRNXxlnx/g4/+qha8fYUS0DAZEWiIQoYfx
chkkZZbxsMDULdR00Pog3YNf42QaajC8YNMhnHgVILhJi3UPkajnEf49m3Nog9h7
aJVobm87P3AO4VrYk42OY+kU/CaXU5XZ8/3LNHw6o+EdZgc3XN+ufZblqUZFFjzc
IqpNkvvIeh0U5qHUmSOIWcv6eUEHxK1rB0wD44iHiQHkqBlqNssvGb915n7PfKka
DeWo7qTa0Q3N/ll4qclZSQkc6DRjdFkJZVklThWNJeMEBcHaxfNaWvPy3GDRaUA4
3RR6r8XCdrMnyZ5FVJ+rqLij8stJTB5F5iXB0fn7/6OFqZ3fuH6sXRIAt4UZUrFR
LyT5LfOYttF9KXsyYSrk1bB49l/aoU6xh6ZKjookNTyg3NJ2HU6V9WqLJ4Y5+Nix
5HF7gmjntEI9AU1tWyrkoymHknJ0EiLihp0es5rxKF2klMkpbFEYXf/n8Ex3CaXm
pqhraGg013ylSxhniC8xL6IhJyW8pYH1Lk5N/9nr+g+81ZXqUdA8rCZ+vdnNAS9w
V6SfS8k4aZyVh8R9STePRjqhM83LZtttVej4n78cCc9DKcI8MIsiHYBzR9J/uNvZ
1wMAhMiqyzIcOzCYM6j2Y9KkhZnb1285Y8DrM5O0eckbgLnOJPPoUWTX3IgUDc4m
Lgxxu2B9JlEh3DUcMVhCoZdltd1pKZoaWYRGVO6w6YvyBFGURIW6gjpdShPFCgaI
uDadZzc3KPpn3oGslI97gp9sj5UuywsvjM6N68XirfGfA5hLU/LjLFb8Y67bVBQD
FyCNgybnvhX2X8oNHE1ifzbYP3oFMQk8rCtbkdcnaeCYK1N0CE9GPzry5Qn4hNRY
1OGd2+zRQBhdPnzP7oq2++9VHdGj1ZpGvf2R19EkTTEW4UYHaleUn8y91GNIW8jk
hruCoVG3c4r0AAah2Qnuo1W09uL7ZWAkjoYdOHkarbEetS0rVp8njthbTMxbPdcl
gh7arZgiXUh8qdnN2Exs5/gx221RKKUWADe/QXJ68QGmWpFLj451S9lGeCAMpN2R
/pArWE4GrunM5S0+O8pnFGWnyYugV9IJjkZEmlxYEyyLSuAKY/rHog4onMJQappo
+c08q22sMnVMr20zgZ8adt3P6kCxl5RhZJxoqXvyah/sBvyLVmvKK8WcTaGYIXqz
ufxGEP9ZzQXLZoLPqHS79d8uuMR7EgRkAC0rk96QApUwYtItV5uKDs+eM33V3jqC
NQzNQnEJf+4XkEgKr9GbYHyvftkp78sq5m7JrFlK/ASXUn+ig4VzowlkvL5NhDSm
Zj5o81VxyhVuw0m+xd35X1WYyUqWCvR8X6jL4yMRY0rL1Pb24XGYvl88mSIDpfrI
DKcA8UURRptxDjLF0ScNNqsI4SxFuc2N8yVZV3miw6dSmA/IFS/f14yADHF3Ntkd
EZbGmQEE5SsXmFrGaIt2j7LVOAneIE7FHb2eCIgLSWAujrFEMlLZdpF2f7dv8cmD
1bFNuKvaNcBI3CRZZ19YlC9noNfpFwVCvMiQwIF5Psft0a8JcypgHRtlJjsKzpgY
gr5Z8V5J0imLOb2EoFfX521PA7O/vaUBHBNiKRITQ5i/OziZqyFBckUG4liI+DiJ
bg2ySbwp1EgVstmsVQ4AOV8uGOIsuN5l4J+nd1dJPTJYJBkFKw/UG1wo3zxZYv5R
RQvzbuw0AHuKpeyhn8PXlziaLUFj5FgRzTaAMu67iTTOx3BXrCJp2D+Y6yXiMasb
K3Rmrgc1WqRZpaBzLnRlIlgUppnZTEks7M6jEuIb2rSIVQI2BqnAkLJysutoachH
AwO6+uKCjptbtP3jsqele1nQLEgNyrdrKvt5/8KS7p0b6pRJm7ZRllQpwXB2xxbL
2HDQPddZ/ZZ6iOXPmmPWcn678Wy7yJaFSOa5qt1schoEM6t2XHRgywEnlRCQrVxl
idc4nsr3NkAVWAaYed6YxvLvqkDNLcgA2ia/k0xJJYBajuKPiC08cQK5z5GB6rJc
x0ItGaW9+Nb+iQdifcSvuir1PputqbNfR+5/AwAuekiHPEp1exQzPFE0tp1Ocqey
45qWkUL98ExjrbKRvTgU5PNopkfaXU1S130hyoRdEWnT2skbl+nQvKU+TtWRrB6O
yoycykxhO0JHkw99ypdoY2+WFYGxKMWjz8gxVun6ik+TMfJEhGDEiGOwgYc9QyPH
W51JfHAyKjIHcX8ALe3Kt8cDFMAG/DbUN7r8M1mPFGQy7QJbC5M7Q76pJG7LDTJd
WXt8bgQHP/rADO/yGwpl0O3ozMQUpAx0ZYxALHIeX+QQNMsXVjfMfaHFjhwfPkbD
t0iSS3iFMxue7yof3MC30vUnji1bheRdeg9/z1rTiNO9nEdzPCpZ888n5dKkDKKF
dCmasBYE4fbD5F29rAHzC4ebTsJW375Qbd11FnRYlLNaRkoxFQCNTQUDZQRgPo0Z
5wy2lqVa0qPnzyAzqFeztc9xcM0ZWbcC0phQEZ8I/xv5Y7aMWtOmD5qmcUbhiBJb
gjx7VzT9NmxAzR1ESN0ahg2OdhepufgwrcEN2wpjUsrBM2Mht6VlUXRTwKXH1LGt
VaXiYTtGDTcF14Y577HTx9M7/3KVhBbU5roV9XLLeAIoFi0lfz/eFOs7TkdjcD93
8DVLozUCG3Jke3j93V2Hlztf+ZunfPVm1eEUIBMWo1AkhIrcINkZ3+MXPR6JOOmW
Ii7Y3Hpxhb2kdqiWTHZmUoLaCJ3e6kvk+ybsz/e+9JnDbZl71TItPxQntjhO4Ww1
qbnpnDju6OwfrIsSGQUUc0wyn42AyF7Jj5RDNxNqZ523MWEZnxaAIjyGmj03mw8n
xSKgBycapM89SKnwNnFDAo7IIXmudTuielUfraNi2/i11/SP4tYqjuaPABNLIJsS
0Z+EgmR7cLQ+YkEOZsIkXHjJmFGRc/9mHhSj6NAGBwzV96KDvarG+2WjmYs3K0+C
+UXSpJTodruCwZLyVfyFcTDGbwQtewOz+E17kd9t/BXxnvgRHECxYqQ7Cgsyu05o
XsSIJPFspvJJHTFl09qZbG6xN9qGYhE0ywhSrePJmzDiwT0TGfEFH+4a9FRB0rqd
dYP1Z/wnRFqtLxurt99bg3eIC+9tC0l8XVwLzICkTQ6b/RV9X0mXbcEs4tHUvFTF
43xrTOQfYOZ+f6GaR06N6SolM33Zevx9tVnd1eG/PliaJsT7paQwyAbgNQdJRBBo
VRzSrz67hBYLmJmnGJPXTCRGt2WWQ2/TaFhW3kP7+adls5eZri8mFP2FI1w9Cqlz
qsbrzW5YwaZlHm5OB/gKv7v3ergJOWDk6VAUKzTZnZ+98h70UM6ioFseX8yS8Djc
LtEUe4QIkwXjzgZXOS0sVlCjFOcvDVVWUMi9RlXxRmZSWuqy825RBHx058xlLQgV
t5vYfzSZKJF2j2RAbZmpZjj0WDyXHjTWNPGhmY6NSegAFtdi0f+nKnwtKTCa4qz9
BoTYm7+KYB5LgDvUlBfC4VT9748SXSOV3wOo1Yzup+31LOAs6Cd6VRVvY0xdrWgb
Q3vuNE70FZ2kMQXLUOnEPvLD6NrPcSyfYQgxaBQeclllmFCvNKtUsvBrtSNIf3p2
6BfMpjwSSQYQyFacOC4OftQ7RGTs4P5K6Xb4VGMIjNOaCPODnpSFcMehZs9f6qbd
qCmTXGEJaitDClLkLuAAmU6SyZ8yfQLtX9J6Mme0+kCCWO2X00PGr/k9S7cQdjcv
WfXi4xTfwnCjgOOlWR7GNjRWGYsG/wB0du52XcAVG3X1kv33K8wqiQgsLR44BY1t
QDY2ZL3FFxQlokiPx+oyjVNqy4jt1rlbYCj4nwCVukl7AF9bLHUMFkl17V5OADNe
NgdXkWCZ10YW8gmgopqIErZlvuYGuOn03Szre1twdFx9ZHokhqOk08haz/M7KdbJ
DpUp82Z0x7zrYt1TvGxYMu7oFBQ9SK3tegdIuqvScqY23Iv9UcKknJaaldk2m7Iy
XzXUJzy0VknKIbrCVNoRrkfUxOe0ydknVO0XcJiezVZhvztoLMd5xyZCtxzhIFDf
GBeRNoNPCjTRhxLIWpSvTc+mQ25HK3dl7wGTZmIw9BjGdBGShCiJBxPWouujQyq4
XEuIeQOeG10xUpdftAXclVMYAuhItTrx0WtSNDrukhuzWDS4yUmJ09mlKwNkdhYb
icjjj+vZP+OwRLg3oGLETDr/pmM9Yu9mvZaBIgYxBThVjLQDdvzdKEIlCk1q3fLt
An5bG4Y4tQ6vSqx70D1G9+KQ5bq9q0m0Rkzx5HifZmE4veVmNx+R5tG7XRg8d5+5
R0Ydd0xMbJvHuUcpBk9yruU3aVAisB8C5HNgT1aPOqUzRSJYC82G5jGmNgt+0GFt
jG1gNVhbi+1qU/8I45UPEvdX0qiu1gZmU2sBmtIYeYPLOKmJopcA7l0JjOfEYkHt
bbRZX7usqkDZq8ecnzBaJXX1/41/8mC6NYm+Yoy425t3u55VWiTcvp9t4nXx9++f
+C50TJHvtzsXT9u4RjxUZPRWlzZYdBMT4jo2d0dCtNK+fafbvQyJdi1a/YJ2lYaQ
MWJT3nwKtkHdZgp/bp3G83ttzPq1Q2PzGl/OfiYjdHgsiFwP2jvYQFzILSC+aIw6
KSG3XQ7LWuKzaB4CO9ut6yUfWNU1/ed0LULNyyVAqQXqb+VuRxtBp2blLyP9N+L7
GMQ1RPGX+EMvU/x7rc4BanMfUOdt0uEzm5gm04qEZw4RshIqAVV2hkrtBC2EORQJ
+BmEFdY2jjjx6Co3bTZlA1T2iurVId5FUntkQuRpqEHuu1VsGlQsum5yM6zB3Kbw
mybjC1+caht1TVfevPnYYGtSIFYOJZ7iixMRm4I5QqEdjTDAn2BfKzvAeCwrezgn
S7oObWyozkO9R31mJeToJHudao13TrUDTv60ou9cYTNhH/2qvCBOsZjRExDPFRqb
sbE0pKcWU5ld5PmSTPQTKNcKSrO6DXL8B2grNCs9ZjcBougrt8esx/17l5WdHTSw
J/74YxYXIIK+WeJ5xN3uK8c2VPoYdhuByWh2WaCAgOHJ3bdzj2ywZ+nwGryx9g9U
Ew9bFby0tOgLjrAGNSzHrJKLqR0FXNAAquQXAUZkbdiqSzS6mfvrpsL9ciywPM/x
/f0qdWQcYc2X4A1vHHjhscn8VZP3zekR/ARLIPeMbG0/EZmcYWCsNTYBXSSmWDL7
pk0xUUrLdozE1jQhWpmEcixB1LZL1y4sh5A/R01wIPSWfHzoRORzFSm4wvTMaioj
/bMQqZw/XaknGkUfPovbVjF7Ba/W0XA/jL97vKbVMMftJzPNo0WhaEmwmznGw4xk
E7P7jJWNDFMZXfIANsZzfk1NC1TbGVDT6/tfeuc7O3dqJOe5G6wiXcmIIXFm7QuK
5zWR+jovpdHkDWDmvZ3DV/5Tcw06fOUhOYOYaG65zMzNoYPcumPohM+5xDTk1iWX
kaIAb7FMNcejoT93sEoIcLiG41iSCnAtXQhhhEC5iVfEGgoTsdz7uzPj2IJtq9Ve
hTqqdY84p4Ya45nai2wvQZBo/Pf0hdzH+AeqDjEte021F3SYsQWVXrBOtU0L8928
4lqhnqvZFWJQae7uijHM+sf+NRMcQ+3KbMKi/1X0Xj6dekaoJTsR1v8A799+1ji1
BNArz5iyh0m4sHqazdE+uhBcrpxFRFq68OmKpc60chEZyL8lCfDuKKYgbzjh3Ehd
pzdeBPHsMdge893VeKcCda4YIBGIiOV6ZNLcfAas6o0S5vOfL0Sy0Lx4oVIGv/6o
nF4vurjFcTjLA8M2bEb36ooOMVBPcLAAko6W0iIv/rZBR7LUQb5uB1tC03Sz1oI2
NssyZBnwcmN6+bq262ETAEhoQtB0TGQMEBA3bja8eGLvtJpfd7VKpvXaxvqxWc/C
Oo1g2QY+YcXAqkX2Vwg1nrAfyxma1C/SgnLiyPvS1x21tt4+h+ni1Ip1K2ef0cFx
/a/z+yL0C1OyRABBe2DXg+AOzLmjVmzf+PgwO8uMU0b1NaYx+gkzdN0tx0Tp4qCh
shFjO5MsidziBCn4qjI9DKA0KH2E/ZaRgFNGbNox3Xb5gR9ql8nmM2eHQJXZA/AJ
ZSiedgI3rxuxLf2UOaJKez5xCeXLv6JOELW1LuZlevOIt9BRQx9/FZt69K1qxdXU
GvvIzNvb874cHE6u0wsz13vpPZ8AFADDkQQkym5l+oeIZTYWeZuq6uaCRPbjyjka
i2kjlZZ1SbRVen7skUeyImv9n0i+hqTvo/PqoGcn9WBqF72ffL9OI/Jc0/pyw5NS
fKzUwIY3ttolZSMuvn87Dgv8XWL0yeALS4zzxEoAjFNr3qrMo89uXV8QJbQ09ncY
o6fS9haxDoMFee64YNHwqw3xHZ825IikrkiwmomWM/KPtyQMvjAxz2E71Sy0B3XC
AKkmM8esJQFzV88abqZVerkWgPuoKYdMufVSy2ZDo9R+RTMw99NVzmFeRnoRijzS
lPwNMQ/G/ee1kxoz8HrXqRqqvXUX+IsZ9x89JRqNlvsSh5uwmgc77REZLi8S5MON
1Vleg81o1NO/ZsD4yG42ab8L+dkGChnSMm1jxWODbKqZVhr4YQg2ySbm76/YM5yv
eqKoixpUTBqzLEqdh3wmf2SfvKsPXhJSL7/JdfKpjf/FGgofieNInm6Qecwvr13V
BNi76zRflptnJXMOypCtnJRnrAqxI4dN7ZXTqfIrmwvdJSG8Bkf1RZR9zeCC2OLd
AOblmr4r/WJbtKNj+WpzVddJ0SDpOj1hrcXPVUlygZNnunmS5BA8eDW3N+0BPg39
7GE+n3kWmxO0qdcFR30KMxp90WZK0peX2xyVqke2Pt9FDvQZ50qmbq46CyFfe+6C
ETZAcP4jPK87RZgj0S1cmfc9nawB/9bj7q5wtZpLH6LkfXsX6j98uLePTRXdKrIf
JLTTMA6x0cT0k+AQe6S5dXyRISv/7pBmbMWTrwPJJRJjH9ZT7P22G2+HWCCqcwFT
TNMaVL0ii38bHfU226DjRg8NFASNCxq5/RqWjvXscFhuFJq5Wj+dAMzEBvzTdFPP
sas/GieRL35iWQg4UQK3ON9ElUxGxudfACWA5pqcrFF732YtEckETUWdf5XYBdHM
cGiKpUIev1S/rEPCH75OPGEoKq1/ueT9PENE4zCWlA6u2kwYhQ7KOVyxlazu3U8C
YduwbYU9G+8T0HGODKerXGeYK9JyU3D5o68Qbvqox6IuV1Vt+UeKoKdlS8M0wcIr
N10TzkFPVA3Y0qrwxbUkudjjElaF6DGVefePJFnMvZsmdOFeGsZyIAX0HGhz9DyF
8QTTKo8jxj0iPT8WWo9fLxAwL86kvzEgJovgSr9ELct1d13P0L4qVErpaIkRrHCM
CXjaJw6e825eODXGJQGVaqmxfJUgCTJYU9Au+gplo+ScqvLhZrh4CPVnFexXlUWv
dPpwhxsUn3nMHh9W6AFWGpzcYQ9pJOSjsD2hXpVgNdaB2F1m/4XePjzFccZzzD3Q
SVhFgdnsnsU6Gx+yFTqu3sRwlcVb2g+pP9pQrkJObwurlTm9qHjkBxvMY5M2wHZK
Tm6f6M5BSrZR1zrHC1lc9yOSyEjX5uJzsmbFhrjNBVaFrXJeo16SCA108w6060g/
k9WtXxplOAATpHbtqEMyo8Cq3ODZ/CKsMykO4DyKW9hCL8EMqiyOlhOfQy/ppVf1
cm7qSrXoSqnNpXK/z2Ryga2+q5hgCDA+RMthJUO02ZerSHHQfeg1H3zyU/dY320y
m7AekA9GfU+yOetEsWwzDBLYWQtowolGyrmaw6eyjGs3TBSz+7eSi0Ro4qyOpJg2
Fb4B/qU1oXUTfLthJyOrCOSrQV7VSYiAVT0ErWlNUkgwl9cs975lE3l51bl/RxDE
2Z3diJKTa10iXoECdh0oLstQ/hSPzuKb9jhR7pyI7RcPlnFVCenfuoRb+GgdK0Jo
RnZPKRoMyZbGwUWNqevrnvToISlTVfH1Nsty25YXszjyVXww1G5YKuaA28Q84S+2
oQenVKcX/nFbHR30eizBoo9Boqk3kIK0C9YZ9+RhjL+nUKvIhTuWq8w/jA2oIOI8
M6WxWpPxzdClMqMYItnyS359VxVuQpRHVzskgPlOKWP91hW/D3Vjs0ilgEdhWoUQ
nCaxlx9aUTkpUUjMNmXp6hO++j64F+dW0729goJMyuiVHTm3eOjwN0zmoJoP6cCp
xD3pMlgoA5CiRu07yx9nVcGxAqRJr4ZeXk1PRDX3Rt03ccWhW3PY68uTawMbGZ5i
EkrUgkgWEycltwslKRrOjCTmFR82H7leODybU8hByCiqkSXXKPZxMEpk2ostLolC
OAdqtxKTxSoqyM0kvmLa7uvanblN11SXlaynjSQw4sQ2Vvo9pXGF9WhPi9JwJY5R
m9B2+ExKx4C2dP5zBaQYCcqXlowvcI2+YssygW+X4FkUxaHtSnq49vAKdr+CVtZN
cO+D8HhxOl7jBJCeO3LhMlrR2U1RWzSzusSl3VU1yZMkPITZonxWKGmXIuYy9FOT
ncEoNqWbzxqUFV7bv0oLxIEJnxGsdNZlQmrXzqlEDYha+jGHY8CS9XN//Vfw1GWq
8KTJ2o2Fptnn0WgHkYCLgc4HTROtVyxY963BE0BzBsm4s2lVwXU+ImvLGeFTYLDg
oa74C/kGO8slespPUUrpwxDM9JXttixeoG4vXtyZs1hwMXOAADTcQpHm+5xu6Ydw
9ik51AXPxJzz1T6S7fc4bNAVVjt37jvwNc9/pyGhl83vHWnnHc3fHy+8qEHc5NZk
F1gv/c5zmaBsSWu+Apyoe5PL2daj+yuuibDzXWSlakdryjVQY/4nVrTSrWleOUJg
be5FYCiuhtAHcCJEENiHNauzVx8T0MaUu6WsBYcGaMzT2N/zfKjnPrpGhWn/OwdN
7Sv0ZS3Wre4uhySEUnGk6bcqG8m2NQes0nL2LhGNMQcvLfTlHFKCjhdD8HVM75f5
BPejzSt/GrBeeY8LSCOq64HZuN1H6spGspRXkHDefwwR+UqTunlDd3l1Tn1iB3od
vDO7r0zTIEE3bGtocVWIlqCmsSX8P49hvzDZdMV/L9FdxFODkqSFFBx7QUwqpmK+
CykRBLeBZdU6HhHksT4cuRM4fH8EdWLLoQalHbGMX0ex1STLQH8YKlpoQGSAP3Bd
WqVYcv8HTRlEI76U27ll1qE7Auf6U94S6XXBJYQn3NTscLvBIB2Pf/ot+d1ZF1aV
XuwevQaWf1XL+yWUKQy654rZzLmEeA/86279L7MIYnCA6+Jyd3uF6MPi+1Vop+hE
aNXntHhVp0nnnNBlfIxHRR+p1bjfSGb93ZT2A5fQf4a6tSfXa4MCuXwDOBry1Feu
YNmBNAAAxcL389qSuUB6htqYaU9Mfmh6YilbapdaywUSSinUKL+Acy7mOjcOOIc9
xjASDaK7tlkiPS7v9rcoaajCN0kg1L4ndxMq8L8eZLDZVGIGs/3bfEEpQdYUrGDi
rRpx417Ngy0kMyhBivgo50ILsmBUyGOnQwc57WgR+MW8fFutbZ3oNT5SW65+ds8f
EcTCddrKtuGeYUr+sKQ4f47/dtrcSV1grPUXit54h4pXKN+/1proaEBkaD/rWzEB
IT6WUcXAkBXxXlBcQdYU0YK6YIrMdMaDYjibteL+hnXA65meDjo3F3odxpyVLT9O
e5wJUNmAgsqb7HQstWmBoxoDUGwV935lImFKkKG0Gd7xuecEW3rF6ZzIa0LDiDMJ
dIXpp5A9PfVFffnNGl20mW3HuIVXC8dfX0U3J6/fg8ZR/CSG081iOpqHFtGBFp47
7PmkyuaXpNwehVGDN1nlL9gXvvv+xXrosvjQetsHx/+5U8QZxhMXyEd7CPdDTIK/
8+WBTwij08R8HGB4Ht4DtRsrGFGgN0108GkXOxGQ7n6pyiRcCfaNf3Gnqr6tXTRS
M/DUMwUwhTdtLgWMZ3WLnl7c/tv8HBeW8Ig+kVg01z50tWwJZm4cV4/nWlmH7bSh
o5zAeLSloEnCN0OPBEod2+MjbJUQu6pRjffWCJWVOdfUlGAyldL/C8CinIKEF5nl
ebjDY9VrbiWk5A+mhSM9t8qbzIMNyx/HEv/FCTODgwDzNQ8a0Dclpnhmf6uPsZ4c
CtZChL85RlzE6dhUY1KVmvO+jBO0eqGmA03MjQFu4lmoi6ZBqVGCZ62sr+qq4c0m
ZQFLQSWb0mVq0IuB/nA5bk7E/FYtBLQ0TrZ40jmMjSI9o5Qel6SQppOa9HPctmj7
MMT/yoQ+UsZEoE/rjAIwI5VtJNnPVF5G7Yq8zO3+gSCf+OBHlUGX+XwqcRHbX9A2
bQrcScnfbYe2sOn3cDYqUgXFh7Bj0G5eQRUYe3gcRmxSEsdOi85zcNcv0ogcr9Wy
l2ylzrlnrMFrRueMM06n8veN10IcphOVs3sfES9T0wxNYo1M1fymhkbHblr6LHS4
if++5kGIZooIgDCo32U5xjeZb24rjkO7EZnZ5IKi8bABrkhWKfdCuinODJv9Wqo6
eeSl5ebXaBC22aE2gmbg3mqMHEG/hMZGGUeBi1IHsRjMvYbZuszkC7jKDPJ/T6yA
rxLhhsyRe53GPhh6ekTYOtG0ZGEQ9CUE5N4Mrs3FuT4j4lqmLv7PUu9MFt4JJgIR
rDx2Zyh/Qv0iG844RIasi66p15lah4Bm0rvn+CkwskoI2c/GfqxypBBrXiwXisDA
30TOTMMzLrMvYdhQ6l/7723LXPFHCB1HQ/23P9rAsXnzLLl5vv6AqRblPrfgWrZE
GbS72uBQpoe0cw0QB9A7hnejYs0txMaSpiP/Iab2p4REgCzCdXRIemuc1JRX3vlr
q81IFkyClJpZDgIVeTTpM+apJXRNdObB3RAQM+t7AvFD1b4znzth/xEOF0zKwmTM
inwU3Yoc/K+Nk76fcp7/O/WpA03yVFpm/GjMpN2J9rG8rFlBNOD1TbEeF/PbNGcp
XBMS7452PqqbHLOXFo1+SK7ExMyjvQ/GkazDjcfHJ1fqO+COUjluhCc6fuv0iTR0
rn05z/lCckPIAW4Zu0KR2suv2prHyZt7XNemWnPz/BO4K9M/c+cqKkgLj/vZqSX+
0kr5a5r626P8wlMHM2dSCaZIrUFNMQvBdLLuIh5i1XiIdYJTjQ93VJxPPtqWX+U5
E2bvqojpVUuC4xJzAZDuJSHJuHKWdXLjPn0P37p2bjbnM9IGlqllVL4oLMIfz1Ih
R2yZPcpU89eNo/ZU5UrJeRvw5ygqbrChHwBBHJaAzW9j7yJwwr/qjuVEGb+BcpaA
BIk+HgITbNfmO1g77WZN+JKFIPQ4qRfeS0Rq/pGvCqHvdGydY3HJTgjXDoTP598h
RBbPFThMUcjFzjgI4s6r4aBuhP8oF+UwbfeQcbPos299s8HjI7rINgip0diL1csX
YVUP8Y94m6mwDwWJPUg5NHKc+YI1c1Xbg3JoePlmgHsaTeUcP5v/Dgnr37Tal85b
xUS0ET7pK9bcDrht0o4oGDJmMBs47/3xtXEp0y/3KSwWvU/zk1kNIWxFnsjY6CyP
LBKrit1bwQ452Rqi/Xk7CGeiBEBUtXX4p56dUb4LRkSSxqkK7yg5rdbGArZTrnWG
RQtOAckpvE+w8pqsnr43zhLV4c24du6tYaPsK9TwRO+u62j9LAaEM7zVTT/dRVRV
asmwKDabbfw8qQPS7PqIUR6VHoyPsTv4eCCHHXHoRSCR22FcyMVXwVT7eTdhBTBx
WOiJ0XTKm/MDveT/PTvOsH/rjUCOkz8grX20dBF3Gn1m0NDsNRrORnsrp8vxdfsJ
H1XAhwegQ7uh6pzx7+uc/zBvcHYQvpvtT9S4lYU7pHAvTiv4zcd9QalkYwqAPDpK
K8mh+lTOUArz4/WoRpvZr0rEB/CrUWQ4RfSo7nmcpKkNXvNgwE5VeX11jkGUo8Oq
qsXjuZY/LXmo9l3IgRWQ3fnFNb7ecd2CFxC730nYzjbQdxahHW6V2L5eefos1ISa
XA7v9zsX3E/hb5t7r9ntbrKkD28X2VIwqzaCZQ7Ajb29Qiktw652y6TVE+IU5jhI
eBWBXohBdbM5FpIVbtwbUP6F/PwFRR3df8205RBcopVn1xQMicSmvEYwiKI9cVXE
Spnpvpm3wgwAmjMP5JpQS0jjaAmAs/6Kb3ZIbxSYKfgeYpkFxsUphhEP9L1SinrK
C1bD0vETOZBbduAQesla38+y6k4lKyz/8ZKvShdNB4XRZnDZPqf1IhFejtZGEPKj
ku6N6sI3wnjpYOvReL6AKV4B63G46qpYxfP6y6z0jCqkoxsrfCgcGNxWY7CyZtS2
dNcn9Ph2GGzDF99a3n4WHY3KT3e+oPIk3VnCgZmDxymMA/Sf2VG2P69b5HGRvtk5
3LaoIuxIwRNQIoQmS15vmz13Fns0VU8yUnTXZa7dxYhXrYguALN15FI1NEBmoV+u
RRjyamTVv0RjbbwbaCDQA+FQU+59W2T7bIQtS5/3ZtJN8PjA0tSm4SUR8ygr5I66
OewpwqqV/8BpVL2i/s+WCA4uDICGObzUKoSWxKW9bvTVA0oVTaiGeFDi412GIjGV
hzihhZ0wetn8T9+vuEtSNAHLtUHq1s1BuwkauqsQWvKMGnbnRH1/3MRzKuGFJHWp
VEVnTtmb09iwvegHjy5Nc3Lo4tcysrh19akFVk1kUcNIiOTAVbACvrB00N1VTgX9
XZbQRSCiNoTkZKD9Jwp92/E9Wr3jIWdvxSxCxePanJ1ToUVeXSmw720DVx+5ZkX7
KtDF5J3Xx1WXPT/VQzXwTKet9eE4wAOt1KaalDUeEgQTQ/Oj5vaUe3pA8RA7ZdF7
0QoAbumc4TIuKQ2NmUw53qQ4nNWteuCdTI5C+0u/x6CbqU6tz46MUE1hbyfEPPEw
3g3/YQ/BHzKPXSVmTwhbup/LlRwquyFdueCoIFUySVpPCdy0dMSy7RNeYpUYGxcP
SA47RN2Tl7vd2dDgAwIZwn7yH7YtMu1x9IxONOl2VXHvOoB9u1I8m7emP18S2GXe
kgT4/en+djoQtfVaW+QBGI3QC0w6iXKVU1JCykmp47bm8s5dn2hvYvnqpYtMBD7o
ppp1FU2UvutADCBB49UAEKdBry3N2BBAqCEHkd1wJCYhgycHPPsbSC3oM+N9WbZa
0BrNrb7hPYN2uIOa40TAnC42Dd8t07hJIyuHcCHNqkj4UYMp/0AYd3bvZ3O7Zin1
9YFwrUmWG19QKfxOnquyKZETBFOAlm0IE7+e9joZl/1xMN//ToMAE+OYEPpUrZay
+Y0R9Xdl6kNgTgH7L6US6QqpwsPy+ESH/9NV80dtVh4hOhuozo9Ibmbg6GmV4Lc/
eI/q9RSR75xhfwdHdqOS1Aw0T2yH2VOqXWYcVymvy80sEQucyViJNuK9Fw/Ati2i
wCKR12ShOBCu/miP7EN/ZpnGCTIsec5/ICkDcD2TNpAnL5dqisTimyggON8jkWJw
QpZZQI2aa0QYVzHaPSWajE20WGyJtEUpen//NQPDOYrOcz+2A3pLTxUKWrZD3eOv
GId/t5rJICWCxE75MvKQ/+zcOKSuk6bLWjf/hcKleCD00wS++0G7mTa1D733K918
oZbfKjNdWviy9uRr0c8IMEpghQZ2Pt+kknKyru0BvQY0pB7hj+wTZbQ7YK+2lRfK
KpRawok3hEfPMHt2zw/SUntJX9kiFtptZUTnNVjGt2BCIhQe1WnDv+TwQD76D7nM
yH9qIMX6tZZKxbOOySb9W3UKOprcP4OIGxHq7wMypRgeLgXa2A/lMec8ltWbBdGA
SG3xMas4F1E2dmMFzhZgCnKn9+lcYI3F29ws0Umb6DkKTQOkM43TZfp0OcB3pUv0
ysUMxPzB2CEGvvguiMFHGv6+Z5zgKqsiTlTN+0DtSADVceKJ0w0cbhZS4ZBZySn4
LGb/xR2MoWKHOO5mjdwtcW/YAfCo3dnvP3P+TOwaez8v90fA5M6BbPqRB7FsXQYr
9KoAgDeKddjNZp+E8ED0TUUqIQV+Nda/sngAgTQNkrEcAbb8FycOKd95SYctqnP/
rSM6i/gNi3WSvEtfWue99yyLiFAx+kJtZgoq30t9hEdYzbUvxQyygH1Ux5+ZTTKD
scBOzWq44wxY+qlWwpxHn8SImkaDdr8BVEf1jzNmwqHU1KjG6OWaKWvvJdzHXSIV
IMkpdP2ryQkGreY9wZOH7pp0mPBSJl5GRz/pWdyhb0QbbCm49KG0wS3x/PjOz4j8
r4Efa0RqSZEn7BtsqbAXrNV4mA0xwFu+vTMXlQA0s8os5NxDBUpLMr7ENF7tZzKv
zPAy5I0aValN3pbf+WCef/9SZYwmp8SqG+Xhh3MfP1MgGGxk//uw+/L1QlZv3uuf
GrZlRXmFe/4caxTd3MP398LVzRFDM2VzhVdQ2FGFBV6wlf94aoZszicIEUL/touC
Fs3Yt4BFO/p2LrgyZfxgejUPQ5QVUWI9WJo97fVHRFLLjgs+HV3BhKPyHiE/Upob
FYbzeyaKIBXHB9SFgMtrdxJcDGnJinc79jE3uQ6JqDZOhBd1vP1vexkS72U3nc/7
JwF4jNw+RhLpFQZR3R+3xO0keftDi/tuSGjFRxOxvuMLGsyth4LCRMeGv6RzBu8/
scHlxEZnQcRC7RMjorHvG699iC2mo99uDvw3Ag+3bigc2VwKuFCYCMxVgu2Iz3E8
ULf4AvKbfPOCXCHWKuOenf2SHpgMmk2UhH3P60Dgwa2rReNs+69AFbR4iFuw0gbU
bO1Dttwy8iZDQsmeqBbyXD3bRoKqojYNhN+Zq1RMz0y3lbDG2uNPw7ogVcJINtJY
9KhUEY6TUDa800vmaMIghr5PKUayD7T7JCJquVhz6xKi2XUp3jhius7W6815SCZF
XneKKzehbPvTa0B+VOeknRfQQakWA4N08aRToVgXvD1LoxJ1nsiQo/REsBcFmI31
4p234mIHrKKZ1RFBkF0VVlnBTSJH34y3wIdj0+GYWxkQtvoPrvbQiH1Nadr2q3UK
O0/vKF0RE6tOC68M5S5c8wBhbxBgMYOwG7UQyh2YNQ2xQqmeAP0eGpIzOn+jZvhT
NF92ZEXRBttQPXOfA5g5jxsnh2bI/Zc0p/1xGmEuEj5Ojflx017OToCKZ3mNutHJ
t1lHhqhD6aDxzvRSDyYDkQlkcpBQmuZcW9bpZ0R6JU37PoeDcLe2rsygftnkwQ2I
VzcKIeUKbRv8UwG/wxkIDCmRoNDz1P/z0xW/Y/WyitOFI0kvXocq/4Vefb+l/j4s
F5Xx2Oa8nM7ccQ5H7ZVjrt9eKSK1vVzPJODvzIrAAFNcDKMxRJzhB4ep4/A4HAVy
xQl96rPQTsjcykURClT50Rt5WmZF8w9JGjTZifs5K8n/YvSCbLKxFNtoJYaSCRQK
VaLOLxLpq4ZP3gnl24YZk+fApOFnxIAJhETSAf2jbkeb1zoVfGvrKQm8fuwbZn3i
oNXir7TtU4s0ObOZk7Zs1iu0g/PT77LXsTBe6ejnpfYvcIS9tnurkQUKk1zJVoRw
WicctCjenzpOMWjQCyWctXaOu4nIXibOFlz/rNuow0BMUk0XFceMtfA0N/ENuZAq
ReDKhD9yo6LtCcYx30PIOes0IcynuNKCxRipTGUvQnkfxq/C385Tr6gtRmCuUPxD
NKHGd6piFDks4gxBypVCSPZpCl7b8qfY1grFjSfd/DCDL5ksKkCY4fHCQd97NhGC
rPZwGWOWwcGOpQiG7K0fY1REZtdL6MryPNpJJgzHTOxCVe2Iglgs5DCix3vU/cYg
GnHyayoDyn0bzPv600hZziKeh7MoGFUKu3G3MSkXHF4Dy94MyYZRhoRP88i2a2SZ
O/0g7vMAA9xD97AJORsXDFFuFNcwK2drK/Lsm7t/HFQFh1dj6bl4y828JLKbCHXm
OlEpJwKYYrUrMR30Yv1p8p2z80GdHxpmtOQK/5SS/+u8u0TY0oBSBMT2Lm0o/IGs
tFS/CUTNFWbLH1xTxsFZUSf15ijygKXOMxZ8Z7VE0BaqvMHX9tPFJwGzeo6pEeoa
Q4v1Nv3NL43CGE5O4HhN3sDwtxAlm2b5dytzWs+ZCWPMxTEqgRn6kS6rmpK3HKdL
+llZGfesEttl42Zu/RPOpapxxI2FdQ9JC/7UBn99Qs0cRpJQDk+EjoxZ9YEGtHUE
kGibs7BfVgeE7qez5TT7ZfzHfkoU9MDq5Hw9RaeicWXM2w+k6kHybCjqOKiOOaO2
nCwzH41fy1UER78ahjW4+OHSmmfkfJTqsraadC1GjMyY/K2X0CUS79yBW4eFFfuN
4BGF7zDEO68IG8Z365acBlfb0sChX1iNX7njOI9+yZTLOBA50SSUYpfT07sXxkZ3
fJOPJgMSxNrJGyRixzmXgnSyJW0nf2TkR01unRpXTNk5aRTrqGKFqaZpH+Zw5QLF
ksDdqzpdE8BRimlOgQ+QQnWXkq6ipJaYhzMOH7g1jqz5ENZWuYW+2FwTCAtr2NGv
w3ccyJyhWcsFlY0+nMZPcstva/jiyk1OkpaLM6fW87YDmU+sfHoyk6CinXAdQ49G
WuLrnVYTj0uu2KzzTMqKkQs20du9ZWiPTXpuxSeESFFlrmKqSzxyNbwevdj7ne1k
/lecy1lKRvy3ET0bd3ZC5IHyrjMZwJLk3t+hLo403MFj44zjPHrdXVICfbSlZgjK
e0s46ZWFp1BPsEXr5N01ET5eFjSFl166rKqXbZwNAU0bdSyGF5ygNv9MsTe0g4aO
YjP8ArX5EeC+Gep7qliuanBGriLAPsb/GLRGqwgNYLO2BiyD51vM9suIWpL/nzkk
hsNMNM8fX+7+VHeQ9Obmp5ritreGWZviX/odxovXx81HMU81no0HJPZay61FuCcF
19tUczWFGTnJ/Xf7CpqAw/wn71Rjy0rS90xZmKqZ7ikDkcxK5jQCV/tHcZQkDmoV
SPPduycBuBUNlGyLIv1DeKacmkWud/fdTYlkUnJWyPa/8Su6G5c4gN126wO6Oidu
Kjh82K3nrOZjJdWrjeNMGwkFmAyZrRZp+0rxhFaoBuRLbIxqWppnVukhmWCBVWRM
bJVSeCDAfLXH6dRPsRP/zbNpkyjT98ufQq1TnI6IFJYqMJ7TILZX0DhFKef/PsNi
wMI97nw88LO7RWDg1EOUJORTwdjQmSq47K9mVRkzh4I7lLqlsg7qjOoBFvXEdorl
aOluj7idnCfZV4PDinY0Hu/w33T3FmcZQQjLlOxlKmUnueoSyWMErl1g8x/nLtBf
1BxLLtc+sueX6VLu8VWi5ghW8A6BmU7dh42B3rRJTxjCiBpgvliKWybjj/xQCBgg
buW1XGdIaLjcNDO9oDXI8F7Zm6LeB7DiAl9eTAdpB840pv0uiRmQsga7fnNeMXCx
9ynI80AgPgN1UIdZiUffqGp3DoXprgpWs01a9q6pDT/RD2kzzxGoKhDq/CKs4Tq3
KNtj1mNilp5QbJoerqGUxxjtGdWWMFGE2zeg2PGD7Yc9gcwXGpxFI/j8xhkpVcxa
qrenje06eG3TULFmhHAbtDMDPsLe/mYkiTM0DjnxniyXuYD0quu2u5DBAZKL/goP
RXijRHaCiFAubmEoVhwymzZBjSvaO4PerVs4fHHcUGWIy6dQfTYoxjzjAtIlCm2o
uFZba3rYY+SUFpDLfAQbqn2sxEML3aiU7e08s/ueXZXXf+QjoZ92O3WZTTatzl24
Xbor1Ty6HX8xO9GozWp7nOVQRqWaVsR91O6guD0ZQpAVXH1gUDdWV7i7acvv91Sr
s18O6LhFbSsUkSVag+c72hWF16AydKKXc58oLUO22yv5BqnA7vzs3dDgL88lBhGB
XKPj1EF3I3kI4jdF1kZe7ObYUM3PU1GACF6dhWypfQRUhTPdogo9Upte/p+CzdGI
qnnTiPfAuub/vDup++Una8BH2Z7oAeLYyKiiwVP4JQpnVyKLY1ixGsRPUg/Vy6to
nQtu9pXAT0BsiQ7rDH3xFBOdyw/1S3IOc8HkFaEWQvJZ5WqnY+ElpqNAiIIn82UO
VKW+ZtEZuDLTXMdEHn6AZQ8RqCfNvMtD/JChJy8YOLmpoT4kS7hHmBQAQk0osFDb
I0Y+UoTtKNl9BH2l/3d/bM/Dn06d4sW0+rcNNjEqTCR2oXWRypPyNny+BFp/cn/l
YUQFK3wKAusaQ/0tGL6k6n7OLMwLnKCsC0NrHh+Bbu6nkVwatNs7nKVJ4Tc6uekZ
dC2SWHnm+fa+FcCy1+dE4Z6vYwveBouXvvDhBSo7lmOZcAnZ1vffGbJm/TOQO77H
01gW398bFimQIIvUJyznoBdqrKEbrdkFBUx41xVjhD6D/im75cLuYg/OaSRdcML3
tLSjJ1ss61w9PtbRVYlM3UQ52D6STNQ254giHZ+MxarWZCXmlWHBLZxCa7Tip5H1
M7ikqSKWf11y7se4tj/1YfkbVvK3UItTiuiJ97Zq+ZEtXh0lZ5lRz0kUkKMTNUFL
LkKiuKzalVFkEtuzo4zYFPXxQ6nZNuh8aDe/cM+hxkBkhple8PzuatUuMo45rQnC
4xCxtPMaLuP2FnfTGcfQK3K+aswuYzKhr5jws7SJu/2CpZnw11ACXUFNt5Y/xTAF
ifWzlyXgAbkT10XsOtOFKe1Yg1a7V00/HsvKNwBk6X9wD0dV8zKmtXpVd3KUeog0
x7cckSfsrXlWh047XIpwJeO+mLnxQj6n9xAfyUqN7c3dJSPSZCjUw7yd7ByYq0Aq
+0HHOFvFoltaumFa36Ay3rhY3ZRMNpy9kxPAx/AJK2yR7c8Yt9Q+H05C+7wyHYl4
vyvZo57pS96xA4jC8a0bizgGIWvtW0k3f3TSdoQ9dzXPSN+78H/Qrqx26eQ6vG8C
zdYCMJKzsRYyuMalULiJDxk3Pcfu1ZARIooZHs6/Hhsle4Vk2Oo7WB+hWnaeMJeX
k1Q0Q5OeIKdCz2Y6R5aTgsoXM0BhedPi5umWMfoHy6LhsJ2zU3g2gWCt35C3xafu
Ggv2lfq3Kz5+11LXDrn2atKF40FWJuNpLw7r8O1r2CF+SLH61gHRGeReP8jB0Nmz
8c7NvU1nTJWcfYB2eo3K3c6QrhrEMOUi2t+AVxNmFR33iGi/y8fgPmA+DGtU6uLU
b6R+AiKyIH2CaXiijbgW8GFxaq4k7n675tNp9u3K1TbE9bD39PHjz8XIw23gz9pA
BhnXbW6YWbDa+jg6Mda0Xk3flBMrHOp4I/UqxMu5WrLuBV7e6HoiNPYO/ZUjdnPq
Y9vs+TWz1AbMSa13PEGudWKgD0qQNIptPpGCllStqA5h+zZoYsKytIIAaGjMO+/N
NdtlKDSfOpnNsKnsjBBIi5b3LWVXXDC8cifdWKUZyAUGacuInKAULErPV8biNuiD
3so0/49AsNUG/LOW7ZMDS20AEm1h3IUHCUrI80q+ei6drH0LsDuiX5t+kNx2PtTP
94Sj/koMyPLbSJzFMdptMyRRJ/4CwlcrViYJpobxxnYBTOMtu2RVcWi7yWZLFnWs
g9fhIGgJCIKBvT5LlzQ7iOMTqWNsHSCnP/5SyLrrFIPFKG5mnVgVcpGcLT9iJ8UH
SwN84EXfcnM62wyu84fOj54qJQJiTRzdq4FySG7ChqKaQ8MU+JUxf35rtFV9Zpn2
LVtw2Y9W1NQzynfRx+GToiS1TO8wXVbfNGJRQa9VC7g/Jafgo3223JWLZzno7OvD
Wn07KuXSTbmrlvE8h8x5/gF2+d803MIuVLPpOVSaZ+nIMn4QqQTyOU7JX+BOgKYY
MUzr7k3z6yWc4DirfANogD57V9IrPnQx4JVRnxLZ78CMPGcOM3KSGM9mOtWNEWz5
jhMYVHM/iKq3w//O3+9ozis3GX/Oc2zLRTq1H1xQ+a8upUXS3/SmdhCPOigje2vR
LyaKaTzlJc6YAiH0Wexpm3KpYGi8ut5SkA+NLaJ4xQTPmgNPJbOgY+GU0gVBJ1YJ
Of9t7c7AMYGoiyMXRgN6S55nWn7bVYLn8bmCN87KACYx+DH3Z8BYGilfbBGItuF7
BWQ74EuWi58f0zbC99j4xEG4wC4d/kfwk/+poOnBgBHRPnRkOvoIU5r8ksKpMS46
qB3o2lwq0LsHIrtMML6bfr/wo66vXci4QuJOZDpkNAb/HoY86meJjvGrjYiztLvt
VQxhIfs5o1TdvNvG2uwg5wDMuNZ3XnXrZzktTP9ejEdVltLCpjhW+7h7jqW57Uh0
x5Ziuhdux74fXnsmnXCH3KIXc+Tpb0hkeRk6GBshS/ues8SDRakAqhRqd50zukyL
XdEJNmvp8hrdHxuGhnnCkJ+CnftBxvvdDg81oi50r3IUpuEhCPWpVZ/zIviCSxlW
qafi4JZwNZyU59ZgDrxz0FCtK3KMt+xf/v7rHzZfWiJ/XjmTAW6QAxEQyq+wiuFU
Hi1X2iNu/T0Ll5S6v8qbUDW8MFQdFHhIA+72aTy1dJSlvdEIDKjd1YfcQ+RWNjaQ
++QGBZGrX5uf/Jaialih+9dJfcT4rqnl0xaQue/8Efz1EtvKg/xsKWrodcRRNocq
+pbBdrEVeQ2LsAlu/x/AObnGxWiMYvJjbKKf13zVJEbl4Z/Wkd+o1GiOwcz1h73p
TV0jJy7+OBcBnRDa0oJLb9bq5Wdhq4uiO4jNrTN7x5iwqWn85eUdvKARXbBsvUj0
bnNEUiA8ti/iMKGYnsvstzf1JLA44T8tkeG9PjhNxtj8XQj6dEKy4bG0ruwvAmP1
h6krFegujjh0Daq6qHE+eZjwbPX2bt6dCsS3DKAYhI+kW0g5w+tSuklE87+9HXnv
yWBIh5Jui4MVqppjWtUzZ7b+PRAdIb5qCfqjqggjw6l1pqdiwMv4ZOBVSENk/ID3
L/2gM1Jiw0y0TxH+/TWKg+UzdBws5CSf30WLpSZbVpCX6iEe6svSWiDjYjES3d2b
Zv2fZBH91NtyYOoq1gKJVUosaF5z056GjLAF8/3NOYu1zuhJMeUGqK3/MtKTiOYE
/HM26hdos7CE66jq3SVShk+oU5+o6Rn5etBxkxLVmaR4MVkivn+AorzJPtDOQ2KL
ZiiBt78zFMH85fW9y0At1yTzJyohTzSFADlTk063vU2Xe27Zqs8lM8qljurr8MPh
OckEt4PzUyz1lB6MZb3hfniULFtajkQ6cD76a5OZPYOMj6StpGKzCZD11KcX6vqd
W4btemmLUtEBda53ibjmV08W2CJnKAgNx+n8RJ3Gs+/tmh863UhlCMFPEE9kxlh9
2cbGx/AbVgMTJBZnzrFoteJ59nWcoYklUXLyJjUYTxLvfp9rXHPXGuOakjMV1qMO
nVQWFuDdcO+PR4/fEccLC5wfuM/LJqvtOj4zCZog3vb84QPYTcNwQz1kyo+BgLTi
+7JobcaaLrVpg2A5doY3abod33LcSYlbu1VsPvhGJqzJ3VmEoXbFQGQ+vuPM9kfV
jvkUva6cEgI5ZeQPz5OevR9SG9VHEcpmeIROqiUkSxH2QvNkvytXx5lTPn1oiPDC
I8bG2vf5+Iu2hwVT5K9gvnf6yluJnH3x1LshgdFhWmMZPuv60IzR/bi0fRZNMCN5
Hjt9zG/CGV1sIeyKMR7nralhKrMZ+7h0Fx0LJhoF6x8Zp8fApo8PWJOpzle2Tuwq
TghVf4iMcIRqhGIu9dVVQgO0EnmxFiR2vVLb9ipioKmkre63eDGY2wGzHr/yypA+
OMlaGMmD2OpvvyjkpJqlz4vk6gJs+YxQuvkKR0IeLS/6EzVwY0ZK+ae1zpxALJRQ
Ng/rwhEW06LGjcHH3nNHgCyzL85p3pMjmgszCib3d9ivKMkin2AeouOB4K881SC8
iXH19MPt6nQOdNJtDYajAzG+Q+qlMlhv8vZIvVWDMrCqnP/XeA0JOBC42g/yLe4d
FTAeuObSph9x9LYZrHMpYoZuA2795ckwjdb9ahrzHK/f2bC6w2U3bKaB437591ML
TyIjeH4Ywtu2o9GQcrV47b8z82crnRa18+O9TItDaUmF5m6+RIomNl23eMv7rCzd
D6M8hdyqRSkffagw9kIiDZN+wS5QdPjr8/8SRHN826m9rQW8H+BFVYOLUlNz94UG
dcwlu78YlcnDqU2ZQ3VArGPREQDpgJz8W2duKYk/cGxj0JQvXSP3X4sASs5z5P3T
HhGPCl6U86ImIXOFF3pp2W7wXCmzECSg8fF3CGAeDpHxZxHcbEhcqFmKqIyjFW6f
koACANgte7M7hsrOIfWEh1WeoxjyUmvICfd5VqIi0hQIkR+sKVtSx8z+vrPSKWxH
cBa0zlP/2HgQhhHurtpv1a5AvpZpxwoHbPv9FuOamLC+L4tFQyR0i2okNzxdU2SV
3sY80JwjIrlL0ci4d3C3mHWP9lMeLQmp+LkgRZEtLJFdfdJ0wtC+Zglqu9seF4aH
TZLD2xmwIOTN02jRr69EO9i/wno53cxdklHV88TFSRKtZzSSL+n+dZNMw10ifPmO
LVkTwP71ra4nlHcz+ZBaQOiPi0bmcxNTKYGz0XqWniBWE5CCPzep8zvelnqpI5Zp
U3oTodc4ttI37OeAvCotCxQMVCVlvBaanSRLsXMIc8jqj5D6HMfxX+RMOKHrGRG9
RuzBOUEkp9qgZyB188j2zpoc06ozjGYo30nV/859iugW7tFcPP00neVZ8a+ORYwF
YEi8ZA3ss0J8GL/A4+EVuIPE7y6bY7HHPHi//6SoR6yNeN7S1FwGyi4dTYAlpy5u
3/B87SP/4f8PErn0hSbK9tTao9jAtHSSrHwy8dKSXTPfut15zzUL35+Ao08yh+Sf
gy5T1vFQCv3tLKD4YlAGW8icS2SMrxmPGiYRR3/HOSBnGBN3a5iKyPN1rtSYQ2fo
sTygXQeZTStqIvL2KXrpLvIEnmEUEwYbpykOFUfLw/C7G+HSfnJRBJIPn5Uzr0sj
169Ge/M7wkx1ErJhObIiMTmxtVjlDUd5+ObQNKIy+ZptsophtD24XTx747w7IqtJ
sUrqy5X0k/fcaVqCVCT4xrLb5NQ0E9RC3+MkNJzOfkzvHhwQ7eRLskKUiFVuOdLi
1vSYXDk1eMVA74CD8RLGVZ4zOhe3gnoLpZIWVhsoaId7TxJhFyHdp7NPcnZmXVER
8o6us0Huxd91pDBI/MlsoRGs1Dw1PJN5jv1yGsXB+wmPU0pbTLpSARoUnCf267vT
Grp6h/vJ6XKEy03BXaqmRhoFoWtTu2mqgLtXrCvKawGEBgw5JKvgzzZBbQFzH0G0
jrqFp+UXgdMasDvABOAHlVLbfGv64dzGJCeBPgaJZBSSmU8q1ZEQ1/9F3OHkcmi8
hT+UCfHJ8AtjClO8D2B5zGkZCyETdJA+7S+2FQuTcM8BEHMYvvVo1++svwy36VQO
L23fjmuwS2W5cd68EBjNNPy2NBTtfWXejYQt5LttlzrPmMNBLqSmAl8qCWW59xcz
j9wthvuefTGlKP2FT/r7gCSvg2ca6Xe+pTGDrTTq07F+T/BYRoY1bkQShVrmt6jg
H6NUd9ySBYzVcRx4Uoj0CHnfzKxPcTeqYQ/cgUXpUSd9wYgru51IjhfeG2ZiFjYh
MlR67EOnLPt6vNXIfPj7+FdLUNkFVCFTOHLRaHqnXLEs0Vwr6kNwbzY5ueOIzrVE
zdJmNlc7mbjpoKeoj8BoAQTM8vEElCNW1RR3TCjW8rIwMo4T/rejEw8a31D0SiPc
B2Ir46ArQi6LJXgN5y3sYqdNaV6Gr2rzdr0YRKG3WyoZ1ZmUX2FQI6AuM7Wme0ge
haOJ9Tr9ECaTkp92742szJndAzuuSTz9jzY84oIZ1yDk/TAwKp0kdi+xh96bsL4e
+0Fzykqt003+m2W2Qh5pS3DmJ8NNlA5MWVfkBFYulBSTtCWUVxlfuTSh3QyQ9D1E
x5K72NmHp9qOMM2t5b9k9gFEXGJNtA0cbV2lEWPTEISyxXEvMrPcqrKSD+aGBATx
WJ+lYBWoB3uJFE8NOfd4PIENoX4CMSrEBePZseMqhQrz+/zajHT+e1Fsw8rSnq6U
ZtNHj7GVItNMpWGDfLaJw1sjgMIJPAv2vWelDLr2aXA5CJmnjQhcpAo8szlxXQIn
0e+1jVI2kKnOB3eXKkP10rKScN8JEMLuybsPk69YszEufdT+lMDs82N3+7Kimrm4
7FldZHBkSmevl0/PRT2rzuxh1FmyYUFsSCJdTF2BFpVeyzrHCTgcPT+zLqD/3vJU
9N9DDN+Xzy7rq96XYxU2W4wOJVNi0mokiJJNlL1exi5us1Pklo7vCHYy8LxNlcS7
kpdwWOU5j+EYy9+ETkh1S3JV70usCokq9X6C8uVUe13dmJBb/+Ed5vHfqh+5+ZfW
InIDib/zvMce1CoWnOAexcdOlBMHbM2ud4NfUzcxR5cMSHAHB7FrYUvJk+ehzlGt
k4Mgp2wQVZ9mNDMuiHruvMDWmmWETo2czKVifsuAywl2DFeGZtY/Wbv+24Bhji/6
srX3346AwNHM5LUlqPDIybvxoI4V27Dgd1BBrniS1mVl3PIFYNdcL8EKB/PDuIMf
bxb0t/fgP9e2Tb6YOlYTAgkMuy7GrS7/KSPLAYbmSSvqsSdQnFkGNNutoX7vd/Vk
9xFFHEM0T5zNe6nXuXL1WQtbStxk17IYY+yKtfMBTCdftQ4mNve0OPa/OkaXwzrs
vZbLFBfnmEFdQ113eYP1pDNGS3cput8/p64AnPi3i6Ba4qzNbW2R4QwXa+kalNms
XEw2Sw/zujTyVLw7vUOJTY8DhbAOLWyzrM83FnzS67KFNQFap4EzsxD917Bws7R7
yfiyfFb3tieUdJNiV/+JGwgwAYRGcT6bYW64D8awy39iFi5GOtgf85otEltk1zJZ
mw4Qt6fF6fRpYV1kMm7lhvrG12GrYL411pp2EiJvL3rAOd2jQ4rz0kas5gVC90w7
WEP5XHHFTqyT0EsQ1+czUWMThFOUINFs+xD549Qpe2/eA859/j+vKKm6clyBxfU2
0+TnjeWH3RZtGUqSX2H4gn8Jj+M638JYAbJgYct5L9ocC5aelmJdStk0qlShKx5A
xRRf6nPsbOD3Z4Ky6KTcE2X5BwCP3woQzXmiigQwVrS019aIJcw701VHoO50Nqo8
sPhOpY6942CKTgTRo+u+aM3r2aOSblRw0yqd59QNR6A5pYDrqwf7a+rVMZEPA7ll
w+5/0g8B+3VnevivaYVevDzwYQcnoKf6C10nTVLm27YZSQlNt+YAJXYG6qpV4KsV
U4pQyMoR9oku1vjUdnUyHrJdzRHG+JjdqWi0+zGO86J8YvZWeg/scDl6mfhkUbz4
rDG2GK+T1d7hUX3IV0bOMlo8RVOWh8zMyAUWUYm7KeRjU/Ilt0spdcE2kYRE0rrK
r9B1CkBSGEhtM786SML5OjPHvvBDnl7ZqEjcDIOD3LRx57DkTqNwqKVYTLSEsw0F
/eCj9KMlNgx9Tj5Yv/5llcEGtNKWT6cfd0cFgePDOAPENEDC6cfh5ilNPqPrPR0+
suaGaTfhjR9GY/VJEisapMoUD40NCNTn0/AhWUT0zI2954SRZal7NYtVwyMZtMwT
etVVdL5FgPWqol2JNltH6uvKB2L9wu75GhFHQ+lHP9oX1O64GHgVhLXTr699OaGy
Zgl2uPZWRUx2EuD4uaNG3l8QNDN30aMLjzd9Kqw09HHnUf/8Y27ewtGPtsWoZERW
qFWhdEkNc54lxa0hUvueYA0eolMNbA78bt/+oEZ5fDeVymWkprRM0lAjsqRsOmpi
X+71LD/Skb7yX+1JWCf1SeGTbcmMDko6yWsc8vTRDHUyBYK/HvYjHZA1i87Omltj
OrDUHBLZjo+QnpUhbpuXaBHgKL2Xd5h2mT8wcVgo7ZJtGHLQSm6XXAnRJx8sp0zJ
CTSmkCjbhPSSyj30N4k3r7aK/wQ3IQ701O4vP1l13hKbv1Rn/VdVFAPD+W3uwEOY
VN7lT1gjgjEz6Jr8tepkFDAOm6rRmZrdpN3Gqe6RYy0nM3gRPwJN58KfB+24/rWh
JFCTUEiBqt3GL6ChJcErZ39Gdu9H+WsRgEuNGBWn/PST7EEDVa1mBNNFbE+cc+rC
JI3Y1qYUIjGln0CMwYuInD1Fap93cqfbVtktkSYCPsqMlinpe0HSQIReo0BWnPJP
r//rovgARqN1K+Wpqz+nTDoprLN82wiaTtMgxZY6i8caTYZADKJbmugZtpYA6bZO
bzq4UsFpXtqhNKbEJXMoP+AZAATDZWnGU0d6vpkohl/P3UM7t//rA7epL6WiSdal
jh5DV6vOkqDImTP4SJDFzC4/m6siMHfv0aumxznL12nj6RHhnjldy2KidmQheA6R
iVbftX0DJqgiKi7TpAgkr7ELwatWiddgfE0cMPG8q9O5FbCt0oOhbvTnJSGLZ2p8
2aIvdS5jqoBBHH8D5qIlpM3MxUuX2pyQ7plcSy+MuWiLU8UCVRsYp7MaHUCpoZB/
LgLKaCCa0meBtVd+ESZGFzUzW52si5/ej+IKgexIiTQU3kOabrmt81KvQagJwFKb
55dSygW1LtPrcgYZSuvft6tLa7nLkm827YXVJO8/t2MXAhi0+Yyysa8gkIoRfPx6
ZYKtQTabEbp+UPj50Cln306plJWJlLydRRVT5I+cK7LnFtngnCMwSbqV/hHAxJM6
uZUblZ2Wl+aVGAcjOyjI4TIySXge2Cew07mZUPx+Y0PBXJFbIrLG4LHGvDvNY09L
TPTet+YUtcseBkKkFm60HQFLkIJi+wann6Fz20bLmS7cWOOkUNFQKhV/zvjjw7MA
Soo8jNAe38AXotz3ovzHIdpH3r25+1gg+1LKh7njDUJoBlI99UuXfnf4UTsTg77m
OoNpbDDc0HPRCwiZTlu2anEDefYvkFTfzXKVs8wzwK3zIJBsoBJ+T73JBJPMcDkV
mJajloCyRthpulckk3/F2FRaLhh/lzAxwauRSOrhUmXKLIHh3hn4u/UYZccTLF4M
WnxD8CxQ48EiBO35hMsiWdc3zvH4QwNaXltQ3NzM2GhVTQolP4HFb7cE3PAY/CUc
WlpHtnNv+qavIvszMvglub+w0x2PLiloM8yQjwC5isq7fdTfUJbyv9xCrEU2yEq5
rdZCGev6+fcrapzuKOR7xf8C5VPPnGuMKkFCvRMsrhgoVgFHcn7aRRdo/go6mmYq
gL695vv0jf79PDQuHXdbRx+SyGmqiHOtm/KeoezWq5Wmy9ym+Wn4uWlK4EdArzx2
UQhsf93Gz/KSpXYy4F9uiHqap3RsQfmvmSqL4SirExeJQO/l+Sld1CyTNC5KxS2m
qQubBNF8y13VDWzMlWZ6UKp5ybDrWOpQWZwMvLUJHaBQUkJ0q4kpTz598tZwXSrd
3APCEZwS7yxUumSUYfkft/ahCT0VCa/J5SqoZmSxMuiZcZtzEbZ+bA9c2GjNqwSE
qGdaiqTHS67A/iqisBDG0jZYCyQ8sHsybbZaTGZ4d/88awv31hTcHqALDbNirh38
uazkIkXEPvc961V6QqEX23U0txVIWpz2wpkS6sgxfZ6NfkQaMHHidtMWxSxEH/QI
ont83Rppcftfmr6X9U1y75rWWI0YxJ1Ax7wV09yaXtfxPnw1awhRERmop+eughlU
YSMnhQrGCKAdeYibBiMcGLehmnUf6azNaHrtsmL+54CpKJUuA5YGIn1Vir3Ehl8E
i0f8+E7iWLTSIJYJ2ny0xDS5QIEP2M59O94CtF6vdwdI27YuNdtXJzQ2/3taCsb0
BqjMDzsh/GB9Ve91YZOsPc6OrbHKCYuigtBEKTMoswb8jYYQplvd82eAmBgNJG3+
SFEOmT46K16S/N5ovBGvH84MGcddgKn4Ha0D0bGaHV7mpTrhcpOc/ha6n2FGJRX7
OTEKwT98b0bZLqYNa1zHc3GcZRpdVaM5l9A4usJz2kPrMo+1Vk2JlijS2d/LpfGm
5VkJQC4VWuAyF37NWtuNxN2laogwHCqdabZA7fjlBSaRdgegh2c7w+TAgI8eRsu9
DnZc4wbFebNREsInMidWKuLnR4Q3WrH9N9AD/7ryPMyH3goEFLaXBQIlm+HNisYK
rnmqXbCrdQ/U5vA/55+r10vB/xIA6hr+hSaGhiNMWY8VlwNz46+FcIWkN5quYP/V
si1CnNpJNJkLqc/2HhSU6D7gTYPGi6LoGGeiwR6oqRePeaBjPxc/kvbQNUlR1YPX
bUZ1Ht6Qu61V4Nwe4lOnonXY1UBh7r90S0NfESCW7O58R7FwqhVShWqu8ZZMRLYe
nlBlE77P+6SghM3ZhNeoj0ch6Ed3ctGd79b6Ta7MUl7+LS0bvUQn0ox55ObI/0vk
Qy4N0mEkw4Y4va6g0AAv597syxxjm8hIkaIvtaP04rgh6N+idUtk47Vt6quty7Ja
8ZRAlpl+KfzDNT7TV7MxOriAg9mbyZqNojjUHCbNW58GSVI6WTWyJ1vfl/wWuVZM
2YuaZEx9pfUIx2qg1BVoZQM+1rZN8ajg40Cvq/RJDRZRKBjJlV9zXfYWCZX61HMw
xYaIDSGUmjaUCUIVryzUUN6Mfv5FbHmmJedNMEYuJ4I3/ceON12Vs5Db1aQsWQ23
4PZELAoHu4hmtcJfyHsgp6YxETzYqWnn/iBXNvzNLPcj3KgolwU5t6s1bxXKtFf7
Z9OtGZMnm1Uy93CdGUXE7T2RqsbLXZGQNaTiP50Q3TivYaxOU5dmbO+V1KUU5tFD
2ZOtIRCFoHXQ0BO9uk2TxDrs1BLyLsPyYEJxCknRcsiuAcAul0uA/fG1pSo+Guc7
R4xJR96gBoaF5UPmvcZdEEvSJh9PdyzaPhW70XeT4lNzIpTT+jsg2c+Whxn65fMq
3z5GoMvaJq+bJAxUFHOSmA8HzgSu7ge7v78p941ykyF66WUYXvFaaOw6PVuOc3sz
HWfUl8xq7d1eg28S2xjL5LH5geEQwmBXR7MsiHlOlXbNZqPClMUIbvd9h5KMNhvD
iPXl+OPirlZq9asueg3MmQmmfqmzVP3Rtvl/BdzYJc8cKNLz9P8s/wU6P7RmZoki
nKnFOppFgN0mmkgNS+94phardO6WEzLRJqwTn0kLvwSrDylj6BIjb1ZDzj90nJXY
+G5TYzmxAP7B6UOT2M3K0MeW5Ha3/7Cs8H2w612/QrevqPQ9PSoD9mORHatPWegN
C33JVEUGl0njLOyW9YOXnfQPY2Ms5zoUzOMPlqZ7y0cSj5H2Eka3R7ltpFenp3cC
8ePd+WQdJAp1G6+mVFaAe83C11RJDQ4LxZthTZNgjsb6mb96Od5ZG8Ess5cv3sGA
cR5we2DScJmsRZGHpcdnM5h8F7HE5tKzIF5GW0T4dzvvZRI0GxarmWpw+eYrFW5/
BARQJNfCJ8t/gRPxXXmjFGx1HAr9/oFXT8etl1r8XxAxGbTMWEemBJWTvbP+aOtH
dlURLxPp+tpiM+95UHk6DS5B2LrSUPCmT0Qh5ig4NqZUcEemaTyRHrXsiO+ujvbR
tmtA9+7Br3zRvVZ012pL2AepH3tehpw2qmm0SqkNkGHNQvyFnFyY9a2YPClKj3na
nHZL4GcKYXqu8Bje/ajgCzyNoEHmIiV7B+TD5jKN9k1c9bV8Ol+gpdX4jYQq1wS9
ZV1RBQUU5f67drY5CrkCT1DdY3BmD2U3pUMdxq0kwxNNl2Uwk1VteYdb70mDdzlp
U6V8YuGyrMOtdEd7AIjZeGLHxtvpCchgpNg4AO99beuMAFn+qSOIII/b8LTj1Wka
vyQrXuNkO5sQE18xGzDUBpyLsFFODqFiG1S+vRRs3jf/Pa0x2ToG2ORTeiL9F+OW
9zegqBqwiAkcOJYZ44LvA26uuQje1I+WjKt9C1f4KA8B4X3klzsDK1NVAKJ23g0Y
2DjKt/Q4K7ybBhpzh8dI9WEM9uFGxqzXx08rbaFVpV68v495yn4EpB80nE8sslkd
IOptdH8vufr1FsCpNIWO/QJTsxWrjmjA50KLHQzuf5x3gxRTCRhpvWGcvPG8SyMC
CuMugkIt/f41VhgdLFqjqJwshwSzVc7r9B2988f3En/U1hc2ikwsY7yPKnEnUBF4
DZFT3ZV2DsP9qFTZiErZmgF3UDerdJPMwK6FQQ/Vm92DoTiKqnPv10miqCbM10xN
uX2Km+sJM1eqhp6L7q4YI94rzCdXCyqfTfGwWJxFr6y5Vn/0Dk8688viYtyT55nM
WOc91r0xOiqpb6a2mmDxWFs/ySi+VQlQFCkaBURCtg43PHrf9PDoWcw+rPUooe7l
6q0KJoAyou7ulGXttUtQWygVdf0f5ceUA1EbfjAga/ej5VSggTLrlN5QRn4OaOt7
w/dhj+3IePJTBWIywEStzylMBhga49JkIUm3LFPj2zoiNzOmBAzgcWxUqlsU7fqA
7fHV4WSX1HL8hnmMag+eBXd+LgQbTVNJCOe0fMn9nDG35bt4RHcwKqWAZuP8J7QG
NG2eu/dWDfqGxz1K8M75dwEGO8cTOw+WvjHZH6ZHnvrvyihmz1jxzT1wywqwRfqb
6NL9nSxG8Xj0yfAQGEYTmIU+8qhQCwFNLX/D5JEehb2XrGK5Qm/yhMNgqlcNAqjN
TNQo4WZvyQJNEaSDqJqUNopVRTXYQVUboyGwbaOxQ3xvTXOb1alKpQq019qYgpUc
oBSI+K8o/y4+3GuD9aJ5epyqewwqQx+NKXVgWa+B6o3GyAo8w9psv+52/HyzGClj
bkkWXEL/BBMANxQ+7A3S19fM6dsKwxcMOz+mst96lGQaf1nGbMLj71BY0BiIQSbc
ysTGb8ujhzweDwMHB4isY3RER+QoCHaDGz2jNPJN8OXGyX35wcRGv5NaJLczH2tY
QxO03EJwTreGlI+Gj5Kh9ugayfCxBxA/ARDnLfS4SwUJLrpT0Zb7fge0Niemu2kS
s5zAlgg5D5aossQNM4CWIZZkGr23AAK5xLlE6PbljntirObUBJU0TOd6r+ofv43F
nb+EVhpz04qoTYIU/AX7QT3ST8tRo1ZXhMlsR0IQ09RGqUjNARxnyZBv2V1GtBYH
CPEBZ6EqOccEbhMDorwMJXEPDODpYIa/L6g3cENM65cLoFMGxZTsjxxKZT6z/IM7
mR7JQ5e3ziT+QE9dx6WyOvoToxMphexZejhxdzli4vkCHlg/LUoFYixMEhXrxwGg
laD/kpkCspebMdCOlC8MOBehYOXuwqFDsah2OoVBGroOsU+qiNZ5PNYGnV/LYZX6
yzpopCDWsFn6WhE2zOCK2g2+y4eArDGiDUoLmxQfR1TMGj9O5xA4cNRRRHqqNXWi
IM797dA3neRXdFTLVp2CdblhOogu8YvFTC+VUIvZ1030shRJQW7raMwx2XKHx/Y3
mD8ghnLoVySdujXXj/sI0ncgFfD9HArKoezXIpSt/GSeQz81cc4bMUVUxBSmlCyF
lP9RK6RJxcFn6NRhZ4ZWIwXr7DXrsl32tjRuzGxbWK5xUBjy1eOX5ac+uvI75m3d
Ogg9dD1WAy1RQX2p4zT7a3ghQZhvLUHXGYvt1SwiEOx1vmNIGJ3zxQq+bmA+MR7X
8PG9bvP4D1zNejMUi1V11/YLX2nWW35ujyIXIyNGjgw/mn/Mkwl13CBg5aSVkGSU
pgQk55EGtbiknRtJoK6+CSEvCvALWJnM3eT/9PW9H4rTaObpsxj4KrvGuywyQDO9
W6H1+IIL7JRO4oD77cEs5YVrnX90IVT6qoMiAiEaGz5v8KGS7ISzzLjcreDPMZ++
QwjeYRPPRWzeXy519ia28lyDyPt6TaGZ0MZoQ8m68014VA7kgXB1ibwvHaHO3EJs
aKBJ444LXA2qmmP+YJj0QuHhRAX4uUpX1JaT5Q4JyZOvCOgblho2ecJajmECdypF
i9oN4T2wT4ndwnXkKH47Drpd2ctWGeFKD3TMHCG5inVtodsiTm1mUujpYnvhADc1
icqPLjoXaE+ifTPaybi3iWEkGuYgD7i7bDnEGfmknpRX/gEwqECzuKin50cLTrhE
fFJaYFRG9nWszjHp6BFXycceJ/0mNLVvoEEWly2hd6HknQ9XKI50AmP6gjBz/YY4
J5L7ay6m2fMFxGS1VnyiXn9IiOhFo+SpHtmVpHPwrZ6zNvwfJ4A20j1tLeo/2zwb
679/HrArMhP/rIv6Wiy/Wpjsx/JBTYtO4PwCbjKXuhgIrtiIKR6KeKdeaxxm4kBS
4CCEvASeY2HseyQJMyx3mb1PkdYAB6dcqKjKhAVPgsYPXftMej2fVK2qXl+fDseI
7WLOZbPnv+aigLdo+xy33YXL+1KkpU4Xt0+C9l1VRFY/ELqHr1VBOlGwjd/cW6cZ
5NvoZFCDKxfdwOmfhYOOlguaKRzyxW8Gh4c3E2+HvvbHspepT1u4BR2YPkxmILnM
jU122O3VFM3yK6r6dX3MTJ1QE4hkI19Ux2gXT5267lTv/9+fXWEnmGQObFh0BOFl
hO6HH9yhuzE9Im+V6q2gQHjZq9FUPz7iQ017rsfWXRu3CR5KC1YxzV6IUaFcC2UQ
0sTyBfm8lTbI1m8yMnjO19XGZgMXncMA9yx1OfEr3pYkB0Wcy7W5ym9M9s1OOqSt
/DLRz75xYSMsQ3+512xNPfTkHvorK5JcGyCKvx1hsrr3N3O1fOMt+h5LBqrvI4C7
cYdt/tUv8TYCwtGfEkHHjAC2t9PfOqTiQ2yotqhx7e8ieWBUTEojL05u3YwLkf4D
b6ouJrnxKAxXM2Xepj5zx96Qs5guTdP9GxxlAl0Juzkg6eZE7UHEexnD15yWBGME
8qnegJ9rHJaAA4E1MhHDiJnIpWv6RYrTI2JzD50Tkt9feshsVgSdm35cdz30Q2dH
x8FWnDY2NcvdlFkS5J5Wz0Dc3Lkm7l1B7xhlqchL5z1UzdLJD4odtBMRaXRN9aLE
PXm2hIAgwZLiG7X7L3iT6MTAGBLty3X4ZpQTkbNswAFo6wx4X/VEfI8lXg0cygmT
lLbQrVvdyDJ1+6VM/y/uIVdNMUsyR4sqkskMoLCIL/8Ki5bnakNIVno5GADe5RPP
WDtkm4q3CVfoeV4gPR9380ufdWpTX4BYdB1ciP6dubyYKYGabP/HZtyKgJipHtGA
ix5IDEUP69WABjESbvVAZt+IAn35EcgUDIJGHXJC3xqFi7y8YeP3L/h7miLZ+UwY
PA20+RQ60J2ZLMi08VAAnke26jsQponF5NPjk7wsLkBQxImrVIvclmdmkn+FMyhy
mEQ7hm8MniVOYRSzp6f/zYo7oufrtUWl8RSWboSti8lb3uL+1EdLuL4I6lfaJV1A
JlfcJ9j6ZlCNorBmfX9SUmBfN1J6we/Yr4VPa0AU/cqaH4+OclNLZtzL9Pl46h5B
AUlJtGQ07rcP36VxcRfegpFtnj/DGQQW3mBPmG2XXSfJT36gP9wt0RboMnR9CPdv
PZgzIURF8avrkQOGl/rYb9vSoyZXPHAXT9nIsE2mHPLHY+1h9MTgc29NfHcQAw5A
RnFK7WCCALRb2Q8hDOZ9yRtpqPzyDE2F7vza7L091HQ3Z3RaTxnZQfU0pcIVzAjY
soMks7LJ0/FiUA7oLgy+iphka5HhpTKhl8oZG0OFgRmhgnnn2tGUbXtoYZWODmoL
tuqLY8wUXohEIaV064QlfEdEKonm9n9Zyg8+4cj/UBGqvcesH6VrrP29x32abMzx
Q8j32dMJM/RHIu+3uYLm+Sm5j40qabIq/V7hOOX9nzuq9O8pONYXZ9FvjysXMzLV
GjfWCyUCgdKvOP+2L36TJ91a0Dl6al8mLiqNltADBOQCjfKRoUCKGGe0FgZ+wkb9
I7Mk3kU1erLveb7HgGQv8r1upOgj7WIazt16ZYTfaHzQ7VgsuK79PgrPUGV3nPju
Ut/qZSXFBPczMCECMPfQbo3orLs63Rh9M8wi+XlaSbONsWtFrJTxLqkiSNX0BYuv
voOZm1zYRUhyiBuBSwV4DpDHJkNwSI7Qgk231Y9H8qYnbi/jf280Q6I2wy4Olinr
JVkd1YtybsOhlMj7WoQzdA9h36i/es391EDRYzhIMJDp8a/GY1/CLpxIQbvKPkh0
5uqiPokpp+lERyLMI+iEUVdmHg2/GiJSozZaeDSisgwljdWuTwG+bs/nAE8k3Xto
zLLd7hZTk6q4q5vuyNoB5nrBeSY/Ak1GP+ruz70UoWqvJzBEcaOsk3z8SSo+AGtc
GorLVzPE6+UPO1CMS4834MPyH0T+/qBTw4BW5prcL9xR+DZddpFsOdegI8vaBZ2i
MHtotrGjlaGJCdnkZISIXjkDbXEcD5S8zljG7Q8zDTE52w+K65U1kkYrI/D0ql48
wgDuRYdwgpC7dURxaWo5FRIc5BDFxUOq1Z3VegNCZGJmCUPzp2m/V/aywESk6J19
IT0Ue0blDOe18y+2umcCa+pSj+XpH87SyfDVnFNsOoabXEZzMaZ+bHP8Q0rMmj97
3OcckCs5WU0DNfGHSTYaX0UPvjd5o1xTBpkQaBNkGkd0Y+FHF0EVgGf2eyPPPUgg
TuVwhGAZCe2dfInCUT741SsgztDBZnhqTpPfMUr6Ey1ZrNMDlwGZZQoYU71f5cvR
FSjeypP+JNOZgKFegcShSCozmjWZQ3vGTtqGCbEGVo2UIAQb+adrQpTVoyG5Cm6s
GerhX8SlY+EbteUt/pYAV62YeYX5j7EH+lXmJJaEbir5v7H+0sx+9WlVuFbV1Ow6
dxGffYU6fsn2bzQocHPpsPU3xfV0BhBfOHe8eZWztIH9CuP8O4cKvU23A5JF+BN5
mvsUQNaSZ3kkuUcycDg405p+NvVAVKJu8KbMIRZ81feXBq/W8MkzTvtJN9BO5yRV
HJFWkw0vR5GTr5tYzlo2eCBN1+APPeq5kPIqXHoUQgbhUWslZ2r49vS62bcCx3OU
bQk041HOileXLxkiPXhzRix1X8jynn9BhgO/uE+Ufv+FevL+dXGwvSaUEgaYhiQU
Pbafp/LKy54ps1zz34/51kJ1Wy0uCD7hHKVZzsQthTpG8ayFdE1NSEjgRGQm9nrQ
0EDW29kEmZENDYA/iIp51QEh5rGLC8XhcdhdHtQQjM0NE8IVWNwV2YK47aN7dggj
h0CdtCaCv3zBak19UpSC+duswCOV3m91e451nwpZb2KqGtH9vMgL3vx2ZMA7eKZX
hSk71EnOvsxvzqTTrfIZkfv01rIFUzJM4lz0bUVSs5GXwWiyzpM5UE9zhexByoWH
2344Bvg/p3ToD+zI3zBz21bQN7R9RJ0uZ5CUWakjLIpQKbsZkN8x4NWzVp+bkEgv
9Hh4EmLKBzqC1dUBvjjFaeprLdAIUIq+8azUtvfUJowXkXBaSR3LUGyPcl4TuCX0
SgfJqU6JMTeznoLUvwt694x/zWvmL3weH0vnrwZpDvxNXLydnpufQNdfWJG/KNQ1
VEwtncXOlvEeDohfhAbA8pfqfTSDKH7XCEfZp8KqkKUzifI1yyfvH/6693TpUd72
ycRIoX8ZFeAEF2vNfqA9jFjCzJvHeXJjQetYMoc/3AhVUcl2XsV8i2oxdvi3wpkd
FYCIxTPveMLWOfjujq+PglCOPr3+0aubkv800No3S3hvOIJswFf711DuD0bXaMAy
0+BYUyqeo+rGfH0e+mWsKuXuJ/xYSco7M2GFZI+AI8sj0ULW+zebJ8IWjx7nInWL
AsTy6nwm/gUHD9QcyE8iZuto9wEo4Yfxm7yM6szVQEOmPNucSwAPmU63xvB7Hd+t
LSYh2oIX2olPjdgctXvYzY+Fs/XZP7p9h0KYv/6r+rEkbVzgBxY0QzeTiSZ0hTxV
1uQ4QRkrv8JGNVCrJ5UBKyX9kSOkjoBVWi6msUq1scDkEHtGchU+Z2EwhlzQB9xA
aSwuyFJqGJsupyPMwV9yINZhZoMoKPOWrUOoiKzOHwd9LuBjYhmTzidVZ4CNVVPG
jc4D8SOZQxvk9viJZDtyH1jf2NU6AIIsyQr1qdVQDQw03ZjA8OShGSV5gX+veMc2
01dQ/9nD5F6alsYXAqkcq24ba/3Qyli9Vfpa0T7BSZi/5gwWnGyrraUbEGsSY8w3
tbyhZu1ezliQWLriPSsuQZV+AhR5WQ0kGmT4Pgh+Z8AS5Y5kT9/3ZwBLNzcjUDGf
PZeAppa6ms4O5Kiiu2/PE4jGbOZ0x84R8zNSfe0gzMunEi3BO9FKQ6u5m/EtbVvB
R8XysN7uAuTCs9/W2hgh9GPTQ8pp920a2V5FlcF3I4faTogrKYdC6nEUXzPxIcub
CrCt/eMLCIRUzb5np6yi/4Fw4dU1munhmQYVI12CESsNi/Yuj8CpBEDqhDeXlEOl
FDuqzF9lo5GPWAfcX1YxzHMHNe9UzSMy8G72cL0MalqGRpfVTcIaldly9EqaLyoV
PtRaZvUzDkoVy3rWqvPngK9VjGfDIzD0nuKj6A03eq6x8dLa8+uQrktl4mr6c8WL
7DGAuHvZQjgHFLdUAwtJmdDHRuRCuMOX9y3RjHePfTioQo95vZADjHyt7yZJ8+3P
s9KxwD81sENvbQmsrxM+0UP9cKfx+bS85WcF38hFNvsVA5eLt809pLqLN+coIMno
8IZ1jLvN7e6zYvHeGa8wouR5DJl0O2It0F76EQdMlTPKZbulACHMHkML4eyvXqF/
Rea2HgZHXwJUxlo8XUhBRpNx8Kcsgblcd46fSwMJ0pWfA6en1gjZGNWia3s5F/bJ
wXinNxvJ9s3BKTUjmPEEc2Btn7Q760hcrgiVt5f8bDb8JROLKlBeX2J7fY4432Oq
hTGex21TSo+LWNz1z7RUi4vQAO0bijs/UF8MXH70mAl2IVHt3J0hqH3tDo3BN9WC
l6AbhodOQFZe0wMWkHCt2AbJQ1Ms/M6VfLX4WBE/Nrduxcr0G0EanFXSmTOGalJw
JaZVRpqqG3/fsoeSvVRWlcM0Sr11adMGnhIZeOJOivVh2fYoH82wPITrg8eXe/BM
HmrlWq5TCAWwVc3dPidlYPYWtSMUhvOfNU3AJvY9yIxlDJJSsvT8XZBs6y5qAmwB
6CeQGTpIsULI3023lu9wSlNRLu5iKbVQHWrhfxhkbp2u58AsnTG1oCPSevxoCROQ
dHB1Vc6z4pg35yRSBrFQuoqOCjMEWbrKDfnN7/vdDtK3sVYbuoebBbG4orrLxtat
vbHoAoVTIOnnkYFeYBbhDfiAHflGYCnIOpAep7WI3zC8zIukr2Nzy7fdbOWci9uL
ZJR03Fq2llcHQQl9e1weX0H2//w+DYB0sBju+8qp+NKVxC7WDg9O+wWXJSsJM8Ko
hOvuH59KIZas1MJ9PZqB32F5Uc4t1yeWsrrydCceZHV3kebge17xAPrKhBZ3kCHa
Pa4xARLgu78Pp/TVgowpOwxZYFfHenEpkIyHSBLMMlsMJ92Bx8r5nIz28aYqwRIW
Np7A5H5rgauHTKeKyuNxbSzT1HZhm2gigtFtL74S5oN4CYZvM3MbJ/VpsHCUSsUr
cUFh8RjmlZtqgGKULKv+iUzNFrCifjSsRoHaq0CoQTwemzphYyvwZk9QBorSjNdl
4m49Ta1L1NMGaoiaJyDeA1k06ZSYpD2nTbvqS+6pFc7yc+2r7KVYyQA31MMFarkz
miJfPTVD2qZAl2KLecHR0rn0JNXVNmxzMbOpAnV2HAHNedpOrKHZlGJzzNG4QR6A
9aZRHCrG6CImeoFmXOwxaEALx2jL+T+lYgylxmwPafVeu6KWn+C/A1FS9X/IU6Ei
+tgDC+gIspLg9UOxTEiYkrB15R+loGvok9GINxYJRg1/56IXSuHhFnYRnBy340fY
Lo0TKodvfPg5C9jc+F97f81jNI4xk/IlRzBlcLGfh634z1whhMjhrXwCqc/YhtLW
BlwrMvKVFkMjhsQG1yKcHnbFITFwmW034aCKqwz7LYWPe9LKCNYcv8YIVkm7/AkG
z2bGjJ2Lev/TYIDZ2ukFQIhQ61RN8yC6gnH2dh1WZEZBbteu/pFtBwlhvdWYYMKy
tYhKI7HUAgfrY29VMf53BFtf15surSDMemkp6wka2osctT8rZeaVsd/OsRGKGkX8
KWX/Y8R+7itPwGQAAuaZ3bCreaaFStZ4wgHwmjC4ykL5NZ+THQsM1xNiWOVLC1Zv
A6+N3VVFGJy59JUWXmEe4GQCrXftLbkCpjR4VZMZRsFdtgh6thv6OYy9tVBjuQa2
BiZGh49jkzNv1DV1n6IOQRmqh9BLUnB3fwx0tp7VUpV6SI4FH3xqNvDUcxXktUwb
3BXCo1vft3FmdgdfDRIvAAngr8T1flKesf6BasaFK50Jz2IbvOazbdSLxyw2Pr3G
hfmtp4g4U1mpBAebahZ1TynO/nbEXnS7QK3sgLYePlh8Xmk8hgGyRyaE8N2RP9fe
CUwhsViNgto912ndyonMBI5j3PGjhop/K8tRH3FgI34u6i7JYrmlO1UbsaarAgK8
xjn8EMR6eFSVpSZedgUKbv8OhlW2e4MNwUR+neIZIhq9wHis+e0LWWHwS6EYSmkU
n1LYg0WAznAfOrMEGPkxE1CeeNbhK7H2HqKpxFIjYIiq+26Fic24XA+gAAKYjdh3
aKJwC4TYZVgAKrWYmQXN1H83Nkg2oo1MF+6/tU2lP9wphnv9htrx+0iQXsvtDSQD
Z/Tfzkwp7B6P0+lxi9HTYXGm/kFsbGG2Zf9u0rrpnN9Yj/bYygJrs5AB1enYzHO0
02TGpb8kQuTvR0/SkXWjXdX50r4OPBPweWm5B6nhWdG15K9ZJ66aHHNPfqsg1MyC
T5Rg1ZexaEtumEKxYexC9DhycNziVwOp4/jW06M5z/T7ZBZLjXm0Fngi15FHXnmx
mXEHraaHeosCIJeQUMzjd2fcwaxQE84qnA0S9UNGD9mtOXPnDVzYyL8Mx5OJX36B
nUbBqowNs4Ef4H5W0ecJ+SkS3o7N6RUWvjwDGMZdTvH1iD7hgT21zA3Py/ZPUbah
9AaLtrADFUyA6vnxolWRPYkug48DA2XLC9cTOMPwscH8e0ooVGXGHnhhqc6kSKuR
AouIyglRO1U3Fp5XpLx4400srvDB2gZZ9vUkMgMOQplxefNVEyFbEM34WefPl47V
FN4yel8kkH1k9lnv9LNudjWndzMmHaKonyxez5/tKlW2r7H7xMHVye+UrkaYaf9Y
UsmBny8q22v4hzSXy27hZfFZLKIOF+Qzyr8letSsMTjZanIZbdwOlgoaB8dkF2Ll
rqbulHmPBE2evqsJIbUBq50/s/8w+i9YQ/de03ltBndKkPcvG1Gc81PdEd4OI/Rt
qfoAOdkiTbjrvXtBNndhzHLXKoPn1EHMAY2LumPSbkYpZ2YfRRBGv8lV7WJYmc6Y
noD+R2KqT9LGxQVOLY0BT86H4rTQVnxa26kIlhVPyRj1os0Wz0HdoC9mgN0LJMu/
/dJhhOZtgCdXCuKMKeKXT9C7+q24LeWEIHI6Xu9x3P1sT17XOkj60txo5kwUg9eF
KIb2/KsKbACY07KJRyCgHYp30M8YTeh13cTCSm5QiajWSL7Qv7un3TYZR2lmu7Q+
i8gpFDPGKr4vD3r7OzG+Y7Rbv5YuTSujQ6X3tZr0s7wO+Z7CPgmkNANbt0PqkYEB
iUgI+ESgpJs96l7YD5tq6GTxa7F0Iq+7YYgya8e74UsXySdPXAuvlFP0QwWFx6Bs
jk7NaVdvumDjtRfTandP/JrN/Vb830NNTUgC3Tzhp2OsCQSwo2p39LsaHwwNBA/p
fUXMi0smAKbPCQlTFiauBjsfGl7dpbbuLdQ+zsmw7SvIAJwJOr0opo2eXT8b3WXg
Bbvi8DHguE3dgfdS6PfjJSf2G6BmmcUts2T1icWZP0zh6O8keIfD39fkTnlokvtY
pgXy3S3RrvjdGwlYd/bLsUS5dQMU5eR7L/f0d3lRk8TX2ai7qF2IfvGKsg1LmvyQ
NMikJ1UhYnuEtJ13WueHPFNhv4TtF4sQPKGNxZXwGzg/dT4bhjnoAV8cQIpBu92K
Bhhx7rBqwMUGU60GlT5xUJbotg/DOX7TYe+2ImunNlZ4rVy3A7G7NvBCuS1cu9Zz
u9jeP2w9NfH+zZaH7TBkgx2Vyd/sXthCUtGtSa7fhp+aIR8VkqxwTy60iLUu+gTY
6aoyRCBZFAamlo7opd+u420oswdiJcPEJV8SHAsqT3P3d+qzgo2XuM5Yj0jZ51bo
jetF8Jn/Vs36CZGuq+XSm70qNrNX8fOwmH+8xHe7EGHAbkQMB1HSO8e/AjjiGEOL
jLJ8u5SfSfB9COQNvpuS+skXBN944/VK+X1URTce3O2KR5Jms7EPfIANUvyUuKrD
uQ8A6SpPtZj4eaxD207jUOopPxNEB9mIQSdcNsFNKPhGscyrOcdCduzNfLnib6eU
J44yyhtbGpOpr6R6LugiezkbZWzRlH3E1ezNnf/KlS4TQKcb6lAWVU3EjX+sTDQS
SNYsz63xEj9kXT6J/61TOZ15NWGjYkrAZa+Tbb0Uj1x6hJqcruIfvsddb+/ReZVQ
veHH3OaurYuTql3J1r7F442k6lGYOT8Urt8qPbl2Fc+sP/WNtiXM4KuJWm3kYFcq
P1W5VEpmugZxfW1bKsBC3G9EBJIxsczvxW7lD6gUNrvrLognmcMQBuhr3ifYEmA8
2s0NyD6DWMqyiwOh7N+9ViIc3UOmi50QRFh3hSJ+ACJci9wJA8VvhASs2cH7TQdZ
UFV7JaiyE8VseKmBgO2NVCv+AZ8jnRda41Z1cpemn6qu1nRfQFI0jnakz/HO0jEz
bAvv2wXXuuDEIqX0Pr+iFwJDdHlJfHelUpaqRlSRDB7uPnCNh9jrnuV6hhpEIO3V
840up9OGfi+87M5OBOrM7hz231fMavx09Ny0Jc/Kw0A0ksmRRZ+nJWdHvvhFGcF0
ZFu3xXQrrA0zPg6msd4IjS8bByNKfsEv58EgTNEN1m+9nKJab8xPDXaFD7etp5Zk
ajaIbLKhSgNk5Ag+8XlWs4v2fd+Cl5kCfuT4aCGJyXsV7w2OnTAZrGM7pmtCI4SZ
ZqXQGjBnmfHW2R3eBxkHppmUUWOmxsthJKukp4i18L4njPellSZR3/W1GW/xN0Cv
phZhwM9XndIkoB6/Jfr2BN3JLZwRAOjH0w9HHbDF/KKPueVo1H1OtNemnmIm+Ju2
WrCZELF1p1FNk70gUEWjnRoXviZjYKIwhKn9R10M12xUo/YF37V0udJ43sSqnZqn
h254YXuGuDOgWRHf93rg1+BCZLRgFI5B5O7E8Wnb3NEXstcf3WGpwdcVR3/UHxdF
Gih31APkGx0rfQtVGmoBq2alnT9a9Wj+pVWyBevvGXAuxJ+6Qgk/VPGcxrGWDcrM
EfDwhwj8glsq5Fx+uEpGaYjnpW52uYwjPTuKM1eMSTM5ZOm0ZsMkUrz6+hfdbrdT
HU8CxCm0jBT9C6iOILrsy6qlt8Ysj+RKVd1cENiC3vZKiobdnyMvJ5bOIdbZ5ihU
PtaMgpgtrOAxjsvtNkiEwQARaNOCPLE5RAkMwRKP1gde3SOsX/NMdRSoWjFcklG7
AdbNxoX7HApAQXs/iRj8HiJs7RUqrvlmn2mQiR+q+icgrBGWmzJbS4V3jskvG80X
MrZz4yKhs2XMVgTRPW/4RzCu7qYn9GS183bqAYJkKFOEusxZLvh4QyeYAkjoqSPC
Oz1H5gWiXvQBUFCxXOsneJSeF5+L3/jBHd1gnYB94foklRAByn2OotuLRNJfTyyu
+jbk8ln2YnfpNHPfKUql7qBRTE9GvEWrgHwoEEd8CsVCYST1WyPy+6p6zbh5O5Bn
09pVB5nmYGUEZAxUSCEWPoMGELeWd8pQ6rauAiOmRP8mXjndQPM4PpBefO4lBgpQ
f6UanWa9KJZ2LZXUxQYWsQXvXxdEiT6Kv62yt0It+sIIrSzaYu1BREXNgAWYyXHm
A1MVwX98WHPhDR2RoF0Nfuz9b7Bl3hW64EPpEy2wZPzZyAPXGC+jWGVt5ikj3d1I
E39ElcB37OUxOp9szkEClFoP9D/rSWuK/sUxBX/Ps2ACfwujISpphNtxr0ET51rY
MbenjG4RWN4ojZFpkSTbX+2QqfpAxKUkPPz+eTonWtI1rBr2Z+B1IS+FRzichfov
OU37ud/HSi7IpDVIN7ctCrRlKUS4WrnaoUCtkpilnlE63hKZoupZoZbngUADfG5s
q6rg+CkoE9aUnX1yOHUst91Aq7HqYefWUMYvHUzjExOVVUQDFI3pk2ApTZoG5/z4
zzvv2S2ch5oC/aCmuRtedIfvMEoezHnPxzzBjKDeB36wSJ6r3p1d5corL/I8JeO8
/TMJ+DJBlSO/9nTYPJpUE82jNDl6uNMlP2njHQo1YQO5vu3F1asl/L1ohlIpPG1e
q/UucLpmZMM9BweZWh4DTEml8FAGB43TTCg4RvXjyCrAVL+gRRHvMzgpN1d0pLY1
Kb6iEtGPftTKG9QG9kCMnUHN5ZnznXPJnAIxZMRVNq17704Yo8+DU+luAjaYMCXi
ciegS+Im09dWVR7uVxPunaQrlL6OpuFIeZh3KQjzqfUPSn1tpv1kvV4D0e6WlJ1X
OttlczfiK//1XKGXmf7Y2uw/K/87sIJmkhgr3mWsUo8eUukzpYHIw6oE9v4MQGkO
+KEQzH/jFIYaA9mN+Odby7/JnRMI2cnzM1+dHKQIyFpSJ4ArUJA/fMK0XMiN9nOL
YjFua7rlXFBIljP7luiF/kBLrGugPT5s6BkBUyUhklw2yLKptOAaIIZotQSqIMIb
CoE9tpqChvEhKpr05V7HKK0Po4eCxTjcQ3ZdhKua6kNcLm0F0G4cruPBP5eJ1z8F
3sDR8bCY7pkhHUff4+Ejc/mma6ZrlUg0f20cBZBoEG0XTTXj5SDt7Atc+KzSmsa7
hv87KWK7pn+UFZ+RRBO1Zx8XRAxXtyCVWJAo7D5ccotLeH6nzhzvuEC78t9Z0heK
hP5Tbne6q2HJAcVe0Q65I/NeyWlUtbuk+lf4je8+xLyEIKG/ACKBfvezb5y5JYCw
QNmzS2emH55VMui/ELikjRVMuvGbUIWs99vDaMVfnhoaPIPdn5e1HqoTsHp1RXee
Cnv+ztP9Rxs0Pen82X2S63G77KvGtj/6UBW5V+g1idvpT/9zHxeD4127i49xB9YG
ZU2+Aq5Jzf0ZOTH3l6TnxMQHeWytAYC798p8entAlFrWZPokNXSI2gwj+90J/vBN
rjZZlGQd8wXTCKjO7hnZZ1DW+/0a2HqJmifpsKklMk0Z+KlA6DkDhPETdWtMvtsO
PPiN+hQaUbK+TbLp1kF3NTNVx7UBmmKRnsvbaYDINXocjODkT7zCAjXPZUVoiluB
TGFmBY/vyI46Xs5UVDTEciuw0XCmIH6s+ZCmNAJC1fny139E/PioOOdt3Zfmzv2j
RhxlJgET+G6ktBTU3EK8dRKyDhBy0PC+tUpFTw2w0BC+LhgSsKpZvw4VY6BF7g/a
KKkzAHMVU1ngMbSib/jEDyFTPfRGLbm1rZkm5SwOWcSBqujbF0frVy/KU1HFzDS5
GqSa9A0z15k2iB9szFbCggQ7iI2hkbiCu2HwY7mTU48IQ6y+nl0vIugbRNOEgyQy
78Ygrf0c0z7V2oAA8nPqWXnmhdAohYqXLt5Rk8Yr0acMsleImfUSVQ8jxAsGO6Ld
G0Ily2ELnopu2snCK5GHCWt7N/Gusfob8bu0uiDtliWp8dpiD2YiaEq8gu7PblBS
LBPQGxowwRcqsOvc/PYWxXlCt7e5hTgHKO/3cUl0914vMIkcZO3zjz2ZVQDwR16y
5OEi7FPgnmZL4CEFtMcQRduDGbuMdEz4keAfGUBg6GP2EP1LgFaHeFnJ2iM02JI6
dJOUPvz7fwJjJSytzuRa9OeQpQUM3yeOxSghg+xx7fj9hU0sb6uxyxxAHTdUc7yE
HzN8OIjOUOXJsS9vnIu7b9ja3+c0rWHG7Mmii8WeqB50XDnLGDvfFkUWGE0EHKl7
F81oYjCl0pms39uLMmIlVgab7C8uyIA/AjpiXElz3D29oIWOYyK3hd0wR4NiWk8Q
Ah6t5ZzBhP6wO8B9M3WPh9ChRl5rI0MBmiSe2UeAl2gxr4E0EBCFgSfNdAQIZmU9
RXm7yJfgMVraJ3BdO3hlLrs6DfNz7/wpctvRdaN60zYorcoadV0huqP/MDM9kGEC
7jCTv9hC334KwRbV9L2tfmrvGtDJh78rUXc3HpGYXl7L+Lj8DdQ8cE7Prft1jEW1
jWTxM/nbCByXMpbyyHbp5kehWZmouEsm7Rdka1YhmZpGtJmURl3nVhRGzTKM1/ET
c4BFEHY559/s+5hLeWrvgLRf/sYyNybX4qCT9lbY5T/3+IadyIM8whjgufyUWPJN
RxPC6N1/FVD4RtzYdYafqkbB+bvmyOMvHiXkaiG1M/hGacG3vFUTICEC4Dh2foZT
Sw4CSusHR/iZ1rb86l7SoXK2+iCm5h6iI/3/80/cbdTuvtCjxKK1kkmbDhTkqw5l
tFIu05kbbMwJcuqnrctMIoh0fQeK381fvc4YVFzlt8GvUdfiqJgvykfRJQ0XVtZ7
L2Jj1rcT2Q4ZmhaNLY9dzyPeR9bK4ccFSevzcWpGd2jomwOtLc973gDMZASGQN2w
kAuNmOErSoMP+QttAFUUhsUGW3kiCA8aES4oh8RjVqiWpH7Ffcd/zfhEJXI2vJh9
6pGj1ymTiTOEtBcPC+9ZpVn+Qya8+QlzpjSXZtxziW4U7nhiK1vymvSzWfXSDxsr
VJho4PTCxFHo8LaKA5auGChB4REVVWwgqD65D9QxvBAMgQC5odCdRkDaSj3fdJk9
eVwEgBskLuvFx7XpJiohjDfbTt5Hh7tvvJPQt7aPDjdMSZavr47JngggOysYKw6O
ubjB+/bLzzFlBqbGtKfvFgVisAIsNp1Tr/GO7lTfNHEVjCVH+D6jVnax1O+WGzRX
iqTwfWnQOYn9aP92KyylbzVBnpKhp8KNUcImqGLhOz1LAZUmj6jr+ae2iaJvdQW5
rZyC6KPuihNvFjlT/6sPf/0wuYCF2knCZMtP3YSzPdBQuuhcWBQLBlQCnQSzmLNf
hEo1ar4k2CfPrxAFDmOE8OrWwMu+nvwl6FZUzA3SgHdQgNa6Ko4LOe0mzeEKBkO2
iK+WEpJs28VKQIN9kAiyNQDWpNOxhuvnZNA0VwAmx11K7RQ+cpmXuwE+S5RxZ9HF
gkhabKcaAqJRDvs4oIqV3vgXvNc191rMEQyDR0PwkkwIBDPYdA7SB/upTFh6QhHO
CdsU82xONsFY5NwVajaeIBp4R+AlFWtyQloMSSG5gD4+H3d12YoshWCYtZbCg/Qj
c1v4QJHLVyIWpeA8e8LCEpBOAw6dX60qUfxbOldvSyyxZAfJ73OANF/TF9vslss3
JBSwbokGq60fhYB62LOv7aHTbPEu+0P3tDsKY2cSCBaHBtas9IKxH8XT/4IzwN6P
5ioD7Xjyg8svsovf9K7lknvKz6FBEHAxjz7ZkYzPsdeTZOdAtj1t9S3aKlMFHuAT
Cx4i5DERJTct+ZdJ/IM/xDjhRcIV8GXwDa5PJEsrMK/jn7CyZSBriQT+WcmWvBE+
CWx7weWnbn0VNlQOCL+yrY/uVSf/I4FhBHmYJB09ymivKtk3mnTgB0Vkt/d2w6qz
wt0Vz2aBB085pyoG8v1lSC+O7QmkUVpqicjl3deKezhlQyJaeZ5FzoPjLMlXHY45
MbLMc96U6lb8egkoSqbaykfFw9lQ9z1Owqmz/g23/IlIfIgZxKNQTeDu47XV1QV5
ciByVfsCmTNTOoLqwao81jMyqFZZ/pni4VPeE8TpfpEKJAZc4zJXq3W/QyAsIHZv
wwtUD9uUgjPKboS1jKxWky/YXNc7IyzJUsCK/sSO5WE50PXQMa8nIH3KxVzAaVh4
mchV5P0iYE+4dqq+gJ6THU8B1sYZxCoQVeVFI2GgLOq2Wuj64BbdIJlhrFoa+WGc
Q5Z9fyBB7sq35s7fRWj1zyBX3T1dGkcw8biVWqlh4MegOgolydbAsnvO6P+HUExE
LdpGF1gLf69FyiJX/pHglUvZgYCrTRfF+inCNykxwa51dqPwTSpCrFIwT4FE7F0W
5+TVm8Em111+sZA6miodc9UjEIcN8wwIMlSmSck1bXtSVJrFG/82lDjpU9M53sCy
dI0nuWvhTNPubArd+NswPBu85JkDY833amPA6EXBNtQW3ktsYDY0FaAuCR6IhiGD
/o2bz6cSI0wXpI/TeKSbZTa+JD9gD0JqGx3GCIPBrho+PI8hq5lo9FXKDaDnlZ03
FoQacC+M4boTHXghXYP+oEHiqmVDQYSB7k6WGD7uZcGXe7R4tHxxc11jamRGcHYd
bChSmFbLTde6ym9ik4NkFi7TdU0K921/j2wx/BY1OS+S8BartuPYzcPjeNi79EHL
n2DlBzJG6IF/56gHV/IasSzAmw0n6Qx/UqnWGL1SIaukw/B+XK0CdRoxnsO/IhI9
luIIyPHAd2/3TRrWkACnodP10tkqBYBJ1fxXXDtx0lo+q1wzgYmWl6qseYivI1Sx
Fj78KcrABJXo5K8Car1kjjd+6fmpe6HLWE/LG1fyhjmjdMAgCNPz1Xj0GNgaKQZX
QzbYWqlJH3NyE6eVGDWlJs1m8ZSBizOGqpR3A7NYDftAwqIQ1eDljmLocBXj+i0W
vb8rGXPRqgebB69W4JPb/z9an+I0andTRziRAu7KLQs7etG8FrLSwDRZZHZ0GhGw
KWotUzTNCp2nmGYFMctq/tIX6AqF8Kl4B7Vt2RuhEnnYQ+fL6V5oimjAk4KqCNiU
hm+xJ2tcIVZwZAJXbIJ3bjX09R+mkejt7Kx+aQXqveAw7LBLYkozvnWaLrf040Ke
w9t6RTtcAjdULIPwEsMbCrX+c3uWBnSez19+G88RewY07pOD+j7k9P3i34Gcyn+y
HvLyb0Aj8Oj2sUpAsRnunl77Jcx76HAZuuqrVD/v0ft5XDCcKgBSdgr7WkcYNnk/
ts8lM1M5hPIb9H4fbz/32VrGcRIa2F9gEUt8p8Fi8mLULKaVjQWsaSGmknhqE/T0
+p449pQyA/1ylqCCYdlvyfrq939F5fFXEyy6o1usOWpqquBWTu2KwUSkbr+KQVW2
qGIX7ACyRgD/Cg8IAbQRJeF+/38/WzMJPHtV2VA6u0sTF9Ltl8CqL729VPJ05RMp
YK7gSEaMhv+bShyVHqqoI6AP1MUdickFVrE5376lnv+UkVwYK07ilWVXDC/TW+ch
IYHe1MDZgkAHqJdhs1cXDEQqlzX+X/j5+9cSXoLd4Q2tsfqKFjVkabsJL/VpFPV3
Fkxo4kBI+T3RAziH18a11FlcN1w5OahLLaid7OesiH4YFIsm45DHuGamb24rAuQ/
fIgOIfxzgn3/K2AX7tPCH3xq79xLpYjXm+xsJOvUofWaoTEnJaF62dZyBBMgJTiS
LuxDFr8fMXqNPQo8DF9veXRzOzDzc5MdsvVBkOBM3kw5aXYvjYlBKgWkJruvW5dl
u9RMiCNI4ojNdtlXzI63AoxpUfnTQksxnPngOYGbrq+EuMOPqdevsTG6ei6HYzQG
yiG8mH5OkYtRJx3iNdCr5s8UQk8sEWZ1cMXAJdfV7YF5Oc42cuBabK22iGIEoU8s
uP9E8/l+6W9HniBTSzxjAOytGq/qazyS8kDDj38CCMDVGMJE5PSB7begwxn7twN8
/m/TFwTzFw7YyqBWCdhV0jFZlvQx1ThTXnYYuT+ajkY9rS8sPNbsXgP8liB1F3vb
0DY73c/7BMH+ZD0HPvr2eiAyBpHCEywl1IDzeg8tM1tihPB5Mvwej4p960QKgYne
B+shGDy7zU0xy/ragiNOacQwlfXNjtC+kiieRKWRjlz+w8WBUKi/ifTREsPXoNgw
S/2Z8V93lSd06IOPOG80JDKf7CKhJfQEAP55XDC64lYSrQgNut9FKdDLl7n5t/n7
laQwrvQBNQaTYm1Gb9F8+EdA32bxrmPO+9UOLjkP6hU3GJCRoJgRI3z7/h8Zpr87
2jEjwkdyArxkCVvqOcIdCqLIfgSSahk+EIcAo0pC8MT/oToiBLXoIeVUz9KaHn5D
HJiv+LroQq7qR22wVg006hJjvg6L++JAQNczJKoqDgpZKFV4kS0QmbmiZw5VFD/B
yqwlLnww293u1ux0TseHOOIUe4jhx6xFxkdWcnokCZ6ZhPLHNvlLHXPPdLJqfHQ8
OI423o9wrI9s8kka9VdNZ+0jjbfBQh0olxn93IKyFAmQt+hkKBv0FLF/DbCb3bKr
jIBN5ko/pUuq1uvQNUK27SK2DDbnPkBnUJw+gm7j+tTtg+yUStov55T2qOfB1PPZ
KdiRAo9EBNH83e8BAZT0cpuFvbuzumDkUVv3jk0x95D0YwgI+BOB4j0AcaUl7Q82
otn8OGRcNafVRTINl6nZmhEArsBcZz45SaAtUabNG9+7StWZymoT4t2oUN7Xx7BR
rpPBNbSFDnsRkM222l4O1UNN46iMlLnFLIxtU3cLSiV7wFJVhnVtcQVrUI9qv1NT
Ru1hxgxIgDpH+/WtehTqPJkJ+q5jhqpRCCYOaOY2dY5d5hvzVuAZzmWts4r0rhSg
HsMjd1DFLdOOlyTuQBS54XIpp5gZUAleVR8NUaHS3aZJjf6KTPdfUYXdfvZcWmDG
fEU8FSYaB1rtQRxLuTSpUhdyeEZ17PmBSRj2b7IXqfuZIlfL3T7CsMk0lZgvTQB7
A4zF2dnUp81siMJynr4+oyJ0GkSFL85++F/HWEP+cWhAzQlOsUlhxDH+ChVNJi73
qx/ClrFI2Y6M6bLFVA2gnrSsTwdazdCQOaVy0bbGQ6/S7YivNhPklpDJN6v7G4bg
RhxnH5ZxXyGYv18owpFZ2F8G/SlIqwUU5Hp7vL6O0IphGfELTLtUp/yFxX6zV1rh
VOpsATPpHamy5ndl873CT0yGYz1CV74vtB4ZSlm5BvyvjQtraDa948nhXKgiYUMF
GCAj7qu7+2PoGmQq2BWtP4N4J3ET26YPABGQ8b+BsVBcvuWoXrL396lKPFYwJtyx
yV2VbEZ3HMDBKPEg67MkMl42cO9vt6fcZpKxNMnHDVJiOpy/IrT38KOXV4yJBGQL
KWfiauh7wXkMVFQAAlXKoHQzIcBTst/TjISSnZ7E0E72OY5AJWOQOBQA9wzoZOBU
ThcGiH41fcUhn98giTGXX9Almv9UgAaTNQqBIIgbemhD0ViPOHOGVHXA20M4DGHy
1/egXrDAG37oiBuPLhfPg6DMw4hNT9l8dUChgTm8nPeNkxT8oP04WC1NeMQSBC2E
x+ZOcszNjkGFeCAfiMChzRFMvujQVBZ7woBHQNnWHh86lvgZFLsJCqtORpJGZukC
9SzFN26VdQrGCjPndlcL7UFTeOd0dLaXP+93Gxiyalyp1KElbpz+TogOHuS7jTaA
rJCtlFlW8DTNqfZomcTDJX9Xec+z1CUmpxRSaTFnjLrUH3RUGKj+IiSVuLTTx0dM
JJLuUJA1GNsUpQCEWpE6iy6RT8X42pdPRpXTDHoR1+4F5l0LFKKlX/4c6OY5XIX+
z+C+UiOATy9sPWmnYqh6SpKyBfJg9WIPqIDgaIxWhwXqQPFYvq4aq+Rl0O8kep2e
8JaaZRCsuynFfb2qjELaCg20eCD58K09fGuAEZPqvv9uFoUuv7Tv8BZXe1Dee9+W
qEwyJCV7QwBe61dwW9Ln5ItMQ9oaE62ZI2O4EZ/xRVeO/JtMYGv8n18YNAlybZEU
WR1ndYsAVvld127nOKeaHX/qoKW+2tudcWyme6MpzNxQzYri5U+hTdfAtYuKmORu
Ob82VbwZ2bKVqqaQyxSkPJr9qGFrpvAFoTtKMSw/WTcUQhHgNVnCRPBSOsb/VOeH
R8fdBzkaUU0RC7KuweG50QNeOSSnKT/pOIN+SfvtPZ6iXUpdAAXByT7kkTdRNr0F
omOC3wK/mnxSpBYrUuB7Mnvnebs246Cl5MWNxWRO+azaE2sG2RRCkJ1Sl1oiiION
IrQhCtdhQKq2NDpm+Xswq+yE2+lx5o/AWknSabW8whM41Ccp9qy8ZCUR4q0ELgS7
EqH5gjXNC2CkyyR3fuDYW4C0DFeu4Ayctgwy2D105JzMiO0CjD5ICi7Sm0FDP6mN
4GJBQoKxijpkBWmb3VvvFLtoRd9rDSGFcoEiPfNw4E95nfrU5FzEEu5+cDtl1v5n
bCdQKw1w2coFPd26q9+/DkPFsAJ8R+Lng3pQ5/y5FEyxM23YepxRdeNcUXVBHEZm
tTwMgKaMx1VNeIlMQMG5hspbBkPsbwpUIYW//RK9zhAcUlFKB9D+SJ1QpMnClWLD
TjK563mu+KUfPkrYMVfdw4qHRbmRWXLD0k7fqfMM2XcXl4V/cFD4RJCCXxZXKmWV
AaX33pcfTedjUwaXGPJgWOzRPZKVG7S9iZJFD3ItsTEe1kKcM+L/wjZl9fIrZb3U
kQ34OKG9gFXC+m3UKC+aGnSLcw5iEFcmc2zTqAPlGCYELIChR63hl4c3kAaEfO8e
q1xOrSKvQ4ls4aBDIFhEHEoJ66JktptObk9QYsn08TQsKFTNb82mHC6OuN0EBIvz
1QbhZ6krH+qtQq0Y+RoVlj/DAzSaqZ6QVF/fGSU5EChcX5jHgqhmY1pQazBAZFUA
tdWvZ4o9LxVIQFl54VDrQG1SEVpGeWeKPWSYvfRpCJkfWocPPdBcW52qtuZ+cKU3
7hIfIkuP5NmW3QYXOJ5pU9CxOowyc8Y+dk2MEAs6vhSoGY8RVyMvKR63iIqq1jmv
5f4By1AdzRe7r1zp9BZYRSlcaCddpsRfwKxemDwym+F9SokmMhhfhj24ColT9mQM
wdBUo+d9XawMUXvhdnCobLGEKaw9cnWxIjrFIHKrJixNBtJMZ673KDc7dekn+i2s
Tj3nN6nqumE/sHQB7rKOcugd/5a9aQgEt64myygDtYwjaURbjgRP+XtD9ror5Cq6
P5MJb4lK9XYSJg2SC9BENAvMevLezGCbnq9XNWjxobScXNEjupqBqXxd0+u4XtE1
3cI8A/yuwsF81CzVZfrDf77p3GWdglKnNsussJe11xVOwGy2CgSi6MqavvREBeJY
yUMU7cO++UAgKJwAKSbgitF3LRBWeE5dqXi7moC7FcjgIEM8Kt2V9206ytnTa64y
qj1daN5fAKOv0OkENQP9Dl0wtV8VmJI7f7gxkAK6KbR4mIHFzbWk79WxGBTYUI2+
a5ku+jB456dAPf1qbGfTAG9Zl4sUJJrVjOH78B7I9mwu/kxp2mjqatx8CEbGGErj
n9QWKdhW4AFibIo3TsIYIeQzhAl1IS6x4LhIblJ7Z1BykDmO7m+gBmDkVrC7Il7k
h+q1fe6q3sM4MXsvCgiMs4QWCdL+frlXpSmH9hnd2sBqNajXmMMXp0l3eHc2ijwE
cBozP5Rd1dDAqZA1tDos79Vy2o1d3GI+L45Q5ygtVLSt/wrKL2sOe/3Fx9/e5P5g
QIw5e3Odz8G+nm7Ro1ncc1XmVigG4AeobteaTS0MpNoF1TSFhpzXTCwoIDeP471d
0cEVE7gaTKCpE2xsPmGReEdx80H46eoAOGXB3tWUthHZio5g16WQAsBdLnn+1g/Z
347/eobMhkMffzHEEPGg9H0zOF1VUqKFunptqG9JSI456jsX4jfC6tyEhs/Kyqfg
ORnS6NRjXJkwsBggVAEO2mFly6eT/NBb78cW3khExWJrGuFgS+PYaDsSZLHG5vi7
F4PMfCdpDQpzdt0jQZk46xqLZlKmlIUBwRejpICBRzcDqNrefTapEz4JqaJIZYJ0
jEsilZvEBhJx8qWyIQXOt6VlnNKg3Sj6Vjw9bImxBSw0jVe5+9XRYWRXV7i6Xw64
xS1odpeQ5XmKrYugbsb3xAaHu5eLiDWr/cHX4zwb6U6oYltZnplvmXWaM/udEYmy
qKanYZmrs/g4YumX4rcDIpr+tzltgDp5fF6kO/YuSsgFGutn5c9gDXtpqFeIobUD
ZbqjoYDOuII1KIs+FK8UXgo6rWvEXYfQitUe43Ab16FxrHEQ5IFQ6WZ163Tre7wm
tZvG6klWgUUdpQqXuaHaag+nrhAKiXMlj5yO4gyzkETwHeketyISjRp72umBJSf/
niq20HDcu2h3eTWJe7/PYXQbhKYFDZWaLrdOmAi4gpo6b8zgShjsb7N5Vi1r42D1
+9s4Fm/feVfUMrlY1FLt+1VxcriMXCwM61bfmlJ3OrSy3gNOdwdcNvtO+3aSRY2L
G7lRlcPiHqbpnTzUhtewiwH6uPszcPoEkCU85NKl6j0XQid0iTrxbF6YnmcpsECY
L03bgfnWOUb7ifKTDGkroXqN8ISIMhmVabP3PxMMxUrIYQR3kRkPtmQH78m809VB
md3Y0PyQXD5EaUSqUQNu7JCYbTg7RQ0dCmOnNdcqy2bP2Epb+f38CaiZsrMIhHth
5kbBi7rqMkCNwIdgxhelUldJT4JzUnIGyWbWza0sPZJtbDziErnlpmwwbTAKyz4+
xhNpgbbw7qL4HGGK09OQ72IXEUOJovGjnCKxCM2v2crmMbnOv1TPi/uVsF9fRReQ
z9UnqFc9MUnMZp4mM0ARsZdoMebMvJ8NV/spNQ0hM172v/SJUuhgx1Zr8h+gje6O
HUmFRWruU+3GBXNuo4y8raEndTR0q+trc4OSYU4Nj5TwnP5ffRKK0rDGxB2vKmrx
hAmZrRgrTkhYCNSiPdXXjVwdzYYYG89SUZidxFUxWSbmR28gcWXZw840LfIGtVzn
QgdXggOGDVg3XcjJmFlxuvPylNNmXV15ZmJjP2EC93eAmkOaJ0fL5M/+Ke1//H07
PYqK12SSXLDC8UC0LspfRAosKgXkqgsq33vXgUJpXf96276ki98cpwqNJHJR152K
3NglBOFqWJNgwcRSAuqP4DEQ7iAHcK8b7x+DUMc9U06lZEk8YZIuQWTh523qvrk7
ZyzeA3d+iTumYSKXb+b50o7tK67glhIDRk60I7Hq1ALfZp43Fa0VF+3v0j4NzYua
FSp2EMoZ//dsfyl6g6vt480NSVwhY6Ak2u+fk4RSX00o6uRKH4W1c+ou/77kxz0B
PAFuSgIHjQj0zNW1OSoVkpIYfnKqdVMpvBynI7DrvKncMHlXpejBC1+HQ1qtiGds
SU4Dx9uLlzcHhuO0Eg5DuI1qdSdDlq1rnO8ILxAqpiWnAfo4suBAvLlGC8r4/feq
omDrxK60U1s00z2CcFFhfZro1tisuiUUQY/7NELpcxyp04QoYWn+uylx9LPs7Cxp
PYesOq9V+GND8D64MtXStBq6ryotSfBhtbjuTC8NF0VcmlPsDlFA5zxlGqKSGCsJ
HEXI8UTTf6y46VxRwDge9bo11WVenMVlpbpmbaIAdYF6xnCdKUvZU3GVPYQWYpOr
DD9lSkHgBWT+Y0WgQGY+VQq7XvxW6oRtcdFQ1PVDHoL8Oj2VwN9MD8NGMVWhGBum
J4lV5/SpNxnCP5yN5kMgBpw+MssgFFl5ExbVncL9PAYjXtV+YsTKB/4ItHO9PJqx
hMC/o40X1Kh+gDsgThHHiKS+5UEKHoJx028/Ym7v+Dp+mHdfeUWQGYVKlqZYlEEH
rTMG0DyYdxlIVQ73+h8Ckar3ECXW9pNMAMy9D8YkXL2ZHor+AXeuxuQ1Eympfz5o
XBO3nbk/RpkwyN+3StcYHidDWXS0L/j40RMCkIjtfHp8EV6m/tiS0dVfAKp0IXZT
V6islGuq4DMsK3O2stXFzkwSA2iGIDitiKV/waV+557WmYj+YEXzI0cTMLY57OIl
1DZgYMc1sMJmXzI3Br8dK3i1aMtKXnL0lYqRkEcjNzZ22PHstMrODBTYkpSZvYZ7
B2S0gx3ZO2keMI7Sy1BYVcHUTdK58+NqTMU7YO7f3aYotX3Ty3UJpEfAMpQ6rgSK
WVkQqdkQmH59/d3ObsQGjD7IxzT3Azu4fUsp4yUBY3Sv6Zjluk/S0hgp1b65rzMO
CQoxQrzop3fq8HG1t8Ak2CmwyELr+SUnYGXG35C7gV5z/F1i4dStwBzoSCI3AG2M
rzYXWIaY61tMvK7KUIjq7TfTnOX3ChSZengBWERTZpCeCbD5yoaRUpbon5z5uAh3
5UY49QASKBoQHtkI6FadaASZqG0TWSCTYiEdSglBHuHIcqfvEMIma2v7ueE+45BM
eHwB9d/g7Dqk7ukGDp8ti5zdIWewTYRn1h10ULJSO0g0oVsyyDrkFpLgJZCdazlm
F8oLus5NVat58Xl5EdgU7I69drNW9B3OK/+rbZxcDELyj6eBxt9SrAlyq4z0wEgO
9NWJcwdaEx6jaiWeuP/OCvt8x/1K66+beMw4Op33kBcmbapw6elSTKMSQiM6L7kt
hGRmXoSpHFGjAb6mjpxDej0ZsXo7Vnyk6EjJm4SE9DZvigftX/TmHKkVfZ1eXQjz
TfAjIlY0E1u0skQkj7EGSlFKkheba+WewXKLhfWCqHPLohgkHUI1vp2hzvb3G02b
3iX3Ku4qjR56TDo+OhiXFlXwzd2HfQNBLNDlB6kKUwRotQ3wdEdUD6bncU1OYDn+
4XvWlVdw+zMobuwMgRkcpXgJDKzt44zZMv/BAzddmpTFOg/Wf/yART+EelkmE/9b
bTSee/jNhHbepuD3Vg2W12/77KcYS2A/6T4d8Z/g0wxW5WBWJV6mlk+wJ5IYnBOH
EJPnAQ5ce0DiZNpWU8Z8foC8BZc8EPaKR465AjadgxBj+7XB77/JBwrIBSeDyZS5
JQChzjkb3A+isjsxYi9E0veeCOKwt85ywesCwtqz0N5yfXCwWZRj1TUJ4zBAssD2
9ngAx8zfynOkymmN9kqzGN7p5QU0C8j5KHbNz8tKAVB7II12I4W+jGoWqd8DAOII
HCsuPvRmfSypnMwBHD50ZA4VW3oiTgIXCTFb0nCk4hRjphxFX2CAeZJEPGTQlxM/
YswBm62/K+IumGcK9Z6wA+p8tKrY/TNeP/v3DTgqirCngPMPmM+UEAiWU9diamZB
hfyDhaz0u1Yzq5gutla9ACGr1Cnu0I/Pf2b4eAJm3F3Ty4ep6DAoRX22IEP+3kgd
hT7JNuli8AymdAo2BXBNnYHop+zMtvFVVWS1W4rrnIV2HSB2IMLJB+q8OJLzNNVL
MhF7Z++LH9Vz43NgSc85S3Xwf6D8dg/Oo5tuW9k4RW1VDfShFmDmFJEw6UJTgFcy
HwZUg5N9fc34XDcwGKsxkMCurg4UEAm9Q9DCVJZk/F88Cjb8y0FRH+2MX//NMhcQ
TrWkTBCUPkVUGiejqsVIOkchSC9GdlU70bxYJBl2dcl0JDmNdcsD14tJRWhUfMsD
nuV4nFowfqyujDJEMbqorc9aC4tp/pAkx+6tmO5YKq6pNIsWxJ2RtLsSadTCxFGE
Ss+lKq0gvqT6elK1sBRk2/clA+FAqA1O5dxp8WjQXvXE71Ur0+xdd65Cac2SUC+v
oAN1ThYHyJUVjjvuJPH10t4pBe+sZthp3vvH49JNM6+rFto71LBv6+iwOwkDhFhI
AQA2NUgV8Pwgm71NHLt7fZd1cnufH4wCGEFfsx6335smh0KVb4o5QQOpUcpSTU83
kn9aYrErkHhMyng+X9JUaMvhf0zhbtAIZTf2aiBLu6QAXM4rEV5huUq0YP/TVViR
B/z1yc4k505kCfS5Xusn9YDhOfwYuc/Otg05qVVErVffCN23MvVhL3gLVw0VirNn
bsjG61BBxmLpOSMKfPRRCeYDPEeVqeTxOr/8ek8if5D51SuyBEb64MIDtZccejV6
uZoc/zhv3PmZqoNU8RFtqLXF52tZ/LjTWpHjiKWG5ZnaC4pUgwsaC2+PqndWhu8U
V+QGZODwp0OWvqv1k7HlSH6931AJ4rHMuF0iK6845sJIYYq0P8SxvaYwoZA11HrN
X75EYkZdMP3u+BccaCi7wcvuK/UaN06/4GHBb6L4So7R3Fg2kGVBlHAU5JEux8jU
JIDWwoMBS7nBMf5u4ng9UF4w9v17/fYoEXaWOp0FPV/SHWsQF407GV6UqfOVCGWX
RsVtaw7/3ldciPefCQM+qeSoXlxMpsmKhkUPiIf5+D0rAaYobSOunqKwOhU/toeT
1tJC9ha9to1tn8o2R2WGjyOuAsJ4jqgvLLaElUV8LwfWbCSGl8i53h3qJNbEB8lb
ZuDR1yvDizx6RMNagmTm2Ur5IKxSUPUtwqIDU2ZfMUOyJha9u8uELm8MLqRY57nZ
1mjk0X1SPITpoJb+U9h516ilA8i6pDhhjRN/9JKJlL63pFbtcqjw/l/wgTKzawNk
AOeu3F/4ZrLPaycfiCKkHAcQkW+YbJRQmI2c64EqYme7rgiU+DdVDnNzi8Ss9mbW
fBXIjKoTWFgXLKc7K4QyyhVXWqi2kdE5jaCG8NGd63UFk62hSOesnDVmhK9hPkod
BeBZm8syZbspBiGGLzA5dH5vY8wWQoHMlWf42hL/dexe8wmrgGj5ZAJfkRXWU5RA
8laDVDP3ZDYqCsk6TWRvoRixT4VZr5irKMZpA7KRlDUTpxKEkSy9OQLG+K3mgRkR
pysQS/h1zq9jVnYIBiDQtT12Xb3tt6MCR3TJLjtmiCY69RWvnu7Iw5L4gO/mOqL9
XGrqRDBZvZrBX3FjANMQo8dyORGVx0utgdhDnCOHDmItghFdVBBinfATeIXi2iij
9jlOPVd8yEBEiK1A1epZUksGhW5yDximvS9IZyLB857wA/BldE814/PrZM5NBzvo
KUhXu6+fP8vHZDzuirOqAbsvd0vaCfKi0OpqMURmGFFhKp5Nd4qZAgub9YNhIVuZ
jgf9pTA8373FvwtHXANnJkTaX7qwUyHE/pbw/rUpmYn9TUfYruxjZeJTnEWDH0bj
pdANmMcSHIZJiPfdbZ5GQp/HSm1u5yNKUULQsI4yT3HKQd0is9cqDjJ6GTJ/klm3
1UVbvGBqE6K78O7oi2zP3KdBQaGfwiJcVhCzVA/wnoa8Kyc8v8DT3Zsvv+Sk0Zuu
94yVFI/2BMOKCEZ8fE09dy7tsM9LhtXx5LaxHf54J2Ox1zICRM+4rgEMS0Yo5rQ1
7aBcLlwBsaCOTIxqLvHDy09xnCYWXVcBqZ6VgWyndg63vTddX8bto/9C61w9ZUss
+Sd7zGXwoY4okagOEewqgLiDSiA6fO6RVYeyUTcykxY8jnhIwPotqlWFC3VP/qDC
2e5wuv8b3hFC+Lg8lB8mcxtZy5c57UGW7rYxe3i9KA/S4SVQC4B9dh7oXQcnM9XP
T61l6Jtbo0EYw3k4Zf4lVK94AvHAcA5ajdHpUSK34cL5D8GcBkRHzQvP2nzdpT6S
NWjoooHo2LBw/IbDBdQPqfSCZ0xXl8xxa2vDEsS0vTMYLW1o/YQaFNg0zccBc7La
kJ5blVe0DFGa6ZTnonTQ4YvgA4wvEKPqOCYvqjdr26ld2tx6xB0cazm4fIoTFzYy
iGu40gahOoxQAVVeCyKBaxCSav3kb76Ig3bostc7lHc14kKby36fSRPLFBBqyen5
pFVXd8D5fZOFc+GwBOImRVxZEqw/NWeGcPrOtf2egMkDFcaSiQ+FU4pGyyAFLgG4
XWh8KZ0Uh16xWFHN7n5wLl3q2bH8xAvjiUgrrrKeCpvlkcW1aDst1eQtJvPUre5b
kXP8B5j4FkixyoDnv4NF9VTBgKUGvlFb+A79PI+kGrx/U7G4+vAC2Qkq0YT4kdZz
Wp5BypXzH5kZe5gTefqiK70DeB2arTU6u/1cZ2/3SEdlrh+A1seikKZ1KU2U2Kyc
HpAoJO+akiMMjwKm8xnJd3TX2hsE8QEuSZxX8gUj2cEEPWq0pJzbT1VkqrqP2CA0
lyk4wH80Uy6N9uuEl6qQMahtWlgJ0yjX11DyeQyxhQzNOLPpvfr1QPcNJrkxYfVk
bgVctgL1yj9Wy2sQH/pbg8KhjEjB+rvFa2Co3yzYiOAVK9uk4fpiS4gbAXVapmad
8tpauoYBBlY0Gx356MaJZt6WImXvtkBy1Q5lKMPQMrJm/5hHykGClNEbq9oYg/C9
QCYiXn2dYEkB/OEC/SQTAMFjWVFaSwlRWm/TpUjFbtZWMPlJYGW9m/ITmscba5HI
cockaFijD2gIfVb/i0/JCByEurshH/yX1XBGFztnan2/zyNvEQuooLTwzT/RFH6/
TTkZFUCX0pBUnV4SKImxwOIW19Ca0+UnwsejU7zsvfKszNucQFgte64vvcm1SrYN
Uc6kRMy10lrgtTBR+dpsO+AcY/TNTg+ZUeO+xHZZXG5YeK6SknFR2Ot1gQKtgGud
RdkxrOlxv2b2cOLj8MONIRtG65KV+4oVpothpJZ+sLaUZOoM6C/d7wD/V1jgAhL9
L6EU5JHiyqjz/roXPs3AMQEOV9sZtNDt5k1hTElBUBDE6O+xNWP0nkJcNvhbTi4y
z6gUxRPnK9Hf19BaM6uOrkmizJvFlbO6k43Bh/j77QL1MpfFnkPhV2/eL9s/st45
RmqiVNU/SM6lX7a0i2bouy0P57BfOXkUB+sg0I+DW29GYbuXiaXAOsfHxoK6CQL5
wBJJPrxctBGNrrJegPIBcrspi+fVTkDnlc/OE+WenNJR5SHFq15cqUSY8mGMPHhK
3MJMywaCvLyCG8mBmzt+ZwsWVQonsuW99PBkr7XJY5/htLyoP/7VrX5kzMOp1U1r
NvqasxkUmZXHxSYokULgn3uZM9iKl6UxhAcWfI0MunnrB0stKQhLVqEPzJEyS5yW
flIpxU+sG9FGykVA1n46/K/5Abvx4/LxURbVxXEd3RvERcTTNfCA3is2L/6WqD+4
fqoF+6tP3oeazqsHLPaTaYhJZgrMAw0McsoYgX7JdAWSTcmIsz5L4UrUyB+DvBu1
TCJ391l4touoa50Dp+tWke9+XJ9JutNvGqAcLhZqhTEuYYz8Fh9g5oZ9irjoBvBA
+7cQYTO1bXwkofWk3yunxt9cADWflDau6lIJRX8m8YJFuNSMRmbjcwVMre1KA64E
JcCkL7DSTniiHPbSjhuPdhhpDJ05eldaWH/zZgmX8idrkD9M0yJEF3oQKLNJWO4y
R3MNFbuVu2vd4mQLVjV7qLIWPl+YBqXxDhva6UDPY/R86csVBR0fpFLUnPy+XM52
mbm6AH90KU2oQ/4qSlOO8qTsZ9ymvOIHTq/7ds2JvIyXtErHpjLy4VoHQkBPKtqU
X9Hv+uvx+BOADgVtjrE0Vq6nH5iZRV8wQcCYFO/vQ63w2NTR6+e1PCovlhXX0eiG
1I2p2Rg8775rZRQE336uqQ6b/SMEbhfj+HPcrvAkmMu7Cw4lx9xarJl0/6+bAdIz
Cfj9zyaBlS39a/cqykqShq1DYQ5UTodiNHqXB1uiT8N9nRToeVKCuB+KBzTnToka
MCT4gpd96yLrdb4EoiOHmgFx3dMXTRx+Nh36JNW0VsPJ1n2dSjSfJj9E5EzEFlPk
SPpxhCY2BSNpOxiiW+2AHVyrAGUVk8vvhUIVdMsYsGsvykPuFW1/jw+7m3HFunfr
NGT8qF77PbG8xzRiGyL8OHzluopx91+CUMzOYvJ+mPMH7YT9W15KT/LlI3jw1yhd
3L2vS9ZspiJSlzWCZNWv1V9chBl/SVPmnUtZEGq3E0I5bu1KnAB1pHkDzlmkuCh5
IGvGA8R5Ehp/HUSZ3H41/glJTPbQi37g6n481sObIFsBFp7Z3dogeWHK2SsE+jmM
5kQJiWTUkxd+jA2P29sUYauAP5ifbd3Ip6ZBM2vqHJICFlqWCKMmO8gA6BZsnvSr
Vjau6uaRGLWgfJVXUho6YMyJJkwC0H2QudjC/7GCIhWrfZzZKjoIj/zlug/wftoK
SV2N/Kbq7oYk3CFMSAjRGrP9yNnyoHdTWpWiqAUDQy+kUwW4Dgwtbf9GvqCe7xYv
gwP/PPWA76ZYr1gEIlYqQxfmErKKxC9CBNDsLtLGqJwMmAuwbgFs0aysYkSqTQ+B
N2M5g2z1MAWtHh+NbSAg8zGBUzyo5e+AMGGMpN3cgSN4hShKOyF3Z2nR3dXkmBfm
Ub1BAzLoxtOMpZG7qbaKt/ualV9CSHAn8k+Pucdgs7xs/ncoBxm4xpZnZnq3lmCp
ktZHA/jQqo9dgUO6yI0TTwxEWwdE5AVE06DXaw2eqmwSkd1cZUOjcevLSlsGhTdR
PyMAj8xwV0eFQpTs/T/wDOynXNEGMxDxKPGEZNBypwybuMAPP2/A8aU0n4H69PxX
Leu5vSEkNnupdzTxrpeTNsi+7WxItQu7X51n0sqPepuSEsu3nEqomOP02PCgXMgM
MrVN4bijqIE8sW390SQ0D9SdhX1E7e7M31O9uBMnd3g3EC6Mn09vcHqC+2SsoHCL
fTi4HCFhpLoOAPhiObYGZC8PY0oXUKzUrGV8cnelW6+vQH0OhOJtXd9dm0W+OWD5
l+rM+9rIVOlLtawhpMMzkf6nW1hEK442dlLGhyvyU6Q74Q2yInGkQL0YDUjzqsnn
kuZ01D0Y/dUiEFZykX5W5jaGYPhkVVfyXUnwpxlZmuT0C/Z3UwthFYZ8sTnL/q78
aOHGW771RhF0fzkmnMg0mpQtZx3XkIWu9sU6skWt1MbGADZhIuP4ONV0l4bucZG8
JO9+HqFXVTtjcbmAxfp8sOeh+U6NPzPKVhNUfAhz2Et23OwJjrIoYUTOfkPYvGnx
JmRjYetRQKBQiWgoDqy9FSOyx6dBAiW6bQi1O3Vtpvo9mDhLs3R0L6sdYM4pPrHv
e82SvlWoU71TPRuxr+hv3nRbADpFt1Uk+JdMD1i6HB1fgyta28wLY/5Z11UZisEa
3+lAgT2hNEt53TsAZ7U79v028Ov+jpcBRQF/nMBUHzBZu2D6XiHTwAobaS7hBUpV
nQprXtGW+vddMQaVG+q0H2rrhI/cPe09yaiQpiDgOOaXd+OA8CY9O36Rr1J9YV48
H/6QcHdYHE7nTUIJTUmjeOlV9fAOHwDEysOcyvy80PHgCwgj+CnCoqF2cGNnqFSv
0lfBuwtedKP1+MZeyc6CVogF76IID6wqhhVGR+ucC1NxeDabI/w4BqAsjJ4qKEg3
PEWqE7oOfaR5IDyDqFhOPkK8WwfB3tb1eb5QKgZ1xqDLh8XXJOk5JhRfBslTGWIa
O0HjcC/rVyP7/oB8SZlogq8ArUhGfuynlrXptYfefjG+6yWQgXzsvgOStJ04/SsG
QXlA2vGUeVwLowYzMBgWpEhabXGXIjdGcCm9hhNpwFca9WkqtL5SlDvHoTvzOzuq
F9fWTXS+1veS525PgBwnapXRfcJzJQgvFGdy/3TXMsgBseshxQTqm4YMsX9PKr5a
nnMzwG0twaXgEDn7eRRsm+2pCzkT56PL8UmdwSQQRzBUaq9VlYnGa7oGcxaPADwo
2SLdHHHyeHG2OR2RK2u3cRpMCCo8pHrJj5m1EozMzj4XwuLCVDkrxWlUTOn0/w9d
MZ9PZT7BFAHhcGUSGkfUrK+4uOJVCSJDz39M/MCDh+cSHsE+VidY0x4iKQQ0Z0pS
Xmj+ByTmFURjT4FZuLmMVJHbj097JhWhxMX2F+Z2IblVd+iAgcC/MQoyFTDNuVHp
O8CrzKD53gkMY65rOBkxFyCqAF+e3OaH4mLUhfaMDV7qFDONrcamYX1a7heomKf5
65Fuxs1oFomUDoKHcPQBiDE/U01+3fsW60LAXPOVDlkIbhgNGtW2rCS8q92GA7uY
xtPLdvbBmNAg8sZOM6x4Na8hsMLd4UKtdQzZsaedErS70eVHIJcie4vwombpnc/R
LXEHhMnCGjepokA1I0EByrh465DPF6gzA8Sesb7M8vLTQJWFebc4nK8cXPNha66v
yjVIGOosrQN3k8EoxnzevwrX0NKyhOuUMAS76L2XttYJ9vU0a4dnPLHtnYoAPtwB
K5KPn5sYiKT/0CAFsHZt9yO4hUJK2ulKBPhmC2Jv1c8NETSoNdovBkQeBrz2HkZD
+kb29bcxL+EDQI3o8UUdMYGDNMCFH4dogiNyiWPur1DEMYX65cxqp0iZo+lvwPvs
YQ+i6yLBNI6PtX12A3The7R0/edKZBVHm9igo38mtCyvCkMT3piFfEeOS5cMIiXE
Hj2+SZ5sMZIBhVUDacM743vUzTfBp/EQUrIiqqPluUJfu6C4m1O4prQsD9qh+Pnx
hCqIMyJK3bRJ7W1cls6RhYK08PhDl/As55sxfFHWRxLNNLIQzsaBZxKIAq5aGuIe
t5G0bNXZxz1hrjHVLWJAXPD/hiol9H3rMo3bhEn4sAS77ODYp7WF9UFSLM8BcoJN
GyPNt4xL5Afm+hVlTrYFJkfhKWJH7NkGbzkhBrKXYQ4tjckDhOX5GJ0yvxvGlVgK
7rok7eauxYNvX7v+27Zisei3CYSuddz58Iu8O908ZIqsVFaaPIw7C7D73GC24rom
KqphsELLRx5TmGSnTcDGyRwMB0Ms1pxMGNJEE9UEsHF/WX4PA8x9vVhtjeFMge6o
BL3ezzIcAlMaaR7xLprMevIYjexAuiQBPcwAVn7gUgh9mpaG7PPQIUQJucHJ0WwY
HNbH3zqCD0t9gbzAY565SgQA9d5QWVbv9NH+VlQ5teJHzBn7xaynAlGjRnw5NTNA
noKBNV/X+zK2K9kU1V76UFfVW0jcOG5nUQJEmsLK0B916Khwo/bpxJSqHUuOCRuB
Q58yl4cSrJ5htPeacoibpopKhsKsVL8nRrVQD3C/N0OHyPG7pZkyojrHqdFW1wVd
ZWq9JQ3mNiIPvTbi1p3LfzYnFFUcYhiVr3MuU7m3lfvWqVn4MGokeLEI2kzpS0j2
TuiDjb+yb5tjoVQIeOfCIRvyPozSRWl2r0jgdhxaskptBj+e6fJSLy2Ra3Zc5YBW
CqeRE+OQ856UWsJBFj7kQ44lFWsWHOLH4Woxs7eldfGoPW1FzdVXrNQ2zxiE5qj6
5LC1SxOhuCilCXEKm5VR1vkdcd3rMICHvJdGmjDIwitJzcwYiM00ntyTJt9xptXk
UPrOnLuEFTgHPMS3wdsK29lMWJg/iYYOF9qCjG1pay1E/6N46gG3gpbxTAzEIwPt
N0KOdDLn5PUlU0wW88ZEBSFk4DPK4edP4PmkgQLl2O6/dyYtBWr7Kde8cH8Bh5mA
MIbcGK4SXlwGCihK4tnraMJW5P8iatFZa9WIY6JJWikPN7mG+16rBjpT0mXKdHCR
m4LdKAyeLkrGnL47NY4RmdHI0RaS1iVchRUrHt87mdd5SM/rchOD22ePOaoQzyrx
oTrjwQYiY3EeBwI3gXRtPcWsqqeCDwZLM2qls43w8w1HQ5AvtNXl/pkAeH97BTad
NbDz9xDlekgsEneaHS8KOgN8FJE8YCL++n3P+G9dUEPfiYtifHpaPsx8DHfNixak
iwRmYPzJyWRok2pGK+U339afZVarHJ5JnM1mpfjTaTe5+o38yaAO0wAvr6HNbNJK
is7VyiSJjmbtFI9m/kkpUxbIAANiDAmJVNC4SjTbwusEzJOuVmlyMXyZd0ywGGcJ
/cgWf9p3hlIaDuJTlGmBU2gkCwcZWBxL7ku4Ap+GXK8/zvhoNZBXoBYqC8vH1KZh
gLGnh/OdtLE8L7kFaGan448xTgMlZIILastlyF4R0Z5O0BMAA9POUyIR/uRusa+i
rUJRa4mLtcUnXgT1oMfny4idClThaTwG1tgzGGMKfOAKEfAXXSeMTjdGI8JPu4bn
8s2hJCc65Ejr32oXrNk90/s94Emzx+2jITkWhgXEDyi9dbdkNDMGrGJcnk1uoOG2
a7kdLGkd0CU5wMDGBgWvpve3VwudmCzxh3x6L2uDvxqFwyOh4WMX46RCxjJGX0qw
q5AIxx9WyzZj1dmmPRLXaB9RY1nvgnPB5VAEZJJZkMjqgCkrtaT5v/Jv/6uE0K9M
UV3fPH1eZZuywzBw5A9K4/phiX3iTCZTo8c9JAwSvK2DCwL8c4nlEijBBemiPzzz
I1u41Olt5u2eEG1ymG4m00Pa+AU21FF04Si7AOYanp0eRzhmw1iq+PYHVMudqkAV
L7zKqksdF/0weBRrdVxhJunFrX6OTOqMqCn2bQ6U/gtfTVPplgy6GipwWIlNA20o
LqEaXRZfc5J7YGzkAC7sum/l9xXnmHd49Gr0K6LRIu3jixEBlyTOWmVPHjiHYTZy
W46OF/PHOqPW20lB1gE7cUxejbvOCeiCrDJk7kBmTl6w013Bhh+clMAKJAKcZ27f
dTgW5NstWCaP+MwnkcSLLaX3Dqpf8Tu4bEx4NNC/MAqGKJN2JiLObw8LCn7VoTvn
QrcCj/GSrdQrfzaaMaokB3o47SZeqtKXr8x1NyNbBPguOZNVB44XWl2EzlC8bVdN
jZGlbFg7MxiSa9GFO6O8YBPmoSRknmrI7Ut4o5pX05TPh06WzWWsJWT7u1X/eESb
GDpHX3FhjAfqvIqRkFdfxPvMTkSLpFcKIKC2GdZzAgNB+S7xhf55jjo0GGqLB0u4
Tlm4icxK9+BDCmYZkhl1PEi3VKdCGco6g8g1DMsQ9Q3dQntB95SMbzwkvggPgDhi
MEd3eVcVjQkuHfu5abqV674r2dW0vp5tZJf2UB8TWPLuew557N1Aa9KoZsvlC8wX
7eoLL+mCxxBLTLpiwr1MtYwP8/ocbqRL7M5MZMc4Y92b0oIQc4SzbbYWJRU/8vMv
ABzJKX2tVIO7ooUVcTVy7RAvDCmhGdfpckRi0SwziRvp21NseG7MTP/y9WCvggJ6
CpObhlIlF7ugpUG5mqdWw3+ubSNIxRL4N0aS1HKONsYTPllWrWsUS2EaHUMtpzN+
EcJFc9HBYc2lS0/hm6Y6s9xiKP+Hd3ZU6XXo2pqNQzflxdTlW05wKwRIXn9GRBnh
Zgfs47FGvPaTzx12TievVB4xhCOx2VJD7UHPS6ipKuEdom5oZLZWnrrCi2dUegXM
mQQl2b+Py0s85A81s7nTGpMMer3NRK8v/YlO9K2cO6FiTFeJqyXAtbK5UdrXVq01
jITfZ/YxUCKGBvncd4Ess8v4yKpzft81kiK7xfayYVSh3340MfawNe0ihVTZptcw
JV7eXJGgIbNipxa7+4cyswj+BVSqH0b/KisvPvA4NBNQV/tMPzQ6B3bRtEhXNWtD
4YR5bGvSDfKsq4kcKWe80kqAsILKW8E4dXO31RddRh9/TO4qW+8e/EJt7Rr0K4pP
WkllEgPkt61BOsnSlcuk/DRlxrBCm2eCZxYtyJ6Ghz8HNCTxW0PZYefXQAJrScZu
AeUJP2KE5yE39y3MwCOgbbckBbfDmKuRhGv4EKQmvmwy/dqE0qXplHMDU+WZrlMi
/pBLQpvxsU4XS2y2WAUAzp5+vexjfIRa04gMKkNINuEmED7ylf6aWTe4oiaq644k
MMJaR5Yed6MVwl7N92ybeaE7P3HcSS34iBJkr14pcNx/BV5xrAS9j+ujGAhtvMrE
fRe2pwvbol5xjcpB6ShKP/HIThuvoFBySAplcjV70gPA9Pw6+hJtekLFYSVbtckr
BLj43Ko7fmJ8N2NYgmxakQhPYLRvBSXS9MFWQqmgEHu75DDuK7neMQUvpjzNoraS
gMK845AHPrq+ylLoRsv2VH1BZTR49BrRHkykc0ciwcFiccQegSyPrpM42tlPpF11
MQ6v7vI/yBs1rBjuGcR0ey5Xfu5RhbkNRSBeFrM56inuADmDFSVaoEyb0TR1nSrG
Al8cKlu78liaPNY5A+mIpiJxpkxBfnGohxlW4u5QAqlfirCznj73Ic3dTJPRjxsS
Rp5CvnU5CkFJwQILpSqqYk856cYq8fs0yGDfaqFhOQXUtn3E5jXXr+ctntBjNKcv
7YmVpUWsufik4G8UDvcuB8k1DWKACz5WJMzlh1fYNjeS863ilEVQcWcJNkbvymS6
I0JsGSkmfbs0ZarTYXHtp53V6NS9p/MoBlCRu35VdRt8DGldU3NVLNYWE5NeoKvd
OU1KAe8uEyzi/epuvFlZXMJL6eYio5Q+YLBHFxdYjk9mXvHvFwsmL92ZpUkqSTfW
AzfxyYZA5BV3u02BqOx8cjkYOVqLqX96UHfGfZiRz7pAHbZ4Ab21FkdThfskPZXU
ffFqAiq/4UobUwfcidvxKETjntWypHg9H2PIqE4fpiCijcK2ca5sL7DBrMoRYPoW
6rfJyE+gxZBgHX8AATH++R5sAL3aJxTAuc1gTyskxA7vrcQ5RzKVHva69H3QHeWV
yw+lrId9nZOrEB9Jl2sDm0uXuuL5Nb+ThmC37TMWGjNLR+5lINZjHZjA3HpvVvui
073kQn9sQcgXU15rDCaW61ful4niK3kolnjPhMKYoWvH0qKYjg1WNG2ziFigapnr
K49jLhL3diCh0m5r4b+j5EHT5VvB22n35DIHpYeGJHZ/pb4dzrYqPhV7YKBzkNyM
ZADDdVjkOpbwMVhZXJWkRHvoyLHiBLEJ/ZxhIuNU715iO9NAz02EZFevTUhVpb+W
hI9iIolnRrU2XV0+vj2c4arAx86RellNV+/jjXDYqY6ZoZX3/PVYJo4RDqVeW6L5
WuP776KWNmRnX9UMsRzIzDyCSd/PP9u+bG6TquyDqFqqnuxSYQxyTH0cnZzfTULz
He6hyQNdsSyU41xFNUkJHrv1tVJnX6m8vQItv2EyCeOolnWRACsOOQuGYZHPnXn5
c9T9wrzCKh6wChfwZyr7bn7iRzcQLKqXqh9u9dwr+HTDZLOtZagXBkyDt5lBLP+7
Kdipd1Bz/15LEoh56P72bZaiKH1icGdlJhQ1VNS9P+Z6FZr+NpGwPhsqqLoh1F3s
Wn7g7DIvFYNq/WYZ1B5g7mRT/LO4xa8xDSji4qNBOhuSo6HEhQFgV62ZyNfl3ZMD
phf6dT0+fxD5yxqcfe6fPtSwWUqN9fdoQ9F4KMmQKAgB1SQbhdbEVCVzUPUUHL30
aV6v7RuXbfSaqnSjTp/MXibATQ6rztPbqbMUkPBOFoTUrPvT8NE1eE0qA1s21T//
3YO8ByYfxzpndAJOjQAkQqaaZsycQog/Y5QFcTyuN+XkyH5hUQUPChDFkxgCRpJK
tNnym6MEcOaNjY1jFz3AgZldWGhhTZsn4w2rvOZeWhAsOeHyn0/UzsYFJn5cK96d
eYIMhqOfukh/yvIxo+Svvt7BFKzJwUmXriYQGjjXOERjrCzUmczSc0PrzbTHseZn
ypefxyABQF07yb3KHoc7beubKruAjaj0ugNC0LoCEZOyURkGQGuAPBs45lgdtgwF
z8mUe/E7rLYwq7krLv8wgA3xIxEiNTlOpjwfMoNPeOlTN2MFsvQywGgJ+s3w3XkP
OtHFnPj5w8iLmZwlnw/dyjujPynPKfcMKVD/GvECoyQyHhNIZLh0P/MN3mPHNCWU
k4W0ob916b/Zp6u1OebBp1jErBGCfCP9GuyoUDb1qzUO5/7IAQ8w0xxK+MvJ4nxh
PmjWXjHba9KzP4aKhZuHYGgGdBpXJZ5nrv5EmXRCKVtXHypTcQkZMd0rhePgjJZ7
cf+xfyTLLqS5QJ0eldcnq470Zm17Cp8bCjjY0zycBSAZLPJrY0dSF8PjrGLWqi32
ilfqKJlLBBduFVut/VkmWuR2LzuxYxTneiPqd/3z1gwIrhmVQIU2VqOCgJoxIY6J
MsneEZwGsxdfzjHpMIT/kVdp0cWLy6qD4CmPgWjIzRFw/dLDRPWd9KIrZ2Ci2j8J
G+KHBZHCL4kYkZU7rR/I6FGIKwu00vVRa5UFbtj80dSGKCZmHq55Pye1PNS26i1W
9JuIXNcDYuZtMlgnySEuzQtmwKuUEZsNGqAIu1lv4Ez4I+WkP6dq3RhmYkVOSND5
t5S1bHGXhrpnMvWvDtHSAlwLxsnnJuX3dUS+trdvOUBHSA1AyIm5KRa2yjvkpCK7
4PW2SxV6dQqpwEWyYl8st8cqBh14gT0hnPjT8tvd7kOTvBWaralqqTRJoJa2s61F
V5XbuH1eBDZChclYzeft3I1YAtsJzTLHkc1nX0gI8irs2HSOWaZrLquNe07TgIh2
ZzLJlCfu8FObDgucg3jzNcvWUs7VX10DiZnxf0sRQALLZBN4m5dEGpLf2hlkMM9E
KlQLzE4cgsk5NJ9h2cm5MAr14OMH7IvWpkfPXBkmdYeg6WreDnIwWrlxA0pNfs9e
ckjr2tq5INkcH6zlqHu5MidIjjBMFEDryOyCqDYulvAlfPXh5rbk7ZDqrleVcltp
eM/UfiUkBE8e4TaacwQ0J+YQpAx9O3CqZG5/WxcEk7/8E7jB2uzmcSKErW6wtdsS
3YB7GmXG1rKOBXT71oBZNHn/b+aC6v2jwrC+69lNxc8bSCIM7ZAKGd3oSYKF155X
cFBJH9zmCwXk6mvSFgYUb3k6UUHKYfoWAi2htSDhZvHTLAd8DRa6rrgtfHkfwYNd
SsastD4H0XCAwxTViPw3Bx+3bPXRoqxTSGztVhpdhqgKpP+tER6sGT6M/Vlrznqd
cpkPZDZLmlrtOwmtzrPYB7E6K/HYVXtRarLf3loQBoegstW+rAW98ikKizFr+EPi
Fpq7Sf4q3LxGKi3Lw1MsibxD49tVqo/9vU1A7PqWulgWXG8gPXKfKTd0J/0bv+u2
vU70aEjgMPWu7PjG+4MG6DgC/Z4Ik2xXP7sLCSNCaaWZtMyi+D9suARJkN8kkAvw
tCFubKfrTpckBfXLTO1+cVsJcPHCYWH2IsXH51Nnazw3WqGRb4/2o+fNCg3jfDe5
oOE5kgUya0tOp8aVw9OzPcVq77OslILtU1UK6ZVwXw59FA90TdMzsoHl5P0R3l4h
A9sG4wCKgWft2I8mQNj9f5h3E8lgcEoOrUvMvHy5zqI+rDHRcJcGoFP1ConittTz
CP67lzZsZ6aPmJB/uTZ8V4bWW6PfJQz4pq2meZ28xWNHlLrAmjd12E0Gflquxqmv
GhRVc2Muek7wdcfzV2cfpoBBcbFsnoIEAIFGe1p8AhyM5wADaRFczVeFfwZ/plfX
B6V8g/ofCDzj0NXdqikN3CqMTnNYsR0aOBmcbGWDHeCAnb7pg8nYZdxG1fk04rfn
hqiXgHo5kDg0QCKeAwikY1haQ+kdhgjcAAkrX7lAoXQ28bWiAZ79wgB5L0kD9IkW
LGfNkhtb1rvf9ivUSFe0wBsy2VhZDBaSiGRFW0d1h6SfbXADGfnB+ecxq2qwvRyt
v5uAd5dmp2Zz94fF93JH79KeE6Wuk0qiC96noeQYKV3Zvw/oPF6rOfa0oGaerlFy
Yqimkn6T/XN03mLv7iQgR4UufeoC6VICr847iqFcXaFwKMEfHh/Nhniq+GgOWpfG
QAg9FhYXEtQn0VdrjAXDNQTVFVZOikLKU0VVS9xiwfE+dp5FI+9WNRNJebAlz43U
Wo5lf5fPlL9z6NAlYkVqgaFCA04GL6eTwmvcMpsu7GBfCeErv4IuS+/joRKdObf5
p46omBcmfVb6zKkjziiY0JyCzRVmCwYgiXSDRJvuAOLKdJN5lZXNeRPlCI4X0nzj
GIF88z7X8pF4S48jycLcYtRgE0lOz+zom9gkFBI5jWvWgXcgsRSA07ruiQC8ioJQ
JV2AuZ1KQ9bYSfm2px9PCtg7iL5pml+pezB2FLl1MN2MAJA+MSQ3UbrLW7WO0bwz
1EqEvAYxbNp7VUxKAkwqoLrzx7kw5I/zNt23rL/ZL28ocIxPQMVnBiC6gxgFgjDt
5SJan5FuHDoxYP6p6ih9paf0DFS4ik4caGnjOvh/SzyNGYOlrk+WQkE7/Xzfoeup
5JVdpFuAP80tzsBfCn3WlMmJTaHfps+3qfodkkvbZsSddg1XImZ7wDMgg85xbKe6
nFVFgZWmZQ/1FhVxiweTue3pUAE5411iTeoGkDYWhoCwbIVDMzuwYLWg+tV7OiMM
8BbYCkeUKrZrcP5NwahQZCPlilwloCjWHbF3DC55Fe9R8D9XdaJFkQZvLXmqZUBb
tYZf1SH9v76wktQJ4muJ4HkNPBeqH1svJjKmeTy6dZENLNULdp8kh5yfhGqLSTPn
7pKJPujF9CUmyyHC2dFcV/zLT16Ohxx9OVfYUSn5C8ofJWnKZwopoLP8CFLctrLM
B3mXjs7Hbo+2fWoe5oluOQhg/zoHWm4fdoGHg7Nww+ZfwvRbo5uJaxxrD0G+U6TC
kl83i2vVXfy3lXzjtu8fzp7Kyosw3LnWdBS3CgTj/ba04THSuWDF41tZJ/Bb7a4/
VwepDg35kHak8AwUmY9NjaUsRZedbwPjKavJCIG6j39G7VMyM7ItbizSCyv+2oi1
EQFnPqiiq8XVxJ+pyD7gJgICR0AviGommb6tIaNeaoBf/nZuqwz1fEX50GrV+K/J
j/E0w8ogVjHTyjXRbe3H2hKkA67BIUKRoOqIuryCds1V4SYVQbl4SHQEr2/jma4H
uUmASourP0aJy+ZWod2JXF6G6orLsauc9w9KY06yZkkA7nPUaxkn0WBMzGULjOfr
xKvyFXhJ8rAeY88coOzt4SbUIgcdx01socJtrphgB+sZVGWUTQN22RevHpLkiJHn
T6F6oXAXrohIR4V6mNdKwEZpnVP10KMXl+K+S9EXg4uSSigDc8oS9WkDxjzdTf0Y
id7ED+or1koZhcQF3MRGHWxNb6HPWi5c77/Xfrt7trgIFndZcs8IHGFSZ5Er8FO3
UCOpw3IfeSYATOr+Y71dJQEa/2tf/1CEEiGYJODI5JJNtsyOss/ssOrFrm3+bU/g
RBaogLiSk/A3MCi2Gk4aHYjvfQ06/5LFO7HS68iP2aFAgpOLNcA1gJOph0X0hz54
+LzXlcFRS+jdDtfkewEErIFnD2+v5d+DB8Xt8tU3ETrz2JRWuyTHwSBeFPOwRIzl
MPYVnTokiCX6jE1CPfUDfmjmFAfG5YjdD54V/4UpP/615z4kvKf8aujLiPH/kn/4
iUY0uy3izQGAKHlkhc7J5IKhOp9H38xCgxHei1ddtMh/+OHXTRfRkCpcEmITcApo
SZrXSYE8nzXKGRRzyhSAKa9+AuWPJy2Jn2Mq1PgMlP2RZftryM6xCYyqIGrn+lal
63ghxjS1t9kXxEHgGWjHL+MFN1vad2KE19I7EHkSz+29fYj6OXRSXWb3P1EboG1R
+j0xC5K5MF5rcCFkz40bISC37gvKSkyTNvTgSO6u7cJbr0RQGHtnn8CjV7iUCMJU
d41Gqd/a+UmEwjf7QglHx2vic+IE1L/4ogXZ+sVGt4D0jOqqCwl7iwKXbNbhESk6
CmcmfjX4/6jLKsCv6VKwo7uVAIoOCsf7XZlhQYmqLWr7Go10GynMC3qEKekd85HV
TmZt5MDvOy9tnI/X3A1xkX7DNZSpRLXSnZU3ZS4cVDJg86PcdH66T8G4XEvBjqQg
wKKmsOu5OIkRfcWlpkrIoJpTyMk97LHlaIh2dvU1m89wiK/HR3mAgzYEcH4pjisi
QxwpcgLC8kjlEBM8RuthE5RK4i8gzr/aIitGPKyGBLykC0ox5r9mJEZbn+O2hu5F
pPFeyLLa4GgUG0C8dMJ5lRwf5+T95moJCblxrP3sjnTCyeQApfJfG7aj54hhzl3P
MVUQWNg9N4cq/l0IZmoBVWSgd/E874+SC+8l6SYvBomlWftfAp09WYek68I6wwvI
SzAHnavkQDKqFqNl2bTl+9nDNGF55GTbpokP8hock78fF8c5tduKKsK0r4JgdLLr
TDEtjzrd5EehMmhBihZRuF7pBgXev8NrSsUT+8rtMn3Hc3PQPkpKOYinwCljxmiV
msCkeHo5MpuBptobwlNQnOxgWQcvu3jeGs5PvBsbfC6fVMq5P6acf50IQbTF2b+i
6cYypJBkk+Cr6aC/3vgsmaW0gtexVUfc6bXrTA0J3RCJXpn/GHBhnY8zm3U6xBo8
CBE/6muK3z8HC+y2ViFgo745MxEs90zK3DHYLCUYG1vKp30cyG/MiaMxcFUFHPBk
oKFH8kTEVtsida8YiXtfNicMQnnA+TnokJQ4i90f6kX930RoeXd8O2wabpQiCLv3
5MEU/U/UFCVpo3u5QClwxDbNfNPNXX0b/8UiLyv9/yDD+rZqWY9zqR6w3M2n7dqb
wf+nH6hTAjfWtKey0QM1yzW31JsQysHjouPDKdJDMSMrh/zdHbKmYssKZDAeFPBt
hZ4t7+tp1BxDt/m5lUq9AGTfE5ZmO3dolV9XdLtD8reO+XAoKaXHAYC/2jiEJojk
kaS/xEHBKLuAJXraRYHERzd8zPmY2C6EATQXPTJ5vL6Uc7d0dhTUV/YHMOv8TEOf
a0d47vIdd6NZqdXj9mX1Ws7tkK55cElz7pJk5fYR6aVatkNZXtueYHxps7MzFX83
1DO/F4+BigQOJ49yV7hcKRQfeiAtlxK9H/cwX/XtYoMhsYpkI7fKEmdUlOQ5+qVr
J54/Yaeo8BkUC0nXqPNQAafP1fRwykQkI9LitfTysjIhpwJOHYpHmK3LviwgIdLa
uOd5/Agx3C3FeglxEosI1NHsSpX4cexzcMP3ls9RQOQFOoKaPNirfaiKpXtHniEq
TRHy/PJNtSjCf3YPdQ16HiQdWYXRMuRp5peQXwDq+WIplj+qAGcCoRB8zP7LMgm5
mD0nP762Lu+2xlJDStZ66wTIZkSNYI1aXKgfI2+SLybjnljNbatCNAqVUEoSxNDO
9juV1yT08+WdGDJ5TL/PjL0ruixmTiwB9Mw7++87YMaboz1f8MEQv01L3skql2iT
Dghi8aeeIoeoAjI5QRUk/2y9UOoXJOvv3KQOVJQNSnjeQB0DlllC/4ujVIldd9lm
rdcHjTOHCnfbgG4UhNVRSnVtbDiF5lF0Au7h1HVlDobOzwHXjgp0ieh8ULBi8opk
QUWGw+Y6Ir82+UUqdYL3opLeuNhZP9ZG1Vn+/xvACrqID6EEeIQoUvSVQmn5LGda
BeQBTLKBOFZMwH8Bkea/qebBJ3+3AzI31xRpla0VGp03sjF0DtYtLBxxkfIo3ywz
ubR08oDlqr45NKgfbWgsjgzrb/yEpi0eJbpkA8/uS6t4T1GHKvx5oqvjAGMlrKgh
30lLDGaBqTiwHAKpYs7ozHE9ScNjRKHC8EoNiI8i7YoHgGTY5kGxgfQeUnSU4frj
3g2Po8IfkwpMxQ3LcXsC46pGm1tHisVSYGoyttG7Y7I5ICsfouOUoO2/fYBf01Nq
hsQD6ZYx0SavhozDsd5wMZr94aSqxk86x1bXdzPy5ZruzYXnIjFfM6CPqIRc6h4O
h+2/QwTEfS3EUZPTK2Q5Aum+HbSXaqxh36yKG3Er2nO5yYl1goFDRL5+G2WvvLsY
Qmfr+bumbvBdVvEilhqRnEbEx7w3/wesW8kYnKiXUYIkL9KWvGePm6TT1r+CbC0h
+JHnbyUmx1iufOE7BNo12X9RjZbMQuvxUTk3GRDGaOrHkoLmzuzwJKz5+AS3QELo
cycDHCGmBQ0RV3QcD0jcMehfHl8Q/X0fvwpNeROvZXq5aJa517YF3eJLMQd98eZh
0XVW+EsMo5GIjz3+ko1rVi19jG8XnGfoLue4zjJRxN3NFLWIiQmHCDaNXxHnnDzm
JLJHX0y8Mnm9MBrK0FbH7/jq6j1AhS4r31LSOdGUgwC9ZtgeEzwaHXB1js/URKyT
PvUq65R0YFoCksXyKsmo5YbwNcQS5fK9nj2uaJHZn9aaM2xHWN9jW74qux4IVZJW
DfIzpx0FPZjQQWd5H3P4IZkjzSROm3Kc43/anp/M5A1HoysGXHf2yUMIWO2LpYmA
NeiE8qmMrr1jLh9bjcqOyRsAGdPH/euDbANoTykn1vb4k9fXyFY7qysjhPiNOE0N
rgAfakBmrSMMy42tDfMXd4Q9Bz8y6B8Au68KVEl+bY7d10QEeRi7xgqOpOSyRvVj
XHC/XHkWwlSkPlwnuqoXqzwBy+qzYDVkXx/TuximPXoilDMrjNZr1C0BbsfQldFJ
pukMlKvocG5cxrvwA5OeXZl+vtYisSq8x0D3484bfI42rpDZVz2WJYavzoB/aLmS
Ake8eWvzbw4f8vyAXHAneY5c5pHl7yWToxfp+Ko1wE4ghbHgRVpGtcwsivxiC0rI
m6+b4YmdxNYIIYbuImNTVF3cM5xWnVdAoG5AWpnuUl/Euj7fVp62UMtllojXkMeT
BuY5hIYl2WyKlI65hawynGEGR9GE2w0Ai2TdBBU19dXt5ltmbcCusjPOxRIC8KOU
3//YIlzwyWyU0ZI0fFEbjvNxxD4FyXNVpib8uL6ElJ89/Q6dATXCWBpOoHFv2C3n
GjpXV6UK44yf4Ktf4OawhgBaqXE1jtPqbm1SQSp4k+NI+Fdrb+u2//DWYRoTa40g
Dt2nrnXdzQxL2TwUdP5twtoKK1DOyWjEDcm/2GQaqn4M5nD51qwno+QtMnLN2d60
lkEL0Dzq7qwvL/WmmRSfA2ecsSM/4lNN3ZxqmcNliwXR+cdDNaHRtqy1WzdR19Tq
/OfMWUapmwTn4kQEIp8Bv7F7004H8ClgifsfulGNuZ1kxk3kVumzNge3XH0MeAAB
bsT+svN0P0Oq4Zrj9ZpqciY2ghJXeBxiyZkeyvJYNDzkn3SuupXSLPFd6kBfXGb8
eyN+B2BCv6jo+DRYnGEcV+S7/JcPd7RQZXnX+LnRvIUg/FhLC1wlnWN1ytX+xSQz
EeokuuYmzEO7/Z9cN0lnFKMv7Q2W1fWRe5WU6bRDswT+Ty1dtN7u7Ph7ZPEO/IVY
B5TRj2FVcfQwdDf2YWOgcoxszQvGFJ9vhu6KwkE0ffPLnSHWwlO6BE4Gyol+paVF
WtljBm4N2YJDtNWboGUBtXU9C9Anm2HRiooWYSm8hiIITBObrWln409b/ekeSLpB
W4zXIlbCZWtdMiR+MJ8YSbYfN7QOCe1XaNhrPBntVtWEtGMwmvA9xgH3580C5g8h
6MLNbS/5zOJqXoGEVnoYclAjFcajQlNcb/ZhrmafJHtnTBXKZlE7ZGDJDPg/yoRc
UUmXHN4mFsJhpWDc6lS/IF4Fk0iMxDXQPs1VZoin/DKak7Q95dm5y7AMGfwp3/F7
gviOmjYTshZcR3whVRZFPdszJvsaHuepRlsZO8BuHFFk1yD2lpQOMEmqBIq+XoGo
RuWdnbLJsEIV4+MIovdpv+KYEpyZ4RtO45QRDtvjfo7ODK/dPzHZi8H5o4DDbXVL
e6Yd24RX0N2NxfiA+QxRYdYIQgSkNeXgLxNnc711N+RT7svn/xxoOV6xWNyioY9c
PUl/dkclMJdTGGJieQg/D3vvHNt/LDS8TvUJsCKHaAFrHgbXeY3Ql0Ek0A+Md7v9
efUgsI+XgUN/5+Z1f52+sci5hDNN5IX/7rVVZTbTDoM//nDwTfxfAq9Ea6uztzf2
gzgaMqPA1wQ4D+koNK6AWsHULTJaICrTMcPgwECyFT8pMNhN5DkRE5KETxiTqo0I
q7tJthIqzg49hKVePUWuvm3AnFNt9sUULPwAdgBFxjsBgpkmJbr/X3dAzRwEFYHe
zxiGBXl0zBzLeTHZ5zLc8gF5zEtHmbPt6ge2DdIxGr7YrN0zFYvEFqHmx4Oja36Y
e4xzM329iPXLHp8enWeW3Y1F8QOvEn+xJrWA0tyIWcFkLrar85U+syRRFkyFZLjw
BP7JkQvCY5darMdGStLHTd8U5/7ToQVX1KIorVjhoDuyrybJ0owVsLT9M6UX/skR
UuvPRZsr3TbNtcAKcla/1fGrgcJo8/ArxBWeaHMubhUAYccGe7nf2NGf7RWML6ZN
v+wVC5/Hz7TF/3fjyvEwxtfJImfbh/ULIyrYilaf/QmbEn+Ae3OSl82F1nNaAMxu
FWK+Z//HXLJOWgI6EKBNKWF+XGnWScdaHaR3Ytvt0dXjize37+JYZ9HZfvZpD0zc
Z9NEoSoN7hXgsf0RTnzAsYAnGVP53BuTw8wUTf+Q1Q9XgByhIW5hCDirP/tAtU6L
GGgyQnHMAacd4muBQsjGJ15kVRx6ZQ9Y/Tno0fkTOipa4tYqJ2JuKsLIrQTvC3W1
JAD7e4toy6MrhIOFAfsaWrNEjM6jFtjfPqAo+NuUWGAZZWYUI7ARzXA5NjuLCZzJ
eS1wvojU3Onf4gz25DO9KBLpQ/GO0s4Q6crxjNXYWJbh6TJu52m9ooPFckmjn1Jb
DS8bIggILOWPTkYVpDWMxIYSaQ81Xg0PsOZOqrVWkMSQfaGNHZjIOXyvXmyOHMui
/esCAoVJXXGAzxmCsqf6wwYFklSDSfFIbP0hVVSr0DYNzn8ulr1NtPxJkwxJWjP2
vcg29aT8WC++9POYeTQHSjeFjVhfnIqvc2EkT0CH7CbRhpZJV/E9Y0M1ND5tyXzA
kZxtGWFmF0Imalhd1wlNTh6LOo8hXeGnkiULby8jS1z3fYaVkeUadEwBr003A0rg
sLUQ2/e4lDrVM7eu8nDUfWL5tjUZzkbenfX1zDHC8s94PGE6IFwIhtAzkA+OL4D+
s4nATmUUHU8roxesXT/epgWvCtMORAMbx23jYhd2R4aRzSeKKKZsukMHCj7f4EOD
Cznaezyi19APAdaTRxoyNQYq1gU9N007hfcBWAqT1QASxro+ki6CeMZpKEvMt1Ba
az/ViQIHhWaQIR/aB/nNqC8dx6eirfuhRD/2SV2b+Lpd6nk/8bdLeIm59XwDvWln
97ZR9Z/H++7QVXSsyQHe/xW6uK3gsT7nkBrQdo1Te/HrlCIllisnkxrGLvtI3G3+
KwjOp1z9Yg7BaZz3lxrt8IJMNEkSo3h46g1NgHv1wBANK0wQXZ/Bq+f98ojhPv8e
Ah1eB4TzJaD5WWVhLclZgwUJ9EzQi8zTXqV8gXk7xVmcmDbUIiWNgMdGIpGMypea
IpH/EXZqcrOJN0D04dADZ67iK+wRcwqqpokUGzXMYUCIaErdV6Sudql/V1e5aymS
31iGRqbkQTb6/Icgt37tVVEMShyE1g79oh8R2m0mm34UUvq6TGcpVfgMm4pkPH1w
W0uNFatPql/uzmh4NmMysnUP4CvK75H4lAP+X13CJavHv4QjYRaxLB7nEKXOc+2+
gaYHJpiJSCSdEH8ybrsrBUc2AX5VgERbxkRjn3EQOuuOl8wKni0J+TAAKeVdraeI
wlJMZSojUMBEOBlwp+6u7yFI+inEIrk6VOqTxTZ0au15GY4dWGeS7xh7jtvmmoPc
IUAZ0Xb6Eb8kxVe0asT38IuFuMa2FxLGjXS5W2kYE/sqoClxIOMMijZQ3WCp9TVn
Ld2yAjs/ueLDg+iHZQNusWsm7vQXzyWnG+DzejWO6SQ9m2bsN2ZqfNkkUKx9Nsug
Tb1Za82qL6Ss3AWcUY8FvCNtJaOW+MsYWaZ3ja1mwxrsuoFkhNkBj5hcSTHteSAr
6meCxe9dpv6pChXdbEabxiWsGnmGKLmaSZfbLB0o7kGIeBuAHZ5AVQWuENoCf/0/
10/F1QRWUl7c8KxUhF6a6zBQnCBaf8uyGTpG9IOma/sjleC3rvNPBTZwpJaPRv2v
id8z6U3eZHxT4MFwDFWcYMwmeheFheDkg8aIarkhtJxG9sGWP1n/WsfbHwH43buH
C7cl3MyijmrkNRQA8pyduE9L2C1I12kM3h6AMj6CGqRS9RBf3sPbgExALzWpbLCQ
JwvZItyb5mcnZ0ROU1sAyTwuP3kNGpdmIKQd+yfbpi6aPd+ifbRb4jNhPxcOCLP+
OovqR5P6f9E5v4U1qvRWfJqL69Nnsh9q9lBw+SOcKORYFnE3zmBls/vgmo0Iip6F
SdaLUEWg7wSHshUWhRYnaXTOXV4xaDRq24SyuO4Hviwjz1CqrIVI3ef+U1ksrf/q
Z7L6fFmaapGt8s8v1+Rw7a18WFrLCNjU+nHhPViGWoVdvNDwA/IN/rlg4+7EhCVB
DuQGSexUeGPyEM7YavxB/2lId6sdzUOm6X4PQpqyAWTJiaF4Kk4uPAShiRk1GpBT
x60MCO00McpS1/WZbot5e/PGQzGAfGLaT1Hj6cOrsUNXbjReBVw5+9qmyECzmBfl
VZXJ4Fe+pzH1o2HLWlKwV598UCEAvdZMumINxK0ks/EepyucmNJmIrUVikWpC7bj
UVZ9VbmXgfrY7Py5a3o+qVxgjlhQAHCXi4+21qHsLkKJkt683u+3nsL61/9cUseW
9ZYyofUxndDsxCzZdZwx64PVNhY98boVMhZinCrmXwhHw7pjdbyxKizoO6PWhlFs
gPXFwcEjW6NXHxbQIgx+6j0512LQxDUaBTO7XG/BKnUP77v3Ogs7rZ0dAnWS8qD2
fJpN81d0xHMB1SwZUsXSXJirRla0b0sspIBmK/TIdoctIXheSc9hMnsVWRV975ZU
rRerydARwgejsjeloMylOrXikmiEQ3Ee7AZl7ebKjUyftk7hZRRNOtJpgCN4tc86
Eh3DYK4OtuL1e4vFM0O1L/ZX6S6Y6RIuJLBCooBaf8gxeNMZcdPi9NkIwWKH89tM
h3kt0+4wGFAj/QCeDv/jnyT2KWMVSFArhUlv4jQPfOCvLZUwWTmKl4W4lXXNYPpX
pHxoteJf5LJpzvm8yQqV3pR7ZTzLXr2ELUYf9ds+nT9P4kWBGxAwqSX6AI3Wddie
YU0vBNoTr6fglNJf7Rl9E5fFUefABUnnjWNwBXDyK4KwTcsm+naPsEN0qTflbYa8
y8gUM/JX6aDq1s1mtArFxhNTlYXsT64/aJ9LShyMR8sEgfQ9t1XLJPZGDAiqWcmO
mMADzETvIVAJJidp7Wb21Igj9oWhq51crT5fVUQoVbZxvcvsry9H2Hh7XNWcA811
D8QVDbinoHKiJfRpeqZwZ/87XcpG6+blUJO89IZpIb6t9xuLB6SmouLtRlKa7BPU
YXslSRSthKfjh93YN2QPBHqUuyQ95FBE7lIDtw+WF/ANp/BHzSJ5ICaI3WULc4fM
ahv223sJ4s0kJ0LKYXei9MFiY9oItZXYrxjXrDZPSNbSCzoEVHwcVt6uRBLGdqVm
5W5IjTAs/62YJpr9CsFK20IaiCDXbRmqXFFSenMBvNJwsO8L/wEMtHCMoms6oUab
sHApu3xshp5W56RYrZwuGCLMkC3LsPCp9K77yAMiH/upLiQhHwbmKu+Q1kYAQH1b
veIJYF6tIxLDixbNbWjOFcVIxUdkCywh3IErPzzHIEQ/1YCEgZtZpypxgUA5q5y7
JdeQ0YnNroStJE4yfNRtDEsI5pklP+tnW6EuSTWD5bQBiRsxHg6b1Xmgh5bQVwdb
KEGwsEzLfN6EInFvuabP8BWVKbfNuLMZoMNiB+bE6X6uDAxHcwuHTqeBlUPbBtDD
oTyYKiQDDlTmbimyFZo5LyZB5h531gFn4/yUuGpFZ40JzmK5kKFeO8J1ZTNFXYhn
T10DIEzb0WW7YFB7SwcYb5tEh5lyTRFDIHuNgUJXoSMCCOdqt3IifO16ZHU/m5LZ
2QOi/X4AUWc36AAtZ5aWHq4QP/00bRkvPwFUZW9JqsAKt2GtKZ7koclVACdyD09C
vCxTAi2F0rtOjsT0k3jNJbjgQWWSEclL//omFzxR5l7UOfpxwDFtj0VfK7luYBj5
EAHKJgKfhMbzoQhxthw2McYaeEHMOZaMqBNFRZnOFkgfxaG4KGuEEOM1u65uurFg
+j6nDaWHSmZs1do7CPcOyD/Ti3/7Op9sGVpf/WuGzsyAVAffM14LLhdjVyg9KGXM
KScOkbL3dR/O+thEwFIEUzLM+Vbp1gIniQ8zRC1rwFftxKV6vpgraWERjUj/n97F
XiCHcA1OlHahqeEGfiyQFcZ8blvnlnGcm1ddfxi7JtskmzfhfVgEddof1KZl4bCo
whZdXqgpBPMEsEKR3RTy6MEHw8JGlU4371B+wFwPP5J6WtYmmxlg9DxiOLeNjTDv
FlUFPxrhohWgiVJQAICvMWZxMxY4digmAj47/+YHH71+arztmablAicItL4TQ4oq
IkGa8Lvt0xG0ngoBw12CDKGhH8jmIS4jY3tui2lG0MjrKuNnrZmbqtJ7mgtCePRb
0TwLQf0aUmnGWCFOtDv3fEXHEY3rIt76kpKG7LrS2ejHpAUkK1NNbPc1HZ/RZAiy
RVNT+sux1jnr/UhRdgy93TNnuHQ6R8G3f4p+fJ/Cx6MDIYhGtKxRGe18wu2b7+tJ
ev0Be7Lozg7F6uWZwMezEuv7SdzZNHCcAUo5+rVyIjbxC88/tuv7tHPxLPEUYhqi
iBbNDEm+KJQgFgFm1YU5+zKkGCrpQWeDAybvrYutNktks7aVkGUJlXMF5kRgFevy
8ZRARcNn6a7UO23tWYKAQzW3XKIkjQTmThhiCpWPMdfAlrIxDn6whSVRkgKbgsn9
nAIdDunm3N7oKJ2Q9cHyS9TpmTNAwZFBGj/p4FD0gnatYtH7Q7J5ttFoX3AnsGm2
jTPp9DizCXPLYnfCjwkw8L8drjNPMURsNSKj4OSTwEMrCV6ArgrEqfGrrBRMjmrU
YQA2j7V4TDS7+IZ7OchNV3i107Ky74A4jf7bVogzIyQ64kHBlsA5LlQD4081Xbyl
C7F23lEcbOyV50WwmHk5y11fOo5rEqNQUWaIImaoddwAhKobiCB75UpMUdXdozuU
OuStmy6bCF8ffWsWzthc+X9L4G12vklnjXQVHA3Oj0opnxpc+51Pb/d48r1t5HMK
9PsISrGqb/qFoVj3f9CB/AN5ROThfZI20OxXB3Meg9If1QK1AamMSjx2POOWb3t9
QRZwDppKjZMnQtTbKNKv4M+g/60HJMiS3NKIvY462trh7OiPNT1eWn9fzDYkE8b7
M5kfCGKi1xdcdfuntO+SSZ6WIiEZSK+FWF05IsOD9MZt4wF4z6WUuNM9C83V+RmY
mnoWMEdFxwrejLX866bl+9ob02Jm9kjdHDzKl0+85q9J+QhunxfvMF68e/EyqYgl
1LuRsp5rd5I9mO36HlaE615cH86U92sAkR5RJI8iBGK6hhKYo3H1fLXrnjmb1vm+
4eGNkoajYcSsbCZ5E5s8EofSKeWZXcu0JUZfA5Yl3pSk1sSbUG6IA+2x8qiWThWG
qz9wbFvbucvN2fCS5WkzRePt3xpT4rjaNBKxY5uR8RMvQit1T0vlCGoOdmJK+Pl8
gxj6w8uTAvFl6HfZ0YN7SE9LCh/foCIO9fNKFqaoe8FFNrTvYeo4dUSs2VRFJTjp
mTj9rnaef700TivEEWMF28b6utr8oMFgpJsDLaUwBU3n9ayOgHsG3yg8H1JX6TEv
rINFtdwAEYzldjtHIQQuxCHF+fXItDgkEu/x8/NslIv6QhXtpiyuI3bvwXYoFhT4
K44OjviBdFZfY9F3RD6O5qzKS21hn+RGMvCS5jLBCo5We0ZQw+eyDwkG3NynVTmF
dE4iQ9+ovYKeEc6EfHo3pmxCOUWoh4Sn0FQnEMXskmGDf6yeLowZ4z2FiLaC7Nia
xcKiyLhrjtDX8ENLXhY/Jqcwj1xXKP/hL19axa/kdHB9NSupcy1S6+QF6KZswJhd
bYDU5H4NCwX0xmEcnaESbNH9JV+zTU1mIBbePqy/Gns5HLbC97ei2/jLh9Anrdl0
7sasHuZQy0810cbUxcSFMT71fP0hW91YLFr1JI2bpJvDy3ZsFKGjyZeu0i6/BCGK
iv1XRPY3yBoKpXJ4WMgLB9VFc6x7w3l2gvBjtnu+g+5fff+Pdk3o+dghKaWBJYL+
5uJoiHagjf3SfDHfcm8Eaqco9px344iPcPbGJMbFvBoYVkY6bZaE6qnrNrGATdQ8
dWbz5QqWptHBV2+b8YquXuZJ+S3BhV2+LR0Ofnu4fJFKQsLB8LVtQ/m8fSyiKLmt
f54gyvU/JYJ/PNBysdPHw5w9RyPbzCujQtm/UhypADK9itQT4IMcK4ujs/to+pk4
hb//hAleRF2Ixc+Wna75dXhOlo4+dSeRTwqsXzN80qXcwSD9f4ZT4HyQHdPYQx04
iQU8zWtsvV7AN0TnnIg9myVhYvV+yCi3OzODdnoysnd2touLnTbFc6Axhc6Evxch
LHoKdlwrFzbdRdC0JMQ4MVkgqqWUqlqKF4/2Iw58ms6wPm7MuvSBROO37TwecO5C
ZeLn3mCfCJouyKhmQJ0c+Iul8jWc9ROWSp6ZFj1MJa7RUVMyEEe/qeNmRp+92EkA
A1Ap1O2WKwAvW+EfH7rHxWL0nZFfPgZnSuetR4KJdHvX1U3vt53X+JzrjadwBKqH
5jv57Exhewkq53HhKUlFCr9Ad/ulPFpJKxb+btN51XIKYXjPSW0aLjuDa1nGStne
efgi1n8XGF//kMGU0wZfEAv5cbxvvKa7ozXwq1uSt697SpHUb/+93evjsno+HOI5
CiTRdOMPly7KsxLDB1mftfDOl8jbulG5Em6grxNMhx5y2LrHeI3KZMwn8cYeVZsm
qJCEdevECjS9tRX45PmMxiASCFXNMJyJunMV+H9L3Q83oC0w4MMQGijRMoUNdF+n
oDhM7pyrxN9gKair6jOOKTFMcnRv55axo/yn/QNMhvGpTdEwcOd2CZNrjdFsH3Hz
+NlKmj2N7edUL9jZdliz5N6qAjRUdHXM7wuglkQlQ1p1OcdR2SVBAmp1f3esbz9g
m9CT1FiNwldOGL58QE3nkW2tn/lmUi68OtK4JCTfUZtFQj99aG8tr9Tr9gqHCoyl
mUxQthwvpHigg3z4izstLim6mWPGeJr7F+aHBvlR7C8ZliFk4qg24smrA1GNAGdy
3i2GNPSZP9AgOyu7TVbAxnX1zZ7fu4W07oMVSxXM7TexbWlzaccPSbChNparCH39
iVCGgleyoitS0w3RBln9HE8+oW3V2JVlB760cckCGPitgUp4xwLNRuysWg8ehaNK
HfWzzPH9nitqhkZI8xk9cTxGtA2RFNA88zm7KBlBru4Jv4LU54MAxT3CCop4oKhm
eAO5xnbotp/0mqj8q4d2RpVSDS11i2tf/pZSmTao677eLPfsptDCzS6w801dGfmf
ddLTnkzEHzsxFE/uNQHw9yKqdrOhtjC9/2/RQJA7cEHp6HoCo7SHvgcfj3GQl/t7
PavL9T6C7kX25401/DTYEDMUHXYUcix/rNZsEcSqiZWnZVRSXrpHtSCBvAsRLumj
DhlryW+cP5mXy4eVGeGmyEoJLsuerISH80I8GddWIvimwfb0aRtq0JkFKeoT2KU/
I2KcwleoSFPZk6vr4uw8ulJTke8Oy3PP8othUC6y4VJgLoltoCd5FgsxAX4aKDjU
cbW6MDpOkT32pcyTwbswZM9uaj/B/+/A8C4dOjQ3/xOwVOE1jWUDPbum1TH9+cDI
TL63OrJwvfpBUdUapUq9hVTHiIT/d+izGrhUo3g+0BM7KAj3OQMYvweAWoYPzVYp
bZxQDIH1fKf81yzrj199PmtSceRUpbSJco5tbjKveWLbTMhjLI559YQCPH/qdgvJ
HYjjZPBsOF/yFNTmI+bjsZSlhcTjUuZ9/geRVSbmwgtk8Ys5jQj68NOmL8LWtjwB
fzDMF+jaxP+VYtt6RScfQZIMHcDDwr63GQqU7C7GK/seHBjdHVuoG4pfKdwWEDV4
UXWNN3xilDL7cq9/aZXPOE7m+o+KzVWIQpNs2JgjpUoUJSaliASBuwRFRKdh5J0O
KKZhkzmX4+X9XLe7VpJJI7Dq8KDxA6XtT4GluQ8zGBZBcS8R0MDBtmypPOwC/JnT
AqJbiRrYCelxZQa1QV1EIiq4qsaNh8MKMTJ4BKC1BTkEwkg9OfM82vv22AOHmEhi
n5aBBeuDoaJ7eig/8+fzq6K6VzLxo/1JUWySYEauzZFHbuuZSK540lJzwZ6Bg6YB
NroaWSH2De4hSMecoKDEGOeMVcyodNPa+wMlUoAgQ0wIwXjdsa9tef0XP8KCy+2A
+4uC315kVeqTIwIl/nd2NXv3OSqgM8f5Y4vH8kNXNrSIN1E7k0EWVkgR3KjD/Lcp
RT/sgH0sDK7Br4BBorQfswkg/QgW/5s5kB0n9lLwyk6VZwnOe0HZGByUFNLoENHh
BG2rikBk8JwiKEd4rIMorm4jw4uf3Sp7ZvyarsdOfRb6Bf/l8cgC55dDO4BvUES1
/6L8s+j6ZZRvnM0x+65NRudx7t3dPPcQ68VN+CyqlEnnW60vUhpDCEekW11CbeI0
k3JEqhmAXUufdcgL5IT4+b0S0xvNLUERT5pieGr1HpHpT7ks6PXdrwls4YHwzGne
8kgMXmmyHhbT6kjRwv9guZ+GSJOAPzoFUr5Xetnne0SFfmUjggoUstMP922c3eTc
s5cRb8npeV6I7yKOnTe3iHnxDFPSnTz+eRjUOiQYjMdlcqi5Q/yDQKKFKSv/eTt5
Gflgvj9vsKDOpaTY4WhQUityEVVWDGY1etYTlN5yuTuLsxt3DWuHpvIUvHjdUgCz
b+OOlVNEtY8RNWxdNtdRQEp6komPdvrtL+v3Eb/kYhl5ellm5PRDjtL6OU5Q79Gs
aizDKSpBvmKpO04r/yhTJLBHwtJMqp0xeK8dykz7LuXfs/bfm4dn6PA43/6A590p
usQ40IW1SC4CvxN0Y9nmTzxHGFWEj8OTHE9sSqEhXKg+tRKHXDgcaSS12t6wpX73
Gi4IZUFoIpnjnvwgLD8vuRF7ggLJXNwPYNkcsdhaLi+IQpB9m9f/6S6UNfVG4fWU
aapRm7uEVbaQGYAxgAuLN6br4OPfdpUaBC7j08f7b2h+zSsmnZ30x2IUCo2haXfo
3QPlZKIeXmxflcILVWrTb1DdpGxBROZAxgJ1/jf7NlWPQb634yb+Yk9qmneotN+Z
pZ5bSfni3piMcbY5CreW4o10bmcKbNlyqgkbD7TXmuxCrYuPgDifAJdmVZS7Rp2F
SZgWI0Ml+MHnt0cTYEoX5ZJjXbRxNp2lDx/FzCAm9NzP9n1ioy/7z26IDrbB6QO6
FFqbMh1I/TVtPPu46SpLuQA8FTDkWOOJ+rYyN8lbEYUrpGoOQWOkYJKOqyO1IIvt
ompxPXmDsuxZvB1przdpGpgiUc0GfTKyIm+9o0+LXkOH7/E3tlpX/9BrmS4TaNTN
/pM1i/xfZ1+QYeF/OQoQwmtYiyDWJX5PHutpzaO13AYtxOJ629PndKZeX9pjUt0a
5I5vqKG1Y9RwDyl4Ed5ScPP47aGv/fINvQF5NKaHwO/sOuAo2iKHKia56eZkivRo
vq320YfkR0GZlxGA50yOeNOcUmM2RwkWoopv0QzirFh5xU9EMvDTZ8iJ2jyN+qrf
TpFu8jmdCNvjkmUXQ7RA7nz6EvmFJkHQWRBrn0BXwHNMsTCtGl0XBObUEE+JJ+Dp
JN0ulPuTFXLJGPVDFLkaBB+whlVwonHS60tz6YSL6Vv9wum2LRwPIksHOB5PWMum
2E5VY78xn812E5IE8swqyAVqcIAfmVkmQLajy46K4M56n8X4znpXcO/Q5LKvsNHx
jdxV883BlHK/NcywzHLsHtoqwkJGSA0R/eJJnVTcpB3gVQljolv5IQgPtxgkXi/c
AH9SZrs5AXdU0bQJMc3xHklRAb0fN9lggrpJsx7/w+K9hQ75ZeQ82atxydV+Ii6E
VAvfCOs0R3X+G1g1lvrKOpB9eriiYhDXtST0NGya5i7P7KYURtfPJZ1eJ1HZc8ii
CsHxr8ph7YMyezJmuesDaaAEfUvhIdr8HKzCYJfnYSR48YWwUxDo0osx4uARODYD
mDshc/5Gc2kGFczJWSGo/WyBpkEM20iQ7LBbCpH/ZtVhV0Uy4XSue7GCbVGckkoC
1qo1UBPB0FlmaFepaztVJPjW8LaPpPmIR1KOr6LxWJqdKuZehwf1i+G6RnIttFLn
QolmkduhDdK8gLPiz+2E7w4FppCQjeq+bcRrTQBShUWlzoXxOe28nTzrCCZ8C7pA
VoyJctEx69yR2r7PvImcxJDfFdmmTy01ZlKZBcVmC6OFuq0UivHZvisQqdcdLaOt
lqo7cYPP+jjmA6gRjp0xOvvcE7krUwTIK7lKp+gh91WLgXBZM06e7UZt6VYQ10gH
SDxKxeH8VI6q+qpbzHrzYNZhj80ZSV/CZkLcLZpGfTBHJ9u3pGY3e5Hm0vFw/kP8
IkKv4I2ElQUcgiLI4Zy1Hf+qV0lSvDS6AAdluPZkMqF/MEXeFE962LHIIAMQlw8Y
//wJ3l05bT34MEpZLppskorPUWF4eaEmqKYZxy0RQHq6fedE8dzRdwtNwdN7Golf
c3Dzv7KItQTgvCnYhOC6zPjLYdUxqJ2n29E+W18iBQhZ2fnU1QoxKckAQgee+CaC
t6dUCXULUj8X925knVi4f0POwYb2gM6XfXwpiOKzjoYtxuJW8V9SHdKOPbYr7xxp
iS6QJBw9fdt6u0VUBR7r9btbc95fokLrLKR2Ot3p3AtL1+Ju4YdPk93oQmbYaEN+
ENPJfQSyej/tndGpVFcu+JYKDI4ximrx84o4QQlg4XoCyicfjcSJ9b/ZW6Er4ktp
nGp3DaFX3XkjKQcALo0kDorC7ZcPEpQqHM35qjD/nXcHfFbEa5id71mrHkU1rrZE
kRhGbeeFgw0Fwr/VwYDtbeoQZtrETIDr5aTV5TgLJVB2L8Ly5/GZQNFadmdzMHNH
tMC31OpvBUk5gulYuU0uS6j3DUUdgti1VaOaX7qZQxNM96vyI+87CkbHmFjgvhaf
Q8hPPAQsrHfF9pl05HPfgRpK+hcz+oYsc/raTxnf3zXDW0Q5s07kxdsOLj0rBVoy
HLIH00vppyefbQKS5lz9hsN4EuL4D6klXbONOKZZoSZaYZtydHUfGWpnmWKrB0Iy
Dtx4vzkdJ1hEhOLSMt0tvRO3Ry8FRITozsvhcHoQi5MFbEbmQs66NorlwK+FGQyu
ymGH/RfZ+LSG0JcYTfnFOW8Func61xToz0Xm6CV/CF3kysfHs5UMt3qWnZCWLuVl
MvofFfULJk4aiaXont8mQoVjCMr7S8T1Mga6W1fknvlZ0ClOck0qDyX791ppofEU
d+gH3qfM+g1oBHKH8uS/PbAC7UFVKiXCjWwm7NDwed3VMtSv+3vRcYwpFLFjWW5n
NdgiCOQsCgbK6zmlrEopd10NbRHoh+SuqCdvbC692VIQd1u8AMmImQwixOisQOaL
k2qa8aw099hBFpmVKYPxAwIbfR1tQN0eULchLdZ7UDq1H3QmMs23T4YQap6njyCN
PaqmTJUrrLaa32s/ndBHkYqDMymXXhs1Jh04WyUOginzEPgOs/d+qIMBQDhwuuI1
m8ew73NBQIU/SzQTf9UPri7onM0V5et44p4dohZ1gRdLUMs07t02SW6P9UHtkzGu
xzjnuPKqvdm12JmdwIbn0gCPJE9nHiyqzf83fr7FMAiivyXlQO7Pt/HiiuC+sg3m
s6GmmbYpO6FREkJTMn2EEf5EvhxkBWlUSmlF9WGoNsF52T6r3upaGWrrcm5aOtdE
nMKc1s5+0U2rAH4h3Xw2TKbiJrc1JYk12dX8VcrNTiTvOywNBjfQEofy3QsZDZCs
GsVhRDrmnvEyWhQFFYABgzzD+4z095ZPH9EcVfDhYqcaJ0diQxo/Lujh/JW2p5Fv
nXtwTQ2gaq/Fj+HNtqWbsXKfrPLE+ygb1gW2Y7XeaNXPPqfLhMApcq+Pj77v+t2s
WhNanY4rtuloJABGohSk2WXTu3egVOMT09E3hk8TwBnuGV8ni3uDc0+h0wO+7jNn
kkk4jU6n0JoImPPV0f1eEb2rLHH5FPkjbXyKzuBw6Eeg2axznbL+dfkzfaOqyBBL
5/xtOZzNCHpkXJntXRO0i1aWTHBFpgPLQYwQsIBbxXJr7y1sGQAXHJrffayxlIAO
22X7+ht/5jXWxRz0dZtumn17UM1O3MFqvdIf+u16w+2pwt4k9akxcljKBAEAAWw6
S/zzKYedsCeqriuys64jsq7NiL+LcavwnuH+eCtliIP7pZHid8dI1k11TC8lMxuQ
j9XNI+pkfr66t9OngSHWraePW6uAmFTgxGPVRjnbLrRw7ZiYz8LfQQ3Pm6OkQGbz
b0HA5IUqvHx0QQ6r3we3qYqIZjMP0HOVKdQ6F/1YDWzlNzu341TCcutTqfEjcdFx
nOMm7XWsFePIbVQeqRcaWT2SUgHv4LFRrL9da85KB0blbUf/HkSxCplN2iuSrVlL
3GqVOXioe4vQvnZhKnktSkswh3TuHUripFih2BITjEe65buNNbRRrKJEJQvG6BZl
rbPtx56AKCrlWkvRm/5gmhInAT44KFTvv5rTJrSGo7j8WqxmtQzqUAch5eZlq1p8
/SboHcTTn46f4BDstMrfffHVicOObEwfh5rFebrJPzya3yZvgsTwZwHOY2HxySAY
dh8APlxyDB+NH1zF7XnLY9Apo9FOuKWmtPJGh5zgqE99zMZ/oZr8vY9ekxT/EG3f
a3rRDkoD8CxsMRNn6cxl4TzRzNGQ8WGfb88qIvRKhxHNbidsecdHa1Iq9Tqfor/0
zE3Bzj0yZrSsXn2aP7/NVSwSpeKV0hTRr7d4nMESvzK8lxys8uNHNNhQllDNaXjr
sv13VKNYPaCC5dtMPfmrGfTGPxaeGlmHapcXBU3Gc2Q/R2hpAv/uBGbAcKKCDbJY
9FgFMhwsDx9+lBK4S5r/eOlhuUmUapJhNeXterfO5MtMXNi7MkqfPjz9v77eL0bL
JUet6e2NLjxHtp7ByhndvccvnSc+NTXag+oPwjj77lZTJnA1YVRYP7eGg3hGmNkM
pkyx7baVcnkvVVEB1qg9vM0ChNi6K3PMzhmRcLLgq0WzsT0JSoT1aIRW8MeQNSKo
tlUyZuEexrL/JBZwrIG1IRwjbo6cd0Bq7wMuPBVzep2Gh5wf5prvgvn8fOVoPA3n
jtXaER1In7LKej0whdg5VIVTpPDSHcve/fPCF3jf47MJeYF0u4A7MAdEPRtuxrC5
xrMdbkc/ZIH4y2tk7dAhDDHn2HsA7SEy5d0SY9vPBQuRzf+YNJNEor8Cr/+wbWcc
CFog6GyPeEqzEya5mn8BkECpC4OBW3mLQ63hMmousl3hP7ZcKcg+BVx0R4XY0T5o
PrZkVsMk3vdXzsAcJ/aAdXj3Hhgf7/rszdZ0GCVnhuka4U4+g7vdk+rKWbfsMyH0
gjDIYLkLKQ2ZCFGOC57AlpNycAVZlycRv7q8FihjUEqo8Wzn7xABO4xwaEx0zTiu
B+Jf9eZpnk0j3EgvPJTq6UQvwtu/S4wcZ1DOMkkw5XJdHz7O9CKSAPNwRzlOGvSu
bEZXORwxzBaUp8MX2B9Q/iJmQfWxXIrk6sBFlKWcvu7Qaaj8KQn2aXTYpr8uxYd0
KIZT6k20Fz72Ngd5EjSaW8SxhKEQIw4q5mN42j6XZfBrCM7pMw4yRVXQakKoop8P
qJVGcu0Kv1nkulirNL2ps4ywD9lGhrrFzkC6mFC2ZFdXgPamAs7mhNGyFVhJ9RvM
m9QYBNOgdAKYFr29yEanfHIUWCjCaGjvn+LW9ywSsi8nkr0iINGbGDdHdajuRMd1
bLECogt2o90jGdYYTFN88EbR7wMhAedQHfxC4HP27qWwB5wvTjJL7H6rrRC/9NEl
Z7s4XBISlNhoc1ZSS7qQagEe7+dx2St/UWVn2cFA/tElOWC/KAOFQBRtjZnD07sG
RmDULASj4Y3oHEh4IIcjDFTAPq5J9Cs6gsPhaZgmS6+Zc93qLaX67IB3hwl5V2/h
LtvNvyns3avHSzvgggRN1LSGOGo0F4Mnq+PbIco5RXQd2XTWYmw/TeIYgTbJA42E
mEZc2nehmhBeAdqbzGeuZe8nD0zUU5U/fdYVkYQyaBXxGzuh+Qo2AvwWBBfzKGW+
ywZgoIXP1SzPlrhIuDWNZNBKS2oa40EtohvCasW1G/meNgDywG3pzmkQmEwPiQEk
Ih68qtv7/ZF9hOgmSHd5tCo7aTTn65KEOQ+mYFk7jqSe/+QSLhNjTDT8bZcqBYfW
rd2NLAh24/82d4EOnUKx7XHRAgQfUSnzWz/58w5K2E8MuVe+2azW0r0aP97ftwXu
8s7OrJst32io5lXHwmQr03qk3JhlVThxZHsDHl1q4xEOQSDZoAxj6O5os5/mjmf6
XVgymuNWpez6ITIuo5Ny6FJZpOylhmHXeseZ+FA9/dUzXJeYFWM5jo67oT4HIJKl
kNmcj0Kho7SHLoEVlnF1qXipuFWo8XO4V0QjqsKysBONvJ4FnTzzoAKT+L5cN1x1
UxlE2xdRYteuTgKgNRdE+njp5zY8ll1B4HxesKZOFIUI+Lyq4bn3nGM5d3x5oluy
FiFDWhrbxy4dVof/ZOFtWXRzbkN5GcvDpfKTotg80t6bd6U+RrniKQUEMTJGA4du
Py23aYbQf7sMxYVN4p4Gi3vHLsJq318vy5e4dalnAeydmw6qYE+iWJSv8/UJnEHs
7vdUn9i9CneIk2N3lo2rSFvefgtiV/wExNIYupYPjVoAG9PL6RlLmwGAoivwS5KU
zZeHXND6FbAmdShMspx8Wkpb18ItT9lzZzf2QBiRI5yaFf84EqqJ36MJdQV8KLF9
g2XVMAHt60lzY7kOOQKN6FslIfMU11SH19n6HYKHh/7cI7fI2DZtHyMPOBxaU+LS
RqavK1NoI3BoxpMvT2JBHTkIzIdPJuM9LllA5kU04cIBtVcOtOWHKpHQekwHvIY2
+rkBvtnkN5SChGLe6Wv7H1mD5SGs7sMl/a8lax4AsHV9SsYGWBvJdVN6QJA3a9m5
2Y0Ejkca19ONaP7x+pCqyx+VKVIWgJCfSVWm8I7NP8Bannvw683eC3CRNjNATCax
MzOZuNM2ZIbZZ0cpl89wRS6MD+1ePTM/y128biYC+UgPF/7jkfrdZHeEfXZtMIfe
EnkNdRrixsfufFsKotlP9Zh5n9B9zCokJBLV8NVYX+Cfk3cSWCHP0c2KWvcpyts3
B3KJWdOqHDRoslIRTKwzTch0E+MyaqrbKPLYnB6KeZOWkBulPhXxerMqrirMckiM
3hm0vpr47MeaDPxlWdSFxlVVZ2rUWUw2QOJvDOPq8gICIE/3cNmYO1TUyzemKaZN
0GrsaGBfyuPNDvx+vEYtdI2AYFQPPF0VdrOBaPiHrzoFKOOavlGGvfzsJsVXwclu
nR1JxvtyzkBnwAYcvhnSSjvG7SmJkchaHIj1FHlrvQDMUnXEu/IIuOHdDDfOsBFP
H5o+ARbjrlz7+8zpVA5VmYkEdcCuNJPK58x43OZ8tnB94zlu4rLoLPM7lwH/yW9q
ZrlLisHhJdUOSWajIsuJwSsUy80mA9GS4ClUjARlptFHLweSGEDaC1pKZ0IN8Ed1
AtaHktfCKLVSsp8qGN1ahXHTEBtQ9mUrf0/dMGFVQMs1AX7lgP7wiHSJ+mIl6sLr
MK+PDoKrdOvL91YZF6OEbbjzbHZKXSfZK8RA5AbWOjZWPV/SDa4ISpU8DqJfOJUU
7W66c8l+S65qSYQBi11NzCmPWtQxrgpiKIe6AUsCcsqgih6dETWSqKw/QvwEFF4X
WQjtM9kHoV5+3ZwdsHdTCGd2nVI73ZSlRd+l5uNaDPI718jIdmYzr3R3dMi3CtR3
l8bubd3LHsGG2cFLF1H7yc1CsaGnLWlPfl6V46/9B+sLrgJHPJq4b+g53xTIZQvL
ggH2mLoWZxVg/Cnq77qpN5jZCSz/YZ0F+3QLiR9WqlG0aDCOsvjtquHM7WcaO11s
ioDXyuY+hPKfvVgXiuwWfAMP0znLT4Rs6w21NVbhq3c2Xg/wP/watKVGaqLY42CV
FY/YvJZPimkH7973NUWJDD6TpG/VkjQiXNDJS/iKb6HnCtO0hdYkqYcSrqtr/1z+
snlf0cQLYwsfFAUoobrfs2bavqnDbcMSXB2IwP4ItS445mInFnKc7IG2/sp1wmpS
BJwDCgQy5lmnEvS+8R5KSew6PljSRQnK59pY2YU+/MStZc82gTTWNNArHyNGUbWB
zC40e5NduEBvoKTovL2pQ3QSXeCT0MF5SSwLUCOhILEp9vG6PHZaH919pdsc3+hH
zBDGa8KkDf/pJW7mmVjYX7lsumQ4jPlVHL1Zx3mMYcOjFGr0ebdfz/Rf/dvdUspk
pnsoL9P36VIwv1rNDrCBsk+mlxJWEw6J5SmmYZUlE3euEFVYMNiaL/IA3ayd18pS
9cHuu4uY5qAUnigI8bJPcHSawBeMwwxUrKJV2DSgXcOchmsRjmOD5Fg1HRYoEoLg
3/ahHS+DRqhZjGC+UsSAkEhXEKBbvioO73HdGgMLU3qv0zPafAOvik1nY/nfUH81
UHg6Vl+q1sSSmrOsUdThiNkfxwqVt3mm3L3JXF2+c5GApGGBU2mDOszdVPL6h8+W
idoH1WBPF+3kTvnz4Pfny711l2i0+AqUlooEwCZ5PvQ/Sz3EFWciRPCWqJu+QIFK
bjZuD1PGYXDvkYoqPjwu4tky2iD+tC1cUkiA3d64UyC8WYbIAtlithkWrCFF+oIP
KvO9/21tZPldGdLyX7eBhcpbSzRTkm6nxNSsKM+3F7+cZ8VH6RxUFQEVMVJnhRJ/
1/GrENRFyDSOXKixxyKuiborsteokw/EeqY8hHsfDLr+FkqyP6i/mp1WD2YEHf7+
7/vGQLuRItgU18s65Ba25j083DYFpd868WM3l81a7kMIDiOMyICgrSjp6Vwa/zf9
Uz5aWNd5C3Ya+U5UiYc5pFOsJpRhBhubGaOxR6bgxaiXHgdDoXebbUqEsoXP7UDu
YtMbK4OyasyWEWBv84khRKGiHTMxK9qar22Y7s2QBG+nuBgSgOw1r2kNUGtxNTnN
HkzOHstev3zOYojlHWMKTf2fm5EeRdrCxK4rtZAn9AFqHcLNpLdPdS+1iDCFL7Eh
Y6iwvB52C17gL1Cc2m0fKMDpuvcaZMsMS3GSrq7CaQ3VDBNrcMz9cLwBRQKara1g
vIXgZddRj1WXdCn9A4oTU5MavRRIvr1VqJk86uKJwl6apGlZ2ltVyQ0BLzp+qtn0
c7tOcMJ7OvYmenUl8NjVwmBDYarmspP8vZk5GIjFV8tJRNNHIfpu8l9GrthUwLGx
ACwvlAPbErc3RDdmUmsWmi4WrRtq3J8gIdHZPZd0PiS6w19oy20iIjSxx+TPdqVs
XW1bcYNCIitVXZclpqjp1ppz6K98ETfunSjGM1SqI/kL7mTwLyMQZcR2188Ecu6o
1F53jxqztDMl0BS0cX6i3RAWhvRGkE8e/6yEdJXp1dGlVmCQrTxykK6bglJzCPYm
TvXTKPMi0i7ySM+4KgNyScvtab4KHNB+KNgcMR985eDHz4zzo9c7k6sOXIcZ1/L2
WobtmlGLEU1MVlC+0x2JgzOfYk/R4Hl3jLq9csbU/i0Dz9neXBgw2zVr6pmaA9gJ
qoa97VOPK9T1Ut7KvAYv49SsKwP9csEdWZzwaEN5px4x9Ri8sm7KJf1vS89dOwW2
J4dbKkSe4AfJ01R8HtZ5fjlj0IGCJIpTpusOlO1e2uo5Ntq+Zq6S3HSP6ZuzQd4i
txC6/aS9+9K+fQk/wbXAVJ1WDtvXOU0ZhNwWfLxsJdxSAx9whuMN5o7OUkRY1HpM
j+L2THHnNCuyw7XTaprLMv9O3V8zJYPFgro7oWatRo496FKZiVBVAxhImW4gUKWL
aaAflC4URkSNYQ4OekFLLo1oJgp6CTQsOyYTAaML4kTzc0vTJZyYxRhOSHcXe1oL
4Cy8KCujJz/Np3EdEPg3wkRLneRxZV2jtvw1FCx0+vc21FMgp3ADpxHsQaLWDmlR
nUc9dyzxuMwzWz5bEEMJpj658FlnsW4AmFqWa4KCi3whltBRHIxUm5395/VU4WGT
Ayt0mDYfLG4QiFS2TrWC1HbbsJ6cUAcyISS4lzebM2ZQW4bY6a4crJCR4A3ikMrA
NWOB8A/R11MoDoxSct9t7WEyz/tOIqj/oP27PihhuQq9AAiLmEHN5LtrIDKislHY
fMKgY6V7OFrE+s82ghIesiB9pYM7AJvOIEXepHMusreOKpH029HFcPP5uR/TELia
V6FwxW5Yc/rI9gQ0X3AQRaTUdl73lo16eGB/0iNDg+/Ae0fEbSkMbqMC/W2RYVm1
mWZIADVds2bpy7XL5vBtlPr4T58geC6WFNJVFzqsQ7re3UMwu1QPDcKGqvJ0+JX8
QuQiERx2TW1Ow9aENqPudKl51ZI6QY1DHZnO4GWwMW1l5V96IGhQAOp00UJvgd0Z
7Dti6ZSvpTCP9XT1KlPxQ8ndQKLYQAvWGobsEDt22YGHGJYOqwvmDxlOhZ3t9Xrr
U65EWrPc8OfRyWl3R8IJqIVPW+RRrO8MVxxu81FO5hnwfcuWPOUEdeqIUNAtKxji
hE2eyWhyJUC9OIupsYqqbO1yKdvOKx2kd4+VYq5DxbqQfuksjoG0xssiIK5ONNkQ
j6czqLz80vOc09EsXeBHkHrsiVkYRfhjM1GoUpVIn0k+cU+DyhcoCgCxcOb4CxYd
HA99x6qZ/bZQV7q1kDdXea9/gEqAmWU6okV315v8eaBJep1lHjzWKxeONx0y+ywu
qZcDXN3HM0WlZlkW7xNuQ/UryxE9bOsJ+Otc8dfYS0heRzvePp95vsNo4YKYTQYY
5dB4xUEA0LIP7+uknYwYFam8StYa8tFPy6fiyh5Hc9b5mVJHU6MvckSNpcp6fsiH
vDbj9OB2zc9k6E/Qs7bij39u6RMGUztGFyhSTfMWvRhVIWpagOC1ijRhL2juy0d6
GQ8d+dOaxqG6zViFSz+5ZuVqbxRFljbIZJj1n8HPBsDMongG/khR68bpH8zAjpgU
psTzt5mCfLKUsuVh+9SF80visH70S2XwrnZ5CjiMUfDxBg+I4ms3waKDK9kklHnC
d0MavaoewPkVI0ahPLklss3ckw93EpBdALsUlYTQEvGUrGWSJGKFUe6GdDt65xbs
fz7qJosrungKy8ATdJapT5rGxAvhXScjXooNZjVUCerpeHo/VrBKXjrbo6Un2/Cg
8xSnP83su0A5TmmLKXcZ5kLSOYh76FPrXHOkHG94GQ5NHTVJjnJK2WBAfzrdI1/W
uraOq9njOd2zMMSrzWrahPrkcLPiOK1xGDvsPVnsX0z+dVF2/i8GUoqxGffdHcHk
g6IlI9MGF7EWCysf1XzCxcSPHpLj0wE3PNO6Z9MBEuoqJjx113cscbHcsks8wNCa
TmgfRgRpnJm6Er6n/I8ESQ49+ESFBxmYPxaeMM2lnm5vsJc6z9wxFz2f6ofdwKSJ
C5RWZJ1QafpDfvTcBhGYcEQgsydnbA/jnZMsyzoiGuX+wgmPF8wDHeYGddH9R9TD
+4DRCzOJxgE8SGvK3FCYVWvoXa/6W+gn3SuJwnzJqmemfO7e0djA/ixY8YT+dK/n
kI7vonsySNqte2TTDz7mmIZus8HkC5RKueQv9dj7FKx1/Q9C2R5DHlP1TG+r3mjZ
NdoEVDxOyg3Eer9QEe8V4KxKU5NCOtxqmMssqBCyeJq/IH/J5ajEUBH4VJC4NrOV
Zaigsu9NEJWtqTxQwREBfqviJxuA4IOS+SCb2Yslg0c/xNbMwjZvCW6ZPQYZ5yI4
N4IEO1dS44OtRFRoWWXPPOcYNO0LcQnBvfRfKhpUFx3Sw/h/4ohSU8gP+vm70fHs
m2GeZ3aRmoyXvHPS2sSgUp8sXaqUzbY4jEuMknQ5w9YEuglDvDoXPlhHRX+qrl6l
cd4OhYmmz2J7xZu6uIdTetMJsgxdTgwH3Z5qKjlECOBNFePMBfvpcBgOAptYHeQj
OwiHVnGQIr/dElsWOVcygWMkqjKnWyguQsXYULh/cUSJexX23sCANcIzBMHct1b0
0M0Pr0KJHmx6Ek4eedJs50f8dns4VMeembjO8LDyBzVWxepTQOe+Hi/CZWZs2Pwu
lVJE8xkugjI1HNrnc1ANpaiXfT4ifFnIjTh/6Hx1JbG0st80oFfw4xwPW+eWZCtO
8KLdhy6XdwB/lOGVGOB18F5EzJ2H7CvfGiM9QnrryI4Gj3P5hS94oPrRZ8VASmVh
z9zs5/6OAl4QZTUIW8cOCUI35mZJA0xihGtHurf8yZ7PiXk0azAmyJKoeHwJHEj6
gM0J9nZ8Js8mlwRu4+CWoEcW4uzlGHP2oePdQDbTTt+TmuR8U6pqRHsWYCmsM3Bx
gyOSr3BG1ie/9j8wftgyaJ8wPtP7k+Pga8aZDpF7PqX90ClwuP1XulB/o0+DM4Aq
BcjMuqfEv8knYwxyYXefbHFMQpKH8j1LUzD7m+K4Raxf3CXnV2jdrvOLitmt1dUu
Z+UwMGXdevDzEZGExPXo/eujZnbOBcs6r1wX8DujnoDCCGtaVPdriTr3XcPByzIl
r6tor5pt/2PjxSICofISt1FLDwQ7HkVREozAAgZv59yu56sJ6cLNz7LITG/WqtWm
Uq+/JeyXcJKPQ7IfJOu5qIqv8lhVao/uDSg8/eOwEmx6681jALq7lXZlo0bWX+a0
pHJ1SdBWZQoFDabl5UgAvBzZFU9b2nJvJN0mrHwuHwEEfJPpJrIujs+T0PmFCcyW
AbBEM71+2K+K+npEzcoNek2618bVe4dJyCiaF68jSVq7v3vPtJbVoCfJTgqyYTFt
0snG83rzzEBCYL7KHNjQ5WxShO5hfdZXlTYCg3VSpINLYbBFXxLElmfYjWL+uoY+
Gz6bZ/WTMYQkqn26fajas6TtKkyzfrS4GJXcw6ZIW7RtddWOC+C7NrTbXdsOmLZO
uqqShVG9gGG2WScKXfAt9QMK5+kFX4jdRwInijEdJXOop9iYrzT/H0FRQBgLoRxH
R+dEET2tgFdjUvra7uBdHrJA1w+xPNeoUB78hz2w36wcE+2rcVTb9sERRA68mHiB
JWUtYDlbhsh4hEPKG28vqxjBeFHts27VS5JbHMNZaJJKe+R9B4ftmKJt1B7WYgob
ISUKXWBWYwc/Px3S0E3YihS65gFF94wA4WMoz8vly+TamhdorBpWU9L3IZduK3dg
20Qz0CCOR0/XCn/v9vB1uDodaGjhNnk03rLj0DH2Y+YaptWFy3rxqQ4FwLmSf4df
DyyBJtXNpZLXBFSngQvbQ4/57G3eQkPgJTjUSxGmwd32SRaG26RhsTmrs2C89zTT
kdAa9WXbh1wKIdRw2uO6toQdeYvT3zrBS3KcVozNRypR9UX9+JW4xnxmIZ09X9sl
Zv951D0WAXU8BdYKf8sF1SwtyLkN8QrSPtdG8k+v0N3AZJvPTEzJsQ6XYSQ9eTtC
GaDv5fZ/E9A7qQ0+dZIBf9ba3rIaJ789Jkb+07VSbMGkMkye2Hq0QoOV0V54Io7D
pXNFwiKBBetlhLCz6Y9UxIEdBlSk5Ak0EpxtrVlShgEjc+H4n0w9BoZf7BNg6C5l
2svWr9DD+DEpvHfLKzV3ej9u7D0gOH6XgVJBtJC7nPtDOKAb09bbMb2BuqepNdXa
//PK/Jx2/FfGRvK1TjANTj1aMY1sPlMy9GIyiMMGACGcBbPsUZGxAAE0wNv1ccuX
fAyFoPBgEUkB/IwuZXGWKO68jGVkGq8vj3OyNi90+CxrsHm5OJWQ7IgG2Y59jozd
FI5+jFLbc+ftPOD5CgHEmtEVkVkLzs8FAFuh4WqwdNvUfT82vcNNY4RB0MMgrzg9
fmcFGx466nl6SWAYqD74R5XYULurZskkTl/BgmmYsWT+qBiq2V4HBvW2rea1Jlkj
1eYeJDCH/MyV3xg/pWysCjyJDzv7q19qqoDB3DRlnKQG9Kt6ofBSGMwcSuxlzJ5k
zUjL8Z6XOgkpHv4WtFszWbn1CkMA8MUktYXWEobqgrMJVMPD+YFYSVy1yPdDglUm
bw1R0P6PTmIpYWuLs/FmPo2n+zY0UNgVuW1KY+Z02dg8gmEaZlPOdVct9gOMyL/4
xdONF86WwE8HaVLrZWdf9KEf0/TijDtcUhd0JbnQ6gG9P4qLdeefTbawlKDkvNhi
llDVrO5HSNqz9TRts3ETktTcrLBpxL62OJjiwqWoOc2SnIesurudvcarNRx2238e
JCdPmfn1s3W7cUJT7U4nYB+lrWUkfpKVGIo6xB8YxlM5mL5CgjoiSvN4e6RPtYYr
P/+1Ds5+jMTca6GfC5nZBUd2pR9JTTxLgM7tXCdSD/PKbW03Wz+g+/LQ/hNjXb1H
JUQEGc4WjBWRqcSShB3ffR21geTBJ+XNhG3wcIPX3pnS7YsNr7mjhmRUQCNeuuhb
GV+1Xd3yaN4oD5hKDyNxUD2SRerdPiXhnz6GiRyRYM++tmKciikEAAQzJPWIzjW1
VnDbu2Sk7xwjt5tSCJgiIquqWE4OEIbvvQf02tdLesZ3fRxT969L6xclSe8fBBEJ
zOBYXMxuH2Of+QNeOGxb4wY/A7eY2gsKDAtmYnVGcmOBzVGD6o3sYDep1Jy/uM4m
sT59Un5X9RxU3wNTrhMY+SYSG0W8w0qWy68lBHQRAzk/FWNQJGJ1pTvWmXCZCvIG
7UxjiUsenv90ovPfyJLB/l6WmmRMFa2N6jjnyPPPu2ubmC6poeZT4bybIpKE6N6Q
UWRhYrYezB4xtmUSvNhu/lf8zrf4ttzNh8HPZaVQJ0yEnpfZm7wFMoZEjdZGUpCN
dRzdI1rgw5dXwQ95QJ1eM/DuWE8KtgN9yAaI34TDgVwu1VkhHo4D2iOfxq1uTQT4
xqn+0EyUbn5REH2S52UfIZjDzjGRZs4adlTRRiHk02U2p1BzHplqLDcxE/xbZq1h
sTcjVdiZDyfZ1MEKxfCoiwN56a0APtMmIS44AUL4AIG8FR6WC4BbPJ8nQiLzHkSI
EU6tWiol1MViYdSVzIwyJDBaUUoD/GgRzZVxyBAdpIFACYBNB1e+2uUJ4JeT+hkp
LJtOGT73YWgAxN0b78RR2CDCLovY/+PT9SpRQZ+aMG/wGKXfz+7kXbhv2iPf1Lwo
yNjTW9dlVWWxzvdWIKLXJvqvFGOHH5SO7FHoIPRGoAj7n6ci3mkpwx/RAoZZTGI/
aSrle0SkU21sacQ6JrhQ4wdzaRwtOyeVtCksZZAf25JbWfUUpxtc8xzURnPjghb+
PBJLmH8Alga0TXgiTzsRHzI6uk7omkQSeEHl80xE9n3agQb12OC473Qe9BgaB000
OJ8KuvQSXgg5BKbyMDj9AO57xaZYX7NFuiuNxmm3c38soQPtyoAhGkaCzkURD6F/
X91O3Sd1AdEPUMQR18wiRY4ObzrIdkOmysyNtVgNU1J5tBkH+SWbB5S2v67iJs2p
v1OpD9f/aUKZmz2iSFGZ6nRiRFArUv5K8sLgteDxrbPECvXhFktwpwbtjb2XE92x
TxiaDQhsFxSo+gdj8OcoISMUznele/gP5Uc7WaKu06JI8RpgpIKwQWQLh7E1aojf
mgXWOMDkmsFvIT7R/ZRuKewLiV0kfqvYO9FnB4eE6R5xlmrOEjib3LBi70T6Dq2O
c9lV0z863G1/53Z0FeiLdZHA+5Bml8TFupTEyMIGdYpTZLlIDRKIneZ8LizRb3W1
nSEcSHbBIOXhE65SN359WF2brswZCwZBts+Ltw761o0j2eHLkRNNyIBTZ+J1qGtm
ODeOXtx9oLRapdaDpbtCsvfUSwM4Xlg1G2cw7SlMb9F17HkmWGSfrP8U8AM6OjXU
DPx7IMOerrV+H2j/qRTO54K+Man4s5/DowLnagQ7mIYaL+FxOZCkkJFvJJW7OlEi
Cii44AG9Fc6hB5z3YWuijUXyAr93NUlfJZycleQ61kEkWn3Zpv/o7aX2SIbtgxHv
pkLpnqPEZEtHwSXNbVExprYwv1JIl41dvuY8/+A9M3PRz9Tkp43RSpqPGfLO8kyB
X0+I0WK/G8nRBBZy1o3qrlh/QCSr3oC315qatv8dZXNSLPRgGbdLXfo0bYKk7mD1
j2JNTS/EA+lNWH44I1zhPcyC76oGkeU6cGglel2JAaH5iO0+B6Aon1/z8ciNSMx4
JudCURVwXWoOpqAvPFOyQW8b2M90DJk0VSpBjxVXgf44oaGru+7djuRmyKt8qLAv
ktcxqhv9qjfW6Ss1pb1YGFIo2w3M8JBDyjADkkTiEQ+Pcgu3Py8nFO8U3efw43sp
45BB/J615ILIsM78Ux9Hwb1tMv7Ra9YkuXoC5GcW+GIydKaVXjQHa3oo8Ua1Y2c0
KTDaBPma0pn5LnVP6HGe+kKqIt7+o5IlZxbeK0rbPfyTWv+4SJ2GPc8fYR035D2x
zBUhNVlsO2mCxQV+HnvnB8S2sIsrjd+C76B+8mfCQYwDZFFKqFx9H+WfTKX9XSH3
QoB8e3w4PfO40nYl0ZhekO0TZPfGxUNw+eCr96PkS3kSE967IEdUTS6mMDT7oar1
knRW/dD83GLvgcrKXgrqRBwFruqSmEQv4mJkuuIPXvNh2jR05jWm6DR7MJCRMfrc
AB3Xc5ysBC68CK/RIv+zu7TP8hZGv4ExFlKC9mbxa2i6xKcwDcQtyOcmU5XF8W8b
199VMongmAsIbQuLBZGQQSEhSQ/OP37sPDL47Bh2EDnSs6aLWY+1p/2H0v51Opk1
VqboE/4ffZqM5ZPcw5Nq8KK3+78aWBuHEIBi5Ayq5NFqJ+jK4nR5RpoR7WM+U0sw
kk2c9GPYNmCPWUc5W90K55CiKdhyLSfeb9ldwhlD+EMRlJHJx2wh10xS6y3vv+kR
V5cXPEhjPqk7yIQlqA76Exr8TvZ17iwQFvQpegOEG9nKF9wUNgxRefzfULDabHwY
5juu/X7vXt5Ac2DWAPU+r1d8l4zorYoFay5eeuPZzsAu5qclutvmJIP4q5vJIlqO
HEFGWXQ+5ao0TX59QfawFI+5VNcyf+xGpB5lcRHNI2b7zTz8mhGltIfNAda3Ry0+
VZ2MYgPIFG1+c0bmq+Glzbggc8kcGk+KQxOUjW1Wje0qvoiIqQTWDF2ReLakmLyx
FfZc+Dc+JgMdvbCd2rpMcry22kqfnin1xVmtwY7rlafElMlLx4yjg/awkjpoPNET
WXO8iw4RNCfpJk5t4aX/O3A48mKFNm39YbsPUAV9BLsBWKNLyrPkwgbIWLFkP9iy
DUzdZmDGjykRZmyfceOIA1Zyo4I0uN+O0bfycOKZU+fW+U1sHf8HGjfYqiWWFZmv
BM8Vv+wQtuCU54xGiA//jDnGpiQGOSfGvt1oVKZlU0jU1zeh0ay8fKxwLAkUfHFP
hyB30ANki4yU/zKaxtAsy6bly7i+EAJzNodKmOlQ2bGF3gyuEj1DIiS+VieTQZOv
dPMaRR2frKhNAMbh+54IzpG52/LoalEaIZ+yUnSpUGX4dvqR1Q5grsOGvTBydAMt
002zC6mNYcOy6g0EGYp/VA1/1Vy+JvEP5h+bJdCX1vwB7oHw/VyXt6qI+vDZKlR3
T6I+HIsxULQqlJy7gCP6TBtEpl8y/fYD/BzP5psVp+jm63dz1uOhBlxLVstZIWOg
aPz2Dd/8OA1pGOCvsvNyfvehGZTimnZC/YzqsIPz/TwKpPROfz0xnyfjqSxRV98G
omCUKRc3TQResNXnuaOq+JqxqfHv4HSSFXDs4iEn7T7ZAhr8UAjCTCO5d7XCZa8l
lp6FKM6vbIAt8ZN+p8jVt9viUgQAHHj4enkBtuejQqtql2i+++ObqnwcuaK/+CJH
Ef8YP9CG20xxvmUrA94bGVdSxGf1vpyXjM+Rcq4EyycWlYMI88AWt6AelqoVU68l
Jz7hXGH/O7WRTDNSQ5K3FKEVBI3CNIMzVn3KSluPkx1l5TEH6jK8AP8dzqj+tyez
uIzzxbCKPlI9ptuncSeCWMG3EPvNAd5DO7TXJQb44FyiAmd3e3gQLTNhjEDb6lSa
BGaltl3fqw9gv4FpOS5yMaHiwHVjZLzAVaXVsXgxgnYC8DNKWtHgkKf6b5DF4+tl
h2gJZ1usmmzBfkrLY4KB2uxsC4zMR6jcxY4s9LqH5c9lKO8pYxn/CM7qC4UWrIfw
nNxCLN8YgiHNvQHjX22ereJG7+ekXSiPmq6Gp9T1YyXh7RWNuarZndvtzLQR3T8Q
1j3yTHJXtjXo+DZmWl7BthSV3TzPgRNkc3n/mAdIQ0KxNkIzd3w71KxVao/7RNkk
iK2WUuLzb84O5EhziqZH5uK93/IBj1R2Btl3ep6msrvFBe1zBFNDcWt1xXQ0dRIW
HfFArkdyCvlMG9D/biVVqqH8n3qRhbllYBMwFRItGXXybi/PZrQMbRyBdC9euSIu
vb4Brzxn2JzudkfRLeIVlcbd8BRXF/Go177zgEt+CWzP6+ilhWtBK79/9yN6gdYf
WKjZzEnurq/dV9hn0MrVIXru7uBIqBlyjUMKOWnnQzl/azWrFv+Nax5YD3/F/DRz
yHKjfb3oXUTMERiEL4sQpuMqrfeFLU4mdTJrflmd/W+N4x+y7lHfDRehZ+W61qCN
aQFeKs7PFOG98Jyxb85IOWwa87TxviPQTPiaVPhicFQQ1sRhJImW1FqbUfqR1gym
DaJuYNiwihjCDKbUapW9TFeFME38uFkPWr9AahNuyOCTfqgNYmL+naysOR4X6O1/
cf7zsL3bRKOF1jhamSwCquMP9gWUPt60cZV5h0Mv88tjXHD6lRINX566O31exm1A
sVHnt70Q+dEMjCISV4zF5sTOc36K4oX2Sy4L8n/yAg6oW6W6BB84STK1x/czB9dc
muPmgK5tK4T8nhWSVfxrqltHSLc76Q30YztRLoLswgrh48/8n4R8JhvBhiLf08xc
kl8Ab9vhG8pRwyY6WOXngm3XadDKPQg5CA2JIHOdKJLISz1XCmdFVwbxu+mXl0bY
3SMMW8y7QwL4URIsFU6mnqiDn6HW+QZ05i4z9XtV3pwYYMYKtI/32rd+r5Ge6I0i
Q03v0pkwziUJkrQyWcr+YQvTcnN0D4HTwCd+ew/P+7Tmcp7+UxkdwMU98gsztM5q
xq7UGakF+fy3+1lgWM3crjDcPd6eBqgX/0AzcxsM1R9WA/LIyxGI0GpoxQbn0ZcV
P/JJwkU9pLX9bPJ+FpdCI2VZ9oZN3zTOItttK9R3+7Mbqvo4TMtlN714LK4dJY+T
agNqyBmR1CUM4cCdaqB2gWnbeiwkXjLm09J1Grjk76C0Q88SZ9tuPPGwGgL1AaFu
65Y0bywjRtwuQr5EO3QRiW6ZgptXTwNNYixKmMK2tvv6ZPJ9ZMDMYuQ6rnLuzJhM
hJSLn6IVkjFhsmu7LFtrZr5GX8JQRKu7WEpxQrMeclP63FhViDQYDpS9DXHOPy0C
s2UxaV/7EbPnp92lYyYrsmwtais2MdVYDT1acqBoTim5t3m5BWTDHiah0Dgx+3A7
3KAcpVvTPLgJSQDdJjsmMeyVrkLGR+7s/0qvkGrPPJ0IazooD/6T2NjMkJcF56DH
lCwcT2/0xOi6v4GVhQjSim3KIEplmjXxxU1dN+UjEbpbOui9WidkOtHehjJ0x6N6
oDO4I6FZsUT33oq1d/uXmio2dr0vTzTIHh0DNrhVA7XeeuSEiqkA4m7kh1mpXZ+n
lu49Ge+D82j0xshgu+xisZi59LJ7Ptefl1j1QIvO/wA/ym0ne230fj7qpl0iqHDQ
H+szCSI+9OVnL6lnSiPPxJ/so1Tts+bWXl+JaWy2XbgwW9ePgqtEaM1PJlrMQZLV
qgxLv+pJmcJ4eIXFoaKbCvCgBXwhLqX4VaFDeY6Uq6j8a7ePVFEvlGT/RlmDHPxE
zDvoTV+QemXPf+a+XJU2m9cWK+zbulRh7kBnFyCGMuSk3qhgJKyhjQ7i4rV8SN93
Qpwueu/4hgTnAtPB7MVbtw2Mqxhhf6pugVrIW+1QjhEs8WgbN7W4Bj042HYDyF//
QhL2xwwiml8uyhJUt7I+0HbzLQwT2YSW7l4D/oXMUX/Ek2BfAKvmMfvl6xQRojWz
q75PV/f5yKHPUPHTGc94e3avoyuJEKBDS2N1VAHF7cSnfBEPimCnEed4FL2Tegbm
LFgcpHTYk8PKlHwrwPYqoqWKnkZ61wtAxSPP7SWjrnJ1of6xcTgUv7LkLhy3VKYt
WN7sw5LsTMZVJ/YatNvMMfKf/LKXqkoIVTXygbnGB7VDg40slxklBNGmydUW2moo
rdLCQnDPDjfMjJBkbnuxLOvbsW6HdGFzqiG7V2p9TKzMB52hhUXwhTQZX1aPbgWB
UgEiaCLTEWGBUq56hFgKPXkz4G/1htlPI2/tAlCjH0X6//Pwj07VnDiA02IQazaA
XCOW6JBh2O+Qt6V8tPVIFO12t/B+DLxVJK5c5cKtFCn8R6vWNsfs9R4CYzLK+PhY
pjqL9pG/6hYpKg7jQ3BQjV5vzsPD5j+gN1Dkfx/ctimGJaMOA7CgUxCVDGlnZAOi
l68FYXSUJt2NniJQhndkmpvtuE8Offu1wGo0lZNEpDefSgNUKLpB17DdnxQw7a2X
dwY9Td2ytlP/ZLrA43DOy5KqdatajUvDRdX5y4Pvd+HPFI9R0mqhYTiYvNR+B8SA
5OENt21S8NOPGEgm3gxCgNK46zP6yXjCCnckjs5mmmtl1Lm28/0N5Ib/n/Vboe3V
kXzo4GXrRyIom0ztGbF00gnJlXOByapKr5Xw7keoUjzb6noL7uFjm4jnkL23c5xB
ICIau6Hqq6x+nxyLorcYCoajZFdMT/HhL+/PjyqG1ijrBs2t+dtDbZDrrTsgHWeH
FcgaNtkCdc8GJbyluNVuWxOA79hnV0ZMcMJf+EWffGjmMaKWQjxCIRYGnzoYlXbj
a2sbmwNyF1jQ7KH95B2X5nmD4O2zNGOrnd+0GrN1hM3t7VHzLRMjkRQSgS7+2FxY
M5R5jRZ9tmywH3Ya3wOpMUS4BhFplbb35FlZvUAm5OpGnpXF3hy4t+/jB088oadZ
vKGUJnv59laiQSsW/uS9TttetZ1Y+0PjK/XYmjSN9t8bwlJcPPV4FsIRffcc3d81
YCyCR8pIJkZOmemEinPyfym+nUnPY3GSuQPrQaLhSLziUc8WL2hOlzE93DWpKcaG
qwLsbQNcAH5H1Ouw1TrCeiUoM34IjWypj+OOrO2TONcRWlxmQRVUSPq8EqmRT2q7
6U7Srm8BrOZngBOPStlA4wx5JMi4lTMOuKJxqFQGrYlXhFN2yfdQoJYdDSd3Y9Qj
fD878njQj7vztstnOKT1DbbMBvfLX3O4Q2cHUaRxpo4FFOsAPezEzlbVnjzbh83H
KN4ShTmgMK3BlzgYaLl3eKVnP6xfv34Wze3aIbQ9j/UxbcYQf3yjs5fvBZ4CR/a4
K6IBXb1Dr9XhAqpNVkiBMcUJLMuqCNNRoAh7WoY7E58yk2MYcdMj1G9hxIVFqmDh
y6MuLIgFpn82+0u4/03bCD4dM0nUX8GbQ2H+JjKPEnQrIE0nSoOzqr38FF7+LI9U
tQKX2UkzDCI874CY3L7+E7xI7Jux4r0x0ZyKplFwridI5vfgu0F1XqpAjt4pLaDO
mSuqUST92JmAPo32a7j4XPnlbAJ6EjO2eCUwiJ0p5dEeFMe38orTSC1tAMM7IGiI
bccEm8WV8xbmv2wq/okuiec/Xq8JIPuFZ+zKAKvhqKHGvGv2JwdXoo2/ENZZJw5m
80IC92I1SxCzjNxW9HVWmLmE2rv3/BZA2UTCK0uEhVMELtu6XQH3bzUrzp+uTbfw
nn4zCEzKXV+PLG5nCFoH3kvsoNrB1X+2QUha8i69aHFvStvJV2aPFv3CR4DbPa9o
Yd/ba1E4VWRmZRqqrN83rQvGTGfK4EgL9wcyavvXfm33jUsXVckzt9TXAaf2IMAn
A5fbx7iIbPDWPwRbdMk6vfayQ+kWJK0X32mXaq9tKEIBh7cf0i+8b/o7jXZwLSiy
zup3/qUjxhbZU3PDzy8KT+2cKKX6UHM5rn6qkQmQgjF5YuS1onmJDXWKb7fKugXf
wNK2CXy4/DSk2oXxALCn9joOaau5YowskkJsKqDRCUuMsxKkSzRK/VyYCf+v7GUj
O/eSVNdp6ZUbogUdqscA/cgXCHtCvVVepP3LTVUWYWVJIg93R9+VHwcviPdlluFK
MWAAMxmlqHXBaVz5qdCn9juFuscIlCOefBvEfpOCAPwE1KqsutWQCVBIcOng68M4
k6JWIJvi1p6iNJ9EqJ1nNxTB0Nhb8N/tnoOuYjPhMrj+JCslIQjPECv8JkQW9Czx
bpGyp/OHI+e8nj7IFO+bu9YAKwr8KhZC0UcQUatQqTC+U5jUdHudbdlF1CQh11DB
PGux6PScgrAuW7mvKZplA0FPE29HldeOJHVOrnTlo6vTaQx5iHIV5rvKSy4648ri
ZrQUkNeTUB6VwMlz/g9IgIenuusHA8tYgyXeyZ9A0VypVAVGrwdq+pYfKnQhr8VI
18lG7eNVU9tISXIrDgDW4MdmoGVHUrKh4gYylZVof50/v5RNlqFSLKjQCX9gIZcB
taWUuTcmcqgkqwb/by/TtuPk3KbQgDdQJjeSQJ5e6sinOx9irSIS6vaXUy/rpGH6
HZGvZXIIeTc/LwfjAtlZP2UE5Wgpe9WctAp/W3LRQsHowE1CFQuUjOC/VVpPK7jJ
RYdQSbcGWt9ucVXuZvtAZn8ZajcxmhK36fSuLV2G4F6EXGWBnXE7KYk3CTaPtBXs
c64vZ9M8fVi4OFXQ/GG+Z0wVW1aBstDlBgwZq5RYpCGL8yPCj2PHSpYlwG4/W3SS
C90uhRILeXo6yyFIoZNDHg19MYSLhidQHqSnipJbjjAOKJrc3/EptTJQ3/ygwWUU
LjC/ZA0Ta4WjtXyAWyTbcOFEXRcim88ERrupUJ+G8LDlZWlbdcCRJEzkf4hNLlZ2
wYg7qM03OhOGpJrYrgBKMdCvg4F1Rv6v++Ggqi/qPhHGk3UgYF1iawOqNlEXbwIr
+hbNSsXhv/Ekoe5Mb8x6lK+diPdZNaMTHjHe+okyAxfCjI882eQHogeqOkqUsr5H
qCYWGzOogcfMP2mLfItLYoeXH71SrBmI5jw4eGqI4v/nla2Af18zkMA/IXvPMrGq
7iO//bsfr1jisvJNRPvhw0/nCuTTyim/w4Iu9GgnUVRJMX4EThLWIpUzFWV44z7x
zemkAWjAFhSmgZSep6g8Cq2rCpgOuHLBkBTA88CEAkAcGsOIsixjKRJQooD09sSf
PSuLnIYpo9/HqWez8G/1iVKSLogz+2RcsP7ByB1bzffsGHk5ZpOpUYmB85DoM9bN
5KBQCiyugSJAFqjwTGg4JBDHh57IRAkuYPPxDpytGyM4cKNKYpjE8GRDedLssvzt
ERjRT/zwNtnLXpCFiKm27rU60uKLRc2Ptzpv3TGYOwKyLYaPugwlgGYKxkFhlnyJ
XhaJ5jHZn1t1BcFTC7Sv0PrAT/918UpxZvWU+Wnj7bG5b6a149S4esQPAAGbLwjg
xwhIgsJRcaKKJYWn7wnYLN51PAivO4Ca9WG7FlsYkBvy0huEuGWWfMj+lajxgLUQ
p3gA4OCXKLbHZDpU79pIwhxvIQgvnHB/mTKNj4FppA6Cc8ISsy9ATUnTIzDLjHCh
CSllAtRccAb9Y+ry7+hIjad2MlCjscWhjNfJn2op3s3QXnRzF6+hPRzYUu5cLsC0
8rsB9HEAejm8gZy39C4SK3LVoVVxyFo1LKGPskR3kyg/ipdvK2tY5a6wbNstdqA3
DgX2Hx+OuooRWsmH1q0q8RW9GtmQlt/kDvKmzvkHqv7+0jM99/vEeyhATA135pr4
87nsJOxXxJhHGsIA+2jCUjV2bDx37ukc6QyEubOsQ/Qdkeo3l2oix1mR8+jy2B06
VR2yRqobQRhM/vahHP+58Wozh3NKOA2CY4CYIh1hN0K1ItdtNipZoNUXq35iSkZJ
zxFNAYjXYkzZXSgnEvoJFFs4w72185cXl1l1Wpu62FGBlQd8Ctq09vvTzReuseXc
/3VtZ/DDmfZBP9az36T57tVzcxynIbyTStSWHelHcwzdUSkNR4820RgJ/Q0wZe04
j8Syqo0dh1aSb2XKlMUNrArCXNer24b2yRf4VBbn5RJoUv/PW/6011b1n1ECIEK9
1FYRENIiOSM5q3sssx31YacKDT2h7888gdJf2cZqecUhGbGnufIKZIGsHRbRF/3I
j7Z8AcKJRxXXiVimdZNL91f0+MfTuEFEujC1+b74RQczujcLapJBKeFO27ykYLyI
XYgSHuDYBqpwGGwwsh8VEFg2D0khX7UJ9Z4kSxEmsaFUBML76ZjFGauN5wdh5bOA
D1ECOOOAEDfnS5KZwyKjn+SXquiwMJTzNAL0ce/y2Zy9Z050eII0jIBAjZg2BKZA
oLSyYFlLS57UwarItYPzCqQGU5g0LSnD5SKhSceglA7USRKpGR8VJM3fq/2a7+m2
S3a4T5PnXe4EyH3deiTw556E5NJUkbZUCICIq21L92FLDLQ76Iz8nR84Qpb67+pP
14FoWE0xIS20Hu4Vwm+TcnzEjy2XYPOkSfGXth4k9zel5hO8N1AHSS1B/M5cT+rO
onDW48YPZGJ5djGALGsnjmudBkriHj1y9anoJ7w0pbcEDx3Kov1ClbOD4XAv6o8/
E/IwwzkKV9+lENVMP3YUx1/e5N0B3DtbjRg09VZCvdgDE21lju4RJIGWBrF09/Rb
Rp9KKVi5M5TImRaAsQ1arMwweHYpOBfrdp71LGui3MirecrHXynb8CmJSGHd0ij7
+rzNqy0gqbKb0cOtMGKAV35gR24+qF6Bsj2pdhOiJLnvUE/CDbe3Zr9SQrZ51N5k
kY4WYR6mGsW8bTTM2W+MtJU/DhvjrcNSHLZ/sNexTWuRKljx558hQ4FZ10aOpdu5
f7n0EbMJ1RT4Q1pSTr5lNE1/hYUTzWwfQV8uUA2Wokrv9XAXxU80WbOUksjO0ERl
H4pp0YeXGBXlgUvh3IW5W67Rdx3q4ng0ukHkuchLmY3SAKupl7XMRHwYHcAabgNs
WH65dkeJ41WugRGaFjtrwUnFIGMA2xP55bzlT5Z/RxdSywxzdMopeuq3ZxML1vQu
5ySJqSj+jIuuJKksbc4rlPrbxygV2jKxyZeVDqA8zD7ilxG5j+oK3TV3Kl0ukmpX
97+NcG1LpTXfPqkqwIpBVn2sU1PTLM8wFUaG4VSHhK/RryikyizsJ4ckQ0Mf4o3W
A2Fez10Rf5xyVpF75HVLR2bZ+uPHJieOSocNRfL3HGqUIlDTGuyrB6Koz6tBxXBM
ACYhHhSs10Cy6qk3Ks8M0ul9DAWAd8a2wXS2iKbIbK7B5DBVMqcKXdZCOiN1dIUm
0b/jDzoGWAZb+lgZYQeLYZtwmz3PVRxzvg5T9pbziXlCFo08fXGufj9YC+SfaSml
rLFMIAZfRrd+NNEN2Zj1EbcUGe6A1X0TNLYHGYScI7KFlZJJC67tN5rq/1ZhJOCX
SpHNkmjzRuWGcJhHgJicw0bRHUEJlJnWXJ7bzcnEMwgp1SBhNeBhdyoEE+sWfa4M
lRpiCvVwDTLXv3P1su//7ZVpOObLsPKJIW+QX0Ruy9S9PHUrBc4zx2BEdPbO5420
RKzr01E1xz81kIq8SoYmVOkGS+GXhxKi3GiW9W1KOmbZgYT1dCc0JYpgvyGSYqnT
hYNSTgK3e4IPzujH9mE15ASyAnRDtO0p5KGlUVPLjTqdIzezEfMhGYHmu2qXZA7R
KjCwl6Ty0ins6ncjA8U9CmTiR3U0w0Az5kS64X03Huc3Hvh90BxYodf50gb8kwRG
3VQ1saJPC9yNsx3GhRkz7Z1a0DfBk2sSMtgTJTXF4z/qgLifVDiEQNi3mPlecyV/
B7IaAwgJ0v6qcxDmOILvoRUgQV1WyP7BYnN1LyRJdAMh0WsoKBJ6pttdgBflujcH
bewc9cE4acl913kDsdPKrXmefisGFh8dmyxHr/0y1E4dMYEfOgqswcNi+wozYHyD
ICob/kzpA17nx2/gKuiAIhlLlsQ4/75LCsRNi90s39dUmuMY/CJNqlm+2oM31t2R
GkTABFBi+ymsEkeOu9rqLznV93jZkWqOdbJWOAdNQz/tyqC16rsK8EAjjmvt0SBO
HqeS3cy9JymxjaHWTJfy4UDEfLxY0X/OsiUgpQzCQzyRYJ3gw2b/saFdXQBcLvNp
/CmiHb6R4LbmlBRtM+42brjd9DUeAx/wLKLMHxlE2HLxFd3xhajYfI/hhfcmrudl
vvez9oLxYHMiXEKVZjc7byEIaAgnFBmFOriUuJ8g225OrXO5tv9U/mHPS88Pr3Ff
mdoqhAGPukqOB8/kbbx0Mlcjx/hPyi7YGO2dSoO5as15iUPinTNG5vuUI+ZB3Vhm
H8uNMEtTN1LOC4KwZBIrT19eowCR1t5AQOoGt6uP9jX8NQY7fsqzb4h/TgCJ+kzb
8hn8eX4JFlJY604zW2Jvk71IyCElXlQzU//SeBSlpDGGMTEHfuh0jJrIbtCRoxg1
7KH532m3jSUo5TBFnIWcMiNGktUcOk+QKuKV7FooK1RMwNidHAlxDSyThEuOJS/O
+E2ESr5VboPLH8FOFw51HOrEN/pMNovBYMAVqkalUxf7tiU4V5pWOMWR8iE5CPoN
sn24xoJeQ0oWxwF3JsVZL4IjxrAW4ujcQ2NoQmErgdb7HcGnli3AAlJ6TF89uaKK
dWp3B4mU0B2WWX0/ZiIs7DOmnq1ExZuR/2SGtOztHJEqc+0LeGUQ4vmObNRudeD7
sLeHwNYDSb3bOyW0GoGQI6sBtAdS+/2y2QPw483om5lBI6BYxJ4Q0zzL2UcnVM5X
1Lmsi+JAkJGmolkKAT4Lb6J/eqXM3D+eYy6DOjonhcPm+nOMJxx1d5bpx9NIM7jt
sQ4wQeGrUuLmR/ECaH8cWof4bUFNYByi3pPvcSrcGtLiJQlnPchvUsCS9XPjrXrU
UJaIFdOhNsF+ByRMhwMvPUbgI3UxrkiI1N+JmiUMCoD2Yt7dCj93sIuBdRyCof4s
QUv6zC01Jj61e9s7bzcCFIz9XImeIabOJP9XexxNk0946lcBm3M8WDtW27ZdvqbU
aHBj5x/s2RpB9mbNWzni7HM6m/UcW3wA2TbWlStFXH9OjwvXMu6/eKPPzTOAtwfi
boWophj9NREnvGD5UBb7V5+6I24Bw0YF9Dfiew+HFx9X4q0CF+UgnkG6Sy0hugAl
yBgTAREhDJhJETa/dW7eqGUKL9djiJr+tXTbq+aSvREj+ymnpqab6p37Aj0dmBNV
Ld1EBfzWja2XN2HfwcXo8Tahp1ltSM5Z5DK0QWYC8zYY7bo/D0dSoiwSKVXTlUSg
7kZ+JGcPzDW7Z0HTae+ET7EJYUnnaL0imb2QUbBoc5xLQHxe/z/2SRqtfRz6WE9M
pmBVNeHT6ofCO39OQ99LTGVIfBaNol8gB0FVx2NmuECCpWgSsAyFL51iMz7Wsko1
883+c15EVZXTagt7VCoeV2BDV8riIgSpCW4Uu6MbjWaT0Ju5gJfr0f2xJK9X5wpL
tMZHZQhHTfa03xm7lbTdMR5aXC/VQROUtWTzqa8XOtR0UkeHuFJyhIXu1FRggTqL
5UFjqAqFZQMBYPlftrSvG6izDph52kUaDM6he2pOJC7CRBiGdVRhaCIxGtNEijt+
GyKw+cRo6Imc80fW/j/+tv0NBqdh7cFX0Plrm2khvrItC3sAndlZAWHpIGQnBWg3
qO8z2QDB14l4SngzM268r+BNM6i60LsE4FRgvD6nZCzLoj8RcUf9WZBdKVZM+q+7
BFrxTVB8xvxVa1SMZo09+o4eNMK2T31Bg9ieFPiKVhYJrtDhozrv7jZWj3gHtr3K
arCdgLQmikDy0N0GMdlbpZdXRIHrJchO40QP8LA9X80PIBlXalCJATJjq1BUUfxH
ELhUn6LPMZ+1BRb06vENeoywRctZ/TRkdezwl6ZaGrpVKPolQBEmqTOkZy+3EOR7
zMHmlKRDn2EMlt9BxcjhbVWnTxcwXu36oq7SoRmqcLXzn8hutJPHs8X/ANNPRp9o
9JZx6OJHATXRuhH1/2uXfdSRth65Ck2K0DDEdm1RezEhfCMXzxbjzmhMBGRQBH5N
rLNns5kaF74dWhGNDxFM0tV/wk/0vbIUH33qKfJw0d3EaDKfrx1/Gb/KPUkEatiP
rKHRJRMg4f7U0ylRPLZFmwALyK3ka9mQO1sfKqsqw8EJiEQW8Y8oHmh/zzGafi7g
w1VAyBgu240tbroHjHQEvVigYFJeDzlv3rcuppFgkpjpdgjCzphtaJaJ7OxKrGO1
QAVvks/yNdk8RC+f7IqyQu64IbhGhtMlAUWTmSRH0SxHhj7OCB+jnmWYwv4H9xrR
vctJR/LVnC9it/VyhHLRZjHWvtaMoP3nu8eFKMciCOvCfgmiA1sGiOIirnZUbvyJ
JK+xCe0mQFTPhFVNtNA/lYVwAUgrPsWfPaI8jFjekMbNnqqNSMbH7oT+8X0elNdO
q+aqiselXkL5DYlkZs7nM32/RiQqtGyXgkzkHPZRCNhbAXVWBeQyePZjZoSQz9af
/3CUG4U64q5svH1TUYyv2wYz3XxUW79/CFc6xB+/TqF3tlY9JcxHYtl97Ce8b+3F
2qc6Avrb+40/qGX8duliuQxtHzfykjSZ3bOzjthVsnrjRTFCN4AvlhP03dxjN3zC
nS/kyPUaX6Kwge82DCrqMk2iay+42BrgjUK6deZT+T4F2l0JRyDX6wej/zO86ig+
jKhk1/cKf1hrwJohsXqFOJBiwaOY1CBVOWihZs4hbUf5HdthP0Ru06vi07D7O1dS
ar+6wVzPd48U5HtTuIQxUixVLGgVwVtOq9KwszH3kHCUbUk8Y6gM0K+wRQiM1bnb
H4U3jNvBKsB1U5e8WSjmhXe0PeGV3qj2HoEmz/n1YroJ4cf74b9xDUgFDcTLr5ei
OGQ4Y1Tw6D8zJbPebDsXlLz4/Rq3MaBoPJ+nUWm+VV++lQavKXa/zJEGPwbEY5mE
VWsUQaAliV33a10jVbXlyhuyi3B3GEUtHef/Rt/utkZgB4uU6Vln3ZqIDSZCOXyt
Lzlyl1+DLrmH4ZJSwA93yKQRV7JWA1PF+ZUEmkI7LF2nnABKWTj2ZAmt0hOPCZpB
Bm8HT5FUUqXk6su0q+MjF1N6dXxzN0QtetN4+sjbMMi0rlvoO++uUWPP0SgQQUGn
nlEt4vMfHBLeUy6BLzDT6SrTbt2G1mcM/83xJsz75/vokbXOb5NR5jy1BE7Qo0nf
F3BgqYFRvDEGtEqdwGmWRZtFcRYB7vQjOtZDaSum1uzRwDxrwdsYEo8BeLpe9pCp
7xVYVBk6DDMEqVZzkyYcJkz4bzxl7kIE5i1NxJf+kTfs7EiVrISCOWWk3+h9hytH
lPY83njP/0Q7gWz7ypbsln9F8IC2axTFVS5tWrA0sblbUpOi3CD2PFlahQQZx1RF
+SmcYbcKIhX4E1P0UTxFPYQJOo7uyO7e14xbhYsXl220/t5volppovtd2r6RDWYG
c6G9ucQTqiHUmVKAcvx1fHX0JtU1ZCCPf02JFvkm4+uKKbYvwItT2NUZ5tdZHq+T
ZQd/kF9AJm8TjbHwAuuWkEUXxHxEcCWFWOer/tH1dOhLFXq2BkswI6f+A2+jUqyl
faWB6giVuAX+Pyt4ztScz77JMg5wCWTOsmJCgeFw9uGOg45v/56dQOkclg4K7G0X
acVnutKaB04f7PrTBPzl/koa/tB6VBU+gjjHKW+S9JCy4zXMbJqCWz6dX5Sf46R3
ciyCxxyIShwwjVj6ITJ9b0b2okYbTaWLpGBEOr+BMbAJBFbMCfeCvi6Si5TAiFge
pxvbNIAebiKXnZlbpUmIUuL4WseA2sNgjHfNWxhUpWPOIUoZfiQWGM5cxfyquC6i
DRM7oXg1++DFtaSVYaoJKZZLgi+DLVVGVKq85bTaRwu326TTHvWsSepFrx1J2bCm
aLUbaQWqH1O7+7gk3foaeLloIbupDz3lUX8wX4Msnjrb9Ii/IkWUO3XNiKn+ZC49
eCOM17naS2TOqtPHIaQUqP/+lWPxOfi91vY+vbb1x0urU/3DmdFEqTvlM4hfiqXs
fjNqsjynNSexkFTm0BSCTvcR3xUqb7/g+tnaabl5brpeI/6Hw7n0+hfogA3NhCs4
O4lLcJQcEy22SMSapdHk/OVyGSFtfgPYEsYS5uUk4TVArRL18hvOALeKD0sgwP7e
zf9GOTaGFTJ77yGJMOQYDKHbuCPMha9ZnzCarBBr3e0sVtt2ehVlj8hbwJDDLoZb
paA4sgHxk2xigVXD8iqxYkSUisGJ8rok9SHJEZN38+Ck6DpLnNW3Yui7aQsq6PDm
Z462NahaoQoJtI7CQHhYzUpVUu0PCRzYPYzzsjfeKEGj/6WUXQp716rVIWEKesKN
JZtjcIKfqfvIbwcFMvTZTqI8l2ETj45b+6Pgo5jtuxAGwzQ0OJtHZxyLHWKRfgq8
bYAd8/B4iuBdPIMxJX5ZxOuMgwMqlAz9ULz4kfub3fhjGyulsPfG+/0Po/hLSrOA
WxD6gK2qceTRJqlrshnlpE/2AYwmqWzUQS9GdEZH9An8Xqk2m7fmwVA8/VWUifDD
bhyBW55Ki6JkTIFy2uLG3/uyRmctsKv4xfohqz7EydSETlOH0Dg8gMcr6oCFjUBx
iqA8LhqAi4HMdfyyz7dUV0bMfaswamEpi+sDyJ5AHmlNcnb0ASr46c9+hmFv8YBc
jhjYGwquDt/46KsNmHQ79sgAK4hmXfvz93fEFzz739f7BbT9UZkPcb64kkRqQab5
PdVO0J2joOj28gnp9yEyTqm5PfVhir3KEiE1aaBFYwwwgDgMnoFS5GAO9tGNO1dA
p7Xa4gnEotivBdMe27zN3B7VJrXFlqUVuoYBHUqVn1ugn3eK1xPOeTV6rtxdhcmH
Ug1eYP4yeQcu9Vr0/GfK1vx87fuUkWrKrUPr6ctu+P+obAiasV5VwFw+RHqvd656
22g105V5lA2Gmjp7fP2VASFBOS5Ga5ATTVQH2vOPboVCUiuRRS/BBNst27nsmB3U
P2ryYR3WafIHvfsmiz+YyI9ovMYoBxsEkKZFK1hKzo79wJ//GH/2MpH0yH6Hu4wd
QzQLuLdetyD70IgOmk5OnyO2+OyoQEPDU/Vu/x7IdWom48xl0IYEScdkbhib1FPq
MSXfi4QVqz9Ce3eZKboxYWzi0zjr7lD+DjvcyjM8KHvVCKXsKoAHmkEi7y4QIS9x
xJ4ets7AIugvbJFXJXCkPzuuLSMB0D9frBkZq2mdIJRIpZoBR+dPyumTDru7zDqC
tQtGl36njCZP5xNYgcp2FQ/g6osg1UF4yIbpfij0g6GYxOuXj+L8wgOJReF1NPyW
tX8fbCsO5atmdRIbJbMQx/FQoF0tpuUO8gk5mDgyBhMkuluty1AtOv3Fu6wombFj
xeBMYvQkWjWHf+cs9zTIgLdjGaYYFNrRkHhQg3CgjEZ+do3swcPR9uI7ovUj/GQf
bQhac34m6lCj97ugfPJ+9O+xsGznbSsmlET29+0Cb//q3rTGWA+1C4IdHFLBL6if
w/UJORdteMkTECEDzxvfi4tJMra2SaA1PXEtti6V7LT6PCkCOXY9xp+6i4lZ82ZH
5PT7qzoiF/9d+47+cRCqjYigs9x1bB/2iJsAzTyg8okSj+NG5c/X4nPXIROEOhKD
tuZYn3DiU4DkYKiu/iZG3Du8FHIiFnqLpdECtVVuVBYSkCj2KPi/9p9lydy1OdPi
UOxhqU/mYruJSvjSkQUpU+eHj8nII9ZdlDEZ2sOdkUllUPwDOuN7K7+MkfK9fTpH
Y3cPmiPz7IVCSZ9WpfEBxrsVUtSi4bkf4NODL4yn+OMRNrueDeKokAPylUL0nV9y
lVWwoq229/fIrECj6McJgiQKQoHmBRaG0SzlVAkGiE8El85IdRZXxH3lSIJneS+L
PakbUkl64MaestBSDUsnzjpVv+Ag+m8yg7QjC3EUIIdjg8X7SXFsUfSttq3H8QjI
9eIbkz788RhnGvtYGdfxOA10wRlQESzYkruPKPp294gQx0yLmx/wAG0999lA7KBS
C3LDSkkNWaGq9o38xdOgh40IPC6Bpy7wBvi8aNpVuXawVQO4yLlVxTOtKF3pyhvA
GpEXaNY03N5qQoLZJi1RF/DRzazGLZknKIdQ8IfHPdeZjzdWy8m3hOnm0hOVhGDI
CuQdpwYc87B7guFyfU8M/DWQaTtCgYnOB+V9y/hW8BlXBDK3cKqzABxo785G2iMq
0OqFfisly1CxHwf0QwCm8EFUcPMIeKuTrkOXjUzPcBRoqZSpTBPnI2Bl/2Cr0jeJ
fTBBVEXzJd1rR5+aHIe6CMWouxajEj/5oCPCkXWs/qPH1r1vkHTnYqv+kVVD/6EO
0VKOoD1tZ2et0lpfrGqpfPKT8Q82kL6taQrm7GghW9hhfKbZB4gunVy8StFUPQxd
hD7PgG9xUFboTizzoBJG+t/iZMGCN/seeHa8+52O8FSgvpiXcrTwqkpu5wF9ywsx
BWMAFXuRCZtles1j7fIpMWzJ6J3k19GueCGJkJuBPTGI3X2qtRF5VCwNLotfpiaS
lmn7p4HQpM3/Cqp9HMBo8APNQRn8J9CgVkHD/UREpgBJ6qhy8MvB32LXN0P+59J6
zU+0m4anHX9Iv4h/J03/alSaQdxUr5rXac3LcaQGB86stGmirNqTqQwBAgvMY+1i
KoBPOrhvEbSHghNIX64Os5TvM0E200ljbs84cZ2LBa+vm6q5JKODAv/yIzVUqyF3
5uXPECMhfpYanmPoOl/BP7qsnlS8Dg3hD+N8XjPwFR820zYom8TvWORrrDkFkwfe
3GLIDCMcKSyZv5K9XfkyBYo6P6/l2B2IbAghl5u7JNvr95U2xxHMdWc8NStG2UMC
2XmP7Hisj/eyqSfRHGWoxWbAdHA7h7AD6kTM+2wCD+nMUp2sHTq24mi1uFsY9U/S
UEMDs5QRBJu1g08cbflx2hk39Sl+5s74vQJXVkbKEl3Ezk9NScnJc7su9wPDhXhP
02Ottc0QUrub6h9ueRnyv2JZmC60YcQwJK23zFCH+ea9kQUhz1sJcpjIJfHOIMZ1
RBTTyKdXtSFn4PoLSsWT6JAQWOqwu4JKgVnCAmMTtJLAa6tFzqTwl5E7GlyRDB75
TjyXXhVHUnXUTr4usYCCWAUupDY50fWz6zOryxmv+nZ2zOpD5uco09Ohp0tZunvg
eP/WEbY1hePdbjpKeyGUqiB3SGVyBU+rD/CYBULNDV4JjV3ArphsGKaGhSlIYfGd
FqLOb9whYhhA51ELiQlVzx74OgQkX2a/SiLzgwMCqe2im+uiDV6T02SyH/dWVGAm
bs3Pc3ENBvtwl7d1PQpSBsGioglUlm2885He2h5buGpb3wHK1tgg4oFnEeueXJhj
80u0CabhYSRw66kwcaVNcizB5Ln/nn2yELt6ewOOFUJIHEQsNSgCgaaTF0CJUiRs
V3ODFQeh/QSVXo4vpFS0uOLaYyfQjTLoqSsHtoRb2B3eO2sOpHuXnmYZaDT/wVMm
cVOkyQ9yzwx7ZR1VJwzVTXMxAxHbhB9NivQVSQs/QZhjETbRRR+E6bXioqMpaEpz
zVUKnLu3GJDvgCCV1rwoeX52x73Yq9jr/m55Z8l3hhYbV6AXNu+rpQPGYmuSzKOJ
GPymVZCPtV71s6ZuBzmvYopx0HieUgguo9qy/ATWNLXoiM0ErnoxGNH0+/hjM5q0
XLEUEPD47zjMobNEHJVt91RTmqMeFsPslgMrZyvvd0rzDH0Vlxi22aM938EJhr6L
WMtVR8XKyf1Z3WQgNmWjYP2FBPVS8ubClYl3uqJwgtL2c1cUUDAO2iy5EkoP9ONF
vw5Vs3lzKZ0wVUtIz9n3q04YyGbY+kB2fpdcCQJXMRXDSx215G6LbDHd19XXA1QM
rvQF+5nOo6vkVr0qh7mo/d806126Wg3slS2CXLbjLxRUtF/4yYCylnS6QC65Z8yM
E7ogDxende+qe2zg9WNYiDSvDIvI8rH1mRRGDfAd5kxQX0X935JkhFTJks45btH0
TiTiFr/+ig6DIq2A2/Q1xLqcZqCau1wkPGxBh/NeIX4oQMTRQXcWLycvlVz1W6S+
QBBmaAPaus1WKLrkTomn/TogT3i6j7TKyvcAaoBw1Z746dzl0MHuGsRbJkgIJmOe
xTWqA5r3EOIMfWy+lEwwsZweS/8m600Gmjy64TWnp6diUpKQTcRDFb/cRoN9t0Bk
pMKYLfBpOv3QOid0+YFELqtdwS42Ye9R3dQGOzFuKSj5LaJjLaP5fVYAVw7MBlEw
qmU5QwqSwshATzn2OzClZc9pdq9ELN4j40tAX1JEYn3gIrcATAbphAeqk23EXhpO
U0x68d5SjM9I5GZP0RPwDIYnDj8KmmgkHgCaGpJ8GIfHuXS4+hUtjSD8HHk3QUj4
juovFLh6s6FP3psq3ewk9ZdRpIe8+JJD9FU84HDrQiPk4pRXgElzAqdPrmvp+7Jk
HUcxe2BFMcDBjvEJH/T/Gdybtly3WH+5rM0wtKIT23pthyKzmSih2zebSKO8erIs
fY95JcyOXoIAdv8TwRIDBqrfh3ZzaBqYIO3a5Vl6uDOA4cg7NqnmT/cH/X97n36/
4jVSrAh16HXTb1uYE2Zj+/5pxPZPff3xBRnVZJjgUnKi8CHuvUhz80/pQo93A7Iz
V34CfzNZI6qW8zQaSmXhqVpjmsvp8TpGVEURG9uYqNoAW+QURf+xwSXPwdiY4mql
INU87TBjopLq1vQys6kmYMwJvHNec6TetdNkc8z0Gx55fk5xoIdNWNQxmAfZVkSb
nbvC1KJX0WqaMMkwkMtxGdc4o5G+NcpA4HZIeIqdIWayNFrMTfn0e6OhUAsa4I/C
It8QVmGPHjNdrmSe4I3kqiHy6I1+JPEA36PF+lMG+gSdNvN+jlD2F0FSuwgf7wm5
563lYsyxEZ3THWBnis7VWOJ7enkkCONEcP6m60i6VqmO8oG2qxGKOw3dWiYtsUTm
uqvIuX1Xuy7/WS52M3eZDfptJEv0TL8lB2OD2oVfiCxbm2TkIuec0ubGiVs7WNHy
V/J7TYP9XdkViTYkMzLcqueaXuPHWZfQahlDgTfOPeWlQXx9QiRd9RVqVKwhiKW2
eI9XSl8laUzRnrd+5fcWgm4HcwGJiAmqCQX/RS5B04q4zX9C7htUV1o2x5ir9z8S
t53aMGFcyp0Ypi9Qc06fU8J5G5XNPHQehSXt05DsE0KZy9WVyBdCd6GexMZLdEw5
UKxqNWGSHqo0WOhTc/HCLXzQ1rSeS/Cnx3DDC20X5bbmI5wMJ9ejbIqq4uWFVSom
BT+te3seNhjXfFxoWO7IBpiulq1kLyaTEs2+guphuz+/WLgJVKfDIrAIsHWX17tk
AvZ0VjJUu6F6zSo9udnZE4x9xyqu9tqt75yv3BJVNuzxracYMIbcjwOueO3BX4ZR
J68zYBQRp6pQP7PEWdTbrKvAZIBNxGRupTyspI1EPv2nZIqZMd2CD/ucvIuXE186
sg7r1NoBdYOmOYDT/9VdRsBl+AQqFXShSJKRCOdWwYSVgy6i6ubEZDDqpMnXKyMR
GgwHKr/+C4qVqJ100MO6StwiYJWvow/Cf4qsiDYqnki8BXTopdf1IptHggkG447Z
fl/0miZ+lIhr+6Wvl53+xnVrnGkNTcSXxlXovqTtYZwCc9wNgVJUjhn8AQ/djuOq
08CMa1jUxryX37z5QUYy0Td4Gco4WnkyvID2zTdyjSpnwRSpbW1tbB02IQmQOIhq
6MLx1Y+fzybKWnzEupPaWnlKt0baiobkoP7XF0D4O2eB0d6D6vIy5vjRDQ47/ZY0
O9Y8s9ClutS4To55eaNWa6u0/9UoDCM/pg/chQ+9Y+hfL7oQr1IS9DA3TsB6OCPu
eBdsodsxLPl7Rrg4E06Nu17stQcNDWqkc9L10c4+gpE7uY8Xfw47+GfVb16q9h7A
ec2ekoZWpwXbgvC0WWidt2JYpSu7M/cRwxgPb6siVr2XfMqx5D2wgERpED8Wc7t5
oi3ddKFrNnqwfBzg6J86+pPVKKc7JW/1z2YVJyLibF+HClFZRndG/opOva9oDYr2
7zc41HfEd8+pK334rdwlo+rr5fOyJ3Jo2I7kAU4kWz1b+zjsKzhNH8NEBAP7d1HU
yXo2PGheW38OgA0BHrbBg5Dw5rkSMkbSL2dhVs6421AGAtTuthZkMSuFH2LxJKln
vgD2pXC0BsYGtkNy2DFzXKePR+S/HSOyxo0Zqe36HkFo/NC6AIFEpsdh/33hJODb
mY0SxGcdZ2eoUJn+NNyAS8KJxIOVpIglCarjwURLcpTlIkKHo72kcwKVUcca8AlV
v6Xisfo/4M4FqPMqqPbFkgEbo9FK44OG3RMJftA+jFZMFoUEYculk1CszPJm2TM1
gztxyP3iHhYcfQUI6ZZ1LjijnBVWKjHmCzrQx7IjLd5SsSMqbKC+VOaxcfsybYW2
J/qe4l3uicY1BvFv1RUqyNJc1qkWzNQqcspMPoseRIR7i+OKN7aE5AaNMh/iaxLs
qMRvtUhksgExRZlbYPXGnuQWnvn+P2OT0Jg9dbDqyp0M3DDRuHTQR9inT+I+xt2S
Vyf+HpYPvcIrTGomt7mfhi1b/NTC4yerfxu35aFsx7fVP+vnPqNnWMOpbMLtlAUt
/o7N8k9at3qQR1GPoGXqJ+ddhW79dkdgjvWTbLdH0pBOLJknnKdAsfTrSmDW12Zh
LlQ5MHV2tWg2cux5Zf3td6YnrKInARX86fvR5h8hAnH+TxkLGpyTEGBmUq5jPtzL
DFNp0HpC0jvcngJTIBDTVPLnlEfRPiUMT/zXVeYCMa/nm+QoxrnOPlB759xBNrB3
y4rJqDf6CKtfegDQz3C0bIo06cM6BwMqACS+5SogjVLL0z+ZNk8E7YYKvhmFLWLW
igMeg1XEUVQ0GdIdxXxFKaTQqm/UvkLXJBaTKnG6xzyVaLwebx1+Ld5FH0nQ98XQ
JV7ax0soynT58XG5VnKYkWf6VDBrQr38KLI44HhYOhfINPQ9FY9v5h7MWqMAAOrm
Wrz5sXhGnLxd6iXVSG+tPQiaCFme+zZFCTFR+kEcvsmvTKDHtmUNdlspyL05m82b
S2Q/3w77K/a7YhDonkRA+P8dxyToZ6ohFQsT4lqVxYP2aA986vQREMd1YC+PpMGY
6gVO0I831Luo4YAmYp4nO4DXvs3F5xASx9CFp4ow7+FhiNsZOuha/T3aUUnzguvn
SdSZzLrN/Pw3zltZg6ubcy5lBB1yzBiLU1lufRCJ2vOyj7jYofX09Z5/Hm0Owyok
aohHljJGwSyHhOl5az8i7JCg1UIDVTaPBEBP945BmQpDlyBrojgKiLcfp+hRZoNW
NqKB1qalSOgT+wfh5EbBBp3kAJktLS0J/iQvTiadhMqqAYG6JMFoVb4sQrEaEQlQ
sIpAT7Qwax6bCzYfA+QGV3sOK5UpSIbdhsAwGgzgeoP0QShgE7zrApZyQSWvBq+b
9QNlfgZftaVCZG+lBodeNCvrOuaD58S+v4jklF0iBH4duZUuhe6sSXIfB5Y6cahW
QJQVM5A63pwGfYLXzpG9PzxjHp63y2snsY6fXz9Q1zf7v4HIjs/bbjOxyggBPChU
8gPTZgRSwnbRDYSsraldZgNPz0k3D6DSLLgNjxBjwcwaTC/bzq2wpBlJ3B/aDg6F
O4wrpQRhlYlAp3HoJpHheN54DXA5mVe2jPlfYh1QHRL+Jm9AxFSmLB90BQnO0ek6
6TfEYZlVP06wGS8RNbmxDgvBfZSzB6j8E5m2PaygPnd+fuM4MudOb4i3sKHVaF4R
FDGTIPo4t26SKDkYSw1kTwsXT0Id0OqKSNAd5g6s2+EnTCb/Ffv//3TaI+1+avS2
jAtolsJEDDuksP+nWSffcCFCLexn04VFCFG/yj3HY4RE9Z8VcEb1JzB1WuxKwhHl
n6oH8MCTApEiXDLBo4WiPCZU53zmoC03kIp7FeDZ37k0CQh3nUCMRdB/GNos3kDp
YLZUeVncPRcABjvAdv/G/EClbQ60CgmT5AauTtYPQ8QllGsyILgZBxxd9qy4JtIv
jUD/vaD30bS9Jqd2a3MxG7k5nq41HkJvA+lf78Z7PKUc4V0uxpxy6ZkvDdH4jvsb
DlB43gR82+Zb1yEKDzsrQdJU6FMHo8rae+pO1rR0dSP5+Ej18pYkyXZzEBq3pWLH
hP6B4Bz20pZ9gsGdEd4GJIum24p7jsOrz1k6D/fAYZa/Mvndya0tPk3r/KZwq/g6
Ie9wZRV4XfDFFJ6Owpkafx2Bqhz1Rhlex2zffwKqDU3qhiV/kZgrs6bdTeVidglj
4UIpFGZSc/gVuCpW+auEbzxoOlfyXDbNcQKAc1eNHpTHHvfXt+NaYIurfqWzWrK1
scb6rLLM1kbEtlUXxaSXw1P37/kBUM+aZ27ppY+DNsdnh1EHbbVjQg4eM/mAGOa9
cEjAZIP760b4o4rirvHt/OSH7vhEAuRvR4D8oQW68hNVwbWJN058LNx6t5kQo48D
6rM/nso42YZsH+o1DvyonFxqbP1ApwAqdOnN81kClI68jFBUaGtGa+n2jzbqpOdU
RsWK+BsbFe39BT0j6GopGEOZKSoj0fmcVXyE1LYQ6QTp8un3uPG3q5ll0Oc+16JO
rnOaBRO0d8KrMIxnq1Reyf/WXvl8wAujLrT6xnLhafiQR9xH4HyAexjyvtt5WqHs
u5x+l8lJC3ykSd9OuJaDDSZptLULnp2poS78WCr9Ttj5yCJxyByZyQcyQ6rkwgem
dTu8+26VcF7QReWt7NdsNFJMIDGppnUjHdpE094FhDdScf59LBh3vHtAlUvvzTB5
J4C1YyV4IZyUqWPpFLEzk7P22x+LI7RIZha57cDEo35f+1hZe3lRzvs/9sH4b8If
eocrse4nZB6AW7HlNkzcsU/peHik7yMP8KA6sa3cTP0cOeVNuAd8XqY9YdngVmzO
IK09DNq14XrYwtuEO90hiCxEsoVjhZ3JJ/vXFHEGmhw3ptIkw7WLUzy1AyhDNSaH
ohDWuj3lZ0s/3Nm/yV8qA8F/0JuWqFnlGAkpOV17DCoum9Km4PQhHWh+/530N4Cd
YNfzB8/l1udKqIP/2junPiXw2P/tq/TVvISFPAg7R9PQLTeTPiEsugpyfStDbR0G
Qsje4eaAf2CEakCf2yVdXAA/JeDTlGStE7xHJYv+dFsutqhQk3g9gG8cItaZGcjb
coDJzazy6lsqJDefof8hD9hARdRwOutdIBfILAQ1gCt23iNOKONOuNPbCEUFMjqu
r7VcXlAPFW2DSxW7x2G4uwEs+Uq02Wo/kqHx/Xau0y3gWviZsEYDJUAv7NcYbAvk
5tPrXcom9h7vtM1i9F5uEYhIEzzlCy5Dhl13eeZ2jiK5/9CEovMlYzh/BgWCbZjH
XnMM6+OYzIS3OW+OQ9FSGw8P9HDDkb7eBcUHtZbsAd6dBvHb8JtY0kJZcU7NxWpc
k0EdXmhvwmwAewdtExW9h8RoAQu0eelAas9PxbHqBIx7dms2wbbUQ+I043M6/Cz1
fzX/uyQvCGNyzIIBX/k1JwkHmG5/vwtqefHBC4EW8J83qX6TkTBfJw77J8pGMWMD
q8Q5cOG+nnK4C1qmUNTe4lliHKaoQ5hPiE3fi7SOPSAy9WBKMt1yJ4ulQhnOWxz/
07U3048vbyBAmCY7B45ug5a6jaHhequpy3Dwr7wolphVwZ4XT0qhwug/QKgCH9sM
V6TnBNDyM9bV7sDmmDcKHO7+AdBiqpZosewX+qFSmANKGZjq3SH5OPTBsuark4Lt
JckrHhNacp8wKcldVJaBrvgiH0KgXCu96maB4JXzqNfQf8BdlAgSDoMeH3NpmWGz
BBA+MD/EJskmnPc9yx0TtnXADVCiYklK5ngoiwSBweqJ4E8ok8EITXVDi5/4xdTK
ik79Jar4PC5xevJqG0wbk5ILYUUfoEToWb+THyBPnz+OO5ssRRnrULm85mFgodV9
0ILA9D1EPQaJZnOMEgUOSiOnFu+vNvOArL7azLPINya4Wle7/zW1wnwWAIlVXuaU
HtOUEgrEW4j6kuYvYThg0AfZmoaSCk5ewMg4gj1sJ9I4XH+qs3IHB21kt9h8d1Ql
8tsulEVnBTiJR++0tm3NXgrQcvlpmUb/MVRcqbsRfk5XeYwIfL7yCWPQIUPU3iJt
epQmlMiRoCu1aC44iNE8kUngWp7XSWaNhqA1SpGVPdQuDv4q0OCNhqhYRgn3Oq6x
C2PYwh8Ttu187EixHpO2tu9Fu3AsNw4ZgFKz6I61hm/hFU4TTBw31wAPKLWXOE6b
oDtPLJ2BkQSnCwaqJ3Af8s5bDLpMlPRyOQ32od8JOlUM53w4cXln+O+tdr8dbi+j
9dDQ3F4V+SSevHeRnrV/AtpEicrDoUEsMi+UxGp8Q84KjFlPMWTqkg3ApgqsOcSj
HQh+XStQssoZq8AoDEzO2QIerMlwqT/GOVBZM1EKeea+HiHmJKF8h7fc+fG6Z7gc
8NbNZBoHy8QGDD8c7Hc26jVFbb75byr2uFEt42EQsAP9bfNCfqTZI5wY97u2+WZh
OR6Xf2a9yUPjiUk0SZkz3S9nLPcTL0kCOH+/D6G8f2PAHGv6mMAF0v0g7T577cm9
OdRX/j4GQHeuhopAE+mrqAi31fP7WOfkjdWwiVjnnZl6GKe4A9TROBh3/EEyA/F6
sgeS3VWuyten6po5WvnD13hwujI1q77UEqnTei6E57HZqAd5aBPWU7NhDvmcvqoy
aHPDgqFwqc1m0MgG/h99gW5KJBDvHs45yhNRPgcFeBEk7VTL14wzmH2OW3ElknlV
Ag4IQ953PS1MYcE6nwTrEKVR/VSkMj4gHKMlLj7bNggliLzQJoZ/AIlQMe9m507X
ad4ICwagCBMWfHJkWS5DQ99EpmizhafJaFoNFvr8Fc6bbGm85dNWXSIUcus4w0+R
Ii1P0yAPXxXzZFM8pD11o6YwhIO9URh+rfTk5aX+hino9SWD/lTXdX2HPbh2PY5R
eJe1cmo4QRf79L9OjhbHK8ENpleH/x11yNEql6Gc4VjpFsjUKM6eAWwy6qZmA1v1
VMIeTodhqs/8pRwrSz8u4CBY8QapgKy86jXbXah0oEAQUXtT/z14xnsVu/SV+oCg
9/4/VV6qKivKE393P5INeQNb32bcLrTf2bycyJZ1jCZ1Oz+vKT8ggPLz6ZuN97Gz
1PECrZZ48ifnWE9VUHiCuwpim0YEusRM7Xtjs/Tbu1DJ2OSHwprdLydcN5tSqvAS
XBDr4ll5zLnuxQi2q5dmXi/UXnWeVl4V6fOL7W+mIraZlwwuf6FZ76R7OpWDVv/S
WjoGu7ZKFDMc81MYkkRoIK6Hv8xmwequmC7Vshc8beAbNuim6nMpUVPs2htkUrU9
LthFrUV57Offw/Aes0Bma2Nfucy83wKc7hhUql4wOafB/ylcGzqV+m+rWREp+e7G
fcl0DMudlnMZdHGf+keMLYjgrWHFVWp0YZdH1K81e57thmVvQSo7dbYG3Ut3y8+q
gtbjaHiWRE9YtQT1srLckJRLfLAYkX8clI9Qb53AqF7cno7MFVRrCMW0v9OHjf9F
RFPALkAkzlfM5nV7r56AmZUQoRhvRFxgGNRtp2WejXo5QQYKZdS1ykNHR9X2TxNA
kzG4m2DBR/FBJVd1IqW5dZm4ZcxTHFDsN9KdqxiopskHHn2kdCr/4sanE00w52iw
5buuEnVxEm/D9hGDFgt4SjM4e607e5AqONUsgujda7koufFnLbvywSheajmuxIp+
ypa+HhvPvGyuREZkOX9eZ4K9d3cuMniPIdPc3Myija5hlnYQkJLho0I6fJNzD7F6
eg32mizbmDIjRoTbEfqUPceagkLA2wD9uSZRLGwTLYQNe2hf19ZMVWlf0UCzq5es
G0GmEUeRgmLqdBPvUwSxhhtbSzmbvBTpu9OeM/kDhPn61WYjXHIE9bCaSf5G2iw7
wNYCvz71cuqkDnAgJLq4+JxHxsxurW2Iow9CRfKObSzG1QQay1QpcUGiQXDJrNZH
ZqOMv4KVugQfhEsvzOAY1lWADOZgH3bRJh5wGrWJf7HTC/nGLeF1CyTJva5Z0351
I5JNfEeI/1OgiUetIODQ1LZRxY/+FUsndwCm7uyxVu87Kz2gXX9PAR1SqYtXQ7UF
cHGY8G1JFNpbWI4Y/7jrS0/DTaObLBOtSV1W2JB0N4+IPByJczB82IrlNGRAvlnu
Ta0fSm2syqWS3WXEyXY+FmKmC8AsM/84w8vl1924RTOYCOcLu3xNmxPWgraHFwni
fxjtvjsnUUGiz6B46sXxcOLW1tlPu3Hr2SegYCpvS3qt16YZkgc7LpNmZVZ3A4bA
AhCRMuY93E0tuyfvsc/AoDOmH/IMGR40ISxduQz7jSoa+7sMlBlLFoBIfk0ACzb5
5rzDrW50rgP8ckGK50bESzwXBmwKOXIR+96nXxmg0J7JfXlsaHuIupKtoHB9IYnY
rCD9SuZRmMfOZwYuAvWmygBImI6eADug71ZETzeUKjqp51RIvXNpEkmKeLt76CYa
QrItcdvIztpt8MGPlCDjCl7ba/fHoduhhor830H9Otz8EsHsxql1PjyTnyyObjTj
+B1zOsl5UNCDXo+ZL3EnZXWAdGWlIek2+2soQp6g6DJfnyWW8bOtOZQlPNRDTm4+
xmRAxLdzypyKl+fiu8+tW5zmpNf6g5zNP3tZsfx+K8eOB9m8pWZrfAC9zkpzOzYV
24AqSDkHbw9tPyhZBs0CwjPTahWbBAcLXPSZtf25PKaB9Co4ovBoamZM6arMVCAA
8lFTM3OlxKTQ3IxHl+9HrTlfOcd+ApRgjVYvK48fehhAVfj9my0ISVV8dWu3zVpc
WsCZbQ0w6OmXQU7+GWi+RtIS5g7skkdetIBo7grwPL+JtZZ6xENkgnkjz3QGIqwZ
T+G1BeuXo8vLljYaSiEB7/wL14qJvrRo3D4Fm/8kU+fVg50Dk2NhVAV9JpJwCubK
t4a+oIm8VpV9BPwxqMMqrp1WP9rqAaHJcRUut+oQjpxQcdMJNV/gpvRbcFwY5a/k
WOqoIDIu/njVi+zTjgBfZXKhEvRSdcsQmGP+Cye8pGmtBB5pkPQ1TnBolvf2h1gJ
LzgWriuDdda0WZ4AYai0AxBAUu5DspBeg+kR/nks7IQpiyAN6vmmTLrBdynOEIYF
JyHRfPPzpi8/UDK4lR53MBC334xfomsBWTDTH1owIlgYmN4Pgf4Y8FGKXixk2sln
D6E0/gkf7PmUY4j/Fm1wKcPAUaGphlLfOko2jdu3bYXPqC3K8KAhkErKdzmGc6LE
k8ts4SCkD/WgBj5xlznW91DOxO8MsFLHv8T8vTxdgONYdy3gucjt6+vOiIQCcY2o
ERVl07vwmZKIG2bGRjDDPEaaDjvQRjsELNbynZtJrx7F7F4eZCDHU0ir+KuGeo72
rS0r0uYE6yHhPunvZ+kDhWGqqfKc1xbIbO9pGhAbpG5UR2nrecTdOg1GFzWtJy6P
RrkMBrK2M4aZ5H2FyAuEuvA9SdQ29uBdrkfvSTBHxSd6MB3EItiY3J67rY7ILVBJ
Xa9/9EawPb6XQh426/+DdZXjcVkzmkRKDopmEzPAA7E4cLlsGVSFmfAMw+E2i+Ky
9Noo/1uTtNbk9TXBGfp5VxiwbfWDr3VdT1q/pg6C/Z991dyeo8htvRbeHvh6GGyA
neSOVCrotAzbcHdVPDkpNqGM246/cMiMii/V1mAr4dOx9OxNufgxPeJnsjkMq1uh
Nngag1JeIBDFFyGFG5l8fc8PSQT/z7GLO6kHRcIg88mByNN2RgKGIlwfsF+AMYEi
Eml3brv3OXtLBGyQ7/OHhOalXyQ4aDybuITtGksC2BqE4MwHuwfDN747mHXdh8lp
BGppcFydASFeeV+TxQcN4+9swb6eRRspZlNVxzZZvulh9bRxXUu8eRA5YtkCBvUF
a/zvBpvkw/9dj+fCa4ZCm8BbkrfY96iUxZOJqCDfuz6u9j8lh05TpQWpTiFxuQW/
hs5+Q2dXNmB7X8anOMckkYiUFRPHLe42jxZR63oClLZTDcXvgIzhTsC7sGzYmc/3
LyLvzkvDaS2x1TylIUctUqmwlfSPEmF72TOAvGI40TeoIgVlOylloAEqo8ltFGLU
By6ta5NtMAmYU1A+5skwWr+sdN8lDtOmVzrZlSdRpPQ8gn3K7df4QHSzHqQxoqQR
ajla4cWRIosg/Ft7MaSn8UXtUn6rZS/guKtPWFrnTs+qxmM3dCTP6NIbWsXERPP8
16niJkChNlH3UgAm88JF/9k/ud1jG/llSVDW3n2wAv+mXYCR3EhXG/qd0w6axput
MpudVykxw8yRb/CKekcY+m+Se+hCpxE4ewOm03Q/WgpN/9AO+QijvUT5ERhNXKtv
lcaQIOW1qjYQq8yJDfP6lG0lypvm5KoNF1YnvZ7QL79SFZyrVgrA9NOc5chuSY0/
mK0pr8y+LnDZruHEV4qY0yltrvSQvnfUDPmPAhf0zOdIAkvAmSnf3VKczkMqNf//
02rXTmuHXnFgDP6XdOwoBKSn5bEc2/Jusced08+JKtyzyH/bXAG6Vqx3o4RIaG2Y
GL8uMarAwTdCBrLd29r/lzJZGp4m3xzYQm/v7YKqZWG/dWGITgDbyQ4qFMIO7NDh
QTRSDuGPVeyU165PuRhFVc/oGdOXcLK10FKNoAQsyZFVeD61z2pWX4p7kC6xCKGA
Y530vDUNyjz0BCq3MqjY9B0Qq4Tfys8IOHzOX9+FHdJdIlUNwoDfP8plY1SyPt15
q9RHkonDt7CIvjwETmB5Xnw7ZxH9WlpU/t3ihbNL2tOfY6vgODNVf6IUlxX6gYr7
n03/IgRrmI8XPH17n+z4j9YfXmqkWL7D8KO8mMFKQYsBDDPqz9UK4ZNcWlyv9Z4X
0eMPm15G/PSPW1CwMIcFZNIWjtrjOiMR+DOcuin3rV0TIXWCez4w2ons1BtrQBhi
WtFxsyKC/7Uww0meYcgfZMoPFQxlas/r6xXAdEw8r/4c/f1xaM4qeH1Ns51BYNfJ
6eCHt6xgvsF3Ui7b5BvbdP23cWRhCxsfZ7UDGID7qRqVLbzv01B5aAu3VYWIqJcw
fVvphijc14pcu3LWUeE5Gfuu9decDTPNN+wPiVbULkaGzr8AYuNVVVnqlOfMQ8xm
sV+UM238OxovP/fnIhNDV+DW8bhAKjtQS/vCGub3a6HLs3betStVqWSGEsoS7C5r
nSIwt8GeX1Nr9W8wnsPX5eEu2vO8/Qsud+nA+zjcHKEajfmwUgmMTwS/t9d2HFAZ
URxDVzhYWzDpJVNuihcSxqw4TR8XaDxokrJXpcG11ZzgBGaPBworWm8pJpsy9pgo
QCWbnxRQMVQPOxY6tJnrqX/h7lzP19d/lfdPosTKzuaMVeAjssUXY1l2hxnK1n5H
E7YBJ4Yp8lOXrG0swNzNt4msGK5LkHIw8eEb2pNrp/LDq3RxDtid/sggkTxKwicF
dVOv3pPVErQl7guWn/s7CYP+H9/BfTiS4VSJkpF9LMaGyU2VN5kj6ja7urLSfYxe
aUw43jF0LATikbWCjd80hkY11aUfcSsKUs01nU+tRBl5JvqZz5XLsMWtMPjaoWGS
/ozHPfcaU49rt4OzcalJQ/XW2YlPUwZk32PO/CIb8LjMIqgHe7eaENrLG+sMsaUw
uFHg+2fjbKOCWmR8za2ZYJntnMnGbT3kKczumK91YWOpI6AoJfInbS9KGFXOp4lY
E3QsWz2Kmuohh/qgN3FewlRIQ5SNmLh0LHbyxMvJ0Glhu1WOL+99JQYnwiMcJr+i
TShYqQr6K3iE7O9IIqfQe+ipuMHcCQvDcJzr/wyKq3//3UfhviiAHqM6dXdV2XPH
TRnXjfSKcUK1dpQeMn0iJ1KodNlBaUMzmT7R7+69FHQ6+rXEZP8Z2cXxBanaF/YQ
PcL0EjfudjPiolc4cDvftgg3NZz8O+7SA3uxt3ckLnsT5q2gLDd1u0qW1PH6idIB
IP8C54AnNk5FmrSeQYf5/Flp1zF248mJdA4EuMKMOlgXgw2/Kl0GpsQQsuq8hbWQ
DCxLxkMmU48LHfHWHwGDI0SSDK3FfYIZOVgUNUvnXuj4Dr+mo5lkPvZ5smsxrHln
xV0ccSg06a4r+NAn5oM1qxSxnlZmSqOGlPj9qdwdICLHWQrRs/Gl4KpjHBu6pWw7
a0rNCuclO0Lfcpsi5eU1l+qeoZUFf3f2uLm+oFffgEzhxvqeeDNMzXyV04RU42BR
AHR03WlYRpWOi+rtwh0VjcVceBtencAKUzyc9nnXiKzvt8E3CCAadXR7IP4kWwQ8
i+OKML8It4n4MnciZ1MVeEr72Sd+YC+zbVA38ID8NDglZqalK8EOZBI3RKt5mPv7
W8ktGcsZtSg8PC+26YZBTLxNfZM20A41YUrBakEHY+SbXMKxCGMzxvsPEeBGEJ32
FuKS4ffu+oFYEQCNKmH/rVjoEzgTRBLR+dAPD6QPuDSkZRwDzP2i0xokaiV7339H
b4BPxPCeegUAuwmNH4/AEtSZHsbPPKvbY+2Oje6M3BnCTnszI2Dv1bYshEYaePfX
4oDypyqe5Ne2DgHdUuhqrnc7PwFMi6Wf1Bnjxz7h8Yp7JWvexiKTBaaRxb6HZxTO
/4pNvCx2J3nvN+WFfW31Fltz5MOQEvQqm+vm55aPZhO/23xVanM5nLSefUPvze3m
I4O9MUT2qwV4l8qZP4HHRf9UXUkRU40/DS/Ndhlqa22qVOpv3MsSBkUGCPZ9Z1j0
1VQHv0I6MuyviX/ShH009yN5Vyy40/ryNcZ3kR5fw4J0Q0A605ciCIbU2MYTlrUx
xUKANIOX8uAcAW7X2nq8fxDaUDH3epkEXmj2BC8vdL0usxYwbbYkoRfYo6qEQJyD
DqvNDX5P6cYr6RJX7EtqwtIjdbmhzy8rtJw7etMQ/Lb729YlFDHFj3goLD84mCjc
67L96vg5DvY0MLz0lPD/+aLHXJ+dAuinzwtpwKzJHx3igxxlw1hsGPs+AYfFbMGG
bxZ7zCfDLtHYQRX1RDy+DJZscgvYYoqms74u3P/ZlOhyvopffTMY/WxtBjaFbv80
2puaeqvYOv+2wZPRsjAP1ljFdFxTgcKeD9bMqDmACN/p59v1tsplPQPQcKgDk2up
+XxbNZfLeo608Dkw66nPpXq8i/lUvMqnNY0+UXiz9pmBC+r8QD+3t9tcDzejylG8
0Zp9294kkL2UPcJUH/sF2rWMKUVvEPwzdfuh1w1F1xPGram9O0gykFF9aXxyLf16
CJXQa3LCfpeb5FMncNTcHpeVXcCL8dH9nhJYe+LNWgrJBHzP4SdCauxx9SQ/vlo+
gkskd8u/R3sgHaUp+dmTc3e/cXs258/XvmeRiVwyQXh0558+vzdGZE5d9u0h/1li
M094M1tIqSpXYlt/G5+Hc+vofgPAiWN8WVXYQyzA3trs2GY+7HkL6mQwQZ9f9kZT
dkw7V31zoZOwyfY/0Pdplje+vG33dTGbWa96+8+oEb3xTdRxd5e7Lx4/SMb0tZNV
NpsotSdPbZJLFxDd+Cqeu2U9iNPqJVnprzOC7jIT+Giwp6yTI37Q8Y/asJJq2KHo
VeHb+sX7xfyfosyVelIJIEuTE+pvFIeNCkwFf2sx4OGhlg8Ql0blmv72jX/yUZkD
yc+QgVi1i8ID12CGMbLDBY4J5vimP4IBYRge+1Elqv0YR1BwMuL9xW28C+3ClDaz
iC22AgiCrSuDSmxbadbwAkQdtZLrRpafV8slEtNcxdqV3mIvGNVbbkY7COYydBmJ
wZfVbvCHyCEst6oRtjJCATsPdqdYMJM0+NVRrQTZQ+wvYk9XWOd7EIaXbhIaG0DS
0ImgzfeGIp4gHqPJXb+UevN/14Z5DLyUImNzYDfMu2t32CLVMfh5FMOYol0b99m7
V4rCp8zc/u3OroevdnztVdzj3Etc2PC7L7xilwQC9TDOizLjqZCHqZsa2OwFoYuz
tp84WDeeOSv4u0uceL1hNJkFajJvvK+6hDL2M2OjrP6UinV6NLmvvvTnbo2HaABL
I/0Qq6VG7XhlQyXI0NiLMnGsb+2E4o2oPRB8iZpfU0GCx7mTYj2pfMZ6CW8W9Bji
TumXpokOvzsDX5EJh7gJuW2L7tdPhRjogTx1G/dbnYJH5pMloac+7HlBTuYbymPS
KEvgNxjPz1YUO5+tE2/KRZ4FdmWNdZ/j06cnN2ynU26igkfGB5IO5wdd54sSi0ch
JBBjT/tmuu4MYBCxLcbepXYAg0XdmZ1OwZU/7wEI0pSz/QTDIj36WBPr69jTw4Oj
55SU+DguTXZ7zO6qiLqDYPE1ex0mIcE7W5TGx9CN4CE7SZA5TXhuP8/Bk0IS2y4t
PVRVGiHTUQTLJjh9bvXQjOMOzVXkjRhw98k93XjzHUJogD34/kRvX6xlJtyeb2QE
6KLw91YzOBPkVqkJh7zj2xqtuCZowGWKYdZeUGXSvAT3QUcLKh+lJ9wT0K/4ovwo
0nZvJ2ks6VaKuYj3pjUriTmK4dDUkd8dfs1mb14P83N4wa+uS9CdxTm4JZefHr4a
QzHDOKWlnu00DSsCKkahRHWNa1hhvSkFJtZDg2qC4LAEJif8h3bjqkHItypUnYrQ
Q5oi112jxmYaVWfZ82O1bhRYfNQUBOepDg8xAOjnEDeRZhx7YSDIpUwGl8qPyFQS
pdW3TjGlokWeJ8vTX7Hp8lKiKy9fyg/8V0sr0wZei4w3v8ZIq6yL1TcR/JGno2MF
qxosOzKRgbL//jjztgmylMQMYN7u6lEu7XG05v4J/aYlLCvvS0zoW8NI4wdBFQ4l
zZIaikZoU/rvSjgyzRZVu4cj+ErPHGc09wJ8HBirhZD2m1IwsrWy8FtTuZHB+C52
ui7xfDsjTM7UUBsaOZiv0jeSI5taYud/iiF0s0e1WmHRFg4iUGdumJwQH4uKWv1H
QWwvmq5TT1rG/QLJpttvy7NGpHSSjslzeacCgIr0EwlHateLwXV3MmKMk6UybrDU
fm56Ow2QDJEZ6dSmZAW+RI1i0h2U3yDyB3tKMm5i8GYS9qKxEodNY58V1OEld1AV
5eQJfm/bexr/BuBB1nj2PWx8nyoLgH65sfepExJmIcgTiGfrA/xDnefPyl+QbpQ3
A2ZO0E77ROkoHPML0G8XPqQccNeJhFjw5Sz4jFgsCtLwZILPiF/YchesCrvKP44q
ENafOytX50a2J2/xCJN96xtTHZjC63T7RybJ+3fozyTIsinpu9MmEO0HThTq/yc3
A7V6LDDtmGJt2fNJZvfFzlEfH+SCzmK8OIezP00jaDfpumL0+rCo6mXg/qcRnQn6
By0xUWVVTohk+Yb0kF6B7iJqhmUrKGjQtGGQhmrUik7g7c94BVs6v9DrP8gRKRJn
hdg4fICeip0DqjSwjNtHUJMMGYC35RbrhPKBsE5Agn/2Ab4/qkb84m8VFDDIpv/V
Esa7BYzjiImtZcPJLPJ1h/4ypxyJ2X/SC0r0LPLFfmB8mrCpkbDNZWBd7vNQWIN4
SDJLwMvfe+ld5H4YNXFKeMKLm25n6jZ/9Xcf5RCZCVKV5nbBY/3CnUOWiKKupBMG
Hz/uqdycNkHiAMlQ8I3YFGwU7scnySa2tceVswXrMsQ2ZT4In840EAgcr+u58Bh5
RM0yYrDykrAwfqPgTOALeRU4TXPCPdr0QvUndMFDl7SApwoeWs7j0m/uDXiSvFUN
SKJUfbtnk5jefYwVu8/Lc4kFzQwvYoBFr+0K5+gkTLdjPhU3i8eEMzVBE52WmCmH
pb/nwivdbG2G9S331Igh3qYJOx5huRtwk60KonMWquojbKg298qRWpryJWUDFy0a
uaonLjZYra4dRHkpZ/DeC0vSyJEFlD42bbDUH1F90Tu7S4yXo+N+O4aQduoZFcRn
qVrOmYc6YSsD7UL6qBcktDAz54gv8RC9S541fVwW2KyhHqIPiX/wxqwwzFagmUnC
SXCbPhUULvYYxQaKEpqjQA6U5AdUljH56LrnJ7tP+m0+nIdUlCGurUbadFDJS04J
UcIxNhG3jroaK3TftgUejiEkfHqSo1Zhk6xlVKCVK+QE5sYA1/S0bNmsUx/7xA24
KgLUasKL0EO05+1H6Dkhc9bgHNAeGgGVEgjgDaKwtLriVAz8xTcGYq+m9Ntiekh5
k4RW5V+QstDMxkOR04RZ9EG+Tv134BqqDYfw3H1faVSa8BHlDxlbafPLYc5BA7/6
ciHHOE98ypZAhd+BH1D/yuWBfA4OfjO5JWoOsrBGxbw+3/vambXqIo+8NOFSJril
RYCDOjpp4nKuPAIl5McO9nA7BtDfJ/+00JcG1JcOgIdNVaIlSGgTbr12pL3xLX+o
bxq9+KqGLRe71cpxqSTCao16SpcBv0LzL/4Spc4BXJo5gI5bWsubGVE07yOClCCk
cuFJsq0A3U2zlwX9hAjIf3AH5K7dW2PgxHoKUCXIhLulLX1I6qXaoEtbQTHsESyE
PnSwR9hlTTNyptYE9sTo3zMGSPDVoR94FSajO+K6LVK1d+dHf23vL37fBO1DDSZd
fy1lk9A/hFT9Aa5ZmYmb/QNnOTrSdv2Rtvk7MnYLxMwrx96VRXFm5Xwt4bMa3fJF
bZe3Yf+RdWwpE5VC0LFZMJJGk2TqtRjVa/4ZWpe4bNYlwuaPWs3LKQ8cnsQHuqsG
U6UFM3Aw2ge+UNF7Jd+z48ccIGDAuOjeGM4ttvuKTeq0E7grh7LNeJU1B/pZaM8u
v0SA7sueWHLt1tcUSOdVftrdmbSdvpdBIaMsPnGSP4LmNscQk9FaelRpF8+1ApEw
/I+rbiAP0yniDXTUwiS0N+XK8IKL13tw4XPM9wOSXFkHYQVVj8wssGJKI/6gTrkS
vfJUoEnWVKwyNY+GCzxMAZvRbdn7nYRLojgBoE7MHx3IhUNd7XOuS7qBox1pPYlO
uTmQvYYrlSNg7VRcMDuZDQz7pNks8/T6PLBxdPhKb+zP6tvK3WxtDu+vILaaFbKR
7g0ikiummEH0RVscQZJ2JR7mMJro8dXhNakcQBzhqDywKKg3HXf6i3e2CuxT0VXR
XTBS8xRF8lAOy554pTyQhgP33nwXB1gqrvPt3T8FqzcxGM2cbqc5dUPBA7PdbKtb
hdt/+OKIzbQSmh7Q62a0fZPoKGmwekWkWS5J+3zyOn8bJ3mkZvZGtAL7lmSTeyLP
af5LaNhjqz4TP2MZhdw3JH5t7tZ8AeuyOaliPjEMvNVgtKRe/W5ODomCnxkGAev4
fU4X5adbx6j51g9tRvpkYCpBEuZAk7nv2Rc3b14YSjOytxEFQl1R6zuFhqW6YxwK
ziI6e7PkTbYC7ZV/xqd/W7F1Ss2KLSDNXjPVJ1mbCpyQBdBWoQNtmkvDdgl7Gm+C
LJxX5dN+QowLz30AAp6cxEahHGcZ9moixgnd4yvmG0AZOS1sEue0E6+zW9dK8z+7
QHDvjRoMD38OfiTLeoHje/bhru0M+cSb5PWwaa16K+1jvVJ4OCGqULSIdH37pOO0
KYdMfn+V4jtJ7aCSSQ/ZVllBqucaR3LCKFd46KtI+5Q+nEgx7/JJR5Cbb5+IBSrO
X0xc3b+oGthiEH67gD9pzrOj1TAkus/CPRUAN8Ij7GjxhRYyacZtVI5IJYv/dT++
i+KhaEODxekRkZLfxE43jBFOGzax8mSZzBTBfvAPJvvwsNw6fmOs+lci6GDTABgs
SLHjffXpJ99EO03jdbGxbDjLWPK5KNYHL1ZGtefjiu92oPW5Trz4Aba4FjPgQ6Jp
A0yLAfjgI8Q29xR5JE+nso9eFKHaBBaiW3ytvFKbFS1RjtrWG50H1uHdgJ6KUtIs
9ADZwKiuizMTsPOTdpcLRA6WrSe8D8aD1trBZtdwfvPMLePsjkA1kYxSEE2zI2OW
TjBFYfRDZktIMkcdugcGRhdpbD7/IwAN+I4K24/ivWjfRHKcDjOYBq5L+tz2gKXu
owBqmbXdpOBDtvwRrYyShnuEsaW5wSr0JKUh5m5YMl4SDCWaXAcB2duwGZIM5qe2
4VD4UTlffvQ5xmJA8MEy+8er2RWstJWdfd3pS+yLqTu7Sb9Kjf5tz02aOy8cjC+2
bDAqjdLlOPQghXv1hGMWrZ3J27pjC770MtUDHvAWDuzqomm53mshGJF76oAT2fHh
WHvLrFJty9T4UE7SGQhMgb3aaCztf/p6PubnF3xhj0NN1xrfE0g3JSyiT5s+uOJb
H8Q6N/O9s/bFfYlQrVgPWvPfHywqmkX9ZYZNRBsqMM3yhL6cj9eNkq/W905q+Sz1
6FWo8p1PnEZaLslZRv1XD0z9DJ/PfUvj6HpqOUYppYbPrwZCabfrnFqpgWxRgA6L
kLi8myZ0g/wpy0/xcyXjLxJLATwmt5qvg4YQTvDu9uZcsl8BwKg7oI2PL5wqw2HM
4ZEgW5jpFuZxC9y3Jkvj8SFBWy4cbd8vLl4VyCaUZD217sqeI6HTHKkp3p6Nu25P
eEZjKx+7Y1otFjhaqFrKR2Yv/E9xVR6QB1PwdOrDfLg8TbwVXCYKdNTeuODgt8DT
1Qi6RdUTeqn4oRqEGt0r9raZCcqzbr4A/v91hvutBNSuYMD7BSSglTb8Ar48a8Ou
Ex3SeBcZwD5VoVED9uKydZh8EXieL5P+jXBH4f5gJLNnpTfJbtFlcmFv4XHi8LQ3
EBr5Nx0kEPlGUCHbE+W8dD5RMEP+mHcXcNA93HsuCPc7465b97UaEh4e71lwlwEV
lZ1+YTfCH5Tm4M3uRAcOcntkJPpj1MwvY4zn6kMhOpl9XjKwwvKQ4UXy48SL4eu2
wEfD40sTiCllBmTJRkL7pu3P9mwitjybfzNYvEBNdV5q8jEBLmqNeZJNq0+LnCXK
Irnw5HFyO6aLPy04fNOeSJySnW17Kru+Ikl0bzEoR2OMXAHicUTZeax1gQbj8qGN
Kh5VnAlSv15dBlI+5sXT60l4Jf7MYRJeWs3P4MSSDnl/P2AqWCfCdq0Ft9m/PD79
GUvu/iWfDoV2VksbQ5cjUF+GVyenmPQBaNP6j4aYd/ZCGspkjYKa7vEjDt9v55lC
/JXMVM2e/5FCiI0R6z2v1UHaeFKA6BZJrm1zSNJYU2ozfGjV9cnvY2lJj9npGYyz
tD/RS33N40um+3C95MZMFIP6ehBSZQUuLIkNW8MAn2jM84geNZXIXWkqNWD5dXCV
359bmHXXvVg74ajKsvGDhC/Z570uFyDd4KioZ1BPoKzgEdi3z2KusygG21J0NgMe
y9Gpy+T04g+oj6FT+EIKHX9uLz5zxrjSmV5Q0LnGwfJG4LS16s4JkzBorOa9uim5
/QEm5wr2E9HTwjRJvQv8tCsS3X2KQUPPiA9obOQAMOJ2u7ebF85d7GTBB71W44Lj
BJGbO9AK1+TFU7fEbtPGE9h1KL0NxttqlzAv0IYgCM5rIbO1AhhbKMq/pLW1HIQw
O40Ue19SLLHk1zzj1X2Xg1JRbol5CqXH50ygtnggcvN6d+aY2x1ZQPmFzjhXmBHK
oo7plKkt1E2kdvfHayV4AwJLidQbXB9aAemNEVO6lNAoxlRgcu952wY/+fg0Ota4
Opxvv0uyEtswYnRpS4xym+ov1R5hvejQ/eNcCGgiJOfZp6XFsEjByyOW2WMSvJBt
8/wEJqgLTUnG1+k9BbfjovwI9MasABWh7TLFIFF1+zbdpKalmCBkYs3Xsd+zS/3t
XgsnGzu1NeYZT9vQGWBseYnTYlQCZxFWfaVv5Ct9AuVpO9JldhsscbmlQsfrMYNp
9le6APgprpqpRM3Qyp6VHW3zV5vNDoE9VLzW2SHZ63Zr5jf7cnnMe4O2KNO/uVjc
09J7nP0KLhHwGlpUBSSa0hpUyRGKsFVrtT9pK3857mB+VjwHoOtYIEkMNA2nmewc
gMpLrqSsXhPEOlshPQOHkHicqvitzWKuexdaFc4+sGSDD/dNaCpAgHtD3Od+aoZ2
O0NZenUMpYLxxK+0Ity2T02uSTF9DxB+uOiHQ5QrVRvCWmbOooUYrsEe3byxhM1E
4rKm3TweKFLeIYUPmw6ezz2OcHsoZKrgQm7sqz+02NMT+riYNGvwzyfuz2DE6w9U
Q5enC/kyYkxKCxcuZmWzIAyguQ19OxXFZx8Fwz7XXT+F3J7/0KS2c9OYgRPKPJFP
0pZa3YzQ6wpCE1seSHD3CI8+jCDVVLL6284dALUgAM86/6gcDkriAPwfr7h+Fe/t
fO5osOU5a3FHs50Q11vOKRujc0boHsqK6yWx8toqs0Dl0jrBpmsQmzuT7qpzXzQS
tQ8ZdBK0FOYW5OYFLKn7SF2lKFaIKg8WDBDngQtq984uN8jz2KKB8d2uzwU1r0T9
wsIUL9W2m9hEg/xRTjOK8o0R4z6Rwf4naJBAb0up1UpvU+Kj1ok6Sh0pycfb838V
0kRbQ4oiPAJ5y7YadDN4UL407c19LRUpp20x4QgQ2+nlT0MqAe8kqelvlE0YMLHc
j378xqNTIvdZA5YW1jRk3SqJfYyURDOnc31fdyP7Oa4PYfmMGq9w3+xkVDDG6699
1CjtT+whKnFvF6R8S20vh7/SZNEhJB5Q2CsezWva7dwuMzdmOX1Z/lT+w65/pl8x
chOp7w8C/S9iN5Z/potz7T4oaIBqHNEjoPTUO1K2997JohdWG2nzeudtsPadCI/w
4ovwilI9q+dsvb3WbJyd7Zfb6bqXCI6tq5J7kb71yrmn3TBSDPJyZezidCa71tQj
jniSyekvchX6ULYPxyipIAyttylB2Ddnw+VVSvLSRiBugxrl4P3W+brXt5yMNDuG
stKXG/g7xL3VArCiWwUALnj5SyXOHuYXiP3Tviw5FeqEEPb/rwFByYNg2JkA4r+0
5Yu7WD8nKtnHB0DcasIj6NPb/0dJOX/q8OkkecRSVDEDlWKR8semb1NiuiNDpStd
6pyZIcKNLJvxZyKHnVXPHSxZkhTxspGClrJxYzM028s+532bAB3IqAG4AAAJzvPH
wqkuNCegfbPwk1pC0GpBjh3ibes9gSbBrpB8/TNwEhCHhKcJlA+UEAhqVGu2X14Z
WVIrcOsvzy54GXiWvzQpIAxKSpxF9Sz6ZbAWyviLCQqGTcgkoecNUONjbQ1kvi5o
8YbU27gHjEXwxVKl0AKo3voNPoG6aLLP0Hk33u4NdlIK6FUaJXyROOcf0rmQTiJ2
FD69mc39rjeyUgA77gb8Chgt4Iqa7d/+5SwisNB9hqxZ5n/32HO8mcJdF8leQnIx
A05netlVSPntP2LvPMZsW52Mez6Xhx7PGMVUx0PPt+hTe/UVL6fTnvz6qUnEerKf
COEm+Rl9NqVeAJ0DshI3mmGSYb43Yf+c4re1FZEsq5WbFPLctFbKDVrY0LGnwFmN
OSESF6dKM+QnEI1nwtxZ+6wau4My1HoIhROXptF5tE/4whJ7hKNVhCYSSl6E3n3m
EjIAv9YCj0T3Jt8373mPn7ba9nD1t4qKZhqNjyPdEvxFaDLZlluTziQkWtM2UUoO
/tBljRkRrM59tukSUP4+fXDu5z/T7KtL4cSKmMMTvAR/O92PtlOPtYyKXDJ5OYyJ
1sHLbwILcCXVI27TCezHsN8kwur2fQOqKPzamm88OVJY7eb4HMdX6hEock4vRAdp
oZ5OdVYRIjfPFt3BsD3csJwoRy8vqnG/JyC6WdfuFlN9CTKJVc+timHEILAVWMHh
Jk30px3iJ2zYz0XCs3fYaBdJFYr5h9frbC0mvCw2mDQ0NYyDXXKi74y+pCGH7ajr
0BYjxMpyjR1YzcHVXAD/FjlHjXxkY09FXLYo7a6D6TIRunJYLPqWs+uQ1q8OEsL8
31N3nbv+mbvya6FVimfX5c0WVB1/JgECVXKDdvRET9x4XrJbVMWcmyyS0EWarqAw
ruWFjfm5BjU1Y1H64m+ZjR7E6Hi6lah/x/eOPLXX4sncVoJBiAN6lE0q82ImLXIw
W4ggL8cZNlnniVi2RhrrUNKrVM5bP2+3VASHGnIeyq5HLMQ2O01Xksxaivskwg2Q
x//7XyqWn32ERQS6ODpZ4mG3VQHEBMTqtn69WVIavUPkJAN2Oh8t61UQVp7KZR2F
+bBHVaEolYXa/sR9NLwx/SrOy4rnWWVMpLdAZHD+pm5QkXizvmPjIejXPoJ/w8Kd
qW5lEoZyt17kvau8ZAQrrafTjW6qIRq7V48lTxuyK0OoqTaTXFUlNgtMApJoFAnF
gbMDKsHcoxPysWOzgyFckVtQEK9Ojgf94ElKxTMvM6ln9rmUqPCQWHE6Vmox94tz
wVQn4dKBjDNMoVsRER7Hl6TOCJU8gTeKtQv08GepdYi9tVLeyzKEldGJutx8P9OL
Tn99fOZszUfUeUaLRIAFDs4Vnw2a7iVzJcHIxQuVPwbGql85FG0nJNuVIWeuEK+F
wLJE0fdH4QTRSP/H60uVaA1RN4S1bbJ6pac2Votr173k94qQaZsg0onA3HcTgFo3
Prk9lVOE43yYpVGcyR3jif9/xdiZLAOVG/q6W5yZi7mBGyPRi8NYybrlfQFDtamG
hYzVcxtnigDRJ/TYorx38UU4ZZXoycflEEdOSkB84j7Mc33hYB+pTqpG2R/KmIdh
8DNPfPkMxdxwdYYTqHhrawhqHC+Cr3tnds1kz4ldPWBPMsc3vl0K++gVdjywwzaX
JZlyhSLnJ+0aYf7s3CzNFLBtJjFxdEr5FEznVyKCvHkSLD1Y7foHznU1s56N/h4w
dAlLw2gYnP+jsvK+Fwc3PxZKJMtxDxT8wXIzu2ZzrTO6Fu1P/Y2FFIltr4wroDGB
wEcf6diSajKKyS89R0ql2umJS2+honu6C6AtWfsZLsEVagizXe8zwDgFzYikTzAw
sBrQpMKeeSwzbB9/nIY+d5Tm6KN6zYsHvxsm3Ymm86H10hIXE6fxY/xdvfSBPCHP
NWG3P/GA7Q61nGVW+9OUhK9AhLKWB8OwRL70k+Znpmd6hA0ta2PocYXf/c0hv+XM
kM7C3bWpMPROmTeJjFiRj4iPzv/W2YCEOnqzdtfNCm3W0NAN7BXpR3vusa+Pp003
iiTnJDyLFOXAAcgpBWctDXMBjmyrn6Mhtpy1rLm4wr7Hq6wulbUoGVBCyp389wX1
pvFb7RvesnflhJ5PLkfrv6KM7qUU1mkJtd9zHZ/lMrqiumQJc+0c0uOegaVuSV4X
KSq7n4Js4TZ60QOPUow557YQh29Z5mntA8OtKXeHCTqiJVNWPhFepPPIDUgiN+sr
jcBARhY1rv8tf28/GYjVKeR4ZeCfwrelgMz1sLpeI8w14xu/SM7CDlS+s5tc8UyV
iAznKgOJG39YGQJ/qCIS2wbV+8Bbr/+CURLShAz6zoeSGWmcHOW7dkXmy3YdxQIL
JoUr0dmRVUxB+AtZ8olfjD2zyokpvYtGbIIS1ke8uhftF4y+4lTu0ssn90JTJXTF
8vh6ltl+vNXK0ir9SjNc2iKcBRq2dqk8y1A9AEcOXtMZcCUAplmBvv9ppwsvWqIK
RxPD9u7aoLe/3Rnz2kg4NDTs5W7LpB3VbYo/1Ij7b760s4Zk77x+VTNic35gYTFl
bvAcuHWIIaWK6jcQXbinU3/QjlQmB/6YfTZGyGwyiyaWdH42hkLcTI485F7Skcf4
l5EjAFxE8IcaAitTul3tWe2zT0DBD5Qe1+rc55sREMg9Yy6aRFs9aCeMS6fvWAdr
DvM/8LLk3raQbWPcav2zNcxqTOpV72nCnOSwViIcIgoUGlnanI8WuDUi0pIFWJNy
9qhop8cKqWKeI0vfb7PUH2FYZjIGjrj9h+JEiMY63Ko3MYjCV0LdvPJ4fT2osrvU
Oc2yMeaLGwNg1FtcAPnxZAMBzS6a63rg6Cpdn8aTk+XJbmoGqx2GnWEDSGWFrFpK
DS+adqnSNBIdlgUJ/UQ/DFOvRnbsZqVDTwJz71VW4mvHAKhU/fwPTqoC7E1OBMx7
DA+6awjJF7/l9C1SQznJk+GQ4iNyV8gJKmwAI6BuIgATsq0f8ba4hOJxfCE0sw0m
3mIqoOKhNHkPkvroUgkqBOk19DaXWFqhHKuNZOXYeTJaBV+zzLXDAsgrX1RlH0+b
NFX8iSkanBem0BqZ03yp7YHC6djwXyznLzoGWJBhksSGYtsxLhVFrbmd90rJsWFr
0KafEvvDB84rYD2qqphV/X+iG6rQvlvNmBro/Mc7bXtliaZUShVS1OPh5gj1Fm+i
8npu4iIg4fi+WxTwHS+Y3Lx+YjiWoZxQFKrdhV0sAWB6AdR9q4nUONzZtzezJay7
psJKxo3cDrW6nYK/EyTxAO4qaXQfvRu4vIFJglhoDK9oJGav1gnpsMxGRqeJ3Yku
da4PMnfmZUvj0FySiSu8nNIfipuZSy+pvYx2Py8zDG3KL/iYkvIpSiT9RDoeViz0
5bj2YQ7M/55NmteXvvp7nIUGo07bF61+7g+1UarDF8HtqjBeiKcbaVuAxeNbGSYD
HVdS/ZAIwPD/iMe/Y2SxEj5EpADF7DKW17p9bwFVLI19AQw0pJcK08cyn51GL6j2
e7VN/W+Fo5aNgaBcKaz+tSik45sC2rlx9dJjmr4klngPOSKypdwVIKRtI9DX1Uo8
ypeHqhATmjpvNjDWchuIrGLpJqb3xdzoT3yNkO/nubVmk7cQkMPC0+7Wz+AMkDV8
+ijaR/FzMwXuEW3Iu/ox71Fy3p32KmPK898ii6BHUmrBPFFUlOuBwG8p0E9YvHgY
x1PDwzSD/G3Z+yQ05XHj/NXZepKMroci797Q6xVU7v3glQ3A269UUYPjqCtv0BzV
OkqWSxGIgKd4ufsdkvQqIf/hpWmXGZcPsVx74TYsTsWD8hqEAB4/WvJN/EHdIQFP
kNAHuvoI1Aa/gaNxU2QQkspKM1GUXLEzrxsTcg0Uluzv0FTGyHPT2Gk+udQrle/C
Oiizn1rQWuIBNEZFdcAZd9iaQDd6f7SlLKI4tAoFTKcr04Z+N1QJ3ivWL5Wv4V59
SiQsTTj9ArcuOONVwChgOGLbjJxn+HFN+ogXREmwi3gzYcwZa3ZhXI6JZfbBs7GO
jBW2bcosmPafBDb9PEmIM7b59BQudQYiWdFdIo6rzEBzCwDc7UipSE5lsMtXvvY1
XpDZmSy5y5qFZ2RXY5MBwBS82yMkkxe53BXFBP0KeFUDaS/8df8dkEmFub4NQTfH
bp2oyyp8wLRrbNFb1R8Ppgld+kWD1fhy38s4htzlW/1yemn25JVkjMWTLVPfmiqv
WgZQYWs0KEu8ewqRuecYOWu0VMXLpuHwCwhp1V3A5DTtcDIgbG1Hagj91lHLAjEO
d3kYGXzO82wKVtu72pRRbTdV/X7gp0Wap0oPgdV0SwLd6XP6vscyOK3JXeDALPM0
5RMrWE+Uj0KRP0W0bxS4jKhDI2CEYLcci6mGFcBQVphImxLVT2N3Ero4K7VJudJ9
c1r98YS+tgS88liS4ZVmPbUZXGPfAknf3fXlkrkKwlVhxR3QiSjY54shD1ldQU+B
DUbKIYE+LH5BAR9O4cdqiLvVRBQ9Makw7nzQlC2ZGr12vLZJhwf2R0zGtUfTGiFq
SDHnZguvaWl+P8o8X2+X64ry82xoKuqCpSiOiEANJYk+R0kcPNnb0k2585KTGgYE
3jgF5LTnhlcHzZi7j/FsbeWJ/NX5VHo2CpwWPRnF2jNxo6lf9WBLK6m8XHxNK2Yb
GCPphGUCUtgVUC49It+i7Xu1GnSazxzUXzQagfcK2DiEDYHzj9Sfv4PiPy4ZqsYk
vFe4irXbFRK1SnyDruv6YPe+OmMgFUGfljEWKGjahH3DyhEvx/NUFI9yNaqfTI/S
EtZ9PMNJh6lEi29gK50A+hsNqCupioOKPqVGoBBB8WwqbzUDOcWguGQ9THvSf8s+
YJlGS8408C8tFDuZI+nkpkLz+HsEAWCS/nrY17nBd/T1rzItvf5ttnEHQ6uk4WCX
arSq2Yvg0k086Hg5JVYPCENA4vElKKpwVoVJ7DBNVelyA+o9EejCeV4V71rbyh+T
KvpNMpnSTs8cYlU2WuB1yUa//O1utGHMxmSzDVmkrGviRlNPQBZUyCvMTHoPe7Ok
K0d5w2TiCb5tHwEwRIw6h64DbnqCZ/6/tTUek0016zJ/UBy3HFepy47dfkQP2Tmw
LFcruJR0+oYztxtEudivF1RdIePK5n8Hm4WmCCzj76iudo+OtCvUBk0JjWegLaih
WB+zflkK8alopWEZZRG8SuPJl/vOgH2ZIjzggh+UQ7a9siLWHSTe0soItjwXvuK6
JVTDCJk0q15UUUi1NXeT0TZqn1nsjQu/VsepJYLjJn6nEub57s1e3Um/X71h7hQc
gBFGAeGXxda+OmL/uAEwPhj/zDjHuRs93AUd3D3Nn8CJMNPERZ1NJhSARn1OY5p6
tcKTx8Jb6TDQfPfv7FPDyTNrdfhS9nfzoAdLe7AgRnLkuS1//IevCtw+Zpir53qc
f/eegqLP1onFNF86vkCoY61f33WNKsyQ/z2s0FiT2ho49JbwLqzzavNm3RhQrs9t
bgbOIN5EY6+Iwc3nDLbSKn7bzZZpY/gTW8ma4lMwkrKw1pgzUSnx/2pzQYvRGwW5
nWAffXFWfZ+UGXRBrD8XenlhEdiwY8DBFFM1NMdzROhmGLcT/mLyZRy4mDa+zPJW
EULjcMABpVGercfY4Q9ZrCkJniFSuTt/tViTj9jFIjggUDvKHPVpZLKZ7fiHItOQ
FmmZJ/GKPpBgQMNWFjo8+LTdhrfgh0QU9+3FSpMsrmet21QF8odSGxbvk0oyVUS1
kJ0CLoo346C9WsDIct8kUeynRqKdr0EF50lvts4BJr/AH6Z4bdO2kdKV8dKpoynn
8EMWCGyoEzXLrr64u1SvoNIFA7CyxE9qLN1caG8zfnPkfFabPAOBbmqZ2eyJ0utn
USex70s93+8QiZ/Tb4HVzE6T5RJBEbdKYNhqDEWLVCFiFRo4AAqfF/PtLmbfSezF
+UWARv/hYk1vMSBizmqMGu8pps/WJdP4aEKg++be1R5K11l2qymgBYRWbfX1PXrS
mr4ipK/0FFO/Z7H2mAuMdFS7Jd1QSnHXsU1WirTsaidNSVW0VjUXQ84jlKZ/GV+t
oRQTMfIu2FuKKmF0LlxTLFbAsUiOsCqfd5wsaLJApFxwd7QgVaX8OMonumo+2QDD
iNDa1jyKtDq0/Kpy+47ebZm+HJjhsobC8mZIyhvPEzBWY467Z6ZehftYI3fUSDov
Lo9rHdgqAfK+W+1LtVtVBCDRTDFX+HLPmTMrhhp8WXqgNxHR2MTtXcrKEkHBxVun
LdxqS4braaKwX+MpflDiamvWfYW9RHDVu/fpcjKN7caNjF9lSe+cFoQE3AeEooN0
BodXkIbDI3TUgEKYbF8O52R8yx3CswdDEG6FFG6cx+lLHRlXD4/ZJo94MZCCLK3C
Q6yUuukf1XtRC5XhWwZb178Q7fUS8kFRgCYduVNTTdUXk0ZKyYhzw6siYNTEGGWE
cRZEu3I0pIUw78A91oFLZkS8R4ycJtGamgyFmVmIhJjPgiPDoMUJ7Mwr92He9TNS
7wHkpVL4eyQtIlkEbiyaEOZzwZ2t70AvwTd/uCiVhb5ybG5kMwmnpg10xOCW89eE
hvoh8u6VOuOcrKRwMx2Zac/FyecR+/dT/rRo11n5l0wZyiEZhMe4v0cD+hsEGXu7
PUHjD23phn6E2FSSfnMkrtCBdradD3TEqo9/RkjeR+MHZPtBxBRBFCjxlsFj0hR1
QSn6Yt8rAguizH2KpjuohJWbQGWGmbvmwjq/YWvY6x67+77PynfUtxSHHnXi01q1
TcGOCYpDD7F6lpSOyLZ03T0/gIxMH7fpNGzTYmIyX0w8KAxfwxw0yU8coDSmp4ju
W9xWs/o3pe/Ug9yXT9HBm03EvPGS/3D6KWEPZA4/R+PQn+dvM/kOSBxdb3gb+mII
C/OhKwcZBCalx/2KrTnf82WhfLBC9K0uzKy6hSQ8mqTE9eF8wkxpgfLUVBs9uYJW
V3/JG8Rdtcd8Q8ZKbzp6yU2YNhzouzCiMMpq0BUkodtwG1WD8tdhVAXRtI3qH//i
48IZfpMQGhupZ3jSbi8/yEWRx1Vv0QAKwFUFWbMBGX4Sf+w7fogUQV8A/z4IAVwl
JNTU+WwB9VvsZ605yH94vOpiUs1npI/yPwF9yg/uQfE4twN+rWyPMsr+LveJzXQN
UoCQOrZ1+n/YKQlQskvRd15QqsgSpat2u0R8z+IrwnXRFl30Lj1W+D97S+b3KcxT
dOp/Eo4Asis20INOfZRJSBb3es5jl3WyA0sqELxGbCp5PX2ccmegaRZY5gCJA7HI
c44lkZlMJtCR1z6gCmjun0UQr+R07cH9fMV2cNc877EFY+f1TB0JQcLMIp9CbBW6
0afktxRatnI0C+9OBahwX/RwgWg0ix04n+2SmqFq+l2RNGf401gWlbyc5NQ0WJjV
TMtxLy7ApgSK0e35zIvZ+5Aprclk/h4O9kQIopEVA1zqu6zzU1x6ijoxxk/f2Hpk
JRNQQvAL35kweUUELqWANQP+XNgW+CJKYwr89wgvEW0vWHZ1NChnOKpLhtLW788W
2NWcJe4E7NvcasLPYuTPzQMSxBwmsI/n3oXQQC5pJntboIjPL2lZH/2lkoawzDN7
UHRHA2Vxx2uKpv/UT6q+QjM2+GO3myyixCwxa8kdz7Y12hOOMqNBUvGxNVhqJyXV
N6f2yW6c5g1Uwr3Xj+YqdcAdD41xOB1b6MDyKRZEM9GmaWSp5JMJLsZ5CcSF1RP7
RaTwKMnUgGvTO7k/47kPIm1qd/VTBjdg8cP9DGH1mMLsiMfXcuX9uUqo1juRPH4J
HwWNErHKpwDPeQVYIY0GJC0JmZpknHqW8RkeCgSreWQ7IUniec2/QhEi3cy4vzrH
uiHcH5xhStm8bSEwces2FEwlB0jUC0RCCrGX+y/GPNmTIt/tsFMEzR4M+cgiqyA2
Zr3LprXrm11XzeOzln7bNfJGSo3yv8HIj1Z1F7lUyO3r5ATpP03j7d2SwoJmdbzk
0rxAeNIGc1IOpBHeoBlYUzona/sgfn668FyG/eMMUcscDEjySgD9n5jjifPer/Q0
6w/3cndwSb4rPAlmtQNe3DeA2mBBuIiMmC0+L8zG9mcmAVkt/jiXTyLRv3VD05UE
m97EiDu3g3Uj/nrEQRmprpb147SoebeWuQDSj3EIxTqd/xTI2nUoI6BNYc0PNR89
X5cQxXmJ4n+BRsoWEEQvDTJTG9KJZ9rNY7XNsax3nNChtqHOn4w3p2XkvloZTGJx
KhP/1Jqz2uHN06CRTxiTbWPBVJl//URp6uPADSCYvhs0PgD7OmFHkL1M5Y/jAqaF
s4xEKbvRth8nwaUKiYGdE7ka6LVTa71dpJlDLQZiniO/7nmowi//t+X69r1kUVZT
kSAz1A+MGrdEXof/jhx52wJSrsplkK7yUV3X4Mhc9cUDhu2coTt+G7KYdyliG6n/
pX79vBHnfy7zk2oRDV5lYPnyEWvbwXYzDOF/n0rHUPfLVaGVVIfOq9XRMCOylu6g
xe8/gPRx3mG1ouGPLblx5sVSB+IESpytep5OODoGM6CC3ayMEbJIL3m261ffYyzF
+ZsUed384OzToA+A3Sn7jPx0VPVdEOxvWHk8tGfNpOHhT6xzUIyZouf9RlddrX5r
ov8p0Oihzo4rLKJt4j32w99qu47T2MEOfU0xuachHaRYRXfBtxSjazG+qekdbUPr
LPyKYLt3fwSzJNNUz6cojFQSppqLVLIhTHvG4QIif9QjoH5RddSvo6rsF3FL7JjM
rO6iKVM8oIbLSSWmGDTHqQrzzwACv84UJFjNOWCaWLM24WqT3yVhSEG+xHqHoNHd
lzAt24O9/4+7YgZAMJx3S3RksihUqJjED9ZbzTTFNHdsoIzzUn3UFwClKkOWGHyM
xiZDfvBqLeLiIVw9DO7f0E97hCi3XeNMBMDjEwZ7VY5M//UVj9fgaiGBXagNo5jb
pNge7sn1h5Jt2al+1iz1fGhUyAM+x4lGsntM8jIpyaHYMsnDjV+xu/6iSdf3sqR+
Mr/Y1TQNGJFtojzBfXBClk7UWaeemx1o4CmdKtHa1P4fiYe+2ubqL+9ZBYp+vyhp
fPIvdvtMJNK68ZxWNe8F2NJS8wHQZ9dGox9ROvf84i++pdhyBpqf4ONE6ye6E73n
8NzcfPSEqeIPF7S7HoqGf/QYEECB5Lymbo05J80QUWRipnUlC2NpdJ/3O1n+DNNu
K+ErSue9qgdwHJkkR+uzNp1ic6eIjNTc7DB7NPFEMH5TlTw0qMDOuCtocWdCqAbz
c/ijwQfEoyClDPcbl6ph/dP052ijX8eQoiQsGV1+5buiAGqUbKvF+lMboYAut3W0
R5Cmk+tE3GpfarCblOyJ+tryy6x9GMMmBaQSmxxO//vdmOrxWdekm4zBLo9GP2AE
pP14PpoF/sncCTF9110nn215mGl0UAc9J53H2bSkgyKxxeS1Mi6lrd2jEQBJSc+O
UAYtkFZbHzXfzvHKMpxL4Jskz3hK6En0Cphk1HlAsolM2/G6KWFDLKh1ULl9CNf7
/NVdDk6kcce19y8ipssPfWU26IVXNQ8863LGKO2BAhA5DoSwp2+8wgjrZpDgI56f
CvgpOkajNgRTiOF8WXVoeIn9W0mGOKKM52vjS3KpsLYCUJ/iwZ0AYFV/qGMszDnW
pvbjnRdtPXPz3x8sCD0mbmzr0S2FYjoibD/sIcw0Q7ny/oOeRbgkQ80ys4JQYlc5
SH3lAU4AnWltpRJk+/VmKUJPup00HtSaAUuF3xNU8m1QQHgD4pxVW1f58nHX3QwV
isn6C9Hg2AmM0PjAKfoqL1NGUvtQ7/7vTA5UmAF7c0KZjWaTijxVa5o/J8hNZm+F
14VB1U/R2+wrE9zVF5YjVbjcHmd6Acz0wI9wcaSxaFe16b37NQMBsYU/cbtMJECx
YfZljuVl1GBlfM5QK1kj7PZIWvU7vjnpyG6pLGgXRZ0KBVztQgbTYB9qrY5plk4h
wrKaGI0FrRjlv2ZwKilwnX3S/O9jBZEWp0/P8RJEdM9BC5Oymu8ItnyrYwLA3I55
fYzJ9hITZy7x8Yi2ZD52u4Uoh+jcH3z6z1eDASj47kday/U1KTOhOkVZXh2+qUXY
dwDrYORZOwmY3rAMHQIVkjDdx9tPteDVAWUQQIliZ4w4Kzo+j/QCBbxWbZZW+wQK
0+NhSaquqH2POpkovi83c52DiZBdSWaOAu9VHmxw7XIuJllkQbvKbsyIZ7y3EdV9
BFROqBtCt7dJegRrwvIWoQnMZ0kPGM/PsPPG35PuhG6aqqi8Aa0qKTG1JckNuCWB
KsSz3xAXs7541fLT7oGl3EgtmpEqXjpLWT7dc46PGeuAg6Nk6hounO8CxW6PXVDt
OZAwke0xcUlgsm89o0/O36lKN1Z4uYu3stvzMmWqqNC1ShjpRD6h7fDSWMaXR1mi
JPsWag39miTQa5RiN9BXwNwj8vZUCR+OFaacsKG1zhoqbvDTYQvoOOFZZBOJy7mS
yncxZ6VqJ6zmHHf0Jokg0snCaW0V7YBQ9JI868dzjYyVIlaXZG4lzFkX5ajOnH2j
eAZOoWNGe7ruu1mwfDEYrGYG8FiFegcgmm5rmk+eA1uxtHgZZrrmzZnznTomuCTO
ghdQTTNsuaQZgDSVGTPtDVl7moPiQjkXtRo5r+mBt/rImgOFyWtyIpzSz1SxfL8V
yrBcbpWzCSMDl0DysWVruGCvs5E9ICMoFN/9EBFxaoEzZ1MRVj0sbf7UHu1CPLyH
fbh6LGwiFlWX0SzqfIYqEhChXSy3YRQsw0htrr71mfIIdnGhEn+59pMjZjeSAMZV
IzkTLwXNcBM47TI873Q4PC5eFE2Ps8Em+c+XwPQNOpYfxMiily382sNsgH/2AgM+
PsT0fQbteXyqsCDVd3HU+eCQIrqQOVe099RGvHAYaby/bPVneobpyJyv1kZoO6z+
CznYkbhKydClFOGGAOx70IUFE14hBANxo9u7YtmuKz67mYwJ02y04zdFAZA3IK8O
v9wGLymH8msOS2uIhOMafjt5yuuEpJg+BIcRAEABM/a015LQaD3nvRvnpEQQPQTI
cQX9gfjYPNihgnJHxe1AE6hN7qMGnclgvYIx0ASMbWCJGJmKMXA/KfA39XjT+S0p
Us7XwEeQ4lQwigXszCBuAXmgLed27vTEF8l1mE3xonDR4nuCDW4G+krlGE5BjTdl
/+HA2ZnZ5l3ZWNkLHx6NFpOSClaMDmgzvGgEilLC/bXBXLzmWs4WdjpCjbZXSkmD
iasXbPuhLFD3DfnTjIZyZLrlaH6jWdxx8ya+raKjbHhzupAIjvRnOLmFQTMpD84H
0XQePAjJzoebFPdvku23PuTE5IsXpRqrR3Z4JuVAmXywwWM02tCJ47i/+1qqZjLP
GKQ1u0QK11xWpKwXMNcpJ58PetaLfpW+wu/RBNw9xFCPjOVPqXnuioeLSNdAuUUX
v9bo/RJjbt4rE5+6MxU7j0EK+xKBHnXi+Y/Ju4LeGrKeTX0Hhu+EBU/Gqq7vZ8vo
CBSrJ7q1NetHJ82aCrwZi0PQhTYAnT0YXYxzm5bTW5u5uj34hy7vt9geWTvLgPli
tncyEFmk1P/TYEgsYpCau4iYt5HtNMgBCOIvlLJra66pWbABsAadvsWlQHMUzyrp
AymCv4wVXn5GihD48UqSMeTCCVTfTyazERTMv+n3eX+hbEDpwoGzh+b4hKE+/YRs
MYoUDD+qyC0But5B5oq0dgGoM5xwWrJBDldmsIm5UTqT6CkiA/SPOVf3UlGc6j6/
BnbPqxNtZy5Z4pZIlzLAaohFQve3YMaKvm3xVaOUGBPI4KcgBUqqKOHO6uyrL+L8
7W41PFyn28zzugTVm+25zcLoRt0UFH8ZfbVe1C5PKDzdlhNaLWlJnpUkaKe0xIh/
DpKftDYa+SHdQGQKEMAVtoL5pIxQ7T50P4c5yuOvjq0e5/l8J+/GMYG8iuehMZ6M
ArnZqY4oclcVMgYuAXBUitl2P0/kGWU+HH30uAaof37HFFoNx+aqY4Z7Rj2MCbDg
/G2fAbHa4Zs1+41Kk0Cj9uGJnWk0l12Tn9fKVYu7fh6XgwxKw/+quPCDIToyzKjs
IWAGMnlX68sYVQ5058t9cPTUs26xF0fRpMY3/G362MWc+NsC4xGL6p2sFMaubk1h
SluzPf1K+RyjW7tTLiAXvkvkIHDphhSvEd5wv74H5C63FbaTKROMrxtpmTnqDqWw
wxg/odBWjEK76nIEuSGbW4t+hcFaPjnCkKWx4nex06F7ATdrV3Y8BdHyiF6dV355
EzTh9zR+JH4YWM7FAn8qCSsWw8nIxwGawCQN4LNHGCYnxc9kfVGGxoxr0yPClkIS
n/LQoVisGknlqbid5ansQoLlSBb3PI+WJHMZAyVdgGtwSe92DZHtAz10iT6jQtEx
dLVE77EmblygAwU34/sCUDPum4x4bZeog/kmuW+1TODu6ex11gV8oh3qLGx0XeFg
u6PpeD96+rBq6i8AiDnXEkqHsoOZkKRV9p/AjkTbU6LNHlxQKfhq/dJneyM8h0Ri
QIznSl0/lPdKXkHidWuPm7U1zGC+zS3fvVgNFFFGZRCnJrzc7nkUlMMW8YVomLO4
Kk/m4uiM8YhAQJelHHPuGUHdVsbQWeOw0myktRU1208djZn+In+W9oUhrwEzuKny
7kq4KN9iTncmhO7c8BHC2WD/QX1mSdqeS6SdYgE4LauKFYFTScWaB9Akgufkk05X
JoCNBRkUcvY8jwiPhgZkJ8vaH3zGnp3guTlJgopBuU38rMJTa0P3d6FtX3OGENT3
p+f3j8cFf0NNPvo0991ovGiyTzN2Rr8kagtGXr6eU4BpPmjvJ/D6qMI5TvHKv2m+
Ori8v2ZBVXJs3uxjJQutDOCuONV0Wy5cgVmq0ddd+kE9wOjZNW5Z+y6RsztEDzqG
dcYHy5/wzgyEcVOKquZn/EpBlWNm9i5AfYgISzwPNW7lE7CJ6u1RSw7kpTEjXq3g
gsBnwHJEkLXU9cESe83KbiaPxNv3yTISeZG7dFQ3o7uEUavh1oTlPivIg5S63/cO
+2vfUTMRHQJMlyELJ35FkgZcvtuXvWfxGG7qfdSgn/0AigGMMJMbXW1UfQxTXhLV
MQYA9P3g7qp2EApDmHUZl5ILoifTwlaT5VihMxysDTZ8AQMgf81rySaqhhSvCUJF
O/P3vm6SjZo7VbbX9I/jn/7lb+g/oBl2xjOfQSEXcIBqQcXV/hv4l2xkxOFREciW
BkZElHya0KfijBJMyB8mxaormDuTK094xHbCnmFAeXzzA+nMYOZV9eD8+XPbpmci
5HyJa5eudnAALa/N/aE6xyBeIjNfcYIYy1sxOA6A9r3LF6ZrB2XtdkDs1ck9Ptzz
sLF1V9V07O6jxMhLXsAx2rmygozB0dY1GCgbrg/Wvk4Is9W5vAMpJB9L5sC9uzhV
bmUB+oUvTCHgELCURscFwRbuXBgBL85rEh9V6GhM4MJhcIerSjk+vAWuIX9U8oN3
3zdjBXHQLPfHgq/m/oWcFaNdSg+sJiNoO0LpxUf2A1L788vrmWcMts7fbZQCs4eU
gBn1Yw4nbIv6xSJTF8a27m2gTc7Oj52CHDKxzN9VmuH4LDarDAfMTGqqGaqpNl10
pc3K+8ZhNZDhfHA2fuN7/B0UgZNdXRcMf1xHNJ1deju4XtKJx2D4Ec0o3cOqqrDY
ctWhsZcdd7ezwzD+2G758sMeu3c+Hl/qEqn98z+X8wdPPe3MJ6pA3csCxmRS3Bha
q5CYodmQFj4J85ei8pGBkOf32vTZ3HlJNcWqFZAv3Wt+nqy27voWY0VSn2R+i9S0
yo5PzwUVxUWByDr9cWkAZRyaUYorqRBJaxDcUlDtnNTJ8UcoJUqtA0o0rGBOjXda
i0ei5GhJYjQF3SG+0Q8hecZ4jxg0h1Yd+NW8dbhulqf+txXA1zGSGH5JtLCLKXrD
2spwz3btWkp+cs9GtQ7IFeAInhlfdEYOKydi4Ny+MZz6/YGnpFrMM78+ggBsLbln
1aNG5wyvlIKi177PnSkg+LXx1cpHmn7yklQ7Fyve1lO9xhxvzQBTlJu5f/GMFZ6b
CXt4Jf5nGe+plNXzheLKF7ioIGhIHFqpTvX+gkWcoGDAIIJUVvED+XMB+z9TKQR0
n+4TxYViJ7MXMEG6qb7OOKjxu+0KnWYKG7rwFZiTp9VpX0VwpOpBmapzwmsvKIC3
F1vNw2CMV9oxzOzPJ0xpXOgLEOR3mG4wdsNh1YKcCllb1DJVhKlnDZc92DWU/tLf
1A4TIhAwGsf47z2rdFYg34dL3r20zgY6mH+/kAPM+VU3G0nl3gLMTUNDtokLpoLF
RRJ4/G7vp+Wvpi3YJFCvOYP3w49n1rNIYeR/7HN2SESwUWys8envRbVya3evcus6
aTgDMqEgQq9BSPvjdlvZTl8bAFyGg2Z5uMabugBJtoY8IB75I5v1vi6WpwPRY1a9
Uowu+ZuIqP2ApxUo8v+ijAo8xLGj38+oth8Qvk2gH9uGoRaFWL7fPvdnQPCRclk2
lfKwq1qdG0hxiRHaGpdY1cES6vTaxa95dpCVjoEVEfzDFT3nAccCEe/iaQSaqVoc
Goj4eq2c5R2s1816waBo/qcvwG+QGShTP5EjkEnL2AWR3IWe5hk5OxYtxFvbAbPd
/0RmoBe8wD4H4/3U9yrh0VlP/wCWUXXsI6kBelQ0IZaafuhs3DwFsNu9iZDhWe7J
tnEGcYBNi9CHcNCmG7lWTeU7mTzVJs76VzJZ4jfG8ZLDgqOCWlNelTVR2A5jUmhY
sqia2fmPK3BBVo8YBvlcurYkP3NFvY0WO2Y0Zk40CXUyg85RjQrBYyjTtrUAIecE
gS9DmEcfEjoXYIZRMjr+Ws5ZppFvC+1PL5tuVMvQ0yjcwg4lLLLWKbLZsJXuLWXK
uti3zEw1FTIGjzlQFRKq9hePli2S0NjmEhfavtVz3XtAv+M0taqpe5iQQpB4p6ll
WBX/3k1SDRZpnbiZrf8RUC1aArnEoDT5VZWNZ6q+Se25j1+xYBftOj3ge0dw7909
capYESQN01WFZMSbdVwot9ticYk1cxcBoJYuXSNNuHW73Xv7Xqr/pp+t06Oxxi6k
eGvZtJ5Wa47wJCmrJF4T1Wlf/e772ZheN9p0AW5iEK/Q1f3nZa0qNGWLqWAwdGeb
3DpJdfqJiAqfvSVNdpkCUJImaLEP2l1Al9aqe/dk0vKbszeUWKA3ywx0Mkuwghit
YNf+aNp3ywZwK73UetQ+lzDD+IOcAxTQeC+BiqdmNCBvDLZUeQmlp0HBj115EfQu
Ox4E3BGrnbJ7NPRvPR+UBK+1Xgizus2hN3I3CUasTkP5Jt42cmI/tOqk4tlQoH+h
8ySM5sTyVxoy7eJsAtXT4B3co8WkyP7gQ/rxZrjVYd7eAHw7CnTdLfoYGmBluJot
b1XqwP8pckPvBC/QgOmoRyUnkYOljco2uJfsA16JAwl7NNw1gi535Z8gFV8R9QWH
8uXIeZBTD/eUWSjkELL86lu8eC2eDbZS1CRnn9B8cFSLAM/rmirV0norVO+EXNJ4
bclFK/omNzndIbWTU3WJhxQPacOvn0YtskVgx2KTF7WXTWOzIK+YpaSDizAO7Dgm
FHdJphYYLC6JgcOEOQaTnK/OZ6gU6QmNQczBsgFj5vd3Y4vM/ByTAkC84k4zpSZC
O+ata9qe9t8AWRvKrD1dYvzSDUroXnLCqdlkFMv/pvgIK0vKQOQ+mBMWBhBZu/TD
63bATCP77weCOLWb+5ji96w/cdUdEzN7FOdx9ij7A4mxqrJS7PFxRi6WqINrgPKY
SH3NpnGG/dQF+RNRrK7KWD+NAGtcOcLA5nvxPy816Q0JWaBgmdxMMyEVAKqSJS+Q
ccNeM8V13Xvsh2bsjRCMxhQurCtluZHGePP8i7o3fid9J0HF1ejZ4RPIN7pjO1ab
OCYgDm80PLX/VANN31CCr8ooqiAKKVz73JEhxozO8wb5RewooK4PcEkaUCUESwc7
Gl0RR/L8TW144iCfQh5ikWjL01RXvNhRk9gKAKOF7IamcSWM7H30slPAhC6BLa2/
wgwxt4Hys0zXpVLWvHeKmGs4E3U4j1g5zkKiQ+NB9Bs9CHUyfcX1ppkG07uKEoww
GN/sX5RhHtko00O7kJh3GuetYwBw9gDc3DqpciAFN+0Ar+mNVibPwZ4V8bwrRbi7
nA942ZCTsJF+G9lpfyS+JCZxufXvFjmShFCr6ODB/yB4QHMNGYuG5iXRajzikTrO
Mw0PWEMFJcZk0raRfY9mkiPLTQB7o/L6pUfshQmi+xvZGzPAU2lle5Cz8yZE+XYF
3mL+fm+wt92Ike4XeHJQhKKhgUGaeKeUG5b0HsCmQuqthaMaSRf8qJIRmgybtFPa
xWo/MUfBWTp0norDR7yKNeBDz0KXwtuC3gm9oEeT4p0rTPp1GsQGOmYTMqKadDgj
WU786jXK37hbNBUp4rPMrKa3r2fdKR1TUKh7eFZ3M3dmyF5MTVTNKTtq3Hi/HtRm
G3uan96eUxG3j7y3XtZvSh444N09QWFLr183zhyPT91MP4AVzehvxyUnZI0V96Rr
m+B4xKOIBB8jT9lcD0Ie5z+p+ceAsiDA1DqP2pbuqDwvdYzj4rqoBG85FgqFkQSp
ao0kj569e10xBDevL77tz7trKR0ORimTJtWs2l/iDpl7BI3zP4s5Ua5MRiA/eWS9
xfrOoqzzwn69gV/hjbtc1gnaKzpwAcXtxy2JQIUzTakbGOv2VRtjTeMOEsw60r+b
n/WF+uYrprDWYr6jydagirjXMOtJ1P9+1GdeMdf9Qve3XGrgACj1JCGKHf2vKajW
bL12UIb+Zg3gTLKV+rbdr6WGmn/WdMH07Rhf2M6PdHl0J4XXOpHH7LkIi5JtCeN/
sSrKoeB4wnV7tCR5YmJVBLfGmOI4GkXw6jkA4uwe6rP4lYY5XA9m/MoyYiLnesFX
R/2IjZU/dAbVJJ/S3ibPIB533cxLHLHts+oa5+zudJkGB0NAmQGKDapbpXT/PGtF
mHjoveGRvDlUYXKw761aEWjSJJH6cq6Fss6AyF0VaF1Yjj1BBe8WsxeZUvOuMjcH
ObiFKHAaJ7ax3lFeouB8aFxpGlI0MShscfr299J9eikfHnFIgj6FTui6z6eBMHTW
FyRV5pYIB01zizRDl/JJ5IljikbYggmZNBP6DbFykXEDOSSiBl5tNOZGu/kU0Tpi
QaNdDiHT9fPcXJPhGBfQGvx1618ikmJV/seAvHCkNTdh83MfHYwhHQiSG377X7ff
5+TsYETRsw/6Q9jXcXGDCYTLfH7L+Ea3DWv4xc41vuU8ll6249i1x3fxwZZ73cKr
3HBthByE3/h6TsU6GiuAUnDMhYTXZkrBCQZWvfD1u6d8Bj0wCcuHTV66flEfFDJK
KMo8AnYCqZT9Drp3Yngo/c3WKrPQwLH9YfCoX6eXIUf5ZHHW9ToCHV1mQOQZYLS5
aFnZDHov5oMzTdLRqt4+ZlFHpU2uHcl/AfIryMWUNdMQPJ1lfK+B3kF9gCQbRRyC
A+MPEnny4i/QbTADcCw7cytkWGR8uu9lx0wHYuabrmkIhxiPzDOJidkZ5DaBasYS
Y2UfOX7kMSxGEHRr7q38vQtqOWNbpnnmhsGGmH++keIzyY62QZKxn/G2M8Yj6Zl6
M9zAFDbQ+vnr4e2fiEEBDUHSY4qCFaovfpXVVZ44sCMYw/GmdJmeXjIWJsFRSo94
+++EdUNBslTYHTX3o9nog/ryeYJ1dvg9W0LPI6Gh9B3ZeSWkINM3zKQ5UkTVLMlI
UKKD9tdBfOvIR0FojdtIizfx93j/2TwBKPFNHYGtyDjswt9ZyZrms1WwN+ZqxKxC
aUn/94Q7iUfbA81Sh54RyJ+pQS4CADmtfjP56J9uOBGpY+t8oeLicJmkkt5Ct6JX
NIZcGM4BVMQa3ovhHpsrwyOrXGE9vrPYQM2vs8HtPb3ygiY+hdJJn8B2loY6fcuJ
TwNrmYb1XMl3EvTxwQKEgbGTUfOdLz8J9LqIjufQ+DDaJA02XGqrnK4FbURx/Oms
cmbWuGFoge225QpAKTLaDARmQ64eMcCbpgJUbvoznm3t9pSth1rKqjOXhorXTxGb
7qjyFRp94CbaotU6CrMbYV52XfaCQQz3pbf8Df6T79XtsX3NFvbgSsch6fsTEEHE
9qYxnbjGTQzapGKtQVmjc+I48/JFpfh1uKL5zWHSudKWz6JdLU+n2yHGUJqQv+Q1
Zzwb3URgkiF5bg1yi5p9t3z0yjIlIk3/3pQfAQ9mUbk5XxWPPl0hNvatNxsPOhht
3+/8tdhG5mznJCfUKxPjkwRmfGQi9KzgtvRNRr/iuW/8WuWnxjQ3jiY2N5W4Mo0K
44jv2RVk+GRhd+d6s2kq8Ai9owxDje5Wk5aOKAZY0un30uUqxP9KQF+YpSH8UuKK
/GtQk5SgSKXuFZ9kXOqqFTsiec1YT0oNeYh7uxQDsY4qA1GSnQB2qVZERBvkFefq
ZPb+4DM3KiGz8JP+LCCIzIY+W9rVSPlqHQwZEvojQ8Xtpfmff+zmZV8fibSQP7Jn
3T6MjL9fKH3sIgqBrmDSGApTFQji5VPSQQWvOvPpJTlq6WCXsgG4pkWqGBKwklxo
sq9nnbo0FL2HvEBJ1JE+yvz94zCkPMitmlSHrXs/939wRriIuihUVuAp/QJfTfxd
nZJ1gfugYFAJCiILoGUYQYEhGJdIoGzuLxzKZH4peI5jpK5bC1BNOqUmvY0Z9MpG
uTiMH24iE/3PbpZXYrQ57QE84puAE5BwBpr3pFJUo87CW6KNMmTXVzdN+032v0pf
qdRWcRlZSc9ntgN+QqsIz6Pta5ZnA0JU0dEJb1CHheh4/gyUlfzsExOHukg/WdEd
WInLer9TTb8fyhllecKRhEHC5i8r6fa+GYNT7hJF/8M91e5wQKVCjrFXVBShoCWT
2PyJLpQKdZbra+gRpk4h8hzYUyW9CxfyCXBKwYA44Mm7LxRg+ACcBATerJg3EEgX
N4+8r1sWMvzw0n3OfrGPS8ZkovKtiO4X9bSk941uBBiPEJgyNZ6XJb0m7dZSS3UW
Gf1m3TdunOAXnzDR/ZjV/JzMOJkoDkuqKxtxfG0rTbL+zzo6bwaZ1wsol5PLAS0L
ruPPRfX5wBajc8PHd4LL+2uYMlvEMsX4w9LJPFUeggNIyrFdaK5XZaK5EWzWk8Xv
irU4FfA4pJPo3o+YXOG/8K4vDcESXwwAwpN+F71n1qasAHXjVvVeo3J0ZkszxYfP
vHd+E9oG7MsbR+RCNNK4PBSHZySWIOTzZv7J2cLrpIzcaCC/4ChJ1DFoK32OapII
VeR+JXQizbAk8wq11Ro158adVce3b5eEp5J5YeuWjLU2MBP5p+M2r2WLP4Y6wkMI
XjToYYs5sOgE0knBJUVYjVbnOB25Ahyd+l8HwWigkqNXL4q6vQlv12hxs0Hl4LIB
3TTAElivhAvC1/l5BW7NvDH8lF2b39PuVNwMcxj6QymeZt4iZh5jDubciSyHJYHe
zBzP6VDUXh6H5LzG9xK+MCXO5ccj4GlEeAG9jVUtuoGqpdS2HhIRrl1Wm2OqP/bC
Y7ksHUFn4Cwkee0JdLHRcR3hugo69vw+izI040wFXqk0ZjTBKTrnwZysKJANqSmR
duJmiij6x5aKM/M205Jzyaxvf70IVesc3tPtCF7YPJVTEDRI/9/QorM8GrbY6qrX
PZxUJ66m4HDkEHUx7adHNV/LyJDJWrQbT4G5fsl+zxt5QeJQAK2xBxepwRPyaUjP
C2lWDtNs5m2qQMqcaY0h+jEEPU99GA5/SNRA6KWJ2QKS77pErGleItKE8Qrom9gY
DwiUm9Kdk60D4a+vRnVCO1MEtooWFH6uwos63z6ZfWClQFg3GQe3ogxSswMxnPay
y98qZauQ8TMzqDMFpZtxqEQmq+wnvHhuCGePDx9eTQ4FHs0mE103U6xEzlRkrhLv
4o9fV0Q+8WzhlnO6c5H54qBYJ+S6a8mvWR2lRWLd8TxT3YMKM+LSDkYVMq9VQYMy
bdE55K2m+PxYKLfok8PYjDPpDdCgfzAOXAyJ4/WAvhnxyElAJD4c+pjn/CkzbV0h
Uo2KFPvP/R91Ru3mw4LW4pzVwbS/hyeidL/8ThYZhAc7KNQeQW0NobBwNbhBOAzz
nAhHknSYJxXiSqMr0mAP9EiMXCagpE42cy2EF62TyeFGzj2ynWZKvGv5UVphPfr7
skryr7TqSSfa24vlGDmqTcPqEM+8E1ZjDIqmS0xNPyyFWDoXsqYUDPLO901M/9P0
gBA4uvFuEEiXZKx+nGbOyiIoV7FX188J8YJP5WJHryf3crmAfbyAAJRm1UGXNZDC
dFcBMOkLm+pxbBu/8OSQhP7BkYrIZ3LiVo4MjDP9n9IrhvFCROw4GHUqhDKOuMFE
eI9Iu4nIyW3NUGVxVuozCOm2qnmFuJQL6apoGQVQ228y1ODwPZkXkchJCP23wyZi
PUFN/2S0sTw1hJbQafyv8eoRQpQRftRK7bV0QR/qsfoIsxWhbLTchuLx5Rh06ymh
2Hz+iRTHqQt2zO7pR1Dy2C7CgbxmEpna+c2xuatTsswHYbsZUOrTd2OlYgJ6f9ts
fAIu14c/1Fjq8RGrIxkPJbzrMhqXP6u8BIbgK7V2zvkVmTj/M35elqHM/1pwzGe0
6EbS3mJbMaM2N/4WwOiWsCVCukSTx4armTeQqBZvnK+RrQxfYKQLL2LTljBIYBuJ
YR55mEVl2dPPP7CZC1GMIaM50AOHCQf/FkEMmE5BHYrQ9ruTQEbKqmc9tuFC8nKE
xrlC2Soq0bh8f5pLa77p1vBKLDqkcg0uzlLW3vniFjDZgWiIQT7BDeCVD1zLA+0Y
DBYgIzJoAc0Q8P/xCrIjkAiKbLhJRclDKLJvyMSg7NF/GQzjaVnFb7u0jNmooyI0
AsupF5B3RaOjwiMIZC3KQx47Dwx73dM+uAsVc2H17NAnBFvVGkDc7sFu/0HfnmDB
yE9LpNJdjQ/g+sWpyZmqQJkuIqetMqVQq+xXNlhsWzPGmDan5OD45salWecDVueM
TXA8pylDQFhOH1PksSbrUHFQxnFn2AsKX+IYWBb5J2SPJz4Czu5EeYHHelNxQ3ea
1TXw09tWYKWr8pBFKq0k9XbvTCAc3nx1dHBoyRGxWpiw9a7WSvGS+LhxocR3a26r
L7cPQaix8iwMok6rGqGTG7iEMEm1TpjN+++yvL2nynGFUv6bPFdChUjNFqZfO7uk
u38AE9GqUvZOd1KxktFSGCEORWEYYgZWtfHdxw3yB2FhjEEMN/uDF5jLJhMaXwOw
AngFYWCCQCe16yL7U17SI55+J9tey2rNqBobzGUWSxrDNPFQ4UuF76egMfE2p280
03ZALRAbeE8UWOSlwfgjxj1LavPSNtIu6leN1ZvZnkt+3TZJsK9i5RIiDJ76k8xo
FHgS59j/fjRHJigPlE+4ByQqYY1Gq6OqMQr7MeD/jxeBuHNHciI7DNBjD24WlVqf
QJDwG/qZjUCauZCzF7o/Szb8P46vHitZgK+ZUmep7RLcJ2DN3JK7lRMWe3vXwZi5
cmS+JN3DWNGdyRShhvK946m0bk1GZHpzXl7JcR1rZzmBEefYQilIewOhwOWNiMwa
KEsLDMX9V4MZA5iIzcgTdMPdZPcRXd+7D2T5EB7A7ZX0BH7hR9dyUjjUdY0N2+jV
+xaNjacynnN6FHr78mcDDzplwrR6a7KX8YpfK4g5MhLsVWzEzS/KBh/UutEW7/qX
unYLnrMzTOAKJkjirBx79l/Iuy18kFdxxmdcSG07NU7unEw0s/YZ2KpokiYwQqph
sQYEwvLGFQ40EA6gluRjQmzukFkdk9XFfHFkmekIpe/o2UgjQE4CNtSoX/+Z1O56
gqA4gTydc70wCvMOw5THo5xAo+XxTmESQJZhXvjIjXuD0KJEt5TuxONzpHG2s2hl
353DIEi3yz9UiWRdSDtlwcZw1F4bjbBxWJW1xSbwQQ/XKGD9WnXcCG2f6+e+4we7
yNgc+cDRjH0GCDUVxAoOdYgNaop62jyj2Txvyq+bbv4D6uIrI12miZ/E3qqeB+QA
GtGhhxB6x6erTL/1WhFqp7S6PRu0d7OL6OrUSruDLtfvE4sBWEZLylK3e2pzQT/P
o9uRywXnSm7xfWpVvL4IubUn3SZXhrKhjYzPzfyaEHwTULcuq6Fq7lWsffsop6h3
DRGV/8TH0GfF+pY03xwrfLCMb3a3o5B/r/JYXW+ueTec8bhMWnTGAakOLw7Mxt2u
pFp/FrRV1GQDE0Rx2294KYb9eq37bWEl5C8kcFrwdJgM61rsjcX3/PPCKK+90Jnj
hGsxWAAn/mWKmwVwlJ8CJkHL9LLwwfembc34HBhXy8GU0NDIxRNZVuQZRUMnc68Y
XbTzYjdjLWIb51I8gqBHonYiSbMYfAZRTopDShng/Nqzzr1ZO/Psex5pxz+84emQ
uCQzzQJT0vD0LloHfLwE38H4kyz1bm+Zv7DGDMhi7KjvZftHDS9wQrzjd22vTGlI
5D1jyOEnC+KJ3W8ILOAPduMfhrgADEpQhXJqUemf8hlMMMMSXKNvusOQVGKz+wtd
YlzJto6CugO2wnpR8UT3/8y7CddHz4hrpBhtetPw5eShTgU5C6tyhBHassTwtEZZ
/PtRv1vMez1iGc4dNuUrcdk11dp9rE/hMMtRV9BVMtpEs6Vf9CY3F8WRC0BhThGk
LZ3vja/4t9AWPJ2gfRPuhr1+p6jnd4DFjh0nJrjmUrzVQpL6+xNh92SMSsp/KQfn
B82FASOqHzViggZsIBIMUUCc0VFNTXsqQMcqPo1jWZ485OERdQqZUGBKyFAy57JB
eC+QxtmZ6Wo0cN+ZR4ZP/7SDxd91CE6R7njBAT/VEHEF5SIVGf5uB36I1hfQssoi
U/7bkRIBVWzUavgin/buuBHcpUybp4BNIfJjIM4SiD+tMzepFy9PCmNdFSHxh/eT
5eCtS0CWdWFw8X5osRIP2P+ROnoMI3zaocjDeEhQ6aqNB0+aakKRDg/TxyI0FIB4
ytmYmnNiyZ2TF3br6QDlQT9aF+CxK+YmyE8Tl0BRgzITRJLnozDk5gWDHnFIaL/z
lK40lLupbfha8O61tZgQa7gdgWz8hdDnfcd9hfnf+mo26P6liFJ+rEqn2rGj/alH
cerY7ARgfWKj6xLa65/ogoXf2UBGeHFVPp3r/K5tJI0q3bV89G9jDG5tXji9SbnU
eId2QNAGqOHOF8ZYeUp+COIP3uAzLmclbTT6x970xNz6DPgQR+ePh783MvmyQWPg
nUey1wZkejspzLTQfNwvktGVbQYDG0RVT4rprUD+h/SKDOQbjXXWHsJEFQgxqHSl
i5ymMTHiNm4KOSVC1tCqTa6D32rSeSI31uV8e0jjyZx55N/1kLI2DHRLBY6wZpMI
pVDKQub5+oyuII+lPQB7aQUHBqcIRuhM2pKU/u5OGXjFq7CbWlJs4A6BAtnJNgdg
12v/eU5KeNPl4OuIHHJI3eVH2TpqgBltwz2s0gNFgIXz5H2VuScXQ88yaGx1w8Op
twpTguzctvLvtn9YDhNJNiJC82XO9E1mEREpZpP3CSBpi/HEpIHkXtumPL2THWbf
Sp2kV95mY9UIZs/KL7MrPZrIshUnEEGV4bPSaAIILuaO9rsz8MLnQMLEzxYIr8VO
W4HwSnMXKcbnZYMe+uK0hmOS5mttqMrYcQuTmJFzVP+a5hgKsDKJ34tO5cLz8DAK
9pbQLow1Eytum/Wnh7syUUSZU9Ek24yzVMOSw1+HcCR+i4Y1LkwERh/rtIF3k/lu
Gc0w8SIdL4kxJ4pG3itU0QzwX5IZPkVbDkndgNQ+jiiBJlvtcIj3Pd/dBp9Xk5wT
+saumF2MWA3Ih7WthTJlDzPwVfBomm/CYSNDZ8bplWlFnmhVIgAUJWGRyWtCI1Dp
+LlQtFAGTUna8KiW++VKRXKS+UNfT/KXjHzf+Bm9+c+AXfUHXoQC3Cq4ckYNaDA0
ADS7ZX3xam67Q3KzEUX7gFO7J1kNRLO1lSOxJDg+nbVkOusTQE4ZuJWSDf5OjMYN
asdAYFxHGf4xGdrfrcEr911l/g6YVLUv+LqKWN1PNhBvKOxdPx70quZd/1kz38OR
TbffYCzVBBLASozuHSTQ3CELl6ljnOJxtytjXOQR7s8JyOljd3XPfp3Z4e0lBxjx
ms8T8CAV9EBnL4iZyoAE7lUcQZZgXb7fomt3FhJacnkUGkymMQ73abpJGfkB6jDo
iIE9lbLp+bwX4pyYMjcIUb61KeVgJQ9GMJpsy0uUD4mTYwyLuZFP+EfIuUYNo8wa
9riQRu57Uyy5HWXKcJtOQShWMs6vDHEw3HtXsYg93ozVycwFWfL4kLQI+UXUaI2N
e5qv5qob/bNZMWQeAIS/iFRRxT5N4NZVlW+g/2v7yajqtfj4HwQpuBcuoOCP+i3Y
z1rGn5E6UNhAwwk8aK4cQo5k1nuK543pocT3PBZrALohGf9P/NRqfz1yZGnjT2sJ
RbXA5SwQNXPySGaTGKsi3KkQtmJ4cos49NnTRH0cDj2TxuGEFW5nF50sgECJDaAA
QruQnpYpdKJvlaTFBjOsDfqQtt8GK+MXNV4qoT1Co1cyT66rwcyMtp3QUCd+VXz0
H07SiGcAdqAcuehLsBtL5ly8rbLcDDFoGuAEOc0ngqXX+NlvylvaeGAJeqSOrMiM
cNAlbobckDQk03B8DBeDkXIlOjUOY4v6jcK9E4RRq8kWehbyv+pwQyjsejsO2Oc/
5FTKbUiF529VoMg0cvI09o4anS+fZ6UxSsmHt8LSLTmpTSa+ywW++/9K9dbcni7I
PnmaMF7Vv0EIhhrYwxZBjJSvViHY6lPv+3MNnj13wAVDORwpKmZoRenDG6HyLbVK
/6x9nimCdxBgNsLWm4UxSLtd7dxakOlrUDVvRZ4nhIMyUvYVn9OyKHFDTtFGI+3A
HT4tWhFV2AHqsEFSw5YlqzndwDf2olG22qy+Gq22nl0VKeVV2dBcd4457hiLbcww
sSf8FID58O49QllXilv187MHx8xMGqU8xevDS8Xnfm5vQspioreBDo+nULAE+o6a
Dm8YLA9iGGLLBF167RWBNrll/mEWk/I1BlQe51dseO7xKXDSwCCWGNmqIwHCiTo9
qCzVDdmrIzJL39rpwOxjHP+/zlKK2B+5vJukft5aZZxcDnu37e0iytEttV20zFWa
+svpE6/F6+AS31G6PkLp6DJQaJY9Jh5ts/CqG9yK6PG6ZXogmDU7goosUU7X76zF
ChKncrtI/ge09AhLD7ZFfr1hIwzL+/mhtn6kKMG+hzwwT+2HGHyQQ9d12XHtP37i
Jzg1arcdhAN5k/UC4PlS2gZatOhufj5kZ+wPE5FgRF18HOTOf4ZuQJo6IhOcn5C0
FOLncEEA1PZDeV2MXEJWQ3GxQNA1RkNF/T6dt/3QyTyKA+bTQcJ4j+MLHNdifMxP
Qw1uGFUAmf8h7UIxGYTTtW10aSpBp2m3uwjnuJs6Q6vPsjmg4WjOQIcrsMoBy/nK
zOe4s6WH6fnp8qqrrAadLxgK+J4/VYw5hwkj5xp6nuCkxqqDBMwbuP7GEbma458n
bolBufa5wsYd1k8u6Lg7Cka4EKQSzFWxiZQGKWC9lzBIYMq2N/X36kC9nlsqTq+B
DmevV7EbyN7SLA2pgeUHTbgT87igxLjSErO8TGWUWuIeuYbY5k6TXPgD6P0pCZU4
ytSfmXURfraCVi+GNaEhjL3gIc0PrATZLiVnQnrpQyWFpXeCstn5ZBy4/h1W9GfL
aBejpKMLIPCm/wwM1X093ehr3pYkh4sVa21nPFUBNJAcJHwBI8AJQM30kaQD5r+4
Qa7+bBT5D7MHyyQNXJcq9BU89CklBXdtUcSTJ7Lvb5RtIXxtv36Xn5TV0XFobpAW
QZ4e/7p0TSBk4PIbe5gMDa6b3jyLIUrCP4C9+S7iIvTnvk5S/MCSWfrvwohfHO3q
uVQT6fGy4qFKW1fHbMOvYITfLk6Gz2gjf9mD5fCcgzp/FYpTvS81vNYYf1J2uTCC
2OFal3kq5wdUD1OTOqGM0eRlcrRlHn4cWClZRa5CUp+8xzAX4dEW6vrK+549dY8l
VmlZ/fwLT0FvYwBj7XhaAR5ZcV8Jek/UwqWAJF2nl/+PR0iv8QpvAZe1TfihnqY4
2j9c/cVopu7VjINB/W5sL8q8GvW7a0TyYOuVqN2Xnc4R2lWL8s2ULPKCDYC26bXt
Q1LR44u/O9WuV14VBlUh3KqHlfCvrOb0Rjlugvn3vwr9SGV5RkuZSg4YGqJp8lKk
pzOLNRuR/RedSWkjcFmnVDecxnEmfSaU520bflyoSHZurxZN3Gx5PvaZaL5d0YRi
lb7xK4IrEKfyDzlt8VoffgYHuzJuGbMpJCRotaG4wp+yWlDABmou8uNkofwq5D32
It5Uta1+BDkx6Mi50/7pKe86WrS12SRKS12nk6PM1td4SBhG4TY0X46Fk9SS5SaS
eMFbB845/2rWUttHLtRR7I700qKEt0NWh1pO3XkM067EJG0+MYKD0k34Ni8yLOpT
5VrwojJBl/jm3v2eU+sKOPl6EtnjP5MO2iTGdsbEEu8cDtsztIOmre1J3Q3eIY9A
ID+3ErCCrWhhzgpU2lw68yOpSk/t9lwyNXS35Af4IMvL0dBnKUaUHO6ox9/sVGRv
Un83Qskofttt9INpQ3kz0c4LsOPaaYdbLWLbhoOSaSek0CMoAAIpJuNLmw04PkcD
OsXyZxiQHPXWAWaxhWNfeoKPo3S7IWkqznKXxDl1kWhaAvS1sjUyDWaLNNg4NY7C
aBTLZjp0X6Fwputjn/Ta/7x6kEK3dujC+KMrqq3IDA+7GdItbA73yd+WFZkVGqTQ
SihztxEas0XeNUruz71iuzv1BdFYtMysrgtGMiBEgzR2LGhgCC8eQhEytzK9aO4Q
1vKn2E9AKfJMP9N1fkUz0h0LGkNQ5ZEatM7lJFC9fPEnGXn6OgLEbE7h9Oy+KfWe
2PBYLMulmDzBqY0lMq2Y03heASg3Ef/+BFgWNd43lhMCx0vBHFuwiz0xjcCC+iLZ
N0sgoR0lI0LsJ4Zm2qLN+L6i5bBF4UXoYGR7G6cvswoeyK4+NB/+B60Scbj7UzYi
pCY5e9bANYe8DRlSL5J52lI4Z+FjjvVS8CmpnCIuA2uM1Fl5AmR7nqZzxAQe2Kwo
t5Bs41Tbc+JgJkWZwvRcXbQGHcn9PCeLgJJhZfhZoGplD/5OP43xF3S2ZclszTpu
cWbbj1FAbD/CI0b6FJPtfJUy6NMACLgNTFDp/6I6rJpkDYuFC3uRkUF61jAxkSqG
/F90Opgsfa4BHJ3g4ZoFXlUKMZJdDxIDyMlq1sU+8HcfhddEnC3ghAguL9/GCyfE
5dwDoRqiIWgLtaViJUTnAAfW08dS6/e+uviYNUvoUw19Ej9Toe3UgzzxSbyg7sxH
FS0Mh4jyyztAphV+DCutFbKtkfI1iqWg7dTxW/7HdwnnsWszmRzOLueHKKK3ldrj
Vo4zXEhGrpVwOEwJH1+f9LWi8J558HeW+fm6feUd6REFuvnYQubs01I7K8sXovHU
KgFYLZonlFpyyNz+YSwdDz7EUfQ34DNgJvmAgh9WVxGHQ9x8JwBcJ/P4Qu7YuHh6
XkMqtJ00TzC+ol5WKrUBi36eTM332lavNNmhni2BsFjpVt5VuEL53wbzZYBwa583
8Pr4sacJKfACzXxtOwueE/4Kl9IoSZBXSqDYoDr/6yhzyWhMHTTPWFvK5YO0llil
cf80d2xwXP8FjI1kl8RVKtHi4tf9Q7FCCGBSW9PwrhA8nA/d2E61Fj1u0365y1Vj
GGzc9YwvGAfXVxFjGhnTBV9U+ejLGRZtylluYblALjF2shZsZ2bjFB/OLACc5nZe
XDXWk2glpuk/IkhQWd/VAezOeE63kqCWc1yX00Sr097AQNNSXuFhq8zEFdHahtJR
i1iUV71AaYPZ3eeg2pRpwJdisTj/+4PV385tYQREE1F6yKGw78S2zxrJWgOJbS5p
qUMoC2n3rTihyskJHreSfNe0NscaZtA357ndcpvXyzDPP9y0/PsmTCUolV03mXrk
At5GZSS9mCu85iwbIKVIH1RORgfCkbXZharMjhr5mFiZqWDsyyqX5oLnu7hBnEls
SjFeKAqWm8xIobliILojqg9J0GDdPwn4doUk2xF58eFo4T6vEllQncNidFTUz5Io
3SCAW9zHRkyNhtDVQh+7Tpok5q+TzY6KwoYUh2L03ruSWgATpvrF1EltY3s0poBy
AZ7K0ROsLef/cldbQuTZVlcyK7uzvwnPNQ6kzMblPP1As/sFdaLksjzyQ1PYy4Ba
GinMLegYFl8czsjtVQNf2R9K+sx+uH7Ud8xgELZ1v8FwVxH9V8dSqdKVpFTbQr9i
H5olN7WIwfy/W6GzrmJPJH15AwAYOselLkbsKZ3EvuR+jTmkSUarwyV9Ecr0nBIT
D47WjA1xAYAP7KQfWpYQjsowgPbiDK0J0oL/lSDYFQMzGJSdzmK0MJNjYkgGdNHi
uTjUJNodGuPMe142MPg1NBn/0ux6DMKcskIMp6xhJ8pfBq4WU8PrrPwLg6fVLdpe
4/wz24BxqSFMiVAiLVHtmHovN2/BDXHtRYXvudcfouzJueidMfe9v9u1Y9uQCwDk
B4M2CL+lcEgmHJI+rrDI5UjZ0hEQJuuaMe3NNRnmzu9kzJGCbDXS5c+vCV57Na6y
6jizrsuFERMusTRp6RD3Scn4tvgL7RBSqs43YkRp5QWGIaJbtUAmQlF9v3xAWOc+
r4aRzr3ZkEDTwwNcCII+rwNc/pLHb8FO74FUxvLrn7e4rwUB0M7QLCDxyKW3pN2o
1jzUEDVIKTS82S+xg0qJPd9jOe0KSu9LhoMMvfD8tQ+0m67FpDZgJGKkSMA55H9l
NGI2T0MnQKjc1lW8ysRYxvz7me7HNTzNSRXW3e7Lry+fVxR3zLxf8Nzj61JTyzLm
P1+2BdueRRBDw0u8cANmBOrMmXs9QHS9HZv3UQVOY9EpalwBb7pO4IAcx5cCDCjW
BcH2DuH2PZKj6PFJN3xcmr+KWV55dGGVUfr5rT5E3GXZW/IgHviOUiM0GcfGYEIb
5nnzxOT0Y2DqnEXhWNtuTAK55ahialaHJGzIsgzGHjXoKzlXzpoiZaHrNfcLElG6
EsjJwapkfQqLeXtYNIUvEZ3N58NV0MGY/xTT8ppM1Fuxh4V0BhRbLh/v5cMbTqH6
4KU+73WpacSzVkTQUBzXHNzMuj+JjlQubKZ7xnpA1lVc/ovPcV1YLlnthvSZ/vmb
9VeSO/u2RXokShQbqyd7P6XfmPri9+tN4DkBbW5WEmKM4WktqX6ns4zlLWf/XxEE
Q1EY9YsPt63md6B88leJ9jQmIxwfBh+5np0zrSQrir0ssKZvXwgvg/8NcL6riy7f
7Lm4RPN4kNQCwHA1tQXZPwjbqQdzjRx6grR7xdgHCGxOugtWrKjPOXltg39Mg4UJ
8y1psN9Mat/g8woniGUh1QNIka6itLMmc9FA1Wm8njTDW6mfoU5q35LH2bDy+10i
tUGrewwevuwQLwqOPHExIf+PdxC57ZavjBB//l59CxqT0isrM4NUFpxUtmwdvjn5
67TnwQP3CzV0aCObjHHRlqbNIrJIT2XlqYRAltlquwzYj6qpfg8lOXbgfHc1YR8X
FQuuUYI7y78Ws48wYpbe6PiH0XTU8a7wG61whbgptGF2u80wBbVw+w4BSroU9Uk+
fqIEi+IMiXYopEIPAxczr0qIZ5ZtAiJJpEOINliCP4HhX1XKz/fUe7UPp1paKSch
m891DXJGTj4yCojYARVNfVCCNB006bnHKaAh+ILOzELMkAN7pzXS/Q9HxXqtsIr9
271JONpLRQXDXIPEJtbZb7LAKrw2VX0Xnyq/nF/bCnvl1bf5XdMwYqaoeJoOVF99
lnyrVlTES+VkbC4p89KhX6rNFn123zqMglbQYxIOyxRXaABbsqhF0CPcZNyedC3H
L2pAVAMYI1vyT8tfe8MyOHG1td3je8PoGzYdrRGHn3DFZBJLb2L+S/k2SUMTg1ZW
E3Pp5OkV2czyY7Z6l1iGPdaAROxDobbUfLRuSAHA/C4P1hkEbtnHv0BAX9exCqom
vl6Ya/gCX+E7K3/cfZMsIBax9z4rHjEc3gH1E9So/0HF3QNO6s4fwgyZENKJmqaw
JZIX2BbPKfyPfzwZLgBlXO7/PmTlQMQiYg/H2zsIDlBxbcWG606tmLHXRg5OXYbP
zZWAqlLiMIOScBqu2fEVNxZbB4uvlJWHUwGBIs7PyMUCTs66kkjsulXJ6/QktFlf
MX9yIR0deM8gf8MwZEtSWZrEuqQRM4UVi1g5Eq4YzivBnPJGtLXdZRabyRf+lUtr
qJHBXwf3As/MbKjhHp4WMUaTghnNXPZCXxHCdX9aiJaKxXDdFn+fjjZaLnNwHpHL
lr2I/dP4MDUV1UC2QmI7V2WurVW/YI4iuh5KtMHBHwELJFJ8HaXxNj6GI0BhgLA/
YjE1S5HtQEbdLgRiOQxoV0TNZ3udpXlfIVRa9huocDBg4PwQwxNNtqy3sK7Eb9h/
8mNSuZ6l9P2VOhncRqxiT6RRbw9/DAMQHlN+8xKgQis6pNUR1tpJTqS2tLV/eO8D
WPPbjCgPhL42DX+MeWvk9B4zGwelufJLFA9GQ7f/GNCgGk1Rg0x0M/qe7RK0bl7L
PKv2Zws8CeIC8GLHdb3BOsUBxXGA3DDCoQMPPRa93V/5Hj6qvfj63diK9gnkHIfT
C904K4HoyG+bfei3+cro5x2RJjyiw7dkkLUA/kMjdvfr2i7l6l66CTCUzakJOy8P
MlwhGDvUxnjzB7m9aX3kj4HPYpIZ23BcZMKZ9DG1tBgDYjt1ZT44taRdWUZfaE9o
HX6DAnz3hOMdNXZrs1htP3O8Gdko5MASqg95kC4SYtq2S8/bWrhPM5QWiLG5NtCp
c3lX41It1MtGOkk3CzvfVuPLseYjhJVa89Fnn6uxtlXig5g/M7DnEpqJYF/PgW43
OgzaQ7dd1uuYOOfc68cVV/rutTlG36iAa/1C/7/5p5u79oS11lw5huwCydWd45iF
pP9HlCH1ezDn+JPN7gZ7OcyTIvB6M2AUkS4c8ttte+/5SnK5EO96j1vzpbWQ4t6t
r6ISogvq9T+2D12fAUfsn/D4pK8evkfwLHnOausgeKeFas2ZH/wysyvAF8GF0CrA
+cPsvZmpV9xOLOm8kxEvs4btTAFD3TGOMiXR/CKAXBTVJ/M5bmw3QyPb7Sr9fvdK
v6DNELIHzthh7OeOoyfdx5yAGC6/A80ycMfEikbbsJiYG0gzg6HsZO92sHlgAO0/
QtOx15EkPP8DiqHbbyeg390BpWffuusliMeNSbxyDgoLHdtlc5N9sZOUMm4FA6XO
5FShWMo8tCrTCgLu4rhJI2MRjjxCZrGFFPxK9LHp+9JG2LgK+atVURKLxgZZmVDj
vnevjFsth93E5Ty9WjnZ3Dr60lf6YTZZR9kWpsJWcysYWl+KjOf7pDERnQxhTwdq
oB1FoaGpGmna4r741BRjcsqC8rTHLt/85+lLu0gzZgTgCeWzcCTsPB+g1m8WIfMf
NRCzxIdaHVnv0sDOuh4JponNL9+D4Jy+LzSShsf+pAMPelhF7Q3+b7S3muYbckzS
pep5MdxogZlDci5Qy+KRmIm57S4KR/alzwhsHNJV24zk0PC+9ncTZI2UgK0Djz3k
X7LWQHIcgYP84I/mQ5btu5n1K/CID1AZnYa00/qQY/FgwEAwdL/6g+dGZJK1TEzX
aUVdjZZBSo9kWE6mTEv0yGa7vvCT192bXS68zqOUoRSaYhtsl1dRXxDOzx/QGpjm
Hxp6E1mukBZ5NRwe0THHtGBLPWOvBi9vY8EizOZ2wakpdoPPEHsUxrPWvj9A+Hvp
yBvXpFJSfbZpmMD2Ld2hssaHZL3VtzqEBuzvm84wdvPNj4wcmi4gTLvEd4h3ER3E
lXrQBkPJkJkmDiTHjxRyc9pEjW49XIzPAEtankdS5UF/A5vzm+L9hNBwJzuZoIpk
tr/vobwgDmTQiKJdOsDp44+QxeYhRDy+dTr1CWwKJgnAZZVPF6ORb9uhBzAImTyz
Cd3gmSkEG7WpWpHi7Px9Nln2Lrz8GvZL/X5msBvWT2xxuTbqipWrNSahxYfAn0zw
bGY38SFpK9uLA3w909/pxFTyqTr0rCEdeMAjAqKVpHmpmJE0YKWCYCTc35tG16rO
pA3kcvDadmYSz5f/B8i6SGtUlf5xWXAotPZ9W+kjqai49IRQpZNZgWpzclVVgqYo
eq9YRT2hAbnBjCCQeZ+/BHOR9TQQ5nxXnC0X09fee2hlPtpEvPKUJGIXklmTW129
v0kW4gIjGnXchy/DaLz5iPfI3BqvYPBMXTuSB4EhHUWrLiQClKW5yg5df11gxYRY
j7zJCPIhRUN+BH70bCKcKwZ7X/FWTX7/tj48vYpZiG5SGA2gZB+ysY9SRBPFyukS
b4NdX52xU7zECOX93X1Ysr7GeDy12X7V8EmLorU+WzqZkdrtLf72XItqemhfohpd
Fch0nK3a5ulqbomWD4H5FeJ6Y9RuM/A+69uZxJVHns8sLwW/7eU+coDjmlt2ycOV
6+/O2RLM34hYym3oDtrcbEXlOU+Juei6IZXCygBO2FYMwXCd6jAp/HRwb3JjY9jg
GQgZ1dwai1j0sEU964V0ILzLxOtq2yu5yfdmhwE6adacPv+FdjmhpZzP3/JjTUGk
ApcFcwJ9wadVdcckxOjSSIo/h+/mWcuAbQQkpf8/zDe1RDpM/VDLEkIrdyf27oRv
zjtbrfPqLUfDjOAvlsLnPMt/qWbfg2896nYyvNVW+vs/RZ7GXUgCOghZm36qXbwl
NRtzDyWCGhq1fBusguAs6bF2DVRGM1uPkjpapAbtOSKzTYrPKhtCEdRGwSG/1Agg
NNFbCbp+/zAPqP1VZK0g+hV7MzaJNUzIV+HmiJWVtWyjqD9cicz/Za5cee73vNkt
S3z4oOye+dK7f9iS7t5eVppffpyyRMUhGNIiDcBF294oyER65CMOCwIxP7pcxSeC
f6Lpjcp4GDZipCULM0oNKG1zlCvlU1VWJsluX1h8wVeAp6W3IuLj6PbUX/MC5lGd
VWQgxyA9xJpPP2tjefi5+pL12Cc8hZ4nbcepzCFUSf+6OTov/ChzyrmZsU+SgFVJ
wCrJ40Z8HMZr0IV+AE3ycxM0B++tVgQShZXgN2uI3X9TSuBl13suz9AULB8D8P12
5Dxcg+1hIARuqOFtdrGZEs9j8NXWhrrlRwQNcDWlvWLQgbbZRGU24HmVXGuLXmD9
CIg+uZDy7NZm5vrIXnMtCB4Jb5N5bDV5ejyRf2ldrzartragv1c/hEyOTcrYo0pQ
e8YKOtK4SyA/OA6XAKZK4pMXkniu2gPuHlXfLzvulrfuiQRH0qKlE4GgvJSTxbR/
e28pJTBmIS43OsVbKcyGlDaQE3cLJHzLzQeV1gYl9OnUSG41R9KI5RSNcOIdeUjO
hhCXh4hIebZqozbTqJVSBzbL23XbQ7/h0bIBWe5N3wbX5xKJ5LvSwFhMkgpCOjfq
EaR2ArcPXFhy4oTpTaxdKJ8YUMxOGASNw1bcmCk8hajjgEGVIEsMzcsUCPi7Spa7
la9rcnVUytsd46PUr50v2ZmSQUwsSjMUD/fvW4rOdim343MDFqUMPrNnkJlX9m/5
E4ku9pSlDo9spjWkN9p4HzHHcybWFkF59Hh7AiwzafgKPA0RdtDeGDZ6RMl11X1X
7+JdXrCJdTdXzUyILYtffRRWBZwLdfp/w0zefvKckU7UXUXDBagU0UbD9mSgo+Jx
/hH4qa3f9rpQrHLE6fdvPJZoaWhjEsh67Sr0Heaz7kpdicPLscEy+QYJHMHbssFs
Q285nBtTMzstT+i73N58L4A7VAOIo+rnP6vxRKBbgJaSGRZs29LtFDzjJxAcKHhA
9VrSP2Pc+mVj1Ht7nh6qwX0ndYggmhqY+U54hLPvWC2uA9WMudeKPaQjD4fsiW4T
SEx2apdZQbg0RaigpOAzFm8ZpZXWXUa0kN3WsIFFSodXp6i+7HxRIh58LzpIfw+0
fMQVwtun6QUTSauKtKwslECMPkDY8ROaAYZn0ip7dYTmwm1aYFTvMkF/22FhO2S4
JM/p0KJddtxJDHGsvq0CIZnTapua4k26P+C9QD0G/TP4TeQddWFXo4VkPT5AAWqQ
Rr58Roy9B0aFYnP9P0d5vGazSAdcb3h2tsgYGTOeppy3o4RH1bwL7JNJK8oTsgQ7
Gdwr9QUuWe+HlI3NAEpeu/1d0UePmJrfHneWnEC6nb9BQ8vxHBIXRNnBK5eyarju
Oqjb8oLoQj5Nkpiu4iXVF6jy3T1MMsLt0dR++1O3yImAWhR2L0cMHKSyzrPvIMsp
f6lv3g5jkhUw+J7U/FgvPucuzse/h2KPAnuKkx0oaKpZ1XkpOq3Sg/L67MA5Oj4J
pZz8Ulw1OLI9mJyVrwCaqvNzEIJgqtoRiszpCcc9xQNcI++niM8pgcx3uaPKCXBF
O8veqpgj5wLFM74yWKcylfHAYFBoZIiKIO0aZikK0GD20EE2WhNfqhswLV/mYv27
+kjs7KyzzZATZRJYKFVuMpcViOXqyYiQHSzfkBzoMLi3vs3ymTARtFiPJsWVazny
Z0HdP3mF+pwPSiCCEGBWK4+jAqC++k0rTRt8EZteGe7GOjnC8JYPxqxqYV6bCdXX
KLOn3pFE7FpzKgCnwdAUMbJZ06yt67xhjkWda2d6I7nVNsFFIjSr3ZnsETeJXz3K
Me95Dv97bLnBh0ZMUgCxGQW7umy1HyW/LBoxu9D5LKIiyiGoicQqCV0bgXRQDWkM
E7JYh7Eee0AgqByEL2QKfnbVCji2pXX5nkEaAHVJiVhYWYAG2ZZnSfO+6oFYkbSv
5jc0VBzSPW7ZwAcwwVHWra2XixOqOgMG8ve3a1JR1IVJxRMMcZM4P1pBttgAWAL0
63QzIjxHNe2tgKLzBV7R8ApsRi1Jq4Jaa7oGQoi+7cDzb69gQdgYbIetpUDKS61B
l73BFk/qGsd24z4g9Rq5d++uma9b1tktH4oqG4HYOAe6q363zuzyh7Hn+L6S+To9
/J4j/Oidp5/gcC0M6AnoNCE3XJXq9q7VOEGTF7VH/9G9Ku7hL22k3kcOqBsAMDl2
PSRPzhzqH3l0T3vM/egZTUuorbVVcE98j1mzJtVPLbc0Hn/Ft+FJf3AvnSqRwgve
2nMp1hZ3trLY0A9+gCJVMManJxJ4PZCGyVLEM4EjFpW7yM8e8b8qYMDHLRHfjwHn
F889hSxx2X3H36mZgZzmywbwAUvFQcNlN7hf1dXCy/FJnF5ZD1sm9AVnq7waZ//V
BsC7q1DIjXHPB3llcyAVmpBFI/CxnMmfUCHch9jRPwa1F6gW8C1AxK1o/Q4OGxLC
vJ0Fl+jECEzIQ6PW5QS6Layn0vRUVOPnyd2jlydqDItbKj4bUVjV0yww7daXThkr
DJTBSBtH08+uC98AsyxM3SBSAfhPbWp0c48K4Lcf/sGNanXIO189tsLWcStNohq5
fimXJnIpcKkFmoDQJchqbKlnGU0kF6ut6m2zHEbvfT+vyNANjvPfE1Sla6QStRnK
cYECertrFw4nlFZqNsddC8kPqYFKy5WvYLVDvYQb5L5MUt9Ofh0p7KEV0LoY7cU8
T3WfCOtpMTFQqN5NA6ZMoEHDBiR5LdsJL6THWqiG3PBxngC3D1bq00YrJuBjrmGY
o6a8owSLEvYxSWlU9vmhphsd3rYXdgZePskssqeaNUJjGqmHJcfVGfmJ+hW0GpGb
wr77p1tlmabNbQX3Xw9O0yjSFt0mVJ2bDdfrYyyRc8xbgwxGhqMhpIpPsch/auRe
3PGMtvwITx6RlSyu/XlVmQpkDjN2vIL0ZAveihesdAJu0Qq0uSEVGRnaRNcC3AvI
zYPXJp02p5UxlKoVBFmLQgC5zWfjDoOjbVcomguL3OpifjlP0woW0PXSKjqsDqzt
AsX6RePy+XYl5eghThqmNAdWhz5tS7k8YhEG7npvNbzbhDH6vIwZt4y/kYjdxWJL
0qv+NdtLebQZOCWDn0LvJA92/g+LJvuwZ1yr131NKAX7QZYuvR6j5GBE5X2v+gML
wuD3WA3jns2Cva383A4Z258RNQrvbfntuytShgIjVijwi4uATBhqresYww7Dvub7
bVUQUsE2cf1+ixBMlNyKJhd3dGyGw74bC9wSRKoDfI6KaNc5rOu7mdlFdIRNPwlw
ZqCgkXl17kKgPxRTAGDtrLShoT2P6hM8iNLKcMXww3QYkBiMXpL4ZUs5Qx9TW/QO
LHAjRQpZDIobrgTDdlyqTJeS0BqxFbSE/qJ66yAQ3w+awNzc+An1RwMAzu3T+O/Z
EUOxcYzYMxHI3rDrPwNtr1TjVZiM4P4yV3VA6tMQ5rwoczigu4JEe79XovaIloly
t74wREIZYK1EXA4lZcFnMpmolelVL+r2YniwfUbcusIigIuKlDIXYkxv8UJ/X/rM
HLmvKTlTHsaa4R7J83CZoJZTJcexbt5vaGYmJOzZzn8u5iZAmnszNN+ir4AbEN+7
O8eLt+URosIy2jlLrN9J/tl1acyLS/9Jm6MN/t3y06p7Vcrl0wu6oKLuloXc6VYQ
BU+XJO25uKW94JwSLlUsrYHJgFs+5wsZgT070XQ6Z9wc9Tu95hZBCRBp63I2D7G3
+8VgCmdoGwEJhevmG5dPG6rhrj1Y5wR9l0u9Shn32HP7ydou01tbSNZTtII5iY2O
6zsyBoSXY0O0Uz/Icep7HYrPbU+cxHr449LKbCTgtgZYUN0dqYY5mcSdvAxTuLtK
oOg/ZIO82Kkw1TTMNIfOjJL5dAuJKZulSC9rmLR9Wd0vEcT2mwA4C+/+0KR66Rvh
NPjrsBbpXgNeMy+kYKJJXv+wc/Lz4w2jjWYbtkQi1V11h7ueyDZLYxJiRsqxOek6
LDVLwfdpGJL5cXFnJPaIPt/ieafxt+aCVfLX/5ZvU+YmWXk+RRBrJgvvku8r+2Dh
WvJapnl4PsZhiwmhm857jZf25O6i6DA+jIhTo4Z4QNDV8fKKusWtAht3pYPYrQr0
qkoE3egh3a2AsxQt6E0kxN7tx27fdoASBNZKjVIMOWpuCf/Gxv6LmWpbYiTq1+pT
Jn1ccprH0TUtWQdFvabT+cyTAKzXo5ZUQoO1uW8UThlYfsZliRWmCDRIVf0zn2z9
ezZRnJpA1ODA5++i+P9i6LcHcBAsnmpG418jcy5EylXbsyaP5WUUcjCdgdk0/ScA
dUXQmFB49VK+hBvPHogdLE9aXHPctgUnENvKftmUg7VE7um3Fv7EhQHBCFC/Dlqi
Mg6/1Qzysm91VPaNb2O1NHqvTv4M9qunqESu9+NZz6dlsw8nbBP+eaS5JJ45gUmR
/7vjTrEqBQsNkU0Ku24M5ceMZEurKsOvMZyrVFE2PkG88dvE0batUyey6eqWA5iY
0nKv0G4+i6WiHMwnp0vG3g4yneet90fuQxmsMBEzt5cQfDhQmj167zRPUsBWi+3D
w9K8dpDaOAE+XblfI6bgLWEzHvcWdBSuXJVadzw6+c7lBdQhinpOLd+2Pd10Ej+C
LwmEamcXgcyTpZHlNlL/k9uvm4Pjo+4vKo5l/lJa4/LDmdTYwGZP1TK3NfTodfEv
nVjotCkxDaxcrwNG4DVtfZ/6GZST7GycMwPi9xbt7p+gOBUXhvuPTTS2ht7kQ8b/
gBEbqpCKyal8O8/tzcMKXd90Wf5uLL6cbrstCpqaeZvqx/NgTHkRXvjBUYr2jMqw
AXPekEa0DWqh3p6bCA8lIQSywlhUthZ6xbwhpwplRk62DIR6oCWZh/A1B2p8w6yW
KQn/kgYDFY+28jYnkSFWoH22DgTWZdz2gI3hrufRi2TsyutK/wMWuQDKtdKB86e5
W4bSPIFYI0oapcfnIU4DR29cGtgQzqSJ7akl7+MXROn1XawgPlK5Nwq5Id5EpndY
Js7aZxpiq2EfF2BnXDMiQvhBMfYi294pIviOCz2NdTq0wU0IgPdCK+HZnvIbkaDq
YA6cf3gfm+HN8bLYIKlWi7hcZoYSbSKSy3mByvYPXyneAN0uUsJicJDBn2yaKrbU
PUcPtpi9T2B/PBwrE7przRsMexg3+cP7ZSG4L8EFu4xAxfBeiGIyPUwXy1rwAVnA
UzvQfBAwU8KhUhYOgK6tO9t2rtjbXZlyLvkyUILAiN8h0df8btzJmtgq2/mlFc9+
RoT1sY1aPw/VdPG2bl2ysfx+WX2jMY1LvoQQ4RvyLcn1evDjodeJmPVhZ7EJRm+e
8NYruok/5oAi96iIMT8reBzAD/PzP/K90XK4Iz2sL0H4Mwzr/7fxT8e08SPoDTeH
PC/VhVa3W5Sh2FW1bIKr+P6iA13aBE/UxZEnNasxTiVS3qG3A3O4NoA1VEAEHL8l
Mr3HNhFHNNAHi8PAxHYbUhaup0j0XCdyqUbbykQctbxF5Ub4jgtCOlrRZowXTo4y
RCb/dg/BeZhWXOR31iIICDeu0FqnmLEYZQj7ZJpukvXhm0m16+1StIEkZhd+brLS
qEJm/xbnzXSzT9I8yNDj/G+qZxhxgqTUJ19rcXxtSYwDnjRFTDJIG9oF6GGLSFSk
oV1g7zUPUdijZIhVdIE2NsPFx8Ii51gwzRYuCqrkpgp7pGvUGFRps+AUytxSv6dp
JtBXbqHiKD5lwmo4Mn43+EJbnqsCueYVd8u6fahrcm+rlFHcFzCZeT8QPKjDundB
gOQ+/zX6hRJzgH48hoxJT8zoKCNL3vEalHwQQtuGcBYAworfcP/fL+7Xiqj4Ga2R
V2M2MAHnKmfPvzjDoUMDRCzvB0RxKaoVIlEERQk9HIPjwg2p831x72nG7i2iFGgK
mCd0bF5kLAN4wE8EB+xO7w8VMgk16g+pRb0I7QQYYBIKCvi61GvWklVfmDFHwvkF
+2D8UA8xLxyI7Ubeouamc6RIFocr8mqMPf99bPaKPG/0q7dG1+cgy0vcOuDsTiRz
Dq2BVG7V9WUNgq93A9xoB8t99qZ7RZcA14rD92TlUrspWjHAakTHdU68E8EeBx8j
GX18WFVif9T7ze9JzWnFVkGcLdl5wUcmei26/nwPbpJ4s3AqEF8r1Raxvfr+kkM/
Z2AN1PC5i4v15g1y+mrJioa9UZ6ZCspMMVT9pWYO3usLUkuMlgpHVCvvFFFYg0yq
8UO1CtUYK9NTIr0uYulDwur87kXU7I0uv9FsE20eUo7vguKFOMXrYa2AnQ8Mnp+1
V7nRSm+7UZBG30KUHNagkpIZnS1onnemmzoe/PURKNusswWYBFAabolYkvQ/O3DI
i//994WkbS1rV+lqoAIbmS0bm8Z9OYbICy5lOQOP/A0h9DgLZs2higl4gN9x99h/
Dzqssr9jaTX50WE0PBU2JQ/DdHRPJGrfidG0Ij/rUkDXIwRsfqR2V2LBMYCokh/J
EdJjiB0TzKelRW19Bxv7cU0n+EHnWtvs+uKXYue1do7eyA8eIyRaCEfvruXNENpN
uZzeDiNO47lxiz8x3/z9YS3afoGCEsCeuZdl/xPox5OneR+ITsW2p5Xfk7nzSnYu
iUWWHotV2I1sVV5xAce/6EaqmDB7xyqmW6E6hcdcCmhCgHvWcMBR7i1PT+BZ7fTs
HGQS1T75i3G6utQtHfITu9is3PzdIOkiyUkxmPXC6HQLkGDCwdosq6pUK+IvW+z6
gEo5kzmMjcZLcQROaUKGk6D8p3Mh4SR49eaT7zESp8xthxsqBg9rUBUUjf0aNzvF
0ngK6A//4HtFx064YVxkgw+vphVeBQ3DJQKmc9Pxu4JgKqnYyQoL7rBQ37Wbmx/l
r6sApUxVc8LLgZZBJ3AJ0yshajZqYh9kuhbeBVuGUQ1f0SBcThiuqktGXh1X5Ae7
1yBnK3uPVx+/c+2iNij8yKH8UHXdzi2ozdJ7o8NXdttezc/LQ4bHAetYJyBENSqg
AE0zYLgE0xrksuKgPeQoOyY+tHD2Fq0lV8mIVqjelcgmm2RpjPoPwak2CR2oe0xG
Z/jeako2CRwmNOkey9hPjvyT62rg9WyUzTeEEzXmYilkimjLVGHbkYF0sc72XDQ1
Nc+pjRwYxzIuNtpWv/s29Z6kdo7ihoNETlIBRl0sIq2oWpyeTRF4FB5ooqp+ePOC
fDvH8Yo+9Sto7smbe5898DimzM8G8GcH2qX0jGQZbAJqg7cbWiQCGdMjyK/PfZh6
U4N5ZbCU9pet1mcYBxHEHt/OTysdscX/VX9QC+FEi/bVfFD0Bh1jbgRc+oPgLZEN
tGS9DM0Rsn9yxQnkQi30nV4iseKSnu7eh+VFOoJ2pxdih5/Yb2ttpUJrkQYMhile
W89Uihgod2YI8AqUvhBaRVKogt2avaVkCwdq7krEIOThukJeKmBzgA2Ed+wASeDE
4C+zTvh/lSBY/fps0V4KWNI9akT5KF55vULLZpTn67jKEGA0Q4xhAr7GxNM2aDuY
nzH0D//Gz68c4D1TZNdUoYtX00hc3i9bPFhDP56gjyfgQ+wYKMBNGBHk5o7PeX5D
plJg824oRfFES9erKUNWmcBLsm1XujLVu1G58HBhnuL6z+jpk95lV1ju9vbumVdX
lympYPDw3WPRBDeZJV1KcdZluRWEQ+4OTMw2y4SNoDevqFq9XF27omuPWJz/q6bD
e8E3jiQr2TB1SKadABDm6tBuopzFdILceC2JUBCEWFeN//Ge2HdTSbnYI+m+nAEw
u3HUR60eOXcJLYpwZUOGgf6VD09HWnmC6+WVS3iuNr45sOcaC2EwvgLqTjz2Tjr2
UFxhEQWrl0hvakQfm306jggohLNmGNBRGc2t2F284w5pJ6BfLfGr5cLhEss8AL13
r9vTqKBOSie8RzgPORZGkeALa0dap94Ki6QXgLXOFD6Te3yuwcsaiQEc3TSGXemA
73Of5625905nV9lNdWpS9xWR2Hz9ral5Xd41wMJQ56HNRXfIlNZD3O2vaZWq00nQ
DdCHhEGvqZtPADg18zYSHD/Az9OfocwOWojL4S/8FNR2uiJuGfx/DlGThvJcu3EI
KOd4QhtxtpmYvBvP+jjjib7X4rjK9XthirUOlJZldaWBi5eWOB5reFN6PEYg6fCT
CvUSmxxSqNvk68llygIAlTsMsdi+gSWLGUp8sOGV506qZuOP3dq4OAprQjevTsOB
Bktw7SlJjIoW6qKevYpGpuJ48cOETudsGugWduvLanmWG7Xh5fAbfxMU5MP8jyEH
Olv7Q7eQ76s+NzaM05n3IOnRNhkZqDgdsWXFhwlbO3CwnLWYFUSxLRui9N2fm0Sd
Bu/bnKIw9IvuiMqSCyL32vfTaWux5F0oZ1+NCZQo5E1aY3tgP4qBglS4flvVri4x
NdOK2Mdbmt1CDYVNB68IyYaQqgXZAtLkN/zlQ3P08hhNEmtbQYomVkrFdBsRSpjU
f1lHm77L6PqKhf8i4EhriepE9MJvbhxJM2IaycFpcI7+beFPGkYyd0IPmOMFeLaa
PSqTHl1HpI7CUyeFN8+sCsI1ZSeDj6eh32OCy01f7Sb/Bg7DMsGKGQQtzup8TXE6
dlfxJFH4eC7UxargRaHsl3K88Nv6AqWOuaY8gMh6XqQJaED3MX5b7mNEchjja7NG
kR4QNGzdOp/R2B3nBYdVP3SXFwvVR6P0wkrEgF0++gkR5+RtNCIuTkwbIOaPIlnd
LcTG01RVnPBgTey/bJhLK5uGz5ECf+NmJQHdTB3O2QFcQxlgKT5sLnMqqlXSpVHC
4rqnqJEchVhxL24Lo0v0paYodmUljP/tNxGwSdB+KhAukOb4wOBackLbZ4YriMrG
WQ4vNv7qzXDin6VQDa9oWnr4uUtmgfqyqaQnoVQqXp3wRrsPUEdrTu0/tb2YapZB
I6Y4x2Njt0LVtBjupyUsHrmzXdug5cnnZvgXPNOi88ByhmXg+QsJFfhFMnmb27aA
QA/w8ZYbSdg7tgigBGXUEs+WDWLPaprL0v+sI1U3CqW3KnJYcwqwBdFEbpeshDme
nqbgKOWkKobs3hfqUjHi4fuIUJ8JksK39quVtTXLktVjHkFdO5epLwyRm2S7Swmk
5H4cNT0IPVNZWmNs6KHEuaON/TDGHnwNDnAfmyaYiCZXBgg675FPZ7Osm+cpglYi
qWLyaP0aqyRoHCRI16zK0rl3WRi3BCLilZcmA2Mf7cXXi2NWmkGB08CdOsCaMTXL
4MLRBmwH2eSC3UnVadvCBuLh+MHLnQHV8JkXZYCs5r3KkiwYJgfnnu1fJ9/xtGGT
8izDfi9tx3wQsmXPyysmLuZrqBB38YLeI/WvL+AnX0nsES4NZoZ+f4o6gCMdVUkv
RTp8fOTpp5K35n/Rv7PXNrHBjB7y8QCLX9syTaibmWpDBuMy3NLlh+qhUAj9GNYy
1yLzg+uiZLSSSC6cslFIR6viGCEMiTJdGMN0eHZaD33XxyaAnmNGA5fQTmDrqR+z
C7MGjKr01ofDsymyRvB5snVCKNQoFWQNznilrme3WqQtxWUozttfSDqkvYYPLDQX
3GS5w4gpeTXqTQme43vRju7ado/P7/9QeAJoMJASpdcezNH7O4dNu1t1yeWhe55Q
etAytp/jByfI7WklAt05AWerGWICMBJDHA7JVwvyJVCzLtE5ows35rtAEgUxZLId
OvEXAvqvY7dgsoeioA8D4GWw7YJPYVGl+rlBwlQEirR3j4sYPxhvpOuC59xeFQ6i
MCiKk9H8WQmeVO8W1M+b0k9UsYZk7BvgOJv7bxGX+sQF4w8TCe6hptuMuXFXVVTo
/z6/HG0wg3UwYMOWr4yjrjO7GRTM0K0BPvGLN4dGvPBpNYZOdMU7YAHfU1cjTLXg
94rZ1bYXV9tFcQ9HsmJoafUE7dA2XRisYlQQDtArPoLvAmDuhTbOXK5mapuqymDE
qMkR8KVsns+khSInRSIoFm43Ww7WNjoNyULjjjdCQ1xNHker8f76RvZFuvoMvLDY
Z4K+VYAzLur6K+6Lh/8aPp6ZHhJut07bl0VSuEn3XxVHxpL12DQfVyl5AUFaiwT6
qSMS8il9kTSfugCekrirWuNmZWD0kbJQ49HrHA4G62SQLyruWPJFxFkOb/z79gOD
TEvhAUY+Fx0tAIKj50rCJFF6wJMijnY63PO7BLPMSj3ZTmbLNbU5izEi6+psPzPN
qfrU8AlcQ6uoWS35NrkXFPOlhe9WKg+kW2xXLAMi1w3U6XLJfnHInZ/7QQ5H7Sw4
hAL/whtXW0k384gZ4P8Q+MBLeUeJdqcoOpfQOcPYQ3NKt5HK6FLjLmdnqwkkbLF5
waIibv7X9p9GIc4Rd5qQQGb+e2ue1pdVZSDlI2hBy6vbx/mq6WMMG+2Tfzb5OL1v
0p0bzT9bchtVyHeZJwMTVlT4HNe6l0GeR4Y3XHTwIEWBMuPiae72bcQvfL9R1rEi
s6yd850/305YKZI4xmxIjEfp+Toz9V/0mMkiZPMmX908XqF7XKe4HjUbP/2Ob8Lw
DF2jWzKDZxrRx2jAnkcn4yreizbQzkM+8rkcRXTVvhdKbod1rMJA+OAVse+RtnAD
EM89YOZhVogYbp55CoAZRYT/0Wm48TOduaRptLBha8sRLap7C3kow9w9VEEG3Hrx
fGicCdQjC8elct3MkSF5Rp0gnGIabBv4cfo+rB3pxpupWEk3106B+0W62Nmgd5z/
oajopN4IMNRa1iFrjPYi90rNlbWWoGGeWNu7psbthu1WhC8lSnIRLo2Ft44denL8
6xf/njWUaSMnA8UnWQ1Mzmkq53Rg2UpiWq1Imr76jdm1Q7e3i4a5r7DtpXJd9kFG
vgDx8zwu64Cxyby9/uqI2WCLb+S4l+tJ1KzQCph+n+CgI2M4s6Z3vC9Xr96JJuvt
0jGNPk2k4qJVofYPYJP/Thq1ElKzB/LqnqOHNnSWzWJ5HkbpAfog3hi8w5zWXZZS
DudsRWTkAwbCVf4Bj7b0mI2pLV7f66H43o0FRZJUNIp/ymkKGxB7+u3mEEWHGCER
XJNATDnoW+So/VIjSQRwvWNJc7V50llcWU6fc4lI+DGIrsRFHuYrvEUFQk4W+eBH
uOw0AGjoLnFyLfUFcnQkZOPYSORPQhV6TkqcNSk6jqI3SdvkZmcGRVEDQRCYJfE4
rEamm//cNksqS1weTKMbSoienNhiIxOUm7bpbJ9o07zgqlegRSAuTveNTvnzqdgF
uLIv1NQwf1A5cTn584JA/0NtvH9IRqmy+Ibf0B+0Vw8bmVUD98UCChkoSKGvwE/+
4efVVos7dsmuvRlVCZmGG8TRyj1YtDp+ZPXYSv6Tps1aR1n5CH0Z4kUKZFWxQv4M
S9jEAhQH5fdyc9XQmaZyjB1xtiTndJX5Y2jxL2pAXDV3rIKj5CNGcagrGDhV6aTd
EkNga+9h5INnJRTfb9NN9XeuYSGbdXwAehj6ce4+4tkOJLPdBgnRqQZDjca/PijU
tcUn1PDUAPBqHWkFwdtoLvrggttvceq19r23OZ8F4Mrd5GeKOfKLwyfliieE5IUk
oUUlZrUOfSqYjVEENHCYPoq3SYiVZaZKF5ceEv0HfMUYKVasGqhIb4KoeRyaRAhS
1xaUT25R0Vtd/YlLRG/RxD42Xad7FiAP8awC5sf7LsVto3g88JLqLYxeGMs8xwnx
9uqW/dD4KzdP4YiTzrPKIs5NnedchbpsLbuk/ArTyTaan7NN6RsvgQwZbnrnmVrf
SEJo2CMLEh1eD6lsnlVTukX6TQQC6ExWyPkNSEcUdxbOW0Ea/0NEJi+ABBr5nd8h
4LKPKEQg9wLVkK3/2eVsboXPjo2TbTdpEUX8vE3GVsvmq2VBUnArHjq2E7D74ILV
LGs5Ns0XKeV/HdqnGLNa6WeOySpXIZGsOOnWPNSCt6Zdwx7yOqD3CPIbtSDWxTRp
MjwjSSrJlf1h25wJP9794zGZV+gnwP4MrLgp+AJ0YWxLKud7eU/S3D2XQ9ziV8oQ
4D3z+U9z89OeAG0pyF0i6rYr8tJnwjw4fkEq899XuCzRBx1R/PBlsXDCtdBt8A5P
2D1k1OPv+ePyUXo7ZHA0e2QNfps/18QIev4q8KhB3e0oE7Yvck1oXzIU6EiMX+/k
EzsH/nBBOoDnd5Jr2NMI8/e8sgGwHizu6DAvEXzj5Mvoo0eK3Nec3mvT33Ma5AQs
dTJIbOuIKG2/1MsNXZ0t/XkzFa9fEi7fpmBTF0VrvF6QiLjlKhxV/3ezk55Ch3yf
/n6NZ7duRqRfIkJ5B+yKv0eN/dZNb8niYfFL/PupnbAc7BYWj9SwO1EqIryvw/ph
GeTN+zeBh5k7HkofVtLKcRpwfwIAIc0PI3L0y9BrxEIn4QSVGYzXl3uFCrvgBEW6
ExR4I/91+H73+kipfV+4fzFZ1mUc3QTynY7NhUZC1VwT1RfByNw2w9/JZhOvFp/2
g/CABbedT+N4SbdjNhXes0Vxh0l0ZXzNzV0mW4SdJ3mnZtZOgUYv6EI8MG3yZIGl
qfFIKAVlRTJt1EE3EBDpNXizmaeaecXUM6vyNbvNvUlIUcHYGMSpIIEAIlmxgnaI
O70kzDcflsCszk/R+1P0KsHn1N2ntWZ4KHJsod2pS7Tk+coBlKvreBbohTTV4+e+
lJTF8BzcchN3vwLqRbGo/iXpId5UBgM6p0aDpMutP1WCFXA3u2KDu1hnngkELDUF
lwoH109j8WvRVb2wBpurUzBdTiaj7Kxvq/LspUsnCnDb6mC2LUbTjmeA4ERX0/l0
lTeb+AX+1IjFnrmERDmF8BsGpmemiY3E40Q7EJfuLS7W/IYt8TYuLO4kuuO69YGJ
3KTL1aIpHF0gRczpI1Ofy92123Hy2EvMLvpKeGQqCx8GmnMawoHdogVkZlDKpZls
7x2phxnuhpdg4oXOrk3v9O1yiMsiwpyKc5l/ymxjisGyhxtCxKqZPymt5QZSC3Ho
CRU4ql0go+SMCEDu+QH45LzeOtW6LkrkhYceN+cSUGHNE1FpVIInhB2eaQhPPMbm
oRqUi1tMhcykEn7VrA/6E82zCrAITUYLpPkt+VjQ+MP/PTIPa0Yt0GAYIyLlGUQ1
RoZq8MI3502Db1Yid7UXiaj9m4vuZp+kyrYFGC8sRSy/1L0GGqSRcqsgk4mdZD/m
BxFY0WvmbShxHnQmhaGwLT/8Bca/3XZQzurZfUncGnUTqyxL3+YoaqI7FFO90eF2
mWC8IRGQNyydefWByihJS1z/LQtLHCyIV/U2FEburyoLKam91g5xlJirCnJQNiTX
SGxFzz0GhAnTTvhriH5mQRIobWZG7po90g+TZTS+YKbnwNERsvuU/lU8fqU1vCKj
SqMbgcUPqETK500JTmpSFlEX5EE1WIEGb1WXV+2S9nfPoYbvVuB72NaCD9z11b+r
2jnrOg/MtaQLeH8kDaFCNFf4JTi2H/S8hJP5YOjavlUcCU6SiN0GPgd67u0Ktgcl
xMLwK1tZ3SXsQMXidMFrZxrrLtUiuxQmVxRJL788kzixbnRScT/kl2TJ50cCoH0E
7fiZqdRFqy/MpDHByR27+tqbmkbpRjT+E5V/o/r5X8Jb/iu84f4u6hVZ3up30M2V
oZQtMBJfTuaxPv6poApzwt2HclNVI/e90+eA4aD8HSQSehFNFucwOpMWe8j7iBJu
M57Fz+sUe+LI1c3IjyrymhGxYWj2oMTqdGIvSm+mdMgQ13c/xjTOJ+swndC7jXlf
RNwXIhI8cPE4xOEu06RAVEABW+9v/tZ636dm2zifFUfbOC8MVP2wUumLaLD8CcOF
Pyz3SWLqpSZusnLZlhIf4VFCvTsX/Qixa/z+wbwOYI4xtRUc5AVqtDi4Z2pY/Oxm
CJdtd5wAjykmtcx6owLqhSSk/NVPkTvRx0xeCMn9QAZeyEm4Im2p9DWwJ3nNk/av
ez6iMj4S6PfnsdAeBhwJck976Mc9wasVtjAf8uWA2rSNbu4sRvYMNRobUhQ0gE/Q
nAVMn/RW7fnpvGqKXeetgTAvhipWpRxr4bXABtIt4UtvTWdl19Jo4AhK6RnB1SnZ
Leh1qRsrlnfZHggn/EDuFmCXy9/0Fm7oClK1HLspF1KvSpOednfHCEXuyaEOCPkT
utC2PK3Y/5UzR2BJ7r5VAKCWlmbUFrt7wUGAqyB/NRJnIl0XGs3RQQ9LX91qu7fL
UUH4tr+c97j8N8f7VmcZSS5LIX/lPMEsxxnBQyhv/Sblkp3d8mulh2dGgXHYVFTc
Lhg3Hqrmye5lyiRvxs2xAzBlnct5E2kRFAxCH2uQIAuj8V9kLVZwphnG//gC8cYM
7DWZW8Xu6NeO567DRz8K2n6lwdzAuND0PW0bEEK5nzI8LDxFZ47o40ruUeHjN7Rj
To4YIo2KhsKxtXFReXKKAYYJbex7UpClrEd6jhpcDcCD5YiE/KigZMFKcSQkWRhv
RDPLimNNfq+Lqr7/5qAwBJqIatetqozZukLximeSuyGgAPjXJuxSmtwF4K53vRcc
4XQyb7gm38p5NVDY62VVItgCOZOG2ZvLnk78/77dwsZ0RMVf2vEn0KtZNh4Rzfcx
WHnzS0CReSCgpiLxvhTo/KNsc7/yWOfj/mQsLikF8yrfhK+DF2mhtWBywPWTAXfj
11Jdpe+LIrE9WQlX/WkiBjJ8w/Og4ExjUCsOJ7cl5YVzN66cuXdFIPCmliXWIf6r
+hT8XbXKvjH39ch9pjh1wtfh9kj9QzC3NVjLmQSVqe9HNwFU6/6v2mRCAFX2EYTW
vZfOIw9HYUrNmKfYAPW1QPjgv5HM3id16V73815DGbGpjJlKV1L+DP2QyuX5aCUB
AoQYRFjHQIKT9o+k9ilMGs6YgbRwgjnP8n4yZ7ZnwAFp9bXRtyWLlYXSd7u1W4S6
JstJ+9ol5KU6mZ/2P4EJVyOf/G2grErbgMRyqkr82MPgXSamIsSA1sZmAdqUfcnG
n/qtvzXh8ChZ71sNSM7GdWgn/dnwxzAZxa0hFxfAUoudKTVU7i6eJ4JV+wSO6KMd
I/SjrZsmB38M3nYzWDFpLdo62J4ITgPRG6IHXt+yjg4Lq82FjSYkfTMGM2CMurb1
6wdMrujPa8iemTsoT/SDrZJG0H9gJCh493nCWmvNPc//kz0NNpX6lKFfds0ehDWP
dC7RMnL/efsG4Fj/N35pEU5CUVkKhxkDAcHsF3Yc6SF102t1QL5yrfeEOuT/Y2J2
MP/LQIcGUmFd9NYpxHIZ6/lodTDWqxYqS66h7GhLs447UaUz/eP/kdYsrbVAfV0O
aDG5RowD+2m5b1dfYA4tRDhBiI5Hi5Ln8geaKdI89TFPrjHnuVuSCd7pNsfsFGkA
uuDALOKOExOqzZ4lcmtzL4EwLXTt/53CY8fe67fWv5zRJVg3521dRWN0Vn3arVNc
acjajqcbDypnAgMORb6xZu1nU2zSMhnV6PYr3xDuP8z4T3BKr/O+OmqoPyxVnb/P
aT6zPnbA+I3fEoP8ruiBCDQfFV2Q7A9zEVWBbVircp/bK15mHW5eaiQcrc15W5bD
mBFwsg7QRYWFwASw7fn98ViSKxePAfhogjOZHdjWzvxJKSV/d2lnYGW+KX4qoj4x
z9Ij1m8DSP/cTYY2UnH1nUgDzvTG9/78S8ptBr37GZXYdD9MlXz9ow4UYV5jmlJ/
ImNp2WpkhnpvSUuN2Dywo1Z+4XHA2gZIvrb0tv++flv94Wwrw/KOKcMy7p9gvNso
++O4Rq1EO4pcoyKl+LkN65kUfLSq0UsQXcdT1m7EQMceKCik/CwF7IjShpHqYjTP
OGK1mOgsxDTmvGhB36yQo/aJp/Hv887NudkzbSNGNnXY3v1gUgC3vrhw03IaE+GT
0pwynL+nc9HRiTV2Z4W+sT2/rC22ovAxly2wJwD54Kd2QbSCy1zrcBeT6IY25eU0
Q17LMGAFOOXagHCRpHd4trusr4NibZ3cVcwGbeKCs5IaxCcfuhb7zYloy6uEX64G
bI5ok58bTjcF5MadcyWOdYSvuYkCI2pLOdfgRL9mmOGl3FKge5oozt6pM3ysLqmm
2EnA53MMFyu9B3NcL7gZXUWk07EQNQkUT2MugF1V3Gw1D045a4VF+5rDSOv5znC7
iJCZKSjMg9yzZofMhZdGrEdefwM0Tlr7OmezRYp5ba2j6Ok5abcHQ7/+S36cboZD
o7GdFu9ZITeaZcrJQS5dpByL69OZCcWVE+w0a034C5jPRQdTEe9gG2wDEBaVWu9t
OCf41Dx+DGwb1ttBKVglrVodUTfPlC+7XM4Ugno9bu35h7yXfOgaAEYuDfzealGw
nmHu9Tn/RDY2YQ0jRHV2eyEjYHQ8gFsDzzhaZE5eoVr//XAqMHaP2WUg75CedHvt
+RIDCNWXAKItdo6OUre0wMQC9Mz9PkfXFob1MdfpAovz8QepahjHLodmhXPZMBV2
jM4beNsbU0Sr/3pYU+v738FOtjRRchSH4yRv//o1koybDawdF3jtFIHdOBS4ylAh
F9Ne7HDQ3hOxYUleM1wUpbJaQd3k8vCCciX3TqYC2vvc0AGu7BBlWjuQtnYqi0Hi
qm+4dZzXd7vfaxKnrqHFgwGdOXgBkX12Zxe5yLcBOVVCiJruPsXSjpvQCdzxT48y
UjLOrjWt91pJ5fMqpE1CRWcTz0oQ2/ja204u1XbLYh70yoTLpeal4P0Gb2ZudpvT
uwZHp2C59R5WefPIVdgy+XGAij2Ts/BE5fYnOlconKT3RfEl/Xp9d9gdbC0VRXmR
LHeH5SyEm4iQ3WYkhI/quz0Oag/heQmobpVbBQTk8NVDFkJcN4ZwclGnZpIP4Fdn
88Q5CF98OtR8UMjaFgMdWdCcFno6iuCY9oprlo+bgyGbvMjw4drT0KPnk486tk5G
Shg68qYKfIueAvunVOlCX73H1n2k08VN8+Z0q1OJd/g0vnjYmMLfJDi0JvCw53pj
Rc4Yq+zx6yrfRpu2NYQHKu+YvOcMfjoFvu+l+g1T/7qGUCZMzkSAAgfUhAPg0py3
r7CFr354IhOkI7gkzsOe2uyQg7emrxwW4kTxy+GdAerVGvdrM0foKofi/AEQ6fpy
NWlPjEqSW/wlXigRKe7s8MJ3qE0/51p+6ORriUSqBTyhoGsG/gy96oN9IdCtebON
aPld88iWYVBD+SdkH+ewZ8vBoXOQcQrKERqrPreIG52Y4YZvcU40FdRe4Zbb6jhV
qZz9b+eSYHS3v0oNBt4oBfkz7UaTlO+fRv6Vw/pbgiL3paxett7LWagYojxV0W6U
UE3lnwKADs38+SmfXHMg7WFHpfjvkVw285ZL6GX2mVUvTRvt5hSakhq38X8BLt8/
yFaUcMMqqdKK+QhkZ61guuTDljMDs52oyw6dC46I0aUOvVaNLGhV/4sylrS7fgid
DGy2AMUQc+rhyHnfZbX8ywKeJVRmxEnWuB6Pj6Xm78XWeaxulo/NTFhXX0tckmbW
qrXOinr5JFohfRQOEsBcMFENNV1YNI5ZZ6gxXrljaAB2XG/MyFNYvO52RBOj9XPu
3XKCUnpK/T4akr26yMEJN0tu0VLZRGV2n7wyt/BBmuirlvrdK7D3LIm+J5EbO5vo
D3wotIx36cKJK6Tzmt4pmof3CvdfmcEQ2RIYfqXu2HGO0wZPvAvT9XLTygjZ9QiB
M7uAQ1puQvC+oiFlZYzZNrpnHvIPywK+t8bZD57ouxBAMTqiQPQCOjUH8InOKltm
YKyUgJ1O1k/t6XKE56y5xTsdgCAslv34z7s9HGZ0QPXv6JYALDWlSSLg6XEV7Cmp
OZPcc8I/FG0wsNUvkWBWuqUHgmh721ZopeVOxEOH9a6Dq5JVS57DMwJy+pO7pojN
qv03erHV/nWQrEik4IPHEV3WIrafXqGh9XGUv0qE7LZ368I3o93wzrrX2kEg+TLl
0BeqREMRf+3oZcBFSLCMZA7e3OgGxapnc0B+Hw4mVUj3DoZ4GQUOqC6w3VBiDIXN
ORuUDoBuK7zUIrVEws7rqNAuUqDYQYXTAsWBIs7IBOJncJS5LGjXN6i2OZdZ39wH
8grXVW+3D6611/c5Dmxkeak8mihAfWF2xJLveV1mw+ncM5lJgz8g1z4lEjWkC/Xg
tKw6R0CmUpXE1OheWMuO0irjPV9Y1Eco/ZyEmeI7yyvFI/2t3X8allBADYpLLraU
nRqRhmx5ZzL7yfOsmgMjpkZ+tPBmaN56WbN2XDETsz/Pjv3s3iB0sP7ygMoyqqis
f5Qjk2asMayPl2TSRW5iE5CDX74yuILVd2CgoPqtP67KUpzKFxhhlBDSpEyNuyf/
Ob+RK4Fhi34HTv/8SPnBfcRTUnUgTUl/OYI9r9KqLsCPeklX5WqlmJtB9WekCy5y
9Zy8HXXwUPKflHYPCChRnKPYsduoIar65D0cN6eDdw96LoQrGaNt+PILj+JUc6uD
aYx58FvjLZEW0cn2x9Rq18Z4f7Nlk45pVyeGf3JIwZwGJPdkJ5qZ68fzUO8UGBJ7
I0+GWG3Ifrxppuj0NS1YbyG8At5dJ8TMBtwwBNERHGJGd4m/x5KSW/UKSdjqMgsN
jVRrLt4D9yFSnJMp7G6KohgW6zq8N5bnufFxRdsezIWzBhn1duVWied/mOUEOvmF
L+t2c3hkj+7ELVxdXYNlzOC8uUP4KrHpgL1YJ2J0WZM9kDfjF9VWUPCFQJtEwCP0
FTZ1toAUHyXr32er+SIOq7M+ShhwnBtn3MipgIi5lzLnJ9IL0QKYJOjdJ3Bxk/fV
inWyzXIfGf9EjvFHu9osX+Z1FMPrewNMdrzyK+dosyiOZdQEQjAPzdaduFUsYeJN
AiaM+E639DbD/ezIEIAyLFqQacPIXrrS/ZUsGk5FccA4d81lrjEtEUK/A6n8OFOG
MJpVZDgDQmwxtVNoFkDyvJ6wAvYK6edt1lrvZqe6WavTY5kOWBabA2691K3vJTFg
1JkKXPY4gMmYTu4aSIjE2jC9vVbxIAjIV4oQtUpObMiA+RT2AVSLQQ8Zjy77oaub
gBdVMYuUlKahjJPBg5reA19A8fPINvv8I2TCcGI/xE8PfjbzRf8Edeha0WuKBAXc
QSQD8Cvi1GM+v+2jR650LEjbWfS7zbVkntBcJSMxevrSd8ykCE3wPN0npQydtF23
SAys/8dJPPk7ONMJ6/A3b6tTS/dC9Eo+HIyg05sIqkuEsFJK+jqF6DNbfL7gR0Vy
WuLelXmcrWR6lk8aCWlgp+ExC6nTJ/VeZZS+JqBxljQjhURORPtK8gbjdXvF+rwe
Kt+Ze+AB8U42uY0UMBqfyR0AMAu/NYmzcos21yBoKeG4ZOjq4hOrsKWtxtILcFBb
0rZZZ8TPZvqs3NKUGXpUGPJyZWCggM4yw8XXxsZESyBmvASY7GkPWVj2c2TxRrws
TUJc4GG12ZO4+kKWhFyTxP21fF40880pWFzv1j6sYEDPxYF5Oe+AwJqIVyroyLHv
ZeoSqtOvvy6joXy1Zn9Awq/5JBTP4ok8REOCLJGPfAgj5cGU0T+8GRhf3PYGleTX
hY+rmVy7gHG99xLJuj/nAx44FBMJH+Bg8JV1c3CPUOSuthECR+pbz/pYfdWv7EPz
f/2jKydLblS3WHVU1VvOJalepcKsDTuW2+Ody61fXZXPgS932d+muDxyjZ22og99
S6vScdqMiPuAdUTXjaTYKaA9CpUl8MII1cPB/95corDPFjAx940xwQyMSJRuosHe
26AI0ztWjGIxHjSkmaFUd14jmb6j5WRNUeTzbQUPdobr132VHFABA/Ed67WsftNo
W9Xo7d+41PVPAbZdKsUtCRv9WOT96/1cpo/mJdJ1ngb4CSXxC81l6ZKxqVDL/m2l
3PnKugTydL86r8FAc/y46JXtQOSvxTfZMqWro6pw22SmtZRCnzlgFxmN616FquI1
SA1fLSNcji6K/mfbK2FLoh/Dcfb6IcisLKX1amtXLXwaWFX1EUf7TJISSRw31hY+
Qt9lABdd26S8Ykvs9mBUFUVh9UgTru3eKPygl+6DgM8dwKhEcKbpjN3N5m20nzH/
gWk+53vAT0SOC+wv1ai5Fqy2Ugg857THa853QdjOT6+7K8tU0UrnQCQWwBVmJqXl
GViJvJeJvr7++MhmrWp6tBoyd0+GdwA5zM7VbrKozsFMsv20GhkkIvb7hYxkUc7K
6MsxbiD41EcLdRf1g+6mqpu4+BvZbOPVNYaaEXylEDfT+NXma5XwqnKwNYOU60UI
32ohEdeBL23UmK1m1ilU0L+iLzEkDoJpGA8Ta/g/wd2TDb9wB3VqeRLnDcoKsEJk
/S5X0P4XIkXX7JCEJ+G8uJMcEMDeB/i0j5GIgkcFCsmgUlKrr9hF1Krx7+TzPMFI
0COnMQRtzacqqP4oWTRp12cPgHr9QSflnKWDOapU6TOQD0eAwl3uooliL4Gq2Fc3
WZNnYRyMJy5PM2fHBG+J6OEA1pYf+/I03CwWSwSciHCI3TpLjSCtPHLMFx7ivD9d
/W/wv7TbbOthdmqLlaRcwz4HVI+0X5nk2a+K0TliV9UHWrtQ9/2u/9i6pAGERRFc
pB6tk38WHSo5ZzR5Z36s+qFj+hMh1azDV8mzFADgT6E2s1KA4j4r0BfnOlnjAVEf
d4kj1CFerjYvYFXeeKKk2lV7bVY1fDxcP2DNbJOdMXe0GZZfbvdnK4T6gwWGdvu7
i1zKSQ8aCqUf+aiBURogUYZMd7H6PAKKrnZYGjCD5sDZmTvOqUpzCeypFoxuynhv
rY8X7/od87ksOtPfofmOBAsc0y1w5aJbAjiNIKUGRhQqKX1ijAmohgw+RBZXBy8F
vSE4whcnpwh9q2pMceCuo7Kv2KCqIENrVeUid6NZtdrkJZdKEyiilSGmBJBcJcjk
4tt4I0nEfZEDeDLwpLDk4bzA11gTWswlR9qt8j7nnauHPRT5R1NFMVjjKgSiQ67h
PS6jLOfUtWUB5c87UDim6gA2VJANeRwynjPMqft52dsOn6LqHRThXskkS/FGXzA2
dOi307MuX+LVZXQc0G01iB1ENezwn4An696S/8cC28oBj14aeQHd1qq+Pf8eU9SX
A/jXaTeJb+i2EtN8U6d8KHQWdnLjbEJaxEadrJdSIDsULzpz01hrNnP5LfC1wiCs
ZshGIDxZpeq5TZRgPR8zGQawpOvIM10kUvkfvFDUNine5DbqIQFTYSJWh1cjMEAf
wOVq/ESgzNVIwedkHpiK9VZtYB1gYLDBCJwo/VSSijmfbVTRzOdOwm7yXGl3H/cu
Ix24i1dg1LeFVB6OzrBz0vhMXAQV/DZNooBNF0FUuhD5uSZ/ZmYwuaY8T7d5A+E0
u7LQC5C7opkpemD2ng1cGG2NDLzTGgBJ1wj+FHqJuLdGGAFOABZPTfTqSWuvBMOV
yI0wJVfyd8l2FvEWYWO7FD5Ic7mdVQjzQePKxayG8QpfSGpZKbptedAvd5jzBhHR
gmPhXU2WMz8puAIThpjhGCVAgPioKMJQHeS9l/4RzuKO6zTR4yExW1rJo5iJuHwS
nSGGdWDkzJwHpcmjjqghZV6llX6iih9UMCeoEbbp90WgSb2hzZ+3vXo2JX84Gx01
Pkl2Ip7UJH/LAWtq+8Tp3uqDckc8Pxta2g+auGzXvbgximmCGpzCGPk2IFNXVMZi
OOYQeaICo3TRuJg2cUFsgM75bsASOb9RvYtkWz7te/uqxZzNhzbN7STlGLtFQCBT
w/r7RSvGhYsxb4XTMAukvtJp0vyeOxQ71iB0XkfKEB64q0PImXTV3Mvgqi0Ww2Cr
57si107eoi4uuxH91f6MJlmup/HRxh2rmWM4dxUoZroPC9xnk9e75nxjpYEypahL
ac8MpQ6Ld9uuZ5z2SZm2aZ2dQVQIHM12XSOgsZh/N4Q4IBMyf9T5nbMEuTMd9Gib
bedhI5OghGwFwowjaBNKoHZE62KEIWC2vSxLRZ4qhz0rvR9CF3lodz+mA/4wWUax
rtWdxXZzXXz/J1BoGg6PDl1R/pRp3x+8+gzQ4I8WqDz9s+4fevVGgWD6QrS08VPF
M0Htdpkk2AF+s5u5adwsx/sNWeb+o01KT654G1NVT8Ak/l2RGBE+KcK7pOmTNl+5
79/6yPmjZ7gAztYR//y+5fLY83wc+yiPMoNBBBiHv4udUzaEcov9oGrDHse6Fc+l
L2LL6Gsc2WqHBKRjE27wtHjrt8cxUFlpc7OMm+Jrzk6/r9wB5otafxQEArlYIn4k
qWfoPhfhC6ju+yS5ZR6Y4c+FONOq62fWOthtR4EOVBio98UzvZMYHait9EZ48u7w
nLpr7F+bMb3Ivc1zzeBZQyvByPB4wx7De84uJokQMKSOeSHiYzv3FmloafQCTdTW
JTPiEK4k07qR77emJaFVNrNgDyZYgQeY8tYK4vim3mB/d8nA7yxMA+w+1b1HZwDf
00g4svF0jPO9VXETcpGhedwIqhpzMEFljHvKyqMdM3YXHjwxCZY9lW3PHlcn+79D
SkAOPYTaBY9qS6MscqSBQUD8lUQljqYO+9plVvfxoJqYXKus4A3ImGJ0PCWcvF2q
UmYzptApxP8kO0vCweKOawqMfSZxx6xzMIT90/CkJJIBVoFWcpZ9NlemOyKBeBye
CPOcuI9pipDkto4u8OUZRh0gepH5V7sfMN9FoJsUTrwzbuRCp1ivr/lhDZKqaJFn
K5gGaVKCVw9Rdh+cv7Pky+Yxkp6FzY9UNbLwSeDWwwtKyOI8svZCQIzK0Dlt4Dfj
kCBDOLVKlPzqazefPOo0wvAjOXObw9jo6KlxwFe1Do9YgcZPryfdtE8RRS5BAoRU
k9fEYdVlC9HW04IAqvHESRXOBK01jnQJefY+41sH3kQ/j7+ACv0OqE63encjjozd
SFlbbw1mLn+uHji2zFq+vlROwrM0YByhDetv8bgo/st9nkKB402gzqzyiEctz+jv
tjWWArvj1s0XgsbBZwUtDIpJ+yq7CMOPeEbGNp9hjdTy6PLTTqHlXoSOAFnZqhXZ
CXwLzvhGh/JHb1FBoY56OYQNaVjC88wcRt3sOH8e/t/AEJ+pRgGzqSlwTh7BnDqh
iSkxL6EAQXpY11dbAfOy/k0GcMFqtEMYBFCQE/XRWZ5A89zv9RNJzFidGTi3vJWQ
7eoAK7fQpb/DBtA47O2Pf4hv9ozdGFYlY9WyZZFQt47JzwIu93S98EW6B8qvzlBD
E/ooQWhewQoiCmULnHhxDn4Fn5Y+TwmKjOu0QM/IYRglcsF3Z38X99umqY0EQ/h9
4OfdOvc9uu+etqxTGXeMvBad5YdlM0AA6OUrF7Xr/7OiHUIEAyKEswA4ngKS/7SK
Kvhv6AHUtD1TlOMKie0uHUFuRHYlkerKAWBhfBWVLe0jjmO2xtgrxiPyceKSDua6
kGBrcmqdhFrFpbisoZCHRPFgA7gphZo/73PNddPETLugIdCLKFdv29wdymO7wZ9d
oHGbRTN//+IG8SaCUpHi8W87RcgFTRZcqBKXkp/dbo5p2ZgD+I6USE+SDkNNgRrR
UxAYFy5zyKX+7W397EU1klqZ/w6BGKfltsC6YdBLJxBDqpxiKli/Fg93ZMaskfNp
fXJYEmW83cadQGQqOiaNuq5CualYcgPZyRSInI1/+Oa/tET5qxcLRwf9ZCuFZ3qM
rY3VYWd59fr9c6GKKKN8hqIxj2n0W4IGNGJBvaamKt4/Bz8nT2b4Enxz2hq839d3
8JchsW92AEgXV5bInNvIo4MjQmOMHVmLshLW7ed0stx0pQC4F7OkHz2njAm+9tNx
FUZz3HOznmD1GJiHE20QcMXW7IYsx+bPdfAaaIHDuYDP1NWgiutHFwDC/GbnOIKv
Tl8UwJx+KhGXVzG5XpIThEFext22VFNiF8h5ygzUZRm4yL5Xa3+/la68SOv6PaE5
QL3zXa4VuMXA5yrZMpyPTsS2DGWRdywxK1KzcbH+YHfNjppKTIVJWKx/8rZCgVMO
pgRSq/WNyWhrDMXVur1ysHah1cCtDDToY296laoGcXs+ZAnsZybhi15JWxOeVBSG
WfJEEYBkgmWdLbAdFViFrlbwhU2Eh5pXyaZ60amB0xpXEXGjNv07kTE3DO3Pcwez
EpxeKvsvoYQPaocq3+Xylt+DL1iXeEJr/zJp5+KVSHfnR/XNC6X6vW7Z1JcL1742
yWAyu93QZQ5UrhVH02XVvkj8qWjdthr0wvPnwrFZW2bFQynyyChr2yru1CVQb/xE
4ay/JAmnpFnSx8DEFGLMCb5jTNt/feTNCEipOOc0nOLL82e3IZfjoW4vyFCdgHmk
YBhY72wpzltq+xZdBQVbYS/VJv/vtq0n9JrBgOCIFRCebHZBHPhME4BSpIR4X3YM
3jLsmSEmHvTWrofcQHrjoyespkJNwKfnJC7XHySYbU4/IXYKUVt9Rf8VJUHLG29D
WSjFU4c+8kqhxdWAwW5Tjq21u5UdfRYuPF3Y6AvPTAJ8KqlZChRCECbqds3MHbYd
zql2U7XZS9H8A2mgnkdjG/tWOBQUw3/teJN3vlbeuNnRWnd+EV3ndIecl/jJbKw7
XV+oP8/luX16RBeiTCQu0p6hi3mKrTeKYrjC6MqQ9uxSxKbDFYnwqDjYYO9F+W+V
kHx93OnyyEu3xRP0JQXtgdqjkkf/WP+1mFczqaBSdQXk1WujfFWnyfyqvSYdaMJT
Wc4ERpkHCvhtrYUpe1O/BGcqidB5aIf2qJjVL3PFnkHErvM3YvNYgd+IsMPaZ97d
49CN87rvTQLdLh48MzqIi3uEeopjZOkrEExgHZdRoiAsv/DeKCLgcbEWTNuvFewF
Ebr9Djp6EZhyz6to9SghfhkhoekEq7Ovf/zwZR9DgxTyzYaAJvIxD0GNovsEAPdN
B1iE7LhQRXaEIADkT0vjSbhMeJ7vZ0K5RTVTTivlnMahzgrMMVydB/hcr/epzUwx
UDgtP55vdSIkm5tnE7rkknj3kklKSjB6OCFYdFvyE++T8K7/JUsBRwDdQVGY8nSe
2y3ZSCOVhol80NWkib9nCkPNWRTQI3ffTbiBtQGMndcEGovqhhffoRFgsR9/f6rq
LbJLtNqNTQsQEEv5tj/49jvDarxWGUFGDjdMK322M726IY5F7BzIJ9JmLgvRzHTD
ntvhI6lgyG80bhQuk9maHJ3HV7lckWegJ2EmL5cSBI2EtPFalyw2TGv00z2n5/HT
s0Zal4uTsX9ncY0+pWCZISQvwBULJ3Dxn2ySvaZr6y3xk0/mRJASgXkm0ik9sao9
oQY0Jh8UcEPLYRtNP7lFBKy4wO7/LbV0psmhmn5wQZPVU86qg6uvbrQNiEDmpJJZ
EG8IrLhAZ8esy9Ta5rEWs3u7yr2hHk7VntI8qYEefqD+akNM4KOvWLI/ub0ug/iC
uznLgUkBwGtAc3BMi+GvYuOZU7OnIsvnf0zsBwShtN+SBr125HM+BTBZ4mtqalq0
A+dQxh7itdEZIjD4Wpo4i56CA95S9fVMIF0iD4rh3q+Gd75TS7d1qYrPtcqB/kXu
VL9ouMvhLnyvxaU/LAh46pYbbg+6jZMAztHknpxMUoIa5e9ng/wTrnmPrKeQkpxB
W179/sXoMoYttDPCcajs5jo9p2rsNSV/35Ib6QVxpqpEPEL7gBp1UwPFLeouTPQ5
zXRL3LdLFygz//woAwl1usALW+r8gz2Hzlrm3XgCFo/jajetqGYVtM3+/PTNnhL9
S+PCntjJ0pxi9DRJIc4WQzfN+O33SnawX9NC90NfC/TquolBju5SnxP3ujaYmwQ4
jX4q1jKKd4EyvuOonQFGmIBTcEoAOZ4JMmDgqYKormuDe2bQPEJdi7uoIFoNSBY0
0UXdcUCxsPaZRR+vtpciXfjn0dDhRFFO5fPCKWzL13gbw7B0Z1J0ase4IGfu17Zh
Y+ax/ezyjny7bn/HGxTvBmTt3gZ8c0mUWR9iDpZLQGt6gYUMyK/siYj66TsUHGYI
L2EKvnPG3UyMAbGdQDJOqaoMRgkE/MncQKaE0UH/ugchj6hoG6ueI4sJVx9GN4uU
C8VH1V/gnW/YcMtPedbCtXO7NT+Mkvcy+y5s6/j/Ib/KXtQrJTYhFlD2afxWDU6O
yZBissjK/FbW7ISnueueLKKH0Hpq3+dSB9Dxgg4GpDIvcGJ9t+2TCyzqF7IXwejm
mNA8e68q7IHZWz+8xtrlkG1Zw+3AFDhTEW76pobIXpgsYa6nM+T4Z7eWhzE0K7qB
6TOYumhts6py1YHWLO3r+6sj6mfUeK8cFhFJpDE42q32YJe165GSyEqZg01REnJF
7oJogaorjZdKlRIIgVugc2iiVy3GwPW79HKfuzN+HNmVWlc8cfIFMUMOyBKsaDy9
ysolKLCwMgVFX+jmRFTONRtPuDL0StXb1AWfv8NF5uLorlYhczCSazI38mjGP3le
beqydKEI9iwihHd0/+QOUEr7WCDujm/2pVy9EfldnjDafWe7SSfQxJhOpMMfa2X5
bstGhykQ96XWn/IARAH4wz+FfkrxRFS0PgyovEReZFIYNzZaABykJKmxW2plHiZ1
S51cckdGR4+Q+bBOaKdwM94I8SeP4GuEEF155gTOSMv5mnNdjQskW68N1r+vGe+a
r/ZabwsCUN9XxIQTZpDpn2qdkLLoiv9YRgSnmnH6GN2d1jp+cM1wolWDPzV5YIqA
GvkMewRuibWdGksLXkvOExdNa5TT+ilRSBRcxDfLwWAMXQ8vzBvi6py+afkBquoq
sgBCNUQtoiAPSKzmCKmld/fW2ED/zi2+Ox0DB1n5+S5JXaeAgLEZQa4lj1EE6YSI
Yo+yDZ4PpheKq1Knxm40eUJaT/sOFTEvbTOdVt995BdFN7WgzUnav+hk11IvS5Nq
1AHnwfOw0TbVvifwbQ6do+XnUoZ17xzxO6mrtiLW6SqfToF1OI0uzjR3UaaBhOF1
JKBko2DvhO0XwqRl+A1NgIGxAjDzqBv6DmeBLKxu1j5HemHgSduuk36Nye6MdWyG
ewzwq6FWAt7DXOElUEVY1LVSi1ChDTSMahTrG+UbUbMLAJxCjaFej0s7bVzXzDE2
ZYWJN4jE4lAOs1xETwrUPc9cBCE4+Zn5QPLAdmRbYw+IYxtmN0amU1axWqhwzrxA
Vusm3yl/Xqzm/BWGD85EpKxFHnN6rzO2GYg2eBWz6Gqd5YMV6y8UjWHzQikBLglw
G0I/6njsEU34ADkrUNYi65plVsXl4r/ss+oNfQbrAmW1/tkoEmpxSO56qdBEULwR
+Gd+i0vN6DfTuxLQPJDgj2f35UUbfSmlkwyyR3Dx5M/yuawlWKZF8xM9bA6e8vlf
Ap6IQGums8aQVDTuBDyQN8llgMvRodrXNX51xs7zYf1Jv7PvRtLCz1BdIgBp0cSF
s4GdT0hbngsG08iWTQX/dfYJeuaGoGqx6HcqAljHK7r/dEvxJDj3SemCNAF4Qfev
/19rlnm3rrLCnrzQswd+NbRiloCmQrHl5vgizVigmt3UeNEW+jTKMgJ3gRHIZT7v
X9DVLaR0/sQz4pX+MNVsUflPf1pitWFYazETS/2RLA8boc5e+EjyedBxkqg2JFNL
DMLrdFaZiCpdAUue749iRqUefCwnHsnBJnK63vFTrk2BATrd2/xqcPI72x44Zauz
t71YxpDxdZXWG/JhWFj0trv0Mj8UNaCTeOBdaBaVTYz1TmKCHjpPbCesA8n+jWXO
akqeVFmED+1gA7IlpnzXIcF6b4XcvTOzRgBsrjzfeCtai1LxoKrAXH46knSLthg6
33WMwVGxHqAglTPO5wbx9oPZjFjRCKhN3Y8KRzdAyLlTq72O1jhy0H8aZQAYHQlI
zBiavNle9wfS+q+sbIM9dh7tAVZbvO8DBFumQKISLnaX0gBxendT3OEE8mMVoNJy
fsRDFu2A8mVOfkgTf3urvdk2UPbHcvpP01Upa5QCNCNAvxqZ1+TFHsOrBNLIvutX
aDLZc8PBlO/px+j9qOM1CJlWam/xGQoFzHYC0QTSoNopIZG5g1Ao5F3gElKocvOU
90ES9Vm8asVHc/CdgKMI55fY/xnYRwb8TmGcmGZEria2hgw5UAU3K2IXHb7uO+Cp
I4/F7YUNc+RT4F7ybehBJ0z5W8AZdp8aCf7lD5MErLlNpLj6S13sin2VzJI9DX9J
eGXHTdSMaFXNP93vX/YdKfVyMP+RGkuTrFlYMDnxv/8Lic7jk8GxUejikUJ9NWnM
eQgXsJgtXnh/K+SLm46xTSDzl3pbkKLCzEkXjJdODRCsi2fTh83Y0BVlRX1PAld7
mghqCYhwqXEe0rzzvnTyBPbx148Rfar5/pYhqY7ddScwI4F2PtEJzcUpExIYohOw
g27LvMDfZPQ7+yx+CEpEQzzWgqMdo6mc0lctrGjnZILu/bvhkN5bUQldyRa892t2
JGJtodb6nu+A7Prwx0CJ5I9RkZRg+MK42cenDN/FKRQY+peNVbamScfhvUBERCf4
5j3+4tjAct+xZ8dYLo4dQ+5MpyMhhNmFCdDOz+OKjNBI5Sz9+zogJqBzsLaGE+LO
bLHvqpyZ6v9LZYWxA+Gp+8Ld5QVG6NOl4j+CqXY2WIp6koSiIa7B/P/4o3nRGVB4
ZkffF8zyGUPAFxtTzdWQ3U302MDIZVKSpEciHExrU0d+c86BvUGx+uJHl8pgLCm1
0AOVw9zAIrC+9p5LPIO/1Tiklya2aA8M5TQx44AdB0BULgBwFb0/pnFK7UwpTLYo
j2bhARzAV9iEUbFBMsmVLkeoGb+aQHFPwzUdwRBERP3r5Q65M9+KZAo75S2krSHW
tehPyHO7OpWshTA8cXcDyVgnPY9XG4XVN0mkkiXHj/VssDYceHM/ZM7jjSviX32x
ifX4+L6Bvup9/L/uiAnVFmaPWQqtPqtA8/B7Mtez5pW+Sy4V5FdY6hHQGozn4K2C
hNtCsvuGP1Be84xXHTuKI9w7OVTp0Ctqk06Hj4Vnf6UiA+ndmtPx5XM8TJS68LTM
K6Yv5lyUske5nJuRhxwkGgclATKo57wbfL/zT5+6oIcTpSVc/HGc47uNwqLZifGc
eeRt6wtViLJZzUWihIPappTG5ZE6unr5J7Vxax3OJVS608DRObJSP2q1ef/1uuVJ
bx0yCeoZK+SvL2ZD+HfNGvY8ksfpO4E+axRP3jsQunydN3v2G/rYS2m+dvz/3cPJ
pZNAAoJ1nsWAZ/9sAp9sbXgcbiWKRtYWz6peVnSvv3DIeCuK9aYarFl82nxCkWAR
otf3ub2C83XgSTcIE2niAevB6z2ZJ4+zpOi7pDy5fm51mq3dRYpawDVuh1qpmdkD
PGHWmOU3rbUteoYOJn4pY778dhM0liAKtDP+8SEeIQXsyQbtOdtHktPLRo+c8Gu7
Q3DvWwqVqlUi58nxxwghNW/lvlPgfqDEjOQiNzrN/4jYWErSOz8OrsKlDR7L0mMv
JYmEOg5mBQvbkeiXqtIjkjZ3h6iV4MXlC0ElAolpZ2IBuHqo0loNA+6n9X7O8gNb
Rb30hvnZ+oSqZdHgrXj1efZtULh6CT4Z5wWbPIgvpHB9ZQ2/8kJuPybO2xzWGXtf
Lw3PkELfj5X/H2M5f3QNb80qqMMg8L7FH35fRlTY+3XtmdhfAl19EeSr/sPtJa3d
1Mvv4c6Gy3XSgjw9QVhyQPjOvY7/xaQYvSaPYrQlOXLqMnCDiyGvPvkxNCf0JQre
HGwABDjsqVcRi4JCGDG4mwW5V2Q+dvoR/qFxIMH+7fUrlCUIbuvfJP/ye4AsL7cH
QgTPfdwdZAO6Khbh3JzumeP2cUR+j0lJCcn73zOczbd4adIMuyzqVUprGWETnF+y
aR9poKDkCFuuNjQyu8vBAWZSgjeSp7vkomb85KlfEzc/ZpQ86JX362xTfKVhbZqg
I7eithzdQzdiwQx/B5WFyGrltCcjngyr5qYOWoEo9DOBV5YSs5fjoykZpOy0Q/1y
3AU6w/hd9opvd/iPzk30+fSzx9JKe77LHP2bJsv1l9sXMBqnHeWPsA0avJ2H/nGe
h3VCqcryPQVypSLsQTfJ74VXQGViahpN2ugdZffOPck5hTrxx4OMmtek+faXVNs1
ZQftNawUUfmX6ccxmVkCKfMyGs/lfIuiT1vwKXrwx6swt/eoH5PLC1NvYiZ25X2T
qTuxXogd82hfgD+6r+4BcAC0TzW451awOUBw/gqD1gxfUxDQJ9BvUezUBBdU1Raw
vmAl3GtblTYXoKtSuQH1cef2a6G+p8YOf4VQHH7T1MMb8Tm1jTYv0CwejuDnBMSM
KlDOdGi4gldqwDxm4wX1HmAv256PAu8OYXj+mENA1ZaZynoCkZRzcxU8EDiCd2DW
U0KUnVzlzB6qrFrucEOx/LHrcS/mHbfHjnlSeFvXCu0a53NyoP+Fytexut/NHqyY
MDZXo8+Ziyx1i8Fg7vbAmXluVtPdqmngnrigH9Pm2WwuIfxjlZi6rfDGyxkzByyK
871IvqPjEFsv6yTXDD3s3e3/x9v9QENMJ8a3xl4A0vfl1I5NHpWPTgIMFkL/Ar2U
kSE/DuqonG2igJ0JEl+GH3P5jRu9ge9jHtYM1ADu9tcQJdimIVkGgG+R3bEtzFy3
FkZcWTKR76RRwt7vuiv/Akg1UClgH51ah6EMMwIBhZ/zrbklOslPX5AQmaop3Nj9
SYFnHpOyfo9xwcaSA+Kbh+csdFnOf3ck/m3+DQA4skWnSlk/dF0CnSotmdYhilds
5KZ/P0GTGOBR+95EBoo20qpcGgiWSUre0WWPgkwxoU0qQziFY6LMkVi8wAajYqKC
uGsgu3Cin6JMBjd8ISRJsFtUm0k4jR+AJVYk15nG3SjMrcTjd0uS6h3q2cai/Yor
JljxawhNw8xREXU5WH2kWv5uoDaBpnLypBzfufzjqz+MBlmYlWuLT5UzwqQRHii9
/mJcJCt4opp9JXcuPmCKPg/UcRk5YWTLLLIPoSX7JJ+Fza5RIpqGelGD5CyIrX4H
+PdykNySNo7h1tUshymnOUJpuVuRtCfu9m2RfeyDOTQvwNGwELNJ3wXaR+OPaS0R
CgYcgcFgBW3iNJODjpm0RbFtPSXv/IRdTA0O6GKQg9rh9clE43REnT/KNnQjD2ex
+IJSePycwK/k5jV6V0jdVGsLohPnFydAe6AZEu1ky7bdvTwYuR+QTPsEHpQeghWZ
45j+FbiX7TEEc4TXVVKGux8uJTndZ2l+74tAzgyHnR0FI/XwB4N4yFYNsl/wIG/r
JwNEoqT30/+JOACB+7MLFMliMNUbacT6WUwEQsMVPO7deCY3fq9STSKrRZpma80/
zyRKdzwY7XghFg3MaZDHjDeefCwQA+kamiUSj/9qxfilZQfo91PKv4DKIMP1vs9m
fXY/61TGVbvyJ8bfaPvMHJiilxicy03UXi6rPivrc9E9vr0sf7PBuvzxGOKrN8Kd
R4xsdBGK6luhDpwjcvIiLYnlpxeCzeqTsqraLoVecYj8lA6VyLQozZuavZNoyqIi
tBnF/jVpeka9o/ZZks0NJK53l/MsWXLZn0UpGBogKel4Sxu3ODBTG4TNME0JIWCl
GubsXZ92HsUntT1vmf/r0q3PkdUA/WG3eImqAXPzUorY7F7Tj83HuKs3yj+LQXR1
NzrgvXZj5Aog5BaXeNTfUhc5y1TIWprqqChaXraFtusqLix5CTMW2XSLuY+pX88P
bgOAdPfw2Pmaufd0JYPJdM73hFkNjwgmneQyAg+QRMZLAhUVpxUhihXzjT9NDL5D
+gB2jxRAG7xEGkuTaMg9wDb5nnf4fd/NKqd7eYd3ekkrEX3/FKmBNtuIL5k8luYR
tIca0IgNllyEWXLxagjnhmdBHoDWALswqmQ/wBYNfDWvYNUypQ3wPMnrFVQfqybm
HlJOVOOFniFCMZvsA/cJsAQ8GkDKcO192QQ37Rf0wtzPSxRV7hMhGmYXaWeF0hgB
fXzxHEy8tIJF5QkVBiJpz5up7s3Bjy2xFVCKD92IMgHw/otFqldyYNBHzZ3BxCCs
tSF+6RCWDKqaVkKwdr+49v9ILPfbwdb7Fc5J+AuHneKOm9KUmbEPciuuqAyK8+G6
4gyVYCoXxBTvc1YXrtk52xuGrtwGA/Z1dCcWTQdIMaEH5WskuhKYqlQoi19rvUuB
EUyrKJJKwf2r/wTmZNpZlv+17DvG5qAmsFVb34Rdk4/fzcis7oLkTqgV9CmNJ/Xm
qH8ME/HaKDnIWL9t/a7Hmx9RIjNXB7NO1wTJeQVphm6k7Bvde04uRaY9+TkQHL19
kvVt3wV0okx71ujFojnCn9XQ72xAnR24dxB1+sS6/5AninweHkcStQxOsTJyx+Vg
Ae5itEC4CVVOuRlFdSej1KC0RiIwQXmBC5qXXzrmH4mYwYjfyGY8UhFHcax5Pmtq
/VZMpjm8rvo4rBeuonqVHKuHVX1YByyzdD769Um/9UriBbxHARlR5sCYkBqQoEgi
we7TzTL13ki+oddKZU1IG+WQ9qpBe6E0T50DAasXh+mzy1m+ySij4bJZU4/5Bg+j
oz+OxfbwaGIHUReUk9GV1UB1zawZ6tbX0CKmKhKylqEx5fjerRMhFoWJXl1HrFFj
rmeVi4quYJJaD8mYsQybZItlRdQmyu2ITQYA8dtkPYCS9i9l8xct++Je5TZlLQur
5xv+Nl2z6wYsOy5SaGXXJelocLQKWkMHWofGphn5IWJE5MmfAMz6Mo2PbEc5vbq7
VQwLmJNPVB9ewlMEaQ6HAEve302+PW1+H9Cf7NXwHoSqBF0c9Ctf7RYXUs6oVDdK
uX+yY1hGbl2lYFNQQak8XXjCY5pLtq0ptW/TtHHolfMYuf1jhdkbcYDPdTWt84hN
VqenXyftw5UhEWD/r8Wo8JtxraVsspqAvYYNkn2C7Rd/aI4teI9XdjE93bnPEp1v
gQr0g0YXwS3bCANNq+D7/4CN/a8ZAFTud3lHrzy+FN/+2X3nZXVLyAegAKtLVvWp
5W3YZ7HttSDIlqIyiG89x4g6ChcWyma5UE7jkmJOLlxB33YKDUi4y8T5P1mbecxH
VUXw9Ugv3qp7SAiuX5LO0ko4aylNv4hJ/teuHdO8lXSC0MO47clFaiU+ndAN/hX+
s4yIDKRIMfu4cd+ZqmouoUi2HhQG4fTcnsZTPdL3vBbwZyP1AV9bKC5vJ3rrWL5g
TdLeblD6EkpUxl7G7YDrALH/vMA+RFhPvOd35MDQT9oYnKU+8KviYjDl9Z0WKWaH
OIdgi2KznZ+iEX7GdFuVdrrZ6HHrjP97b8aD8bUUseA1hce/BGfgiyeqXNgv0eJo
A8wCMxRfuyRkqXpo1YxtBZb4kWpI9NPOJ60+n3hAdgMNqgbV/bGyopJELUoHJGyU
cchPja+s8QGcvo3IudG9GCKMsDHx0LSL36LVV5e8IfDXm1G925Ll37/vXXS8Hkfb
VJCX9cvi7m8MmvovH0tjcEmYEG+mkpsl6+v5BngZ5P7FGDog8V9Itqq/YI4c12as
jpbV65NOi9Sk2WNid4QND67urN3T1EJf+HbpAPpozrt3rHqsWcz7IgZDix/uN6pN
In+RbFWqBmnX2GKBI6CasVodcCqHc9OFer6I6BFyRRenfYcbfHHEzFuDG1VQHE2s
hictZu02sZ6ffrCge39kySnhcuXZ0AxkJ1SY/M1jpYqbF4itkptgRmrMqWhigSy8
wZ7c8khvvORJZKxmFUq8tWG+PQL9SfK/c0vxOc7A7e33qJ9gIdUXUL6OvgBfgY7r
dv89vEVaCpuig09RXdx8vJudgWmUIfHlEf8WcDq+hBQaoSe4AAa1FhClm5/xctZd
1tp5i4d3N3RXdqQnW2bHtJNpcAOVsEChIjlLDcHtNcDrXd2/UsaeJsBKFPDvDmIN
grJtBH02kb9LG9HgefnukppnfZYxkxhsy9dNBW7ZvG7e9undtHjyk2JlyOQWhSTX
EFKdXpgrTPDMw6u+kHWfB+e/a0gwA7gYso2SElntpsQt4n4/9W+IoL3T9bjk+nOu
sXSloIn3bSZCIquWlKsk/LOeiqzqIGESLNOEmEP4MSMjU2uDzzVqJAWld2EkGfWE
+LSbx1iJBUb1eH71Ou9IdUacQkeffZOzwa0xaUPHdBydY9s7IdH90HlzYR5xUpSd
L/R6E/UPben01zkUr+nLpuYT/9oo2/1n3F1o+KMVBRlK77UjGoyAQxibuEKcXcvn
965ej3Ml0XJI9DZ7wrDjq9UsBQzL3Zl26no2TszFuSZGClmBsZjo1z8lYyAgoKV2
7PTW1ZZc/E7Fiq9PGWfxjrhiINrzLjwkfTGin6eZjwYkDd08vwb2WH9dMUsQ4i6t
lvBPd2SIser0SyR62NzCaOPfr3RpxVPs7tFuIWPmx0E+Jfakv7+hc3brAKBygMfG
PxH08j/+Ttp2/SNMxHoFJANCzXyb7uAKvI5YMzGcZJ4yowvik8mJltGBUQEul2hB
NEhmR5IyEKQoBwln0rsb+iiYhJRGWAwLbM7vCtKdkzk+SYmCbcKNlHOQrIPRanYi
siCCoBA13JliER4rIAAbu8eg13oXMxhJAeBKAI19DE8bILF+AyXpiDHzfb3bXnpk
vWZNO6hqyOV0auQzZcTBIDhMIpBJN9FPJ5YzpPWA3KZ3HOUE32aqdrruXnEXGQ3D
Y0CXdjxL8+krUAI2AbvUR6stAbLqMveku4DgB5UBU0+OxKeK/HOPBi6WOm14BlgJ
FuPLCKuN9AE5rzSUHcxWC47XOOL0FaPyNBr5kVBTAKHX/h+6ziI0PjeJy2QR5jjD
p5KJcwXVrcykPozFQHK+K0GyjgWJDxd0vt6Y4gzZXYBhcqnQCET5df2uV+f0Gzr1
R2memIaVJpmW0P0O8Of4npaDIF478Jf3PTFs1wjNKB9eNJ5UZbChWj83Fn2f8mfm
JObzOe2vFPhwW1fe+9HOuaIC/NsVpt/xayQ2tzCDe1YXcGD/kJFMbHBSYuZBZsB4
YTZl/Z2gkndB1A/oG+NuLUYXjjZYfoQ9Q4ddXOVAYFnIo8SwzRleO3seFYc3jnT9
CRbpgrcM0aqdIU9NJ3yYeZC/g0mYqhqlaP+ScxFKpnGzZ22MXhRgv6uXU5rZILC6
BMTV59km9ovetDAzmJvKeymtIz9tWVCdAcOjfZtlnulcXEhnTjLf9GkHaRk0SDJM
3AlAf73Zfl+6E44cRXer0XLZVK01qeiJfD8406YTUbJsAzJvX8HhHlArPyR6W1CV
AIbHouvAzRG+AwxAITXtw8DG3VxdtNjWRIZawXXuwkxkmG5lBpSg3q+/1sqw3zue
H6Vy5B/KjS4seE0PEM+9ttIYYkmoHTs/Rmy9tzB0CB1cZEzMw8YWqzpEOxjxAzTV
eMeD1mmWTfUN1nsxXCJC3hMs0hLxi26nv5P3+aYGzwG4+7yYXLp3OOVfwu8nbLee
BuOHag7Xacz/MnzOyqAIBmMAHLMijFv+4CIn52e0TpD7Unf0wyN0LhttOhWkBVNM
T/05NV789LQuz/E+d8GfUq5BE8rajhcn5ZmXbwNB6eJKqkZlbcbZQry8vOVjiP7t
OCxGTmKJJQ58UPEpfaQmXskM4i7577WcQnhCbESz6Q7VGzZ4+fzr6EjPdL8bmDr5
MBeO3+GkbGjifo4FQHlAvJtMvrOEAt3plvaX7UoA2UdntxP9eT8bTpXqs/TI2zmb
yXannr9EnBTvA/pA83J7ff3HqmPLP4qi0JcxdZewNf6JY375UwHpO5EG6JwSmUbo
gNNcX8rLjePjsWRu4pHfiLXjAY8A1Y1/U3RRBUUCLscXlhqS/Pu6nGcydPk4rCEq
TgvFpqyI7SE0zTbye2zDp3wIRjFOMG/D76xL56PL1sqp+Y3nUW0i3LsUIu12kgnL
oFziOgLHyHNeWgG1eJ7TKMadJISfW4J7rydxTrzmab4a3v3CylGQ06dEJ35caSVi
7gGfBKcULgedwKjmCx4AW4hLVSvA2Z9YOJb8ivznCOlp0aIXp5vwGxBzKtWLm0g/
7x7PUpKDAntitZjASYyJFi1GlK2zUrBealifcEKP8O01BNbEEUJSEP5cKiAL0Zod
Bx2rjcGKy/S5Nmc0QcZc2DQ5lHwiu3Z/L8Jljb5SpdSTXZiF9hdgVEWmECUpFYjh
U2S7xvMBmKithDhU5ScoJid/1k7AdtUCZlMVa3LVkNIrQN4AkPffpV0xA5zmikgT
TM2h5S4ssRblBi2wEfK3pzMsuytgYjNxQMTOCigr/H+yZpxR9kWPqNDLXhHz5MsV
3RhkXN0AEoi2G26KNhFjDxDaozJXydxi0A2VU2lNEqKhRPuRnZREMDRnm85q277h
YqRXThf4YEaBlRUokBRbNRpQIRf01MB+AaMhP6x3OGgEDqD5H88MVqlKNSmGw0KX
xnmPX4RIAZc/6J5HO3Z5oWW2c1tWxFdQVzkxcMmO7MaPnyeCLcYyI9LocCpH8EBr
VW4rRW8XcUVKVE/6QfPoeR5UVd9GktCthoO1K4P3oxhMVjLL1Ij8/ICUP18uU3KR
1qzuNQwqhUSu+jgOt2yqHbFxB+kRIVZQjU2DyNziSdfKfCxM09Q0v6AJg1TaLwmx
BquNyQpOReOwumtKw+iPQKRT1BDqhmFJacHPdLOXOmIPEg/Lxl30xsovvX3j2jqh
a5Kkz2q/gbesTm7gaOvDbEZyvKePbN/q8+y2ylhmIjFqKZ1DdjdpeAJSnD9TZN0i
QG/QmTYJRtX4nkSwNdULUVIGWPOfbq9GjyqIdDEjLoWmB+J6kcqhKvVG6X7nu9dD
j8ON927D0dqExt7P7m4HiwfYTCtshZphzeClXF8VjIBLLS8VwzXA/SDYsyM1cch1
FjDTTd76ps0L7AED9/5Ekboi6sNB++Ft/Mqe9fSwR2HMBJPPma5RA60OjzsHZI0H
F+nnAiumOPZitt87n3kZp3fKox+ECdAmOzFzKgnQ1RcU7Zt55mWX9qY55nXNeV7Y
wDuhdh30by0FLy/19+jzQ99x9TvSvGkoU37lqFx/ck5yVf40pJPHn+kxV+6KmDVh
GBBaFXmEkAEqNrb2tTHXeNhC50tYYgIIf+j5eDe2pgL+4ybhaKuurW4Yh9wzBPL+
ilZnr9Ulrius2cEDpcEelFKPisKc2hUYUsSEOtvzs2nsi01jIPXGLN53LMWpjfk4
HbY/bZp5UbInvnY16LQNB5KRTalVkhGMtZGFWnnQRotPF/nlHpbGuapyHcDORBs3
388aECEWF/b6U4udAUcVupdEyW+FBaBmAT1hoOVQUvSPOAZdKdbPaDKSdPxzhP5r
e+ua/E27f3upInYjA18YA/luSm4Ym+AW8TnJfSQh/cQKSCk1xzLZvCNTrZ6f/Eqt
VR1J3AzuR+cGt8nyzq/kif1hNJQFq2RxHVPemKoDOJJERRguPQmLJcJKOgwR8YBS
/AqLiaFwyGT2Pm+T2eDqbjOSlp1cbcYrrHiPiFcs7RI3Ox3kDM3ru9LdV2cK6XJn
bjTaum+kEwt+s8yT7qLlSa9d4caivF554pL8aBetH8rL5xLaUNHio7w1Qu3ELswh
5yiQ8hvumXrIOTEuKuds2X5sggYneflValACE+PJ98zZhH8bzTgWPaju1LFy7+rZ
3Wg21tQpRhZB2ZKjd5h6XhjZ0RJJdHyzj4mLr+V3hj3z/weSKGJtYUOuFP2q2Zvb
Tul6pflbkEaf2cTCMsqSpAj0U+g+TTBkeg/22RCiE8t++ZCEAsIcbYXlht4apOe0
t6dFqolyAY16PQaQlnJyARfUeMcWHfo3pcr2PhoY2QU54HeFeSLLumYArbPOJHly
DgFog0hNGrr1KheapB/K3owGi5nZ+8cPVZG9asLizpBVHY0/7EFi+qJxXU8eac5H
BX51diTWoHH3NTBcznp+lDsE0Juuu2YIa3+7QYgb1CrmsJ3YqlRL4rM0q2H+IUYk
aH2sZFDb/K0RH9u8B6qSRKgE40pwa6ZfjftuYibsKo3eaajq+eETf0xs90ncZGl7
xnAyZKy6D4BMg+F2DNlVmoIOuRTREQa8V4NQtZ9dCtRjiYurgZ7HvitC22xS/1Ww
t13sHVYC+6NUgCxxnO30KhehbleV9Q7Houz4U/++rsCJbmdNitC3zkKKW0+lgY2m
Bxy9PYgy9LUjNbUjXRP3NX5bCn83ReIyjjISsolCE+o4go4C0FWYSAN7msUVvRg7
ZDRx0Od0dQOK9776Gdkl1wHgQAsry2bDXPjZZzJ5C99ZZc+I9+m20neW7fO6Rjo1
x8U2ljf0Y49nCazgbQGpdAtRABMCmdYGxwxsPwua1m0iDnZFwSjuOztKM80SscxB
fZ5t1XchdibjUzrR+97K2E+j/5lPgwvpJqzKebwAasmzrqtUfJP4P5xq9ykWun0I
RzbyEQQR1j7Rak1i77cGir9h/yFOGauIImyBrzX7/lTgVqLsep+vWplev/sBWXlu
sMBneTqs+JvJux1v/RvhJKITDDI1Ra4viIoZCujy4y+hAeZ89/HNLPyM3HJzOesK
JOtGTvI2fdfoDQwIagHYJ+Pzuo1igl7EHMXvLLHKEiN98MiMY5LiIBh2MrEHgdU3
1h13PwWo5aKoGHtUWy5JzsJsvfsr0Kh8R5oRwV2/PAHKMfegUhhfbKuvbKHM49SJ
iq82J1riZIHxgYsB/ZPTGKWKsqx0uVpRS4J7cp5AbMVBenUMbD2KJ7D81lWNjX6b
f4o3UmMcGCh5Gi5V585Nep4KGJ+vq81v8yjDqI1mNQPEaZuOhTx1e9NiSu3EpvPt
Ey2KozLZDDt11hNIkNOjBol10BrqedxhFXqO769RBf2Vos2Pq16in8Zh8iCYpMwC
CvJmxEEVZO33S+OcHtK4lqkPfhHc6FpfKveDHE8ftTT+oSijPtnKCDN2LhoanBub
6UhZYc+gDMBO7uAlnLOwWc4yP49lwB9cIe3fU7ygQ2Kj0W4YuZCPUl1H7A5YcE7j
oI3pidQafDLDYxWwGGaYJM9stxBFkiyDxIn5sk/PuSGl8eiJct/nUJqh/aLCnC89
IXv+5f3lYQILc46cpPqfPqV1mTMlSmA34ba14hoyf9mPoDUdZK9aHtngimAWyVFe
KCjejBSNuAd3rYZR5N3QO/1brCcdP/68U7DwMHT3Q14/xkWIGoPJ0brWID9EpbOT
Fyv59d9fqqNzAzLFoDfUaA1p37qCyOPeWYmAFUJTLTcGaQK8yaMP4fnY/QaY2fl6
wGH3iAD8XLe3Ehi9o+tOHxg9iDG86MRxCSwXs9ed16ynMNWoHs8jpeT7c2k14rym
t/8xqSVyi0M9+xfsj620JXrdCpOiZIzk/HYcpSk/QGWaD4rGm2/HSF5uPi7TMuZ9
w1cD71KYm20AZk77Rl0iQH5Rs6OUwfiZgALPe+2l/wDHozOp7pdueOXOy3wDGb8L
UtJhqIfIqQLhVHOrqb8+4jRSxV1GHpRGlK6pXoJzo0iQ1PXzyWDPZub3RLxd2rVs
III/eN9/yIgCGo6GqxufnbN/eEi3iMckT1mjSOEgUtxeEzbByuayGlrwhMFOkoAD
/zteD7xYTF78GDuRuaZzz3kG+iEQpSRhqKE2gkiNBGwKE+jsFVJMRcNWslcyRRvq
Qaq0Kq+2dJkKjlAb7DaATqkJwvsVnDOECKgxkcywm2bnoWbNlxgROWWU20mGIy7G
ezJbCYWt0RMz5s2kCVfv24y+8D3y43HqiXdfdH1T83bcMtzyT0ZN0gVA5MQuEq0V
iSV8q3JZ4WiAz6ujVXkEpBjinBaVkKhqHnev3smjDY2updaMKXLsx5IzoCsgjsr7
0xhiOtGeC1Jr73+ddm7J7XPx1MDOpR9ZVuo/pmXk5DM1TguFNPSTFDwF/sj+G18w
XMd9o3NBd2j9sSopjaUqqm8uc/3k00G7WmuqXGOTmOCh1Xpqmiya5qSh3KkhJAPX
83pYby4Hqhlw1nlRPYpfSGhWCTANvSWWb/9rMhaofYBkdSs3UzyubPepALFCG1+w
T7gV00aFrWByUaxt5uO/lmuZnNgq7lOIvBW/abYwba4jHNv1HmAjOhocdoXBQ4CX
7OZJM1fLu7O9TQEG0iwNVvQ0RmNqGaL8O+FkxN+cCs55Id6XQ55tll3y45LGHJFk
7+qg4h6gCiW/9IwNm26MsC0l7xGOqROs49e247igxxKdx2EPr6SGx3AnmvU9+IsD
bUK/Osz89yuqA82Cb0qmaBXRAnixta9Nz4TFNXhRa2JDx9+6T0exYn3bHUlJORg9
xW840iBCUyguM8kZi1VfVchSrmllWYxWvWVOgc9zdda2lcpy7Ffugk9XBJM0W1U4
OZrZIburI+o8W1PeKRAJO7aMORv2+ZVMrO6dK6DmxTvxRg0DP0wQgozFhNDsJ4Ym
+0lc84/hwu0RKFvkag/9cmvxGHY0v0LRIKSJWn8PLPV/OafZBVM0ywXqqeKyWSH8
+EBku//IQIOU226UoPsd7VNzTLPnt5PRgFHqf298SJa3CNy6Iq/K+EveHGdpJ0l3
BHCZWqwhiT5dtj/8/jbC1Mg6Z01Gxk+A9fmGGJfceuu28RuMJn59CaLZRftgwmkJ
ziMG1dSlFbChHDYJDg1fXyS+4HLW09xKAxA7KiQaBmE6KcbYZaSfzKPrTMvqdJKx
zbz93vRKpFj2ox97xvvjmQKvmfJCbkI4PcwNu2PNw2kebmGi4JqaQZpyay9uhsNB
Aj0YywjeUdwNcE94PP02dMb1eAdX3n/l+9dP1rfphTIxtUrNv52ksKbmD9BS/6oq
GZC7o1lU7GednbADOJgP0bSoaZRhet1CJRk8K22KvnvIqqEo63LwQxMm374kkA8K
DjjxZ40KE7sInxkwuWf5DnY9OSMdwOQA9q9R3ZTXLpo2RZBT8AAtzkCv0VgmQHz3
RMef1V0wr+h0iqtBgElT03oOxMw+s9jT13lwjMFaOYiEHmFqXCKv6pmMTRIKidrJ
IFgCG02fEukEZZl/hslHviZna45OIK6AYVcgcg7DdpCnH1W8l7mE+7kX75UQrNai
sX0xvOoQ1HQya0RXcoX4LWwRkODcTiUoqEaLoaVo/a5SQUuJPO8CpVqZtX8ZqNTq
EvmqSc8jQL7nUt6H1m+nQYBuXLTY2rMnJYwIY2bx/ktH3R981M8x8us0R1zHyahd
QxvnZ9RpgC2yPc/dxM/NomxpFW1n7Pok25nZ2yhqF96lEGTA/b8VGzArtoShVCiK
cztBzv95gSvGjws6xnN8e9WuRxnSC+USzSaDl0U3gGq+u1iev9WV3ikXembBaOtL
VF9WvfqsazJFr7zCAiyAbyZVdC4PdQJ4a3TufqDXS+h+iFlCH+3HwghYkM9Uev+5
1phmcsUE+eSLfzbojd6XaUie2MFLCnxIC7fyjx3u8Wq9uUwUEtEW6jI+3gwqMl+v
KZ+cooTC21uTW8rhYBu2gr6SHXCv3q3maCUVzLuTSlOKS/cJzLlsAjspkc3zpthE
j8TkDOMzmIbfP5W4zBZWWGwGrvoVEzewYOip6fT26PBVd/Ck0iQmVvU3x1yjUGSr
nCP8KeNDxLrF0n1gPOc3tBA8ZPXhULGJwaV0+wJasJXbXLNwFU6eElv4kXYcRatU
b1O32DYaLKQSsNZXRWyRTtCx680F0ZFex6c7h82MckE5Gxf4Rhj+Dt9rkmUbd6xR
RrqExWws6wrPNhLtfdyfT9L+67JEOTncbMGKdLXPlGpnHqc9FsGtJuqWNGPTjaLJ
lLv3kdx+bT12ZcVEc3yywtZEQFaCZuLqmYqicd0yt3a6wgml4PQP2NDJCbWB18eX
8t2WzEXHTNLpXqCqxqgHiLEajiZIXZHisRuHBK2k4Rm8Ocpts3vamhVEw6XRkBhh
OXW8rnO2AASkiXBMg6ZVPkq/tiJukJAyYFrAEJECPmJ/hZ7MGM06gh9HlifkM6SL
6oPDwu9W37+PtzO+hhYZYA3iKDu9vOLWl0jDhwI3eYyPWQsWJwfB9HBZfQARQNt+
jjj6fWo/broGyUZQDWqoh2s8RiUYUL3MvWmE/qAkAW53PxL6/zScYXsjORJ3ipBl
6RXAEXu39A0Zpuk6mabAqA8Af/fjm3s0p/N76ytl0fJ5KRlfDGWJALbhWWrh+BQK
3DaksEmdgUZ8o5M0fLPNvkrtni+5ph7dzM8pMCwPxJagxKklUdREoWhYyvymPK9+
5LjMAvvzzXsbz03WIYflA+466PNn0F9FR2Ow+OeAxRKAEutNqhCZtO7SY03DsDcD
PiIb/gfROs48q+hZGL2+6eZkAG1RcsOqLnM44+BMszW4LvTAh2qroCc+qv3I4HY9
P2j/An/wckKv4ZilP4l6bD55hWQ1QYFc7sYPRPyqGRE=
`pragma protect end_protected
