// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.0std
// ALTERA_TIMESTAMP:Wed Apr 26 13:33:40 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
dWY8hPYHo8vMLd2KmPg8vvRhSSprTzYoLqnk1q/E8c7O2/MP5HNkyzbZSTill2CU
C+joWGDeUND2S9aepV9UAO3K8E6lwDgKu9tHCjul2vOIGLQBfxiaXXq4ie/g8yIp
n+OYMsLeuDqT/bpgZEakafb9tukNrKWCj/rz4z2w4pI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 1760)
eWM1oCVVNxchAPKjTQQCG3eakVymaxgGkIJQDaO6vgp0527u7m2Ro/su+joUdXe1
UR+Dws4EnvUtvo8sVchdHUYoFyyOlFibWaaKo5q8HVAQFCzt5LreoWl2PZWwUgmx
bl0LI9I2xLfj+4u8I+ZmjZvEtWNwk53EjMGoHkglU3XmNow93zFuJGbYIVHP270K
I3ayZwezxIsV6r/u0B/cP7+kpazrA6e/elTr6H3npSJI5AGIBdcxNo0n+PQ1kdXa
WuKo3zyNb315ib1+QzTnEHqkXHFgCl992Mu+kAU/MjMfMhqy/ejhDomqpMp+aA9H
PlidB1XlmFloiSqf7Nox87Aw1cqwiJ9E/645rtykrt/xEPZLv388ppxvZsKuloiz
ZC/4PHZxtlrwtgYC/PhLwSZAmxtc2IAEAa3mFAT6vP1XWVoLDsWnmyEtLH23/qyo
R5WWmuFZZlI06g/vtDKz3fgXsBnU+XLOL47L0jepyQXNVRvWrdEOHmmg9BjYJfd0
BT3Ifh0wzwsegNwyiQbKCY3+QOR/MsfeXwN91YsGeS0N3SjdWc0Ihb3geEBw4ikM
00qhZi5UJ3MQBN2iwdaAubfUZO9CHkDgl8KlQls7CnCWVGuDKbz6jl2TLP7H6pQV
mOMWU7Vwlre8ZXvsR59mZy7G6AEwbe5e4SoOf5KWaTr090DnbcE9UeeJmBGInVAD
JJQc4nc/46tGR2CLnOUyG1qBG2E100uFNSMGIQ8TUe9qfRyZv1Fp39eTUrtUdc5w
aAG3zpjRwHHFDBW3ULZzYyzqXBS1y9D1codyrydvKbJLJnRzH12G80sKt33yhsDp
San09UfBMXKieBGoxxQrQyhjsNcj2l1borz6Rw+X0duLXyIHeB8XRLCN1s652bSj
FnIqwql9OvzU0dByLZn7lTMnKfK2CPwulEP9M4/a8RdpmZahKDvxWT974eYah1kH
gDlY0L+4WPN1Z6L/zTgUpXYi7Q2qqd7x6ymWokWye6MxdbBh5ubUb7hOG1116sF5
h7NvVFSaAaDe2ATs3fKtwum3UxjS1oIHtAaX4GXDwDY2w68/ZlWJUrWykoj16teF
zzFySGR1lN1K/9oiEoD0bkz8yo9PDg2IHWRhAQA+pESqZilqQEr0A7YGiFDKEe5i
Z34KscrN9JtBvwdfZK43X5ZgPjRt++99ooL771R05w8xYJywzJNz8edTCT20Gh3Z
sZ2YSvhSap8U4k4vrN25tvFpsI/GB6u3C8b5ghs2ZcRtvViR+e6OBOJCIuYhMKvU
GVpdSmKkvImlpH1mzQfJRtKkzjpnqAs0CrCcrBrBLazJFTSRaIkpWvvCXeSLCzgS
oJuR4gQZClRzK4Xa8kCOWCq5v8YwkgEr+obtk4A7n57eLYSYgvc6MMTTdtDPfkfO
58HsNYFwvA4W0bLRxpl/+MJ9ZwSQlPTJJx/uKTEmKd19XykNPXko9GBFSyxWy+BK
1owiREijKXD9vrjRbra1LIus5d0VFu0NEJI6Liugr+9ur70yVS9aA9RB96UkoeSk
e/ptkdGYnY2NgAxJAQkwlleVh/d04qzz4kB098GCulJBRhVgyIhFWcwkBimURrFB
m/ZK3EOHQAMXCMM50PxrmKAD7lNn8mY++JL31Dud/9rdOtrTMp/XCsrmT0su/S1k
5JvjLJ5mPsmHJNmS7xzHTuyFvA2XLLSpVLi34wFznFO8YhB3lva9vg6wdmgD76MI
9Ub8WvLsG36iMgSotIw2SguLxDXgP4qJ3vPLvqzS3iZn5DRvhV5mViBwVKO5LzKq
EEAAPbuKvqDR/Yd7HV7U0gmWngSUFtDqJtZouZ/svNecGR1TpWlg4pfhjJ0mjeZh
4rkSWPaU8grRk6EPNPBUorhL5ag/kpu6WqCxoW1i0eaoCJ3YcVe9LQ8iRmtmbnVa
7HVpGI7/wu27KLCMSBgdzztK8VnRUCxL1fLExbJwyAEKAqXM3pek7h+3MSwyQLje
t8yo+ktQ1+aR5SrK7HmZQk9mrNXg1+3ld+mpgr1yaLaA7/gANQ+U0uu9FT+NCSJm
6pU4mhvn8l/1UV6QZZyT3Hlaq3Gcm/ZiAwOWDNDQ0VgJlpJP22Vyr/Jv5N5LlIwx
RA1/h326166vp5f8+LEgbIrK4TJunAx7jICkX2OpOrub4ipb12KVtKDjGBhZl+tU
ZXa4B/O3qzvlg+XbIU6sfedczA5GIF8LJ75IC7l2seH0mlIC+8YZXCVHSd+Ea+Du
nut5BN5uOY394tl2iJq5P8RGcp30DU69sGGKnLTUXtFlnK/keCrji2QvVziRLyij
wRv3x1LeGH7WKlaAFczbm5gcpbxk1GzWuqOWk9zOmbU=
`pragma protect end_protected
