// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:36:47 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
qgyOJAdCxNHvvIk3A6D/uL8xhgxefRkDLQ5dBPkcKkENfHc/qnGiJ8/Epa6One5t
+5I7H8po96Wc/7eJWYtvLi6rY9td4NFueuwX8an8KIlACjZdYBwT6nvmiz9xZBVC
kfenEReDZQCSL2s0KQ604DYcgnONF0zzJFuSIcZ8KYI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 26016)
Ui4QsdKNqvTGyGamD6/WFsa5T6Xu7SdpnschW4hO7AhE1snsHqyh3V3G57+xf3c3
l59wZAml9cGgFZD6LXs+yVsq2N1IZXuCjFySthi463giEQYDVFuEz3saEwwDimch
mBC+SfC1e71XZkov0OOE9RPbs30WL0pddkaCzApwgQ9W+zX+wm/1MgllXOYZJlmm
6W1Kb8mN49lAsQQKmC4grbMbxPfXOX+6l/mxj6ltYSVii+Q8mY6zmQheXpTKJAHa
jpJyQbQqqwkrBGTpaAz/zWLzaKzFqcA8GUe3gerijo8BWUxxaWGeObWOIic+72y5
Ay4V+KCFoLdJtoxDYkJh2DX8lJWIDYYIpVikByIl6k2wf1n6aONiN/Gf0QrtmUMf
nF6PYQI5NGzG8gtbBUzXLfXJ+BjzDTq6E088/fqnyekI2eOsAH11qXrD6eYOeLzH
b61zFlnOWJY90HFpkjwPKRbuqTk3J0NKKZuRB7qPYfLRsfiD80nViFu34mqy6hRu
OG2Ggl9r12ae9Ys5Sq/+NWpu4YxK/5rH72aIZ0cm0xq8kDQ6vgtirDnxS8QnW3qk
jnLyOZ/EVFuHkmuB+LP1GSrsV9FCoCYOZWzHH9g6xFJFzsphwYtcIAMRuovZ1dsC
e/xM8d9yQ3rnO7++vGTaMo/R3Y5tuMO7jmrsHoVsxEQ8SkgCnk0Z1QG44Cg51Do5
1xKzRGq42S4Mfcdt3uBA1ODn8z7G+tqrcirhmrFWBUnHG0xoyCjMLkOQYQAp288P
vfLPRjamRfjCut8z/0eIGn//6rGVizNUFjHe9q+rdHMS6YfGMyT8V3a9SmKWAEvR
kKkWTHrNTZMXcqjVL4iL0XXUt/Vg+zf5DgpWpU+GYAgfGW/Cd/zr+aacjXGd6HRU
7OV7e1S1hJsx4kep4gWs0dvamVkDbiKDjvJGAj7u2U18nf0zxfD227Ic080wS3i8
6m28l6+QeZo0STgUJfFhXRAW+IOhYFnzB146Iwr8UVQ668hpnUKTpsQx7zY+d10b
zkq/iZxFjG9TAbkMRq5T6bnnYzN0b1/24cX+iFsuIijVBsnjlJOtBLEEcBDUIjEf
d03Lg2m1gPhrGLffjEnKbwMUV8/n15NPKUscvKXrFd01Wyo6HMaja5KAb9Drd46A
ndc7/QH2KY2uzsNmglCgG89IO8bsjPO1tcPs4uwrmGf5aaXb5HXyLS+OJCFOw/Nh
Mqss/cYNoTPIQiP/iagpzv8RmQxMM/7fJDzzGmd/I9qYf6IVqBUp3E3apvw9+85z
qy1jazT4g5IUhtoK0ptSzzvTn1jKcEZFBz7LpQf6RUojebaTGWgTIwrC3Tb3OXQm
+4ACoO/z/pQX9JJ3e2fbjFbuzK97TuIEvEFg6vszcl1IbalsWUnnRLwmEgeQpK2L
CZJuHTEKeOkWT3DvMc116dkFdEb6OsacPkVDxELanRkvlU0XEVNFdjifoZF4RCPm
ohk0QzwzweWidWlxwXMYxsr1dx7Lb5Low/R6uJFqgIwnKtWvY8gcE5zYPnzXVeMB
Ehx4WLiJVJh5e4n9ZPq6tUg7Lf8CCfh08NkhJnY7JfJGfBWsnBlXGtuhKBnif/k3
Qmq9uy2UnvwW9vM5oXQ7w48IIqm9Y5t+48hI8ihKxHrduSLbV8q69nrTqAo4rp1U
jfNcMbpstKiOuJfafS7vtQIcOqtaYTouiE9jB//j6QxHp9pZMQ2heICf3Ea2tPdV
suflxhGRkM2iElA3vrxQjE5mZh2mJ+GZhZGD7POecHgIQ0GskGEnE99VDGRBRioj
RQbv93Q8wXEuLTP0wKFoV56BCoCDpAe+Ep9H0gframKh+nJouw7wtnc9+IVY8MbN
WpjFuydms3HrevPCQu9c/XVDCT22+Wv/hG1Dov6dW1jeLAph6ObNxC5SFoeTN8FB
qCw0qHU3gS3ucDpQ+qcFi7Rtoyhulik9csLDkBfMHt5IlVrAR/1MdHCZZ/v+uVk6
jbgNYGTTgesuYhBJFXKgQ2IuFsY8o78NXcIMIUYfiOMV6050fzKeefQpSjU0ax5G
S/ND5NdhglneIzkwtB92qwxZPYer9Tqo9rqh9UYCL3suJpwPi58kXOeNjvDtRWNf
ZG8W4agglZLO4o+DbdnxgTNTm8XGP6vEBfSMBamPxvB9mXpohKiyq7OROxHaRDPb
9P1EAtxuX1iEVBsYliTF8+p6SGORJV++bjgT2JYCwTpN6jWabBULSIjYPlJaSodS
MT+Wo3lRfXjBR+WpacvjlUgHTCR9jPT9MzoHYu/mk33TpFcxCHmJX364npzpGCTo
D77r6xSnvlzpCnlDYNTZdhrG/Cc+LVy6hsBV4nukm3zOdydQbRFzksYAINblTGMR
3m2XiykaylJ7MWc9nFFyf6gAjHc0WxIUM+vRjlMU1nq0arCOjbtqaDA0NlF+disS
7twjva80OPkqn/zpf4j8akhJXwLeVKWdDx/dWc6T3sOZgsNFe0KSAXXIfrIfons0
leyUBD43hU0yL10eBC+38JRIDJRRbJn6w1WYLW6EPS4wxY3ln5ZscAYOWVJKqWzX
cCkAYdBJVnzTYS8N2RHQ5q3Z+Px23nq6/mDTudVvNM7RUoifey7+CUVab4oi7Bwg
tdH7Hd2uWW8pHhM8iaPQMtAcSDWeOnXVd0d5MC5RiaFL1OWinX2345+b6NyqJW1l
/iSAa6Mt6XkROL24XrwK0AU7bGBt+UBFSUFPtLmuyX2PzGIUNQgvHOEu2zGoN06L
6WM8LfIVQ4kLLMHtQ5N+wy7qZl9SRbx2SVA4nh9IPrH/KCnbMufQyeX0KwVFBvVs
J2WrMv9934ug/PJehtJ/EhfqgZde7wQbQzjksioiHv+//VpmrjovNdlNt9eCiJla
b+P3M8dz0pVwQbaG2KyoXm+XxoLBKKkhWSBc9Fux3bv9oaifGua3/iObebXHUr7a
oOocIlLdAYrkosyht+lS+1GImcTX/F2BfhQ9bpeFPDLzI79Qy/xA4W0pVLtUMqr8
G+mdUfuNLGR/PEoQFFKmONh0HbyFBJci+CK/WTc+UlKu0/IN7c+2oSnQu3tJOx/+
9OmdEwHphHdSdIMn7se4BFQPBQqyX85LW6SZAjocU9fxSyPOvNl8lZNAkk1dWOgd
fZx4iKmcVECKZ5gAY2o2S8H3tPBGt7hlQrc+Dc8KuP0bhXO+IuPwESKzG/7vIeqx
/45nL8Z7np8zqhP98dN8AJUdNXRJBvb9Wx75WxlGIqZeCtF3INQFoFO7TIc/aGeT
Mcji7u38oGiUXtw2res3In0ZIOoU3j07vzubv2PacHop57bcdvQD5b3KlraIH15B
WInLJvFqfVPAciwuu9DQsxhCI0omf7X47jAQPHtxtKnX85AaWg2xd7sBF0JIri96
AqsgL1VfC+rm80UI6g2JyxgFdCijEHeDrhOuXlI04RKXcFt6QqunXxWvzFMTaoaC
egHoA5T6GpfABAC0iBr5aasb/DYAmmtIpFqz4kp0x6QEctUD05/YIyOgYPdKVVD9
UUVm2HMPMX6ITIqqZwIdUfGKyVHdZBD93+tDsZfuSUpopEvoJkIR8XMJEs8l8zdF
Pl4Zm9LiE0wPP55YNP9fetXr/L8Q0Ss6IFpY42hRagw9oZWfRh3zUxcULYbSoraz
0Txdeo3zuI69KGFsIKG5Mv1zGbNaFDQZr0WYGRXJpaGfowhTLqliKZpRgeKIGk7/
nAJx5V9pK9k2NW1bEBC84OeFyEIOHhT7jx/8GGVIROUXS7CApYf/aSyFBCTsCldR
rkardYTqqLSb7+81qdHL/Q6aCiRam4FNWCpCdl6KKpbM9vzlw6w3CGrZI/nFbyzx
DDqYQcZq3GREiHv7Rjg4s6S4JttJcJXWt0BCcW9rDIDmFLBkRc8R6/bvcpk/oJFt
L436WI3ncUulHEHf6yRCA5S+sLskhT5oRPhhPevma8ViWCvWxPlG1uYu++DZazeJ
ryFn6gjG2k5WoAuIkgR7tlEweW17cG8y0glrcFlBM8b86vC40S6VHfvmfOQQrudl
VTSAV9EfDvUdjessMJcOGvgkUXnuA6s2l6mJ8d/U5v78poLjX+8j8zTqgxqMqQO1
o8UTNzVf52vpfrItCoaCu7M1SHJJTVwSUIamBxp9RD3nzXYOOvdm09nwnZrR/5P/
jIGmDSB/uhtfSBrsqv03m5PN8d8i5Mz+8yJVyl1kW+akZIp48wLg05ge1Ox/8+Du
SlDhT6rJ0vMFbasixfxVB08UZGcPwiMi4sZ80dp8ItfQXX5WD2t6X8Mqs+EIQEzh
KvmNVJ75BYABygGNIGQ49ETm90Vvtioyf3483cf0YXij0UUyeA7xSsDVmRffca44
CFKpB7eo6y8k0LMAEak+A1S2a4pArpPbqiAB94lK6YK97Ntv+VE5OlEpkB9BrZTC
mrIkdkfJYQSRAqTOBvyoH2tw6CZfJJaUaMYE3V8fE5qgPOsGu0scAucHcc9nzp1w
B1Y7/aXEyceNndQVpPqaQXaukmlT529NS0oq/ujDXfF7SWYJQsWLc78BbjzV2tug
xfCXpWqgEVZ6W+4KvSOr0g0il0f4TiGWmIhX+f2LOUavLOmcgq2C3liC+a1B4hBt
LZPRKtxsBBgjjDZfQ5U4rWEpgWWeQkd4LIrz87ZZkEpZjI1Ft6oVjH4um3dMWa9W
LDK/eKTIn3F2byrxkNCc6k66T/Q7fnASEK6cJML/46cEAZGvOu/raxzGfE3X7Jdz
SKW2ql4c19AzD9sUuJvf+ztMTjK+6u9Z/p6U+4O13+7YEicX4oLb68VJM+32mSro
8TCVC7/rO2ge2veh7u+Iw4Q/Y6hyo38gq47AatgHHGPDmwLxeiASiVhTT5NyH+Fa
4vF5ms77S9hCnDYi+CeiPVzxIW4Nu5FUMlU8c95Y1fz1xe13ENgOuNS8BdBK7eo0
FEHo1KTN+DMNYI2W4TG+X/OT/9VSpwN/midhMx9SiIHgO47AHEKJJkmEDPWZRD5o
GT/w6Wq9PnyKG+c6nPJA0iwv+GETZd+WIls9IS93sYzG7Xvf4HYDR5wMmJex9bt8
5u7xX0kSfXyAHMFf8zptVVuXD6IhjezMjiJS8IBg3xJKbmWfxVrqYS6TreSldsc6
WNEgFlqiaBXtR63uVSlQFk+bDtQAMH7yVEA/u4IVs1v+uy10tI0d6ANcaOdSXtUu
G9fzbkfyMxOk0F3mz+gXq7iJs3P34pQvIBcZAMSDZU1asDz2iTzQFb1YbH91myEz
JLvdTA/V8qSGXSQDD3mRR+h1H4e0GBpnHPmL/+FnVJfTVkxQb4dGcIwbwmkQ+Goe
mekY1iTALiHuinSozZ+XVapn4Cpgyx7WFW2WfWB2phxp2+pwkQqWJHHDLmW+Yrr+
3h9ikn7tv7nDfuubYg+c7KUWJ9MmL935kC9QBzs8VX00pBDB+QFxOYHai2LkvAoA
7wgPMvLQE8xvvDab3OnLh6Zr00DqsYrlIvQ+3hUK1qvQ44C40UhEPoHmAc9KIebO
NvyezOif6bG7Em0fem/O2Iacm0RFQg5arJGzaaRwGqloVPKWWshKwEfMXXENPM5n
4xmabpaPyM+jtGUNrsPnJM4AD3/u5zpEikLAXGCiS1bNMr/ugPvvg0Te/hJdT1o6
zicEaesDFqWNX5LT9IO3THr5Jl15xaopQmN9ItxSrAdOBY09pR73qj5y4GyEJTMK
NvfAHi9pwUVs3TU0005KBkKoQ1XL3XmBIvxCxyNJkblyNdfggC0xcypFQA0PzYbI
xnlmlbkwB2dnI3lnMXzHgdbbFbiAtyWdCvwJOXJjcipbvsPKIDezghrI0AZd6q1d
YYQxY7/2rdsxfX4Dx+10mR1ISTDah+aUuFeODcKJmwewKx7QRpbiGJp+AwdQdbhF
r7avVWK/KWEuePmD00B/Osra4/UszB4Z6OcH/zEtKSFLy9vsnLZAuzm3AjcNLKRL
owkz8MgaNXdBfBura3lT1uTG8+LJrKaEzW4YuIVBuenFi6lzBngAXcT9rdlW6Q/S
bxfT/caxgroZEOaQAYNtqWUjAgtM4Wm55NHwjjIkYW/5SljVCDWJmzPNok3PvLnx
Fo/DbY570caLZEwZGAOEvBcH/DR9dENubVaYAgYAigUlx5yyox+XMttjnpIDsXib
hMCA6Q6V6EsVducecGQ5X0sYifpjOuM8z7Yg1gcnVi7XtoxRD5t99YH72+UE1VKn
Z3bJYbFu76Xy6J4r5FAKYNfebyE1g4DZ7vp4fBRiDiSwRJEQncqzpbG95dw3ur28
hIsvyXokG44e4v5p4kBUs0w2qUY3wJZhBInvn+RGPf8vugofkTHeGil4NtBt7Au7
b1rJISPZehwhK6UpqNGIBn+jSP2CvKqlSixG/jw6fgszfbAO2jArxyHwZA5Z/yiH
WEKqAFgHmeBjk+5gfATcvrfyr6YxovMPcZr1mDyFWspY+EknRqjoRVBZdLDajRlr
TEpZG5ZGsl1MdYtzzSD//hz7w83O1+G1+YZOa5uwPTUFCSEABRIG4516Ss3Wt3FW
ao7a/eSTaUsyTkGjCA1Ycn7l9S41pz4dhFXTpP8S31XJ+yprszCn/8FR3bdJAaLU
y4/wHJnTUJMz0gkO6eZJRzS/EMORNIBuxU5idcSvuSB14gBcL9pp9z4SMdnpuI6M
pH+2s4irunu7g9K7aYi3+R1z8s7cVW+bfvVJCArmEfQndHNjvww1fPnDCFPV9CbX
r1m+WnS+ySoKcgDqWGLerL1YD/6X4AE2MmjnOixVfBy0mCNCUGZb/PH/rfJWGUrS
GloLI0CcAEzT7ijmbIEwD0+hBoYgDrtVVPG+e9Uz7cZzMwYm3/K4PmNlG6XrmX16
HmemOK0L9sUh8PN8qkDvxFyxYDeYLYdHcL+Z9TIewOZhTlQSZRUugZ2G9kPwLTJ9
6aqcNIj6JNmvroOuz3r+8bNTiRr3tKHCRrXZc96SRBHpkfhYKA0vC9Zia0OF2dir
1lYYzgpK8mFu2NAb3pPEnuzAR+leuPbAlr9IO7b2l21iNydi9WyfRNFLD1VGSfqO
5c92lgS37CoaoXGsJU8ETlh1NkLk1rQ5ozITm3z3+H7xvOrMrlvH+8kycA5KkCmM
a3CHNjjqo0iuiAm2tln8ukSOxIhn3LAkYCQZ97ZWtLx3Qy6tNg2XqYWu57dZUitf
ahk9eSChnqlYtxC5ITq17Yq/evI3leYq5dFAE33GRchPtlfC1KMx5hZ5ou9wM7wn
SZtqUTPO01HWShk0rvOmhQMTe/8EwlWwqQFpX9+hbD+bvS1J5jdtt1dgsjYAcdrK
6O1idf5SVhxJY3dvxhJjQ3NSIG6CU/8xvRC7aQ3oaiJ7rzO9ZRpYy79lWorWs8xL
4vb4r0hTu1GN8p5jtheJjxtB5eFD2Tcl05mavxNuVkLnuJLuRfGEdawUq1WX5n9i
nJ/ej0lfG6OVGa/r/nYJV8DGrOSh6jg+TsKe7D+TqsrbInfJldqnHznpQ7h8qwnW
AlbhGCYV0rLrakG7dvPZ039UC1sqqlfwtQkU0lojIfBofnhoQP2XmnLuGaVlzchM
eEhMThc6qFlXOhVLLBQUoRgBs/P6xH0M2DKHZs6JsTNH84TT3eUG7n0TtSxFvmlT
iU5HexnZbx4xHPbt5An/0/kMPRpjE4Q8MJYMwLxXoHd1Bs22076aGZig9U8ycjbA
V0iFeYIl+N9DJsY7iL/jTQGxJEE0Bf3KLy6R1VyP6o+U6gdhschgf6hmAxmX4zL1
ihmK1CvV4awS/qFSyqpyxeU4dYLnNcTLhkwHfJzTWe4W4fm4arZzt6NlLqeL2Iww
f/K2K6B6Ik0EsJ2uhKsAg0an2xVh1el3KPZ+TgGKh2NGJELFKY5Ce93BsA+XSiKb
aEXZb01u+9vE5wkX0fkjrWAMaY292jHFthQtdazpxd2bYEa7o0ykIkZjtR2tGB7B
Y5RyObCeAj98sgW2XQzPb2qMBVY46TnJk94/+dvre5HLxx3GZJiHtFGI9rzzimkj
tXSIWqwKthPx/JbkrO+QqXi5ZWkQ7Q8wrKwDEilr4x/fmMU7d9SRKuO+XP7h0IPV
3OE/L45nwcjxjnHAqSTWWhg+v7d96qS/IB9gMcOv4zhB8nBckB628rbhtT3kg6Iz
mHMRuZAEFuiEuj/qhgC7MWh60duR47K0XNaHBAlLXd2PD4QZnGQCfz5fhafaZ4f+
NiLH65/wB7OeLUuP7TDy4UzgWETvkLyqR4hDHr0vvZMDRts1Ghdp9y68f53yKrjp
m4eA6B7nlGHiltKDSWG6EBN/sIicj+05iazqkwU2aNkGxIHC9Q0jXF/xxQv6rNr5
ZIpSbgtpgG/I9RcTjYX3GcJIqhkVyFQZkKR+ZdbRSVBS8o6YDuvzl/p40toLVF/d
KA+43/CHPjdFUFmjpnzSMMebFjTktyLhiSTbEdaOfsTx9L2AR3YciOhZv/HkBB+1
1JNB/Jkc4zAPE2jz0XqVEFMx84/gfxNm1+MfG6llF1AAXkVdeAoFcv9cvs6PHctV
b3PyA7BPThIRtvIgjvfpx61O1MAEBD61QTw5K7i2dxKh686k9brrY0V1/rihqQK7
KveH062E+QH2Sqwx7GSLdDb5o/2fQAVOrG5FdUNVITZ4gcfonkSCNqtKPdGjNyXj
g216rOYhdK19bVQ/XWxhLCYxRzhpIp7n7Rz7OI7SRA/i02/e/gZTM3Dx+cy6KKRU
HTgMTGJ0+i5JKN7Xm/xxpU9Bj80wY1hTwi/WKZuLVpcFmCe7UBDlURzIbcdFL5LL
//ZmnpW0zH+xPKf1lglj/nI0bJvaQpqg0bwz2NE6lRuZE1feoKS6nw3WO9qvMQiq
fXSBzbMBlgP8i060WgBt5d16W4FOgCraMKvgLzeAgg9xSR9iHZYqnL5hH/yB9I/A
9R7oBjmegzM9I7mikbHS6X82PlC3e+XUrUrn/tELa6r29+sP9lZdGdNKdwhdscMp
uGHSl+Vc9YpzoAqaB3Y3PIiQnmsUbfK+2EThPVZQ5jkhLszPuzLQJq1O/Xe/WkJG
1fhmMLdGjXZMIbTZX4ejxX1V0HpNIOrilqGgoxyZwCEPalsdPdTG9Z4xlUKfcOCa
qHJD0jMCCwsdl0/5OG1O9fTvUeFawg1hqo32i6CwK4QTrA5RFPUDourhbckh6oQ/
5hyZJE6Hlk7y0vWqe/VYEj3yVZGCVSiX1Ib1JckpBSlnPkFCrI61RuY3SP2e/G1z
RuOUQcWYnTfL3WforjrGfknHKTlGR5/Hb68vje/Bh1i7IULFQ5TuWapsDu4q2IzM
dW5M1M9r5giyPjXgUbqUavaTHHJdpRGO3cmEac7LALRkLXS7sSirohem23Ug6R9K
zTCV+hg2oHdqSP7qqoZqlq/xCzseVrvfrt2FO7KBZT+hK1RZs2HjiCp8fYiBqxv5
KO9Qdaq4zIvx6/mTqn0wONIhorCpt+VaVIjuBtm1I8TD0xDBQUE5oF7klBoerBxl
FKHapEDxJmRJLjwbwa/fGwsZVypDnVPuAs3CcwtUCfs7+vziAYbayAQB5tZrUnNf
tPMozhsoF+b3g3CSse+9fJaNU76Np8CigbsbZQfjP7cOF+xL1umRVm0AFs+UoBIG
kKSfha2On/uTONd55Q0gH1Ah3KVHURCkiNW02yA6+Kfce9ixgGHjHZAgyhMk0lcH
Zqw9Zge8qD3ZAnqpP/WEq3NgokNbh/qjXf5mvpEYu9iAVCgvHR/KB+knkjoPkUrF
lLqoVxUeixdSVVAeSBhTV2dGh0tG+2FzrbzoEjgefdPGilk1hLZzgFTgT1sJoqXs
WRBiDv27tywn7zyYVJaYX9eX7I63zGgrpFp8sRVeimRgCHSILQ+fBAxrBk8Kcpfj
JXy2/hMGuy1rA4C6UxjCXmSrY5lD/EW0k1od5iL1mkXvgwDufY5Tc1NaaM4428Pa
zhTaTMFwhZw5UKGP7aQeeQFQr0RyyG94u+xYij1SWrgTab1hNg2tqsNGO4+DYPr3
iK4m/ub/9Gmzkr2f8b5tJlKp6Yn9OBpb5QzYN5q6C5M2D0rgvLfeGfbwL5aEymzQ
IQ9ofObQGzlhqgTk18gUrJ+XYiNPYXOczhsWPg3+MbwXr4Zt4AZIVXkTFa8KmljU
C+ZBYAKhyjGdBUj66v0XWquf1rp13Ni4pkok4qdAV7h1UtaHbExHe+XzN4a4RDnn
up3/gBpL74utI9rgncIYTgF2LB+OyD+XJxnGlc1k21gw0OOjAJ0teVOKyrjthtrU
LlgW75hVwj2N9cxwb1dlT2/BzNxFkW8z202fyIhGhFeZQgme32ECxFI5B6KKnyBA
fgdLhO39vC+hoycv+gc3OADVusuJe+EleOQBR1YD583rKFldc5hJ+ibQ4eS9Zv/F
A9GamA/PCunv7tyxTHTNUzU/GUzy74SRYb/hi/ne6vW2EhwmtlcXosROdHsDggSl
cahSK32oTL302fw+sBNDIrBTUuERSzenjhSkAfUmzKzHVW77utM2KLpN0go1u4xe
vfHvrYV4/kC5Tw/sKWL/gveFUXy1pdaB8CpmnhlLQuhqun7IZbisIFyFMTzTroiQ
7D6OIJUA8fgIEszn0uA8ea+jcY/bTl5AwTRJNke6TC0OB0P6hkKj+f7hN//u/YyQ
l4pAC6VNpd3sE3O0MlQd/sFyjxmQHDLnUu2jduAzK0ISyt4EVoESZ/7Pk+Gu5XyV
GMYdqUFWbWhCFdypwBRsXVhesrKCHcy6jItDupXn86LepFeIsVABfBcCJIRU2jpl
LSDyQpMuBkduH4zn8prQAH3bljd4QSI2Xo76YXJs7ypMjUGWrmn/Hifh9NboP0lW
uFq7GaSY/r4VLBSJWtix9mO6SLcii+mhNEzytkukXdZ4B98w2MbuJiROGDwsk1Vs
/uRRpPas+dwUDjgbi5AdrnXl56SELceY83loJ4EwjmO6n69pWfmhvKhsbgkRvbLl
177p+Ezz2mOgy5r4Vw2D9BScG/ayoCRAPsa0ckGoqDy3ZiiJG/aSXnzxXzzMSSEg
y+L6x/YGdS7MRZQUlOkGG85RE+YVWCfI+m5vNY80Nb+D4xbqFHyw4sryor8vOzk8
SuWGCz5BMiTPl+gySXt/VzC8jgIhWpnXCupqXn+owf19k12w/G4BhF1I73a2k+6h
P1DXxFaWQr4qlpWeV7fNG9nWOPhO+29v8MghHhvVJ5QHX6K1/Q8iL4bhEEyoxbRI
5mCnoFcT4UcAWWq48YuZ8pjjGQEPFo3+y9vqq901pHHwrg35jlq3Jf/a+t0/WAVJ
P6drtBhMniIwFdBbJnqn3YdO2PunRHpfz8u3WBLg9Y/4o+X4OhMEurlZoQlc+jd0
YH3PwR0YXOBHYkMUmj+A8/wlKk0n7lXXL8W9edAxNfn/y+xtKO9+wfyOuo35tWHI
QCexS1AhP/qxXt27ZBdaIrulS9aylrnufAgn/pkoMR4IL4V+FsXPPM86nWw8tPDV
NFpqDsKcUZcymokuA1EKN6Jd9so912BOnmCyQDpWPv+MJcAjjyhLpRorMF3DMmjL
naLRN+nwyXrhp4CqR35FG6iiPCN/4VVLXH6Zbnrg7YeJ3L8nnjPFcXctjNe+Ac3m
kwBx3qDJc/2/O2EnLZf1Ui0V5UnyfDZ5Js+6Y+C0rw1l8i1JT4gctCaFgK5wri4U
mnpPlI6SKaVaUAfS0eNtEwEwHbINV3xBsZP9xMZank7z/xqpwvFGWnoirAUg85n2
j8KHYQraAz/ywqLQ2cG1+yeoobIOQGaQS6bQKVuM0i/PXVlaJgO/f7ELudqzo4PC
x+79KJgu2qgh97TjmqAZ82UYk7iXqVuQWqUruw24xUDGTK0xurD7oAodWH9dJ6YO
d4W8RdtOVNu4AKOQntznpZRRDTHlMpYVkmJBzp75vWihCoRsb6Sfg/C50EMBllPg
rJXtfTJO/vrI7IRRbNi0pA/XCrSU5veis1x5hZwN+ZBCiSVI6PXT1NgLXK7s7QJN
N9+67gkRWCdhowawyCdzBkehS7hFs6elhAZCnYhfip9piOR5PsXvbkabH/7WeSM3
Bj9SPLc0ZuSks3Ti+2d9RxOaGkuJAcC8Ip9NhuCOU6rcL/MnlksKj2LXfF9IevZ6
zrb6oOPoiz5Fe0sf7ZleDcOEHsm/Mh2pqYvOLssg2SsegiZkIemIgOM2qODLII8/
IjxcUEE/SSxIyJCvSahVEI7phtdd2hL/nX3FSUQL9AF+ue+O5mwZQcCKZ9Xn0eEP
BCSJNHAC7Ajhac4ew92SrGOMj/RCN0yRFc94fAaEBvqic+8WmbJuyzbfv/bISjOM
7gVynp1XQAYT2bpqMI221XPP6ffPOC3hzNwLIJhjIis0plSEhjImLxcFbkJFoGj5
gjgumtKJTB4FFVbAfgs58p6JM+VBhoL5CC5dDQVgqoemW98nCApzEJKj33ABtXLe
OfBoxd166wpZtSdjIqv1dQr1WqK/hLbMOrAEzXHic+e1kyCogZQapjBsYCz9O76y
OK+Lnf0KLamiHZ+Ht+gX3eLyRVSU4nWeeNXk++wa4+SO3tUbZSc+dmQ0rjrzugLa
jYRUjaBoXMpq5cG5BdEEsELtYGy/iusWunBBYvgsQKuLb++jopqSyXZLZPETA77b
8phvK0EOSFBrEleDbq5dnMufEKXzXVkmwsaLHtZ5jh0uVAAQAKodRX3/wBlc+eCk
9BMXMUwO84CecHN6UpQTGsm5GU3aXDcpGsSWytVaASFHdueXSQDDqwkFT/tVutF2
5MMuNipT6gibkdy+sG9M3xeIbTAg2NvAIC/Vv0461bM6mGshQlCwwUpbl2WQwJdx
5W72X/VutxZvyZrmwg6NSmBkuMXV6SZBDviXG4TPJqHvB2cwDjxjUxq2GUtnuErN
azgEx0DjZWbeL58EiIBJDNGWTihjRgwi7qWLpfbWcdy8nb8YdmNvL3npGz1Q3dTf
fRkoL4ute8zXaFzGluv0T3oYODB1u3ofqqz/hnymdXCVIa187PtwnVmYWW2aGccE
jLzco4NwsM1YlNaAuN/GFBzeq9wM7FSDzc3CH9cESizeDlryhHjwthSJ72p/G8d0
1OCFe9ycPxG5ZgnAb2R48smb6rqv0xeNHnujIuVL8j+9yOQk8LDkCFLCPQ7s4z9o
EWXxGTDN6Zim7xMQ8Strgl0gjSOfqelzSq2QApq2L+gG7tO4uJj4oxSPbOe2Ojp4
jFKKhuXD7zM00z9mPeLNds3dBvBt1lvnmcZj5XoisEca4/Dz5SmIc7fpufGyPZp7
m74L6Q8peYiOj4vu0IA/09k0OC3GLVauUErg1GZJevmNkLednq2/buCMkxd2teGO
9Zv0Eu80k7DM+kZY9I5bdldOsnv9+KejsQ+c46mk+KJbqCSSrprxWtGmixNOreNt
9W61pFKADJRWPRVV02xNM3RawqhsutFjPdOnnwwgbPIQ4Adof/mNBQWLk6nvEQiq
XrmzGni8MmqPbO6Cg6w2wCFYCHzyzxRF7F4Uc9m2aU3MuCOlXf5UuN70OkEfy4yl
4FwHg84XwgA4bGrb0AgFI86z+Dw+izb+1AqnCeeLH5IsK0bcyWsFJAkJjdtMddOY
DJ/S4gHSKmR2j3Gu3JBOLeWhXK3A3FrO2pOqu8dXviWzcsmoxD7moTae3sOzmlwR
hdtxWQcRbeWMPSSQtSC/zxUQbSAOqCG8/NJSXxM5GaTmiVZdAzn1kqfB3kGVKY0V
80pP8hqJgsv4+fTSbeA8v3WSKRZxqiFi3pMF+I9PEO6vjbfakH2HOj65iqQjqeAC
vbcN+FYzrClYahzGYbhEsHihtCz00DfHjTUISETdAGCGOQ98eq5xbHpU5WvoqX2+
zu4lU4Kb+q5ExXd9Kk3QBVAGSbmVN5YV1+RWGyhA1SmV7Eg4pzb3cDLhytAiHhOl
cFIMbBUv89xArDC1XLLyjpZwuVX9fuSfRdEqpreHqnoMPlDPzpiE38zyBcQhrZvM
1zf/ZKZpQuj8N6fFC1H1Zaq/+yy9JZwqmPX9s5qX402KZmdKAu3A9nRR0UdQEzdl
HO3K+ZNDuOCQXEtUNhieXRXykrx7Wmnjl8k96swg8K+PRanh/7FAIBKbZdhf+92f
eZPEnnLrKMRQ+XR4LS/rRPRkXjaV0QsT6eygMhXCSIUT0IcwfOyTxvkr95hHw8zk
Ws84kjixckVTjQ8aPyFcMDb/zmxPZlZvIrfNvtl8OwHQy4p4ZX1652JPyStmpKRG
wlFWXx9zzkGNWE+3PM1yLC1C1bEj9Y1tQjkyqcbUhCFCisHBnK/0aEWkpuNZ3pJk
OQ1CvCzyeTVCtOHTWVO2SrASOvGvR6X89nL3F6bwzpK8K9v4q3ExY6e9yHIzkC9E
HROE72qgmmY+SXZr75VFt00I5Q1FdDrQPd/RW1/Oc3RYAdMBhtYYKGi2MjkTg+35
XN+9aYl+VD6yfQliFYwlWrYGhUf3tG0ChMQt2exKtk55Hfl1obQaXSZ7B1qfGAA1
Fltb9NV3sUzadqIpZ50+IYiaoAdTP5f0JLPERNcDrSOaHtFIAfg0aAG21Qtlmo27
bXHzZyNvJQxNwaFzhKJXmtItIBD27nn+7jM7uBZVuF8R+aHrRrRNx6YrC3g28yRy
rl7A4WRtZ+kNu3ML/hLQ/rRrNr5laqR6taGxggUT0vezimryZLvmcfju6zQS4oug
2g0sJeyQB3XmI7rkBLmLJu/Kq1h/B11KSjFV7zcBBY900qHaTfQYb54foK3iSfvj
Bk0RAI73qUEqq3HLJWbgBC5yvOIpaUUTD1JeOVssl1kCh7IGesyWzhXBbZ9S/K61
R7sdYb8v4GcMuLvfdtA3ICaASODV6F+vDarocVuqql9qkF1dJueFwDpt6+jcbgW5
ajHNuD2FcONZqPg2gowhZl4W+nncIcZWBOPseg7+mvd+72nkpCLmvyssBDXsFxtO
i7cPFQeM1/oWATzlRh46j0ElC6AiLkNRDU1HU0MXAxzClA57iqSMdGNpBOsBrHO8
bEWlQIdKjGIdAqqypQaIMGV5bgTvGLvpFzozU6N6tD+KLxOAihb6MiLYpsvCTNTn
7atcMlaQ+dkWH79QzzOcn8eeWdFx3YEnfNdDq6iWuMbTWV/qHF8cVWJ+Xx1ovt26
I5aoJS7YZWnzwca2rYZuYlW2mCV2HEYuGS8OjvjmLPZOcmfXur3aLW4N0h2XM7gs
Z21+i/Lq98OJ6KT+9HOVae94xqbqS5kbnbEK4GzQVqpy7pPwa0bywvNYvpTdiahq
Bt7ei7MjQSyYy/D4Z9lyzvolq/QkeOekFjhlp9GCBZ0KjUbhfR9UPNZUf4FHGnnI
t6MNI/O85FqZDLnZ0JAs45iynxOd6AWoQMeS9rSveZ2/CU8VT3v0DY2prb5Sn5qf
wcwjZKZ7tm3zncH79ZECVovTaTYs6fFB5b/vTg78mEwMY1UgPQXCGU3ZSZPIarAO
dpSL4en9E+9zdW0tXGAsdSLrI5qDZe8EYJNWAc8TFK6Fn5hJdYNK6h4b4PIp+I7S
XoFW2TTEvGIPvdypyt5iA3o/FteWHNjj323qSfLLQHnYG7HgLDhvT2/l0/x2+TLP
POXf1bqlov6gVBWNL2xgO+V/qDIsjmL+msoan7wEGtk0K2hEjTbye2TolY7zIsCN
3LVuT0pk/vCFWXK86qkUtf5QH1kUXLWiMW90wD5x8p6PqqdgxWJ9OQLw/qOt/qgf
IAy1qERuqfWwuKwHInbo5gIR1ZGuqmLDCSopC8bkwzYOTt56ntiIjcj6bvdBK6ei
arFogLRnprH4EE7mzJRBcECaP8nB1XPaRMgs1M+GRAiOaJctHeM9IT/rulSLaXFW
wON4iOCsJZDqowtgksZ5x3war7ccVFoM/gdbrXtroHCda75d12sPaRAhA+woG+gg
a7noQ3JoFNrhx0DqmHX3s42MNInkw4rMqfiXpjbFEz8uZ/6ExjOsDSywnD3bRbI9
5Vkm4K0pnDBl6iR2auoxL3/1TwzTmzx6MegHcLltJPuhvvekbGvQY3JfB9fJ0ICY
zMdAAVTg5b+/JAJHSVJFVetqYa2JMovOFj3frc0YJC0Zm/yFW0uELSFlSA5K82ne
43C+nL+vNzh5F0n525TcJ7KYaFC9mTT5egZr3cgB7C9InDz7TF9GN3OfWaQUkG4K
MUYiD/ZqFwtLhq1cuMyuplOFHVlvZ8Tmt5LpRGTlA2s7DFoVxY94HgRlmU1p8Iqs
ib6RR383EMypsBFzcGXXqk28lrODM2OsOoegl67Ja1YPkdoO/on7tXLgNjtee2J6
St+024H55dmyJQe06XmWmn1ZU4TRcsr5zViT0MjY8sFc3KSeZHRMExXxYoqCVfAV
Cyv+s0L6lCBNf/BiMz8wOK1zUoGuccpeDDjP8Asu3FnnZSGp7h6ukQeyvT2ucRNn
OeIE2NxG6+kSVqJJaC+XMB8jVbYMwzjpIOuo2i+bYYbI5HhQi8NxEOMnLyUI2zI1
QvFn1iMXc7G3hVOsrjYiQRsBsj1LvGYBiQNFfXip73nP/+OgCepEo+mCpNZ4GltH
AL0rUB0ZabgN7oOM7s6G5latQk79MLGZdoo3INzaZyxZdPiIsiz599X4Ob4Bu4eE
oL2MNZzYIiDUdHdgcXMuZxubTNoaM0Jz1If3FbYXyKzR7zh0f+Zh8Cgm9xe+AQ3X
Jtr648Gurp3wcEeUDvUZ9eZSUooXJLQfLjzB1CtY2NdzeHpKscIyvBJ+abZhHa9I
u8M3nUv+iqPwipAJaB6IsbhSFgJiI+oABy3lSKNqIBQ6wlZa78Ul3KjpWQx3RHyq
gptN6l9pd6GFbMiVo/VjQo9GhqmVt5V9LdGz/3vsfuL26r57khU/FZVIOm9823ha
eYVgezVTB+MndCnywkJ/8Nr24AfIQ9AQT8uDjnMkjO7UW0sGktG6CFtLUzgmJ6l7
O6tGxxoAyAdjNdaWnVhzUBIY1VWRWu+TYXcCrK6w/T15JIYVFAkt6YJeIjZ2dxZX
ZGv/pIiG4SL5KDDSIYWobICUsDALHRifv3jVvtl4ovMf/VKN4ncypzrxbZsPw6ID
G3O5ITV/wCSwZrBls5fhuvWRv4JMPu1tbq1Zm0rtxg62VPXGIwSfRZXDtLNGnSSy
rfZdI4mjdRnO/ddnVoHbV/Ld2xVdE6oJ0eLrRlyj9lWw5y2pYjNAf6cjQ7wzF5l0
thuV+65qM+Hniwd0ho83pdu5fzECfs1GwoRHoBaaRX7JZsBNZmx4cPGcIKui4OuQ
epPjjLdNhkhp9OCFwa4LgvgGGhkc8uU4qg3HSZfwAPFrVeM3TQvS/gkTmyWOfrtI
aa/PDUgDXYuxc9ENsMqke1z3Znk/lhVcRcxt0dSFFsKDMDO2ExKs/aGvq+ffv7Ir
AJKa0UR/eighhIeWuWrWoqx8Og+BAKjjJtrfMi/SOlZwn85tzfZPYujVNNmymmPo
jSfqUBU28kF/eK1HEunPb7tvud5Gr3+JpcOqAtz8RMuGINGNUBTFjJVlTqqq2tnu
dvFNqT7jQIHB16aILJzTzg4Iw7Ck3OADOrJTRWMRwt2szio/1ymySb00p3Mf3C8d
Tmtjt2/5yYnVU+yRiaPmTR8kMWo4f5jjJShlq1kLNoWsk/DPntgWrO7H8xvb3trG
hjyvAQQ+oyyUPxkVtsKl0O6mVCRclH+Cl4lKB1wn95gCJmZfBA/et+5f6sWnWTx8
6Q06/ru6t9xkYDwEj+amyVpv77RrXoFcwuhLv9ITxJKFwXCbDpRiGFsgb7OiAL+T
8WjQVVZoYDLxm21LWg/yoRUjT6PQjVIQ+6gNinEjaN582lg1PehNMoyKSFPlQrpx
Po8sdepiaYo4y9wV+mrNf9Cd0aGznWw8zXdJm4+EkZB96LcUevOryq6YqxLndRYB
lQhSTJnknkA5lTiFV3iVrTpVN2VY5ZNl8OJ9UeNsBohaE+IAmWbG3vJKuSpookMC
/f6fcBOg/Fqo5D04jngbQUz86uaKPRD9KoIODz7z1bqtL8h4KAumKANMaMYFvpsR
HgeK2SBGPtO/G7fZl02tc7Upom72n229lyGaI5ZYNxLewAGd9OW9/ou4WYdUEIKA
P+L53M2igq5k0aclodwO9JFBlyhLOn/CNoR7wNNmghQ+YDYJGNytIjlR6p3V1ame
w2hGIfbclup1t88yrOhFtgVlrncW8qseP6yV9nmpoJ4Kx3N7jJK6Wi0gcgDp94kr
JtgkXwJV/FKv5Qf+Tn4bM4w2LlIWkYrjfX3084Vq95c6CPPur1X+QguGvFzI92bn
NMiZVhIFTuYV4e+rmkN/EtX5OBTwyBJtUkwyGeLUkurOByd7vEWYXEhSE7dx1UVn
q73MOu5q+TYUkWaLpmO7Xhs0IIVPP9B9HsaJ9StmHMW4ydIoxVSDbAEd60mQH+Uz
BndjCFXjDdOOgWXquPdVG0eTiF9wKgJS5TR9Qo3gk2C+WcJhi3oCuABtXsLUCuSD
GpmBHf6dt8rXAhVjKktYnMSv0lbL2isFa0bVN7Y8jmD2gqdrNov7S9gSTBfQjnbI
k4f3YK3tcap4Dvy/egun3Vy+diJennWvz1vHXEqjd/IYpwOYRvghV6kh++Ki+suL
tGRkYlCnp4gZljftQ3rLmTzUwUGXm32xR9RTn25n+5VvuTn2USY059kWXWgfyGE7
HXDj2pHL4ttkcbk7RYsEc5M0WRl367uca6977/eB2kd47t1S2OpBnIzNUiv2BQHF
lTRfRcjQMJPyptKFlMl89n92zy+9XkLFN4n99naQ8uzhkmXecOA9BDp4jPuh33Zo
IDbEKi7NIhgTfMW/FYHGiC8j+xqySJQ0d5TrM202ufjlNJLeIe5ytrIjQe5fMAFx
9QIUu0uWW3uabCt2xvgB/yK1MBaaYqFfs66asyKp8kzkVLecS0R10Xv4dGWsVPP0
lyauSepF1FnmOpkXmrvb1xQrCZVy5GoqWb3MOBfWNW8QjinIlldzWxxeDgysSQz7
tQHWjlCrfXnVIVzpSEJoo76PS1VgIhYnQ+azvZ8oSlIRVf2ks81R0YJgBlYLYv15
rXu2X59sWPeBnLucVniBGfaZEIbrIWzNqRu8TZuGY9Jdk6rwK5fbF/ASVdJpYp+Q
zlOTEkgGjM9swybwMbm5fIym79o4M1P2sgionLERgwGs5kdfWCGAfH2FN+N7xw4f
vray5ZdSwAgkvkmEmFY3QnNNdN3zfa/bW1p1BWz7gVIWqRHUAGw78IfG41QJc367
QH/rsZ67ktDem/4gWrCFYkjkFm+zJFWTYaPsyqY2m81Iu0BNZItq3vw52bCdVCyK
95YnPcy9LUsbS2LKISY83duWTQzKc5TkJ96J+ZYqix4IcapArO5p3P/GmYlmLVj4
8km9OMhUSp6Ei7o0eNPtkRkuxArOSPCX0oFMsdM24rAmWNXSBuEt9bEW6YuEe0yi
od/X/0bJCrNY13gE/gUHhvSj3X8DURxDc6m7PtZQ1uPkmO23S55MbxJGmKMY9FZJ
nlI6/PF0J/x3++QXRAtaL/zwYF2ge4Hk+0Sy9YI0XG4H/HJNPTURyT8ya/GKgdkJ
mlcccltmPSl2/9MBGasPiiojr+jg2Z6Nseh7ItkKKvbVVpRz3bm4rCmozhS8ipWq
VDPmPpwLCM1IyjhFBn5aREoMGMlgxx2W8WZtfTzvdVYCFmnGK6WzYfX8VRnEio4b
61aZzZb7Fh0HV5Pzyktz0tAlnblYEYXufZq8euXMVm5KZxBjyhQ3bLRWvaIwakGm
EC/7LB1A9ceM5NgyCFpGZwfT22PhdubVT44QRmz67mRE/ienf4ZmFc/2YXD8Ftai
pdrhCjwYhxtk4nWqjiuX0gX2zhtE5KIBCvjnvXWEaR6i4w+6yoSlAvBM7hHdNXAr
WU9bGAdxw4LBCTZn10c5FToRQHIOtZY8k4qvRXeT6Iiji/A78ejOGX/QiHfOuvcY
lMSgOxI5wEEEDvGC2oONn89Bw1ZMsTXfaLGVVbVeFn+Z3RGbnSnmy+FeT2ZBXJIV
RSt9WQcnF7o+Vj3CBzda/Ux73zHseJebC/b8ddirSR2qVNLeyHVoi6+ZOeBXLd5N
TRSrzRpv/WYkANAtfrKeaMUT8O3Y6eVyxOhOW3dUgCmypKQ4ZLmrN40btZwJ3V31
KuWzktkUrwx6WaUuDelfzsije53+64ewa//x6WXxSE4lm2HrtRCTcRqZjv//Vnxj
UsPPWPAV2fL8hxEPc/kJdVoVFmQPc7r+t5X2nPhryRpHhqgn9SUuAJY65n+ZUGSe
gFfxzdAAWm2OdXB1AAE6Ivqze5sTl97N9ogMzLpVEuU1kDh/HR4POLaSKBVPqNRh
tDLely4DX4+Bt8uPLsVewWMHtIbcdaGZ5bvuZe/mGO8ukfbeJuwn2pcO56y1yCyA
YksQHi4I2hvCZR9XkAkvYKych37lNuYj6fEumSanPhHpOf+WLWasyoH5vuo0VKC/
rb2L39zK4avE9RP6S2A0+ZD5vu5GQkLhWubABkUJhkGlp/6nWd4kaLMWPHcxzqv8
Kc9W0Pa98imDZcQxda5Zs/LBNVO3ADRLbNkpMToRB+Qd4Bm4CPVMdPXthNanL4oL
9Auh3YUA3pDMDNZK2jcqAZxrfCf4Y6DsMr3Zyt/1YmN1NpatpYu2uIHL/Is3FqnA
oK6mJAjHf17vXa5DzC0tyt8f2U2ZkIqSLGYXQG5mrwHoVR6fDtFdVxuWtggW/Kly
W1hrb5kBmt2hmhKw5MbYBHDqdi6x7dMpcvuEyloZBRyd/Cqen4t1C5E1OI03ECOf
9rSUuy9C/LeQtqeCFODkTYD7iCe31xovq60EGV2+moo2BzCcKL4f4pN4nRPdiVqa
Io9YDD8jsrbwaGQAUJswKJiQbMqX/4DuCl/aglJuH8lwsBUeZFQCfh8ij3lc9YAK
3+sv2ILLtdjtPXyI/QRcdhL5x2BeZEOHE/0mB4UAJbSkjkVcG9Wg3HYOJUAgksjH
0kTuBDd32Jp67rcBbJ8iNb+v+yZAv8Ey52aOBXTzlFV/GzpxAmPn5zRjdbv2j8vU
HynRiT2eEdAZl/b10z9TLqTTmnvh1ENIiVm1ytoyRPgcfjO+NFgV7TwHIeNaGIUc
glGuHugG+6FMzTC0iBhN+WsmTwKbnY9UqBpvBcRKyM0fE3Uw3ohoN+34uoFBDMe3
le5WLwbjnof/3bZ6lONa7q6RSX4uErk6nHRX93OzFeK8j2inzgaDcRKemD4QxKen
hxMo0b7TLBglA9WF36am2myglE7nVtOGqlIylihYWRVHwPXFIU1cHCg0aufpLVOZ
ucrhG6dsqc1lhCV5XKYUnj0OPPJg3cW3/PLFNExDOoq3vTmlnn1V5NSem3QdkINx
Uj0Nq3SUd9+7Qx5xTEefY4NftJ9JbRtkj9WifbcTMIeCqa5xJByUpQlx8eOOOepz
1gLhWKM5zZeZohZ1967icJ1COajvT1aPlHK+EAE9AY4+Dub5esmjDZMM4rOMNIK1
sykIJSjHI05gDaWmN92fzZJue3kbx/9GnLW162CtuHE8VoK+g3Sx9MY3b0yHCnwk
JRXYEYe8/Srh+A8GMf7+MQKRD2raCMw3z7hxCpGO9/HE6oSyJQfDjm1EqFD/bAXG
+hZhZMx8HEIaDIMnzSCdDgWSeqBPTCom3/yBIxed9wMeaZBM+PdM5zpNLCvtvc96
cmMYhuaDB1+HbhsRMr4zgAsIlWG6gb8cAs2FnVb3/CY4LKfhhPu64f0O3iZonQJs
/vAGYHnu1ZQfUNPNS/MtlJdc5SIX/+/a/SoN7Vfyts6g3l+Uht3f9FHj6mqn8SGD
+rJWbzWx5WDkp7wqLvCnBeKdz70wg1+gv84MbLJlLiJdzqNibgR/dWQLzaG7Cd8J
n+XM6YIMfKnVNk7Pis9vh5cAasU5AEw566y3NVk6MwOasBN6KOfHqherhDZ+LDAv
XQbhKctIGUwetQOXthMruzmCogDLdidk9qTmV/rbBJgnONMtbmMKrBRIDlfLg+Bz
v5ZjB1A6WumsfDFo4nNxGzNx22NFx8FqtYUeeAGcxFLHeTu3hBRAZPXDvfwNatgG
bU+Pmum6YNVqXYA1qPwIARTWB1Cvp0By1TiOJGi6My+6TkjgwOTKPu0QmKnYVZ3i
FAPqxCWHfmZnBTCeU0BaYLDqjfBEXyhGXAsWACoRbY91v2cVx8hox8tCDcmIw8G+
UWa1A9bCw/U4wXXm7+Tuu5xpe94cdyuPjlC1hwa794jRFI0X6YCdkhdJQSd4Je90
j1U6/O529KxiuFYQSPjgU2x4FJ+7bEZLkp3ftYneIatuTdTjPbvlIGBZ7ikgRuhm
G2MIyQfhr8hoVJZiFaS0e6dAt4AUYqXUTOxOoqB2VuyxhXuH5XCeaTl6FbwpNHS+
TFsQKGzQcQyBmpMxOuDIyX7HWcwyvE8SpKJbzY4qUgkR6UgMP7dM9mwxVSFgMcPX
De+fUnOs4DHu8idHGelLlczqDU+/T9V63rTvkxxpuaofnnNqBzwAju0kdD+RfoFV
tfpzAbr73odGWU6Pz/8L0bqnIuI4FczCeQS8kJugqClleTBbfpkIbMHVOqf0wcLK
zPoX2ozJL6Z1DKzf9D5B7cEw4N1pVqRJGJsVVXTyr1dqWd29x+kTIHRpLMcAVoSS
4hhiZsypfWj+mtaVuI8yPMviKV/Kc8Qfd+BW8aJs85ALPxrYx1WhrNbdzXQoHt9Q
NK3G35TFIipO0xceCVfQBItiXQ/4w6cWMRr6lW0z0+9ofc/YcZR0I6zDMT8+7Jug
BBtaWn9Z6h7sTVDPL4p7s5/QpoPCjGRBQOSetqWl7p4+DS1aufr2X4Bio+IVnEBN
BZFLIUYY+rUDGQsl7lhk8gKm8aIoy91GHYemh2JTwhZkIhs6+GNWk1xDVkrAXjJ2
h0vng023xZQilAralClEWJU+p48OVGlskxmFxHY3N8bT10gII2lo22TLci4vJRds
0UhXv87oxQmDB/2GgrEldE/J92mX+QOxFNvuByZJ9LQbx50dDwHkD09Cvc3OmBw5
YhTX1e9rg3JT8rAfLSfaphOkuIxwWkhNvTkY1Elu9o2sw+fvNhJhuoUI1YVt4Ksw
5hlcNZrC/gOIg0uyVQi8Ulimr8+3d2MnfTPT7kAxGbLNRK12E0quLQySVUWTLV4R
vBP18/jtNKuRu+QX1meqI8pQNY1JpkEuDJcaQmU49hJ+aJ2nMkthBuijPfGTZazh
TkoCbqCVJYHgPeCQ5EH+TyW8K4qUdi3bRt+tta8HDMiKtoQEVv+7U2bIzgsQyank
zPXDzuPBluxvTAcMmzdpbxLcV9dXKqGwbrC/jaaEfvNuRSbkdTMEdhPp92fxMua/
WKXlb5+hsP1h5FzNnka04+MKgFXuY5aBEFYyhhd9RovTv3Zzo/AZZWupXohblG/X
YtCDDEm1y5SZAkdgMmjY1adatWn2iLuiVKIG/97wVrfTp3AJ3MtgxlEWeHzqhmuD
Oo+gKeGv5/Ler9+4byLTtXd7cC3m6JWIp8hhDpfk4SZ5mYFrIR3X9dsIfvNo+zFw
eEa+Zz7Rg1q4boOWTz1Lqrv9mvaJL77RfOgn8I5RGKJDymsV9iZMhGA8dAos6PO2
jrMD17ag8EdtBqgQ9Dks+0h3GF3ZZrXf3BdJ82yvf00CGEhfwcgkh43dCNUiTdYc
S/tYLrjhsq6qjdKEdxibWoZepRcseFUdNMulnBAj4qNmdySaG0Wt7fKrVrsZ7qkA
odmrAAetxGA+hwShS4tQEsjD/ugisb0tg0y0NJQh/hkYG/AxEPBB8WJp47SJ7oQ0
Ccmt5A51zu/i/lDunNMbe9JQ83aJs+J/aH7rk/powIZ7cnsgpSfu44GYjh1z1HPQ
umkE5+hhNNd3rz8SKd5LtlbG47MVbj7kBzzQRWQwSCEkm69Eb/TIi1TFQhx4htnq
kp4ZGOACqKIVsnXJMno0ygBICqUUxbPAWpdY9agVw1s4QV625LP7ZZbjRPjodPv4
dPaT3ZKxMMoz8iGHujcVWUxZJCYO/8EdjMzFJJbebTuoRwCkOHcyLgSG4lgTZ7jF
4+nrrOHFxMhO9uCeuQbsM8XqQxvl2RHPGGlAADxPJyCdEKXmQ9stbctyVJzjnVDr
T3rgt7PAZi/uxZQzBdBCNZOyCnO9XU/2wz+pzWgjDfkjKOZ3SxPwCCyFZWNJD1uh
gVmx5/SN58SUyaM5S+4GG8SHQvTcQto+JzGbOxlD4I3jL0u2yDxL8asP2nlEesje
gEtmb4rzI8pNmlZ4HacQnfNNeq22Y+T9CEnlAc91JhRgluO3FvlHi91Om9MSQ7O+
6AJTIa7Nw+epA0TK6DurE8KLcaZz4ZWLRmzwdP3XPdrwHaPCpLw3gNZb3Rh2Jun/
LQAndXIfx0nDoRohueRpMHyTx65z5rgxq6W3Ho9JRMe1UUpvdJqJ3iKVgCfQIR7k
c7Pf/RlMiLmUOgZvSPUstmkxLPNVkXDKUXsNpa7CLXnVVc1SIAXB1+Ot2GyuCtVD
OEKskh2rRplHitFGcW4ZbkiX22cNZaaJda34ozSUS6I+gASZBHE6TgWbTXkCHq1P
qsRmqLPHUzO489NHfD4DdsyY2UJI5kGVuXwAORMqewXS6/TirhvM7fAdg5XSAuAS
kk1q3XYi/Mijmh164StZKkgGLLvWwY4oG0FEJP8txligk1Xv6sLpZleoyIUNCvWc
c3OWn5fzHFeDqhlBkL9jTvbHIp30vZSCxxmfoIIxjJfnJ6q036q3cPVd+vJ8knNT
CgOSciIeowD4HH6PjASQ2kMHxsND96JeST8xKNg4wbdFhtrCAI9CH8n/cv0ReRKD
B4CrR0UsI3v24bgOZC4p0KCDzQjfKuShuglufE+8MwDhDwtWFcCBZqGyhP80ku2+
+a3WyszvGbUU7CtYHyuD5AbHqmn2o3trWcDRhnyYtAv/4oqdckCL30FUorOx5VHl
25GonDVv+Ysan5fXe9GGZqboatJGCXiFnftSEhoUI0FA/rMnGUdcra7vTEcIj93r
6B8lbvPhkHTb2TJ6AzvRz3sNICOIRGY+MSdo8aIH2wlk3qkMZhj4BoATN6I5aXL9
tTm8flrvG22K/heE+QDtlt+tmuoQNOXDD9rAhvltafg9nhafWvhOpaG5WGOl9U78
9M8n2Z6PF6W6zZFe8vkujx9ntvgVaZWQHv5umDXyWF2bp/CFcgT24UhfYN+TkDBt
vl0n/pC7gRfNllOm3EBteW+Jkh+sVPuNOKJDDVOHHk8ieNKAW+ASrbvshmtIPl+A
7KGbdJdupY0yo1bcW3L+FiYznahkfND/5YjcYIm1uqwxBuT8bbgD7NWjdY+95fZZ
3KTJWwXiWTRoqpMyc++I5HDwW3NGJvC8CFMsxfr/CrFj2aDFCiX9rrTWrhKhI0AB
Rk83v3yXulL9bU6Xd8lsO2W4EDLlJAKtZM4D4v/UiLzFS2I/D8dbWWiG+WkjD7N0
oT57Jr4ipJUaTXgd8yc30MI122A8lGexTEwiQQaA0D2Ct1+Ne9X028mlqVSjNRg/
G0UFWs2zj5KgCC53eiA77fOjZOaQAGFxU/WTwkuZxyC/ef9yBBCbV9uM9qOvxZqU
MF1YyKsgwgBHLBV928FRA0G28dSg0En3E1AA5EvZEHNZqf4OAY+/+LUVblbprW+c
/SBJOXe1Yq3XkkwKK2Vq6FOz1JJYFY6FHj/HYdv1Wj8Mx0IQJIqydNpl0iRvQvt9
nqI1zYeTegqbkcmCVhEmvtbe4XCkfmotOMfDcmVPPPF5JpOm/Sf4XZefr1kni53m
aTo/o+fNiNLRggBcXjXn3OuO0D35wY0koP2+W3asHuhdSDDdwodkOFerYPrzh/Ku
16YaAF2w3II2XoHWKsgHuvIMpsO7ULSVbTvG6NEXt3BNNQZdIlRRHSlUijM0isks
YNoLd4tIMbU0jgkJwjuy/IJ0fP3M3i/oQLGAH/q70FBxTiINe6dSXn4UbMz8js6a
F/m0xcZqkac1niNlph0tW34wdG6A+EhdUWb1xlDU56lkUM5WjLd2h6MG3QUwDbRz
IJPHiakca88pcg/pAbg2C/T0nCFINKiPx2H+JINSHMgj7S7MSXG1P4E8OlyaN8tl
uf/oU47/5o9ONqAV1QSLgNfPZ6payMP8O8I+DRYqlM0Qbk9h1GpU2ZguLTogAwZS
V/27tDFVtplMM/SKJctMfJn8+j5OBwanHBLO4a1Xw5E77AFKZwZlWlhVa6YgZmCw
Nuq6fNglVxxRr3g/JBm5xC/JE89bFb6yvuCBVDZYgF6fd+leCS7IcMP9eD20lzrB
SovFDAeb00ZSSH89oENrQDmRD4kb50iBseRilSHyfsrZAHhpx8rQTUgt0qYD+anj
ISreoguVkSLUtbxDcHQ44MelLxjqoig+1lnfBxTfrbl4Tf6ztLczC+WpSpFrqmoJ
0iEkfVW+5GebUEZwsWUAr1nfjZfbFuxJko4w1wFMAskTyiEpwn7oqfd1c9e4SjLZ
PGen99jRz6cfoj/0MH96PMIZuP8N8zOP5UlqOHHxq/+Q8cGjnKF/t87AORti/jyx
xSGjP7eHbf4pqrjf3Z8leDueoy90sDbldtZpnVdb7DaYuX34YXkJImkw5xnNWl4J
YWsJJAGlZrW+9kVdriJIkXa+ZNHhlohNoOwIGuWUeF8IJkxh+hdTOcyNR7rOuG6i
N0+S1dyF/wvjT5kD/kCMJOkbEpO5WCT9E66BhzNQqGfOLj6EAWolmYyuw2gqaHCw
d3ggIDLSDxDIsd6sLtZdFBxzzQpbX65JGpHEBYQVP31VvUvVTRStvbwQIsO0sALf
MXf5aEP/2A7sSsd+1q2qchvlfhEeHgbzYiyh7+J6s5ByyOSjPejmcoQHbSos8rUD
AW48LpvvsqREcWnNFKNq5Oi+zrA8yBO5mIBS9ej0ZliWt+mkd31BnyLe285iKSv2
An5QLnFAgwP6JtkZba912weHVW9sFfdXvLC3xkKxoouX0//BtldxHkJ2bVw0uOBF
Vq6ZNkFYmvVtJEKFAiASdJkoS0IkkwZHiQwGTD5sDDfvJiHF9mQfYu/Xz8cbAle+
JK6FJ8ZB/QGHMrTCZUkwMTD5iKHQcorg7Ukm/8zuNVmztrytG/xfhYpitcZlDlYE
w4uTTwQm8om2nSIZUw8HbM+RaTeVuRqQlF94Y7EMHAYlw1Zfe6x3P7G2GC64ABzG
GKs5WTpVkj76SRl2Ln4G+5EpbCTVxGX69QGVT19PFX/o8t5IHP62WTRw6fJJg1PW
HfUfBEV9m1qmcnedn4KchsE28JCAJ1d77W8S0oMTxuPKQcmzHEe8JPmNx7iYfW4z
jEiisBJafm36lpeB57FwyH6tJqYO89B+XTgz+jB+lczH8COMZWkbQb+WeG8YP4JN
QZyZEVc4zxJHXTxK+pEjCYupfNGRE+mKww8HwEB42pzV+9WYuqbxw4tr+n8i357W
Ojweq6BQzweQnSNCBtza9G6xL/kR+UG2x62fP4qWsCfp+O3o0vQFRKx2GGLCBOs9
jofaAmC9OtbXjK7GO/nyuJ58bF+C/LTmolpI7J6oUeqXa7yZhAItkV0Ga8UkUxrY
VFA6Gki6UVpk26eEX3UdMrASqIE4QPDnq8pSpOSGE31PsdJKvYoTp+wEYsGmLfPH
1a0BzA3lC2cVwRCPMcuKHCst2J7SYfhEJ2mux6PY+iCkVkH0w6nmqHOb4tiYQdYO
8GfK52sWqL5AmZ3cGFMGI3/430I9DBpYL/zQgCoJimcj/fBHcgQX7nita3BUrSNi
CWrvA4qoecS/GpzGer9W7rgtRqLMpOsAz8ky5Oo/uqYKSdydPvvn994HYFZleunu
FwlMsMs6n6EjKn2BNpQJaPBblonKcJ1FxfNGRMXtJVVtVzYXiH/ZPCFX7KKUPeqz
rNgKdn2OAErUZG4oSWCLiAia5auJJtGomyPpFxHMIgk+Qe+PijimolKnImSCkFv+
ZZSxdeNXa2tvJmnKcrxxJ1YaaaitVNh/khfFTwbj/G8M0o6Igde4ej2l50iBlVQ5
EB/Myb7aKFRiGDDqwWSP+oNXVHVs5rOUQfqLLy6OMHfyrT5XAlLyOfR9G0e1IFGW
eks+HorX+tUmvoU/k3Kleby9HMi+RwBAd2wwLiDpT8uCzUEcwrBjNCkEpgVDy0Ls
JPQTDJ9JStXsivoH7a6AU9UvwG1Y2thtSVMCZbB9YTn+WIQ9/IVM8+nu67ebAInS
D3ZcIFPLBbRceeJG/myX4tYLGKXSc7hPsRL38r82iQ3eVCaEqnHJeNw1CVtjQf62
lmWcvw6RmLDBvPVCJQ5TcTapj4NdK8u8bZHwDhdoFRhn/s2PC4lV2pmVy2DLzS2P
8QsfSEkeT/BhMQU+mWKopCkEAaD/bd8iTKEHVs7C9Ao+ibvepoXCNv/OfIe+3TAp
oS5QhKGRVZ2daMx59ox/0Rn1PC60k4E+1lxU+og1R0IKUrkG/Hlq3QZoZIkirmYT
qC18AQe0D70l+qiYfHtQocYMSS2vVarG98pGYav9LZj3duKKEUJL4fsSbOx2Xzsn
lNIXNs1WsJFfmbeMrazH5PTU6EnRIN2CXXCYTCH/HUKQ0VrB6rSzUh2nW3HrMwnO
24hV5ZxZxD4xHTOPCMTD5SoNOdofzEqccPqhd489oc5RX8wg89m8bMcgTak38Jjr
GYC3fuMcnO6z7tgw3xCPm0CmxfLjRDH712SSa2xbGfTKBPcvSB6T77Sw+OUEkTUM
Yzn0r76grbhG/ljryMOPfndMQYTCLm9G7lWo95P9ewIZF6KGaYoLIJCaYkt5/DWM
jI6H/8Vg+vUBkRTAh6xAIOWOr9PtXlYZw1q9Rz6qXv5N8fg6c2VS8q6yyJIf7+TZ
GytA05vOsxfxWGEzMfFmYzkOiVo1ORB3Ybk62IdZOqg+ai5DY2QKj2X6e9j5kchS
90O9ulT+/oMqDxWWaDmNfUAzZTXSncJfhueR57iKHFpmTKgYdsj776SBIXKK9ZXE
nAkI331PzJ4p5v3o1JcXFupyIitss6S4lK0bHS40cUrk4HH9uydgRw6glf6aWXcW
wC0EDO6Cdnvf0vqrulRmWX7lsXKsib+8Xahr9eMXYB91ojxAM8WGDIzG1yXv7HSp
2mJ6l3gIuPdFQ+j2InHf6GSGiFVbfkVFx1PYXNau6Bwm1zZjgXtHKWZ9kp2veTz7
0ENbkoPRjS+sa26KGdf23LbwzXRFuIDeJItbvJGhzOC9y5mikl+0o0LsC87k3JJF
Y7GCpkS/Kkx7LmNCUzraJqWEeOPbhvYOkoct4fP5uCYNcuJn2r4vjpoBxHscmXmV
hs0EagmKcW8lzQyzmYMo1+JuCYEXv0pZEA4gbZ4FYdVU/9snVSozbDS+SpoYx0OK
LgyfqZlr1a0ve5YvR7/VtrPmWxYKWLGKlPCCGoMbV640pBw64Nbz0Rf4gTlT4/L6
xNzxA0mK7+PyacVH5uAjuPfxb5t0CsH4tqCTUcN//qXvu28gZyFK9bKjV/USYpcD
9JH9Wl/mLvDGHmI4F+5jKvZlim0oLpmLxfLPgidYLhISPlKdnbU6F1fopsTDc6Ud
56XiCLyO4mWCTtYotRvaqcyKJ7piQMoMDnzTTm69Fwh/HW+BxS+3UBmht4d0fx75
dEzGk3h8HiT66iiQGBR358q9xKIeO+UUEiL9zqGbEAj4fXMdD7/U6lilfBlSljrc
SRW8QTwU4IqIRwZzG1oOZ9v9Ke5f/cVcgtHNEUQJ9iyci9GB7oQj4AW1C/cuZ7OX
zFru2qSvYMgCaFN6JycJa2EW0KySjYWabQUJOvd1EkeZw+gkC2JQv8gdSQ/Z1ZV6
sR7y4t4DCncDDXSbE85VOs/ptPxDvMkXUwtpMaPJZxcmxngcuJSubIz1aQXThEqa
2apMi2ced/5qj94eu/8AZAhsLQO8iR5PUHXvO6n0idISE4g0rn849l1X37E2kol9
clYG1mcLDUXiNQvQCbTxYP2DsYuMUEujSFypOSQXvSxxD6hzvmZ8don8EczEPoFh
cqqp+hb5+a4QSwvC1IhvafteeTX3zqJPuoLXtGWAq462MtyX9QRNF3v2NFYJ4vVK
QpA0tZ5u4cXbF94kTc33VqammgXm5Rt5Arr5rJg5+NiQN6XzFaEZ/rLE+Qhw++U7
ntxqWd+zeG1qKhs1O65tRUNnPSWVqDEYf8oS1Picd3VypD/doL66IndMltl1yVJ0
DtDIyl46YvmRE/9MsxmTa5JgkNxg8YorhmK9Xqt2P9nCLEwMtSCpKM9GD3XQpwp4
fOQ3lZi24Kejza7zrF5TCT7T4tJFFXqhe1n0SXMH2sBTwBZwv2+Qn5eisa8WLEuh
PdMQKHfUDGcg5J1RQOVeyV/GUnZx612E75WB83uAlWpZTksYtpitNmDOU0WGD3mp
LTf08zIzrAVEuvLzcT/C/4GyzKJsN81vQe5TU0gAi4VurqATnRm+bir6CDAlRc1A
oCAuaZr3NuKwFJJttCWVtY3CSWsj4Zxfcgql201yscL7y8Q7fCXWCoViw1aqe1kH
X8uo4S95gS/mKmE5EuBvGg+Mgi1LCJzB0g6IoKqYAfUDnze3jhHbuWPizBdDXkYi
5InjSYxOtDTY/69AUkxJsV7g0ht/eo1/4c+7g8B5JvkPrC4uoW7SwgqF9r4YMBtC
S0A+XVO+u06k6cua4I0Hm2XEkrwYX0RyUlPWk1jistTGMFGU6DKES8cuH6jp2Lcl
fLQiR5v7YB5lx3l+BOWo9v7i/7RZlYI08tArs0MxZRqhUqQ818/tk2uJVZdJGD6c
tDWWuMFzY1xd/0rp/HlISqXtcEk0V8EABnh+GCzT93ZVILTora1a9pplUyfYaSPG
+Dj+jiEVMs/DHjfRH+DrndyTxU6h9VWs6l46eIVTwvgdddI11aNA9J6OoS6t2Q8Z
3v/70msys5ilMtxSqo8zajB0vj24ArquYZJ0MS/F4b0thNYceBYgSIGUTZbYEQS7
1AgxxV1CaEHrgYcIKU+aZtbSpYK95B0NdTsyT2P/MHE/n+h33I3sn/Cf1MD5imab
J16UATK74YA1ctucOQjUhSHrx5v6O5siY+ic3QGMi4BEL0ZokeSuGxZnVTU6FEou
4uGumlkpTLyZBz/8ZErtkkpLfhkhF5gOSl4kETYyAPdEcaLdkzGK7fBjzE5YdQ+g
Ee/U5qzev/5mcJ1rJxJI6RvBgPtUJwzdYG1SrFvw6fyI57t/c8UvqA3PsQZUHAl8
3si4qNNI6jIHtPGqwUOylIqKGa9slfagNSwRyz6XZHSjKuzpAsAROpo4NNwKOZrZ
vA0yp9D2uoVP8h4F3tmeaAPvprq45VU9+v/VgxNUqao5SJ/G7f19xbjugVsi/npW
q7xLYRJV6m+WE+dlL0HUYAmZeaYaG6Dx3E0TXSeNjs9T7TFJy3aa0wF56X558NEE
QDya0nV+HKA9NkAtm5V3WgmgDKt+rKZLl7zYt3Gvbu0LzL2E6XArsLfFhIdiMEJl
zcWFGBIKEeyByio2+Hs3Br++iKlVbrlIjrCs2fy69EiAQoi0mpHdCA/oHqlD0DNR
TiCj4NRiuqlfAEUREV/MIpsiBBgaUOH0pikuZ+F13Iyl3xalpZdIdffxN0qv01gr
8qmUu1RgQAZGzeZFRMKOqXH1HyXSKgW8m2D6Yj01WTp0N3d0YCSZMAf5FccgXlBu
esWT2nhgQwGvQzRGnWZSf/TllpzWG+dcPmp3IuwakGds5HejmuIf5sEo6XnWFaZw
RZaE2+C+3uvDkEZR5XiUbwTB9gLHf0bF9gCCYifWqPUZQdiCpvqvmewE9/sgk8Qc
zt2R7o0Fw63od+0/AFrIvSCOHuewTPkLVc413ldU4eTFJN/xeS4yeKFxjnH0VxIv
n+ygjQm57IhVtf17lgnhNtzbC34sS1ZKa0j5uZULe8EBgGAs3PnMPlG/zVsk+LUi
LhJzYuqzb8GcS2ksIjnIqUiv7a4CjUlDfVe8TkYCovZNLqNdOnBGQgRRtq07ppWc
3zUfwIEDeoyjZsbH2U+uPdMzc+T0XzU6qabXe2KN/kEMB5llRvtx6H9WDrpNRj48
wexjLGmlXVR0Asf/LVZvMpappUksCpHikw2xE2TDi/qY78oJDbrtzhbsUTi/WM9J
rnQyB5zdGDGSgYVyjjPDeVIZOXXYBCrUqztlA2y0YUoKX5XzztHdFzuRyqwULX/0
jpUmzm5mth60ZgOj7cl8MH31+3iF5db/d+NoGwXsK+MkgvUklsvA1qhAZvb5N8Og
luIhQTytkMn+Sum+4s5eoMqKztMmw9fp3kRd9gIXZHz6kgPlng7qW3EEqdikty5x
Qu7pIq//r8fJToPJLjZuRUPA3L4CwUHDDG0oCqrRP+sFFPOF4MrAD2Awnl+UG0zw
XKEmoJiVrlIUvy6br5Mg9QCrJWSOmDrXVodWDRhNwYEMctv95LQlAsLiVQyQrE+m
febZLqJ9FAOJI+fzP/mqItqIUO7qwWGG1hu4ZcT8GceAS1ZpCKTwjT/rwVPBSMWc
m+r0pTZeJrlsQk02AAijFwXvhmd2OQRW3ivWOZTR9pwXH/X1vLVc9FGP2LV0q7/o
4dxHIf6u6m7+oGiNfqdz8U6K9vOyfXEMQBRk62ymnSo3jbXiRpty+6bfVMXJOdrF
nvcibAINFUFtWcAIJllNGdCp8rtkbxzEfng7y5GChbCc1hmRCufiUy7YuXyW+wLb
wz7nMWr46qTjNk8OwB9MK45w1ErLVdbUBHZZe9g+8MWBadKUO9yh+XhPJ2QqoYpK
bMjhXSuGItpL7Dig6jitDHMOcDw76r4P2uqG8aFgJhA8QWwB95wIRFR8j1ucsEPo
oYBxavKxhVHOafvqopnCHkN1OnwwwnePBuLxWyqdgABILRdE4FGkAk7HMJf6uFEL
eCVGaCn2y501jx6951Ne6yyiqoqt1fD77/L2fNpZGWmDkXAZ3odY+amOAFEE+NkT
0CtqVGKXZCarmo+z0/wBLmdqyPy6kD2VBpgO5R/gyaQgNIJGf8/cS5UKis92WGYu
sHR/wEyQuVqFaFFDWxgC7yZH/bo0nx8R4NKlCHFJtNTL5BKg5fmqVh77RZakFQSa
i9+r4eh+XggC9Qtvq7DzJeYFLd1Pz0yoKfwOwj05RbiZJIxYdQ9IcsYgMY8elgGE
sum3H8445gK65/uepDK5EqPwQWysh6hdDSC2mED2CnXMzuirLxvbda0QJeAO63XC
doucal8wJLDvJHpI0qMgmCsCMe72lTJ6GVIPdqRvz4Yma8UhoBuzrd47dVx5BzUi
9hfe/nl+/hJZWG5sfryXTP/9JUIjY2tXfDvIydmczQboHOhHAWbhd4GT1pDEQ3GG
U7QuRA7CjZyL629jW8NGHebrVJrzfsBn/T1WeTYUDg20voCd7pEEue7zYONLHxml
L3zD6g5P3Qphvgw3iFxviec0vK+YAHetNCXmQApQLgocAhvAzbHyDhxvN4NojvAB
dKTsAQ9VCEV2YvQDsF+v+IcovN94y5sv5nZfj0dw4s0PTnE2rGvXWzq/tLCfULta
BlV/El62DJGMXeX86u7a2PE9SAwQgclvaRgV+aKTaFxNqntwSRDfidq+qpwV1zDi
skeEsdNZEkIwF1cMzvPkYHTL7uEtZ6dAWTNwaZ8FHd1KTVUnTV0ZYj/abZjohp+e
bNfx6VgHsXb9gSUhK/No64/HfCyn4bXJBqI8lVoUiIQheGj7/pzltmn9GZE56U3t
U18UmG9NiDZnIiUGsYScHgRZMFV4SXIe99BBrKhPj3dXnTHhiUAF0+SlIn10Fi3U
VehqCab1KhRIDIPeUSWkObKKvkNGoDKU+AGKvaY3Fb/N4m+h/wkWE9ajtaFX9Wmv
HstiC487tsjurQKea7PJgbExGai4g+Q58B0NGFtaPN9+3f1j8x8rKcCa/L/fG8Lf
V6GJTQGe/8RJZMAbdihGhgSxdYbyRop47XKx2PKoTByATmNzG3m8jylyoMEcSNSQ
CR3UIZZnP6DGLbmLaUpqCEElF78WqyH50WJLFiPu6fiM3ZbEC6nFygNGNj4hL5UT
Z1Z457fkaP6XX9s54i29Y8/AngQ96yuOK61L19yEA0dESrToCoJDAoUUmDcl3V32
eHLUPSI2v8YoW7oRo4Kgl09R1KhT/Rh7aaOF39XYPMMTP58KTe6hIvXje702sOwA
3YZu5Vk3sLolyFFmYCO72CCOQK800Ly7xneqcse+gQM4DdnjHtQf91cwLzydJLKO
WYIrkE40D2D0hNGbwyyC0tGx5RyuA5yWx00KxHu+Lw3B5+zF2lcA8GRWRrdulFvs
orZGSXqiMHiwdvg3FBECMdvy/h0Z2rq+vw/Bjbx24mDUDv4ZkNH/+bgswke29P+h
PUoNfpRZWlMKOHIwlTYtLTBfwAocYFnOlTMk8NSjTijhsZdC2EU+FGCuRiFTru4x
P0t+jqPjChXvhEvD+7bEZhyr/bWM2dvLLHn28gCocMkuWZ9AAbGZtgasWsQRTinZ
WmVfMDAcY9MEWPoottwr0VJNViWEPsvcS+f7mGWj3kn/MjkI9/8+EtMAefUnFeb7
8WrfpXCleJjAb9JsospF+XDCkCCVVV1pCJtl78FHHE/LYYkIzIojOMYpsUxo4tfr
8ywbc1rYsWtPmw/Jy3HfoVNgVZAMrV+GZs4ybgGYQzuL4sy8np6jGxegk8od78f3
QXfpwddUNeGEEG+xw/p7PMF0HzhyQATDBq4hNo6D1QIqcZJVVEOr55Du9lJ2V4Wz
`pragma protect end_protected
