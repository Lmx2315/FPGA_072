// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:37:05 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
TIQr6Ne61IS7/wn7EjtxQclF3OAUFcE4ifwC+DNnDevTA+FkmgGRgazkMuSb0nLC
8oWeGz/HqpyLVB+s6BNs/Lqo01xws201rfb6WwhSD7UuwyHn8+ceUnUkHMlVcd4t
GiX+PeWjNpcUrrumFHDNhUwRcobX/cxTkVityuMOuxs=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 21296)
wdlLYjjPHrpBtvDqvvYBp7m/CFeF+BGIKujxxOXQgDs9JOiWmfs7zAdaSqaD0Zwb
1Cy5i+yDdhQITHWeKPOvsc+cVD3V5/dvqTo3+cojK7zfX1pBWnrrz1MScNE4nuvD
vsoY5DNQW1QGl68yLKLJraBeCCEOXLo0efvGJxNW39cjVOadHtjSSCGEtL96X1oR
KCDu+tEkTMPg35K3J8NA4JpEwXiJqtNmTQ0RS8MMs88K0NwVgYR8avHX56H4Dogn
YZJe334z+Lra20Ggv25bWDSZnqWrkAn4aDddwv/4p+daq7JNgLZXVdGGSHYzbs79
MOOozg4SNv26ioeyPLRwsjOOkXi9nKxZ4JP3cwaib2M+tsINcv951dR38F4hthcm
jurFQfFi9TpwDIlNOxI5/IRRlJNG+gSXG4+XjWIrbrg++dBCkroMINLwou5owrXS
s3wBTrJsiXYfHqqWOmGBS3gpBY8vjGjqcpceDVjD6au5WO35MuhyuiWGfHN5vaBJ
DTVmMr2S2TjJv8gPGpA1faO58EQFXdzQKUFFopxD7Dq5DxaLZZmnCWM90e0MTDpe
Fs+dsgy8ZwCfGfpWhEunCAV74IeATCGyJqlDDfqcMOHeAgx2I70xzkzlTb9YmRHE
RLY6v/JGqTZr1R631S5ciC8KPxk7fajmKpty7nABM7L4aBHV+J1dFCBni9asIBrN
/MdIi3ciXYm/1EXPAkcMG+Q4VN93X3IXHZ6e6iXqaFkmBdbsmhQKGGPgtbBnHUTs
Gso9jQExpM0O1LpbUB1sgYqE+oY5akNeuaM+PfcA/VG3SFYXdeYupxbHvaYrbPnT
TCtR36skT62kqFIuDvG5tQw2TyeDSphJmKjBMq5GngGbEnRb45zf6vAAl8vgOnoK
Bq2LqrU211dzHnlKvT5WZVzixyRKrbtsUEzjEsXlDysJ6/uumH79PVLyhxekbe+B
V9UiNgtU8WypRt0tv+LuJJr0HYG9nahQqR0hRjN/UngPCw9eE+4vFKmoXXa758eh
EAndjYBbowJAjByw3vMYvDgFHOoG6axIn2OLNK7BF46Ug2t3YgFoI+Htz+dT3R/l
yTn3rsmLyn6l7xtUwm4rmvJQhmlHxAUyOPR8U27I2/D3zgfNr7S46vBlhtc4eajd
cR+hq71nJhF77sQuGmkppknDXf4ZWJpGPGRTGl+PWM2dQjkdt1TW+y1k/O0hRN1G
cjKItivavaWSDVgka5eGCYuW9dkAvXVd9qazoZsmGUCBAx1nHNbmD3uuuD4B0R1o
jclKFMfMkMYFTFRSkrYx6dcOMqltkdhMLNN/WoLyrGCEnB5ZLlWaSKD4RHFqh0uy
C+aWmGTG4hkoh2zoCaut0El8VIUdH2VV2F2Nc1IwXYK5PXIrETJMDwrVTpUI5YSR
B5UZNu4QBctTsLY+i0CWWGpRluz/aTUV2DnCjq+W1CkptN/ugGc00fUClJFF9Voq
Mgm60Qu3wbmaR74CL9QUMw/ZZXgKo0Qjax+GUzT26DXHHKajKrbotunCGmqdzns8
bQDh1u3U1QSrbmC2m3BBMnmm5a9C2dVrUOsNdplsGq8yqVxhJVUi9O0yCZ3VeItd
p8JL3zU5c4dKhiuXQMKJeC0NJPheBQwpvXXfWSkYVhY9AcF22u+/xzZuwVNDvJtc
apKYDCi16RKEk4cye2s4cRB+iHYEjhGH/WQgNLGXZ+efkyXd8Rg3qnBYqm5rPEQL
y57wK9tMc8NHmhpH33K2YxaiMaYTihGC1OcSDoNAJ32gQI3jmj4EJmCaiWdd8PgP
QvndSCaTCwzKb+1v9txnkl4KfLAu/wm3JE9F79HAHQbkaA7TL7EjO4RkLN/hkd97
R0k1BIS3DGp/c0xEgp1pUvF/OJ4SNt6KqcbYUpwhOS8tb+VSbAMLw9GbGms5EIhj
ZJtqQ5ClZvMucSuPJGfCbttGg+RL5GytAN9oiiqRckRnr2swsNWzvgNsta4rj2Wl
zOyH4Z+CiQxguvssjlYSuCQ1WV8PMn/KCkIx9ovKLvaXx+XpNUJFAOICeXPWKPKn
giQCLBvjxMOFNNHL/Wz7Y435HmdR3eXZd8bRBHGpCh9Rc8neuJpCxyAmfYqDpbmU
SP+ZtbmTRyHJtPJoxC2j6Ofbg/UWMmvWfhLmPyONm4MomcGAj/mT9C2b0zyMxhNJ
6DQ6T3GZO+6yso001xSfgfNSKuMV4dHH2u1LU9UuJdSCtStxMcFzFLHoLe2kkYqM
OmDt+DUGi0X0k6/QyRq73G1bSnFjxxClpxjz+w0FwzffKdlzd/RcgHpdT8Ojjf1W
ZAD4hHwLVAAuYENBHM3Z4ov/L6+mLyTdyw8LWwM8xFOB8tBUDrB9NaIVvxNQxeA1
gzlkp6gWc3SAZUd/NMjYaXjpfNnbtBgl7w4OVWSwGKL9t9TGWjxOwLQtxAsAZBrr
T4ABJI47ErQbRDqWebwkoi+QYQ0JSzPxr+sSDjWV+8AICbugY5wz+JU5zepFiBRi
JWaLGKMQeSnzm1xFYhhQrBWfjE1chUcF/UBtOC5pszWUrHFOwSNwLgfUxoJVZ4Oe
+GcBIgCOQGu2ZmQTq2FfyZWUpSwCL1X/V0W1nHXNNSygbayqzeqXjsYGzKXl4JfL
q/6eFuZdRvLNnPsx8KSgHFvvtsGRi3NlhpQGTfYfuz13E5jdMAix00wQ89uAuFzw
padatzzNYoaG/O7Jwk25diR3AsdertZYd018/EUr6S/9VzvKyCIKmAglIvT/WwcG
jmVl8r0T7X1Az02pA/m+oyt4DwYNio3hQUchk0+ZC75bVxAArFKHpCDOoLbd2pQ0
vnz2yFy6gcP67GVfcoaX/ZelaB55yi0WzAmOCc8tLUHzdDs5mZ4aub5A0TN8Dfw4
axIDJB15Ks0elASMGUW1fXH6vUbA4UWMXz6pyuXt2y4KS7QNLkhLaoAxlix3plUS
GrqJJ6GG2EZ8WDjvWPjyvt+eKtAdhrT8/VVp1e9owdyImPqI+JxERW6ctiPLI1tg
i0x2PzPaDDgotIdXRjkqOAf1sB8z0rIary3iNPyOHXGuqWGXSCs2k5HT2JrFw9ZQ
PyKICpx8zUXNLKnjpnhnDJk5jcQqOxh74yKwI5aGuivqc5BLwsiCQHeEF3DpCNu0
LKtCNKwOS+Brft0LPE5gdOeosYWTd9KhuO2fUeJNYKzd9V8cIUZ2Td9rYxMemIXn
CchwadxCn/6dKo+P71tJ6hkaT6Geb4/2Vif2qqqygnPNGCvNqgBVhOCx/bEsfxIN
F9PgFXow6pd6VdPAgqwHld2D8jzbyXDaPO49rsaoXweVWaVMzye53fAbXvifBlL2
nO7vscc583EDL7+qpGGCfptaqiPMRBgReTfigmbrUU5Qzl6MhC4DQocFaC0mUDzi
8icjfTvIUTP96FENfGrUYGqiEaXpxUM8aso1Vf6gkZAxgpzkHluyTy0zuomi7wQS
JVQ4saY3FMWjiF6SFk4Z4mXQtTr6bZoylm//uB6TvXJ/QeMh1bqlUsp2iJbukZXM
zmX4VzLwAM7wkJO0lJ98DSADqBGmiu6rlFCCT/qZx74jfYzA/GWCGfobuikRg8BR
LiMx2WqaVZ34qSF8Gu7qK928+5xuAqN6XYwtlKHNgWjt3FkOyoPRjXJ78xM/giaV
xnft6HBjQmc47h43xi15NOOVHbgzVVuVBgATK+2hVT0q4IzdLFXyjI1EUHrx2p+X
PXEVpJTE124pr+Dr19PbaHi/zjQPg4UQ+LKSxxK+hNMjGPI6TpBkH6pxHxx0pGAe
iWjZa4pEko88XtDXZURGti0D8sI62hKMYpdL3ieIBz5R0dETBAadXbFow9Hv5au7
KqeyPoqMBnJxPbrrszCMm3s/jY2N4U0wMnbIvytccq5zZIdTSE4BRscBFemzkkE/
V+oK/MneKJBZFybbDrnVPj5UA+o4eYyjNlDC84F7JcGxe7ZjmVTl9Dli7SFcQdgp
fNl3kxthmTds8DUXc3irFS8D3Q16tOgB78nswKszf6jIJ1tVKVSZGhlL3/1EmQWW
BKiCFReMXyn1pEq9W1LlBLjB4PY5DobUH3De2G3fnCZO4c9w+ZWp+VqdrIHkuURI
SMgvj2GaH1hB+Wx0+S2/5WDgyz7Imc5PKdslwbcjd/Bt45RKaoBw30gBP6YwXJp4
ZcZZHgE5sVPTDyWxp8iAXZZpNiIYOyCDEdiB4fJ8le8JN1k2D47Wt1rgRFnQk10p
W91cF71IDIRXeMXHxAG+NWYBumdVP4RBiT6dzOIi+62UBK12rxpU1E9c9Wsyg4YM
vtZBZ+9SsA8mZiLKcc2z3z1nWE6oDaRihmxVhUnM4tGpL1CeeKhFSiBpV8NbSdTE
U+qW1KlunLssaTZKBVkFq8rT44S0svGF8vWR2II5SNoxMneSBfVYohMnOlWabvHY
iJ6hc2lA09LTBBQWJkar9VN/hm9hpeTEUuuKlFC4Y1SM/uKVd5k8vfWpDDqg0WXO
epFuAxI3YNE7PUP+GMTEWts754Hc6IlqiImGkhLuXpaEpOg13sRKirmFd0L8jfGC
oyCKh1LfEMlVYfwYQqaJ9CE2w23sSxAYkD8r0NqyXa423ZQ52RnBNV2vbyaCPcUr
Yd92wa10hxaMEk5tXyZ6GPyTutIhjE/5t/tpqxjU2x4ShqHD+A+iStns9E+WJcrr
RU9kyQjq/Ro8waeF6e28HfDwLceW/HKzDNDYYLNU36HPIfljGVNVqOxGutmrCe/6
sxzUW1rdPmI5xfzvTYlvrepC2MGil5QaWbo5m3zlZI3XuRoUkStRNOBlU1Qy/n3w
ydeWqTK9UjogWRhBY5F9au0Y41EyKFsU/0cprW5PLFDDchGytwe73O+2p2GEptVg
ZFuRRIFRkZaelYs0jKrpBAEn0vya70VElewZN7KEu1WkBhNp41vf03sV1aToeorJ
VTHGscDJKQo9GJ32h4/DYZLYE2X7NxH7ajfhguIhV7X1i+L1i5BHJwW0PpEeeTor
AzPH+5RQtdvNET2FuVC/x/bNyEV8hk6Okwmx9JhzUAxbfBDPTp+paQ9EUEEtcrQS
nv+nHLumNy/Yp7oxHVHeYn6eUFg596UXUYzTB78amAUFKs1SVICsqdYbiP5Xc3SU
FE9bQplrsKRukd9hwTsy6SDPYbDgNa3nhFFEh1rBuqChguKOhq844Z6lgdpPkz5v
gRnDzt8Z5bIzLG31TpJ/HYVwsCKVdwqyFMchTChjbEsMkqiyXff8s1J/kok8QttW
8srmgTTZE9hG4/DFHBVoj7oL5bflqNYv1LDiqy5hsjhIvk5gERqf7N1kXiInNcY5
ixaNxexDia+c/Af8Hvb08E1I/YvfUNZN+WO5hoiOzRTylhj0dwQxboMgJbINaE8L
vtr3EdBBxFOlbY5RaeTDlQw2XCqnGTkd3bEfKCgUVh/+xbi8oqSt3qW0ftVVoxqQ
tngdRDkzKmXyCFg9O3GbPybLvUCV6xcwom0ci8kDpk3cU0ePE0VM5oSWBQr4J5pS
HtUSQAqflOovQah4VBklqLH5AMcBI8utFikdc6v11R5F/xs4PqLpF7RLsTxHdIBs
NfGzv57MMAUUJDTk1BN43Wdx4lUved8TsKrYN9AZk84GYeKfZDEUGJUOLQMOT7VS
DnjciA5slaiaMfzEjVf/Qnfsn03M6Im4q4AlS2qwElKeHydhoLz5qEuZArBW3WiN
Rdvwe0VOQ41K5BTa4T5vqqiALE0OkIXclV+1pRu/WjiVCd75pKo3PbwQCUS1fyqT
X1uyJ51J6Cr2/yQI79wqLDpQFZXTYWd7J72YdV3j2gHTs88/HA8hA543b9sPoJFo
ooWfpqaCrvpySnETQKB3f4pdB5stjTpZzOxHvzheFBNycOMKg8tIfFj1cpD8kz+P
pz+aRXWEF2I3JUd7DfuAdzML+PkLVEA+maw8fEYVjFZK7D52Y02V61D+bJvi9kDM
lPNx5pfk1XCp6QXKzaZ7hZk/TVFC6NP5qsSgpSc5TPOpef5Bi4q21xPpUvNlaLWA
jYe+phYCw5cCKYZI5UXaFuTNSE5pbYwb+MrIN/vsnj1UYKrOI3ZQPy4enf3W6eMn
LI4CMH32wwodKKjQq9uUCvykuiu+vgZPg4/3+8wAi7ZYpI7pjO4N0iCK6rWjYUnk
zpCh0DL1kGfC2VYiplxqrCHUoUYNu2llSZh629QoRCkt2cvNT3cjHrJ40cqiMVgy
2nIrV2nkijTmuYldAiuLJIjJQkY961PqY1kPGMuJTANjdnfPh+ZYBvKNfEAOjh4v
Hy1KvLZh3UGSKl0ShYrDnVmNnLEaZUPNXAY3/z54fqA0leWHyglz6fXszHjlm2x4
7PSYLy96bIO0BzWVMnQZqluFp3GrCyA8fktaylAYiRKcy+0jFfd4hzHpH+5TvQxm
bA8JZ1RWr4wi0Waj9VdVbD1Eka4eeaKz+S5tK4nW/pEr8Lb/3xsqF/S0glB5LkHc
Z74h9KMr5fFryvk5WOxj62o+OVAMK4Crp9uKk2OCBLkoNOrp6ylwdBh64IZyzk1x
Quor4B6Cp1eCbDMM8ulf4Wk+vYK1HRFzAc3qyiobI4CqqFthEpBrWU08uY8bynIu
gTO6HYxMRYFSe2ilNBP6j0KSp8MpmtkXziwG00lgiZkphQo5NnI4FTbvgC937uOH
m5THADS//37ISmxA3Hj2R9LtNxU8AMhhBdlB9VoBsdhbbJKx4/GCwpQW6iOdAY8u
MClHnlPMK2g1Gp5lGc1L9CWXO87btnKR2PKgNgQJJyNWd/BoFe/lgPVH7oYnjTN+
Wfzohqa0eBQtTPwWfsTvrCQw6Kc1D0bnDs4e93jWrbDh2KHQqcaeQkPFHgOQTO29
J+vwh8DBxFP9SFl8RADLHhSLhf3JLYg3NmocL3ehGA3KKFecO/6yf8Im1HVsiim3
GrxAoLIZLOSXNe35OXjlh93zB4Vw6n3XLa4P9YAwjGDvnksBU8AmCmU13Osczs3n
QuZyj4zs+WBHKdgxQ2cjnBvxqyTlq/eKl0ewC/3PmHmmme5gCu9wJsby0OHdSJyD
owcDfLG9FCPT68unzXy7jsV2iL6X/KgPiSWx7ICPM2PjsCmfeCNv8QlbwNrbPtlq
6d5visnYSxFAK8oAFR/3tSK9gRvZLpmZDCz0VIVFCnroNTeP9D+FEyspt0KYHMom
1DMMA6cNuzxUuxUa2eoB/Wj3YOZ2ZbxKjB2zikB/Q7rDoELwQZFjjr8oVQxCsKt/
2XW95FSNkx3a3+JIpSXfjJehJu0mZaOf5MS2O3KeUevK7T9RX+NkoAlH16JlQpNb
aP7l8nKdyDiEF0UANP9zMHfFd/D6OUQc4JLztb3p+CtWKMTOFQE1khZmboTHvJON
kL9NB1Ek4aU0dpxhMPfo4xvHvLfs8bKm8foJWWLx63uKJ1oqogTz7UpsA8vWIv1s
Tka2PasyCCpw/Egbo2CN5zNY4CRvScCJnsh24OsCHHxQTnOZPQoPpc9Q7iBCSHfu
pTBKYiyd21jKlVQM5vKYIiscuVdAjw2TQ2GOeVsXxsUcxNYGHjApZc3JomBvelz0
+WS1KvF20RXQ6bs3KakfH59HIWs8z7Im/Z8Hgh8J/l2GAHgtH6M0tgYt22gR+9sL
ASptNfPCqOlSleA3Esiw2nAObPD+/KXSdotoUaAOB5AHHWa1Atw2D/jTUa0jznha
x3R8vtU8OiLEnaiiAsk2PzP/N+N2x9EOalFnIcBKZ8JE4NdlrRlXUdeizUM3yZwY
Hkk910NXGu7s3L+8hBodatnjiwfRizeYFMgpNCvUXpbSMx83EkPswjX3ncLS0I2s
v0I9fy45+zUqnvFjrIE8+97nKKuWCLoeDxr6WE0XFDW4CJ3TGI2K9UuGbf2TlOxY
6/jIC6+5RX2wxGRKocmuPrYo0k1yg192WibU5r9Q+L72fM758oAv9w3BsrmU53eM
qHw15apc1eFcmzjGiwk+QS0AtU8PEX4LDzMo10VsWhAgt1IarFUWv8dXX0p23724
jcieq7C0zfrGj6qJh6ziLFbCM1CSU0iDLHgz4p95ZSWxClWSXFThekLEWNLQUgPQ
JLtZwFz6R5eg0M1TS5tEgAnZaaA/INleW0yVAlOPlKZtPKZTyXKFFkvdCk9fdoC8
ZySdGPj4x9rqkaNi1wwI07xHy62G2+C/nuy8E7W7VEVp1mmQRAjpgJndWrDV2OLb
Aat13QcbGf8c0Omh4EXXZmFUFuHr4CHrzE9Ny0FlOsf9WwhdcuCU2JastXKgkrIb
hwytkAKYNVUWfOWE9Yn7wfF+xWQyMsvBIGtHpIUec86dkFV9MdAqBp1OwEU+b1iR
5EHI44WBdJF99gSYLR6dsm76uSa68JGp086eicNBWupZteA+yi2Kq1hLqcJGEug3
+pR1qklh9Yt2MLM5tszRh2q3qLLaToFd+0x1K6IeV/9GZYHB5SitloB2eW2tQZQC
ebKkhwkYc76z6FmapZ2fkOSLi3onaAKSE5qj/A7Y+6GMRDmucOQYQCp3sl0DaN26
Kmz+UhhDFzc0Ffbit7LBdjHUbjtR4/j3Lb0pguUsOnWCKFgR/Tbz54up00cJ5XgJ
+dW+rhCgtYTi3kr41mhm1uTsCe63MU/JkIhPqGzLnmDzntxIViXF5fKruzj/EK5n
Tt+ED8u+SkrTF+0azyz2KUNNG5xQ8Vwhm5Zyp13/q26PJbr29sh7NqP5QeLc07M/
+5lGY8+wjgxz9Umavmxu651ARm5hq84pbekl6WyhQ9W60lyOrgE0C7QYuTZxB7Te
CI7lIzCBkQPrkfaI3NIfrhoOvN2wFxEyq0oEiAbq6SyQY+p50F+Lv3xqG9z5MPQ5
q+7hRzsPECgkIil23w/MRQeyZd8BR6FmdSlEY8vMgw1rLw9MgGMfGac1U2u42GDM
VS1LcW6XtNrUUd2++rH+mOHF6i845xUWjBiHKHeJG51UTn6ACPUOILG9QzrshyYt
FwCii/PMw0EFh8J9ryLQt7UBdVCUGMRbj7lu/fgSuGQpt990U54FU1vlFkWwiaY9
QMK8kzaiWUfIzUSPgXQRrtApwYcuMTNbBz2RlZxdBtrw8w/9Opt1TWsV0FY/oI5U
vYfFaKLDEB6J9Cu4fudJ/9oQm5EoA313t3u+ztQ07oVqnK6PySK1x36DIBpV3Lyw
nlyLC/+QneA7iBgtRjFamkzX7es2jlWgjvDpt5Ula5+N/hR3ecyR+07ltcI1Myvj
Vf2V7VBdtgHpjyTgtc2SjIzdaX3qRv9cEcoY6UUouAjpHIDXDR5MaRtccO3RJF8l
wmCqPCP+pztDaSAZPa2UAEkt9sXPUseproR5iYTwEGV/ob+8i7HElKKxfyPe1CVD
c2NzVnuGoOOJID5ZlaRaAiJ7Yls5OE+ySPGN/+UK2ogMnmbhDNvxlNekjPcNJ688
9+0e9AZIXwdkzBBl/xkh8qLMgk555SzD9u4IKY73S8wsOuEvEF6sJc1hIsk/qtmH
dk4hoCGE8F/qpxcDCuCS65+nTLTCydRteIG+aPi94E3DiwC5aWE3q5zD/khBfHaV
+Pay4dMKYop2pNH7/Jj7SDRnv27UglN1zRzOijMgZZZAoCa43wxNPzyyizk0RXXT
tp7mQsYTQk+o2Xgz1hioICCO4yI6pyc1V2QIXiWOOfaUt6M+dtVCSMoYqM+HhiKO
jLnw2fruVlCbG4qrsKi0c2Vk5kP4Sp9WQTzVpyGXw0y4i8O78DanEL4ve8cx4Rip
++v66ioBUOAncSuajW5//uSXl2RhXVVfZsO0h5bD2jugKFLpQNm8/OP6X4v5PKPX
3UFIfkSyk9XI1Oy8nKUFKNZPcUhJF0iyfjnAclZjzjaKCfisNGiA5Bc4XdYDnecw
0rFtI3BJO9XuODmkPJ7LamLPRQXzt/E/wkNS4KvL6aEWVo+xhErFptuoQAZEmNx9
ub9nv8CfaqQrvY6vRhy54eVJTweCfbXhCc4sW/mHmCvD4eTnFllpIoCHpZ0z+a4i
GJO4ntSRcvEhSk57AFTVMskJRGfCMsV9Y5cgeH2+5G+p4a6Ni6pge0eq/0gI/cAk
NzR9ipXQ0NB+lcCOxbOevMqxGmc3CrDl/64gzj02MgpND50mNsfKdTarmMullL+L
uaccshpdhMfSlluAwiNfnJiFYbHtx+5GdfdkuHKYQ8bsIvi8BxYx8HysZo7RD0yZ
W8kmQ57/WLJPjx38JIamCOEySa63cow0T0e+gBp9nYgIQvD2c0QbuZdlML/3HlH6
vC/4AMd4n5zz3f9QVTx3Nzk80zPuzkXKgpZVvk0zZDR1lAX0FF1Lsozj8BWB2zMb
CVU7i06No6XwHWxu4bLIaxGkqU8U7BrpSfHdDqPsM7d7K97ESxYgpJZyMmyC9xN0
G+acLq9tEy8yigE6Rc0ruq3VN1W/3UsPF6Vw24/z3rLDJ3WHALjRDCash9QFCaQP
6u/oEDGcF5M/+TW7+D3pOiLjtsObZ1nl/XNG2uCmcLqcrTZ4DZK5oyc222nMOnNC
nBNGqscGGZ/ZVorxQ+Mdn8YvLxaTbHrt5KRiKrHa6jvbHjJFKxA51d0SFubzG6Eb
73PsvOE/t04EkIHC+94eHV+nkb9w5S1tXa+ORkYS1tdNTKwYeZFSpu1M9L3RmNVs
2b/cfXDAPfGY6gB7jvvG2ox8NJK58u08fohJLlCB7lO5yl9cSm+Az3qIXkUE7wZy
7gGW4eUUiPNTbJLhMxuXNfhWU7bWOuxjf1LO3XSdo1ICrNZF3t7XQeUIGai5nkLM
XH90OGPj6+W3tnX+1se4hi8taT7Ds1CMZIHGSX0cFvMz+H2wm5maUbUKiivFkkO3
+oXaeGcMCIK78+BRo5J37Q8VOmADAvYcwNzBQA3c+80EKBBEWElxeAW2pmEO+HBV
ra8xJjvkJs78nHlF1FOJt1oQRHEzA/QmTBhofvjrrhyPBrec4x086Cl+0nNQE1v4
xvQDgDTod2OkRCflyXlDbe3KfPRGdlC6K9hqrbaYRWf049Srl9pPyB4YuDuIBJFT
ZnppE3qITbUd3hus/skbyghqWP75KPSdnx/H5CZznuF4WuKrx5KXptXQqaZcBl91
KF9uoYqwyFNvT2CFg9MEixZZsOXzWEwW/En6FaTuFbtCgBWPFdp0ICprw1q5NmRw
9Ksrr4k7vU+XWvKWQMs7UPIRAG87Hrg6O6RjIeO0st9z69EGDEWwasvqVYzPVgxW
4vv11aNX5aw4f8e20ksKY8dZJpoNvvO089pN3de4QUfoGsM1wAG9jkPpEZZrWIoD
L2IDOVOtbeouN5EqBQboFXs7SGji20isFOsDsqWHMGmOoXv1D9Go99XdpOebpb4v
oGTgtvsPtanDKnerMF0uuMcSFyzhSYX7/MrZB6PcQiRFzj5+jkUiEreYwiJzpskw
eXgh+rTEDlmG15DiJu55zlxOA3tG+RU3U33E9ota8oJ5ttv5v7eD/0ZbX26QuEtf
vFho6/gLOaFfg7mlJNKINkrW8pyKmzF1v2PMAZgB4GtVuriJZrp94yJCYCEnU+w4
HAv+oBzM7G+jzoxUuM+jyLGd9hUfJlHNNnmNNT/jz3msGrnVVoSNe2nE/qt5BQku
mTo69Nzzmlxa4A3lcs01mwtCH42tC8FuLT7SUDdZZL6QeW1xa5AxpCowu3WLGFV4
Fe5tJ1QQD24uQ0G1aPMqXFIDeAVY2ISSnxlNNf9nhiUQfmWFyiNTqI7SNefRl1J4
ffO6LW+10HoaFydgUpjeIEnICPQi+JAez8mPKAy0TFRwdMxaJ1VIW0qcHnjJ5IfX
d5D7+k9Z6nlInpxJ04AxPJwxo302TltE6on1CJI7S/x8RIGiX2KJJWpImEdALLrc
bF2e8OsquD0Q9AzSpQoTD0l+GHCSGWybOtlvH/yuBS00aS17ok17b6NnsyKbSf20
UonuDNg5eAw/wglNYf7ussqievQbwloVm9dASh811FWQoSS3j6g+5OXK9tT6ZaIJ
jNf7pm3/APdRvnbo8dHu/1Xr4iL6Ty82618qEEMga5288/yMAO0pyBtyC4Xx1f3v
vWaCr7WljljrLAht4q1/98Y+FWm9NUnDhfZ3Z91pCyM4rUPJ6N8Jl0fum20eWYJh
mZ6jkVTxNm3k3ivfgCWLWkl7I468cWzns2ddBCu7iln6TdSZ/JaR2gPR2uh4BGd+
93DkCHPWwtvFVeMrg3KvoVhRGpM1/4DrWsJuR/tgYU4ohJeXMyLsqJHBosJsYBP8
mPR7bHqdXCEqW9Q+2cCpCoWf4Qro/dcsaOAlhXev3az1NqFQKJiB8pKt2qnJsUsq
WgZMAqihqsn/HuSM5XPMy4iZB59F9ys77ti03n1YSkz3aOuh8JVkmnTWqTXS4IbT
bXsEam/alwQ6K+SDIVwymSm4S1G/Fc9ENXInmITmUlv5gxTgmMAabyke89FF3JWl
Bz/Naw2ejQ7echAwgDxNcMCtcMabUCCTkn9+UvEW9AVOwXqrNYfB0tYVLAMRbf1V
G6kS+6kB5VuI/ZZTMvEy2QeWSsBUAc+ep1DpSpB8ogLO/ejKKbnHgCGnCV/k6l1T
CBisgE8JsPVh50Vm3u1oUXCIaOCxLNMsrKdVUZLvaHqZOqDW4ZccLXpoSAgMxXKl
rf7dKmaRcRj9a2nVd7eqwM+BbD54OJAMpd+aStd/6oG77Wftsh6mJ903SL1/Iff6
i9Kmz49q3yOhb6xE79PKcOI3sZNzwRNbj2qppoNX9/Wt0BVV3UBMwvUvFnSbcNYP
5CGshVS1qSnROIDYAzPwWsW5ucvk8JoobKANOkDyIAK6qoTTX/2OfHJpkkgoytA8
66EvFQCMZ4B4yNBHT6pb24QiZCXzyNr7M9yc9aR6Ht+NswFVS0fuNEk57Oh8fGTi
6rIiX4bgAzT03YEQ07AuqKw1i5YzN/Z5+8tUHpx9LTqzWTxBVAaOevWoKxeEOwrV
KlZvC0M/J/5Or0hzSlc/xQj2OloX314FIPpOdlIad6l9tOwVRhd9AjYfH2jgRMl5
I+uvef/QvTom/DKmHfY03oFdAI6oBXIvdpVyz173vbVPwh1CgaBU5O2pOg3zPe/N
TgNpMqWH2StufxxXYfwFS5osrLG4gMb8XxJbZ3dA663pivUxvAsAJN2tpncYfA/I
Zf2h/PdMgJBwBLI7mgFVJ05FfccqR3dDJsziQRyDSE4oLmf9uF9fIqnMYMT/VaUJ
4wmxjvi6lAK76hAJJwa4B38WDjWkkBA/dvJm6wS1ScS2EBva195lukt/TVmS5pGs
Xsy+wz1GyEmsUAmynQTqlyecgHBuWA6JIii90UMXlz2Jc1eiF/Ihv1BDu4Zo9fUJ
TlUiKc6qGLotQhLzpeURAGT1xhDlWLpSIMphheSROdStFCk0crBVaceTokmjI8cz
DP/ELVt8n/H3WzsJvna/QoKk8zZ09HiQt+i5jCf0yTyNthBJfnCXmcP9byAcUoEB
ZkuznSKJwloxuIK2qkRrWQ5uMFTQy75qLIgqBhNX6mSH5bXpjAAWyK364pi8+h5K
LfHM5sKYYyrQKpBXJG7rRtxdmnBzFm8SqwrnZdfGP+I6HaFcABVRw/knsbKXe4yd
m1n2l5izSKXNUj5tzrYBNewF0386XXbCZReZIztBm8asTIoSLY6YPdhMaoCnsMNs
B+Vt9ZVR9SfEOzpsboxhP0wpqKilDw5vs1VpkBpZBICIoL4L6ggdkiCUhALrVC1G
OmHfyMKeXEJxyWJCvhjglvjZM1GXZrW+gyl1Y6aLthQQr35yRiEh84UBRg6wGemP
pEOVxjFFz0YfW4j5Ey5i2j9QgpeIIK2k4AL74MBR1AjCgOeUc1pEMrBotZ62ZXpj
o2CgxiMhOrBT4J32aoFshM225t8Q3rYQFktGctVqfuD4XVBukd1gQ0kdxx2AK1fG
2uPpHqG0B3XG4SVEqzJpx+yaohgVlDlQA8/DBD+L4KD9gegs7seOdl0QD0wiJC0C
yFMLakfbU4+Ln7c7kFHC8QzCW15NWxjaYG+NS44xE33ZIzhSsLl9HUg2uS40krMz
I4c5Xpo4bGybwA8rmKoR+cAS+W158TRZFzJjNLEI3WlZnfaiu0KxzGeHFDy9176r
szSK0MC857FdkNqCM1Jy8I73wC1qMrQr5+u7ef1Yctk0m0ND9kHYIJpPvj0r3EaW
6ILHRRRqBwe/KAif++6P1w3FRi6N5B9Mwxcc5Ycqn8rb+7rjP6nGPWquZW/FSqbs
NVqNBFDipFLZHd6T8p68KsDabCLiCLaO0Y6XJyqVYQituAOcbHvzZWg0r128rrft
/K807VwimCgb5zUohRAZjs2bj32SGNMvyeg+l0pTxBrxDRhVpmJhxqyGkJal/OK3
X2YcwsZDkDclREs94F6Rdv3pMwItLbJ15+y/dqHjDUTFQN6+MDSrdjSzpZ+GXWEK
cVmqYFTJhNNZFn0HMJvIMqZUyHL/UulEFRHkXAh7soh99mk1nrP/5etB551DptCa
btFv1OO6QgBBXtjMfgebtH8qAYutEX5FTCko/KCQNYXcSOXQKNyn0sB7HHyFxkXW
6VQOlp+uR2QA4lNhGOQ/KZ+gaZEsawZiDFWk4W+GRqDFfcOCjrPCBDnnMI2ib2bj
3FA0cYTa5B5F6015R8nKTMMCfhwu0yiodRpbKYfSBdnbCYJRiCcr9y3GgA/xqPJ4
alQ00Rh/x9NYYUL+tnfRgHphNtdbFUDI1ZU7fppa/Ld+As1MJwWFwJ0TJSgC65Js
dfUMtv8YkDLZEllbro0b1LHkrf9+EIIkuDixKX4h53b0bQQypzgaMTONtZ/kGg2e
2ZC2QAVp5YK1O0prwdsplVUJsujHgLmF2mm+4kbGNiqcO9lSb+n1w9XSV7QSYj2w
MeXGwhO6UNFbabXK7imbUCxfQBPUlXVJ9giuPTW3ySB0cNduHUrXI1gqTnHWKSZa
fB7VLL5Dub2NqrOgjjpCXobKTGxWm+Yj5LO6h4Rc0SMMUlxKrcEiRmaJ8P2fKcwv
btDazgjbjU2SIxNEA0FAqHncwp99BqHCWNlW1M/sCuhARyKdJNUSZpFHay4clTNw
vNvPx2Cc5YlIq8Jly60+0jOFAr6LxNEEu3ayWaus5EY1mvkfYcqPyzuiMKW5udXV
5I84KWb17kh+feWR4OcchZW31Oqer62fh24FhDmKUPHyOkO+XneN7R8ODBaiM29w
73T9HMppMWSPS19Ex98qs8wl2WXbHPY+Ta9mnKKpGQHolyAYUkMB46fMHjcXEPK6
RLnmyEyNfNh3IaYBPydIEqjgdUTMCMrlIPGBNR7djK0sDRwxvUe+YELE2iO/kpNy
HPZGRWVOQgtcr0y8JwP+Vhq4XoMwh6IYyOrJYa9Yz6JLAojxT2T2IgTAT7PFrzU4
vd59LzXXRTK+VV3OYw6kJyhHiKXLz6RKYmeMaPxrsSdrC0Z3VjzyTspPyAFjQXEi
1ONGOcWx8Yv4MsNsWD5TSDc3owgT5iUWooCRpZ5JElRuBrpGKjASk9zgK2FBmR4x
kVVDObb+2mFUsw9dGPRayXvYWXoaaz5OtXoZUAZD6CBsoYEDe4gz7fesiu4NUqhL
hA8r6nPT2I4d5CUymccWWOZsXAG6y1hWIopcXdZKsKWcoSn28OS8Fv5QTHiViyvK
voDV6cQW76dFqlNwnikUExB8CWYO5flO/woDJjRlJ1cN8184J5N0t/pN4Q/QPrfn
hbUO/4/mh7KPeKaUNyJUsuI93SJTiXMvsS7la4npCA02dsdruXwftTzA9B5wLe0j
gZnzhtPHV9Pw8QVDUwfE0ibZ0OmmTGd3WEv0ejixuc2+cib4gBN9Fe6AA8OXk6lJ
GdKvH05OdcNM4ni8Zx1KlvPjEV6RnMeCour3/1glYu8WxrLrZRu8ghvjWpC8KPLQ
V1CCJkPra4+jIvtPJpnKdIPgFFwej5ky7b4UueFQOzUEjvrarxpPKiYQQFkJBVqy
6UikWX2fw4+G8wAMkH+G8JkV124QA84Qw4yRXUXBGsLWkqkHG+3v4jtfpgaJ/jAK
K9PsDi/oE8+FSuuCOwB0b1yZUoEzYYI67SPrc8Z3LbniJCL7bcWKLvLwlH1djnBa
fCPI5fYCr6EfX8kZsUxU5NhPKxlBfpdBwuCJ8iSUfVw0ZMI88/0gboNwJNfvyxgg
Kj9LwHzx8P+j8w+wLNavIH5lBdSDNjqxrNmC384S2QRE3+8Uz067XU4H3HOHRZNb
6400Y/Eit7CoLi+Gy9AVx60PrE3HgLI4LjfP9tmryIC8KdmcaeB9HLSNJxt1XBa6
gCsbMUtQVGwj4YMy75evgc+/xyhJhDJwD6p3R3IuI9QrMqyypsgXHHIoPFAPFhYy
ocMf+bmXdjtPRpio8tNkmXh+EMgjmv67j7ovTncPieYxuzu/VtPQVjZivCiUIi1B
9XzQz31w9g69UKQuR7wn5h678+bnJHaqsEJ1RANBuulgsmjqPn6QtWeAxDlMxy2M
2XwiF30pzaSaJsxQkMuGGgQ0m83rg4wvzZNjGn4odtvrVDjdlaoHRLdQ8B9LzWz3
I+KU/bcbOQn2kibQYnu5P09dWabhIGMAV5BvbvS7qIL9j5pUq1CHsfcv1PcOydBC
Iy8dTMaE4ZsUv8vC4q+WLSVP9lydj7TOuz9KNrAQXasVYqB4+J04R/DRygveREmH
Ir1KD4yp7liRHJMrIhN2GX1UafetN6AN5nYxRWJ1oOzogQJx79Jg/iewgDXzPjuI
YWK47n1wxSlElk4M1/7ER0xPcz/wZNAd5HX3773fd7WRN8Igb3Nllj1u4isnFWGu
ZWiwgvVm7DIxI6UB2A/WpK9B0R2yumek50bcsGYzjkmf1r/S8yu5JkEZmABXjP2e
N/G02bNFHigm3NLtva/W25oS3vre8HG2y5z5IE5L919MzgEF4mfuCr3rnitZdefY
ttHHv8zknsyEXPy4uf/qNZ5oCSKOCxD2+wVD6+9V/KsECTf5E8FeIqLS4+CJfKHF
rdJzwo0j53904UuZekYk0u6fZviNs48ftAjp4Q+jr2eolS0CnrDSg3euzPjQ9z7o
6ibqN9G79gUXaKK8kd+2vpII3iG9LXbm9JXrBCDzrAixTHA2d7nStqhAyJxCLr5q
2mN7H8GN4wTkaJa85VY9YCkYOGh66Suu8pgLFIfIH29k2+dyD4e8ofVze9fRtiVM
GYmZuvAdPUtHzT8vSu49wVmWSyXV6UfhtHKr6v9PhHHqIA6HoNykqxQE6wIsrg1m
tTs2rGWUvb5dDZS7xdBAoQvp0O5M4SYz3lPzsW36gS3yobeI1l00B/4bAjJ/5Qhj
4crIqERdS/Ky3PMNVjMa87lgcV4Wa99KlRO1P8RCZvVUF3QVpf8G569X8/LXLK9Q
zEeUYk+p2iBtQ2T+tpXI5FcjeP1chMwmftaHGjYOttwmhVseaC5yZfHIs4U2uroo
Fb5AgB6cweettBdXwe1puIHBHY1QpDGDhVlLlXKMZgk2p4Vk+vHv23MpNFbXzncN
0VKjV9jalNiqUuXOPb2MD9mUDzwTcoFO21f05UCCywCu98oQaZ4cpIchLDz+7YpS
NMX4W5e+k+sIsCQ/+bBDKvuamPzZiXmx6JzneGoqkNUwfJUUB0M3mf48nSeAXBYj
Ah5kzZp0CRAdsslnQuX0JdZ0uIE+K38BhlOjnFK6NmZXe8Ecnvg5rY35aEKdRjXZ
7d9vzDwBXA6BO8KivQgm/3wOcPF+Ch7UoiNmrW75pf5smZNFIkaxIgMzuxoT0HU4
pEidN4rwcyeNrjY+MRQdsPe5a8wBaQMPduJUs9oc7URIdJO6gwt4BWj7QBxQcbwg
NHFHGGcwTw1YDB55pT9+LbUkTQuC8MC5/HHcnVyxUkhhg7ooIB0/lOr42781CjK/
C4sKiFEN6rWktl0+klshmtp8kczW3W4WzvROceCniqqdG07lf0qTFstgNlZmyW+C
/RzI73TTbFdaXXk7QhItsDidGcpmpaNjOJ0QLov67zdFLKpIGlEkeMMHYL5Nsl8F
fu1F6sc/eeVGQXkNezVBz7BK1g4npgURgX16rWEK8Ar7qYyZn/lNT4D2jMXX1vxJ
M9M+tstZxjK+x2afH4v7RxyaFhTX4qR7xksqY9Q1rpjB4A1ZQBTXTJ7Jfrcw24CC
TIWAw+ujgDRA+IhCsrRvneu/UN6HqGdR2sJcE1nkRxVHpIZ0XkXbbdxdiplk5Oe8
NG1NGlAKpkikiQMIH4sWpUXbutqEUZUkRoOE6BIlcJQZHnRJ3fMiiD+Oq47x+9sj
aydAi8EqCZwov1kF+1gg8kd1QIbp0Yc1yZVNRO0Yu+6s4QGmslE+7SREMxlirfF6
HsgBV2aoIbeoDpjABZWtGvqpzKn/0UDs3wKCUkbz32TKU9ILUQiYaCU8rMmQ0QEz
/I3Vk4zB+eulh5jj50CHq3SXicfkT80uuDmdqNg1FIH3x0gZx51KOc9U66aaEYy0
zlD0J/WLKgDzbLcnhTrCPeQvwL9jfXlFM/hLU9qvA12YUaQINGSVWjJwW5e4R6VG
cTSONop/7AEr3w/4RK6P+No4IZIATIR7an5ASkA9mWrvnhSmTdBdJW2MoK8ideRz
4rQPi9OKT/bFQTlkBez5WZk6v174gAUpbRK7LGhtso6axurPGtyLzc7goDnj/nfZ
hwJz/af5gNMHFdU9EOLcN9WW3cEWIWaCWU9bVJJmB2ftZb8+V6Y7+UDMirES34Zq
XLQ5bGZ2sVsk9eTDVIt6dEjXE/wSodAeMSKwPygO4c5nF7IJtn1Ag+x9WdsD9HVB
7HY8bnjhnf59vs57u7Mo/C9IeKDSVJAhWcx69FG+YlvNpVhuosHDkg1UTU2P3X+T
xHbOZL7WiVhUOpn3zcsKOawY4vwUYW6x8S6+iryC39dimFtXnWFmRtq4m+0Sf7iw
JR3EDjIJLc+V1hrvY/pxqwy7c5UUmCxXwpg0r8Yz+Lstcb8ZulGwiRN3gY81fpfj
3fOHbspxytcNTvrhxptOMQMQr4DO4s1p+O198kSOL9X9a35/CsLAKXBKWw+RC5TZ
Y8UD2vUkZrGrUMb5MvtCcZA976pxYZXdqi/BNhsxZ2QlsTX81OEVoP+12LxXuaUC
1GhO00YXGccBpqxJ9z1AVlEPsyOL4W9VELvS7ATZbRs/S4vaiT7TY+ZU3u6bAHja
2rOKEJo8aIY0QdL+LZ1CkgeYkiAhr7L+oEzjDLbc+n8LIkRGzXTxFzAwfhTSjV8x
cgEHj8wmYanbiaXU/Q14I1c7TDPEPP+ejtJtEIHD7kvA5akn/qoRd+3Ae5i+fDgL
ItRBgGsbp4bscNr0DbITDXxGBZM0dkxFgZxXQk0oMLCSwk+NYm5bgEpFUiH8n5wj
xsT1B3pHuR+0pM+NOfhN5BBFvZTf9abdEjDzpaUiC8tHTMZO4HjI6nEkmthtlCqy
raM39O5+bXZTXCGTymquuDeEHQ0oaS3nMb5sYmBmtkSF0USb1MNyJduX2eePyc+s
LEJ5cWZOLyDa0Dev0GEPKwxbb2VkB6ZN3F8C6xZEk6H314rhWd+hDl3ysM2A/R+W
A+lDuAeiroNUQhtfFrlalzzhg16dHmDihK3TMgtlAe9XsKwFXUm9AAq4AB/gxYJ4
bP772en3LHuIte2qjhRVscpt8uQh+qC03QDoFekMHBFstdVaK0eHLzGoIAGoYmoh
hVPdg5/vBeE2Xl5ecaHHFP3dDtsjkcgRezrpM6Z8hd8TRzG2evCFFscae4OBpoyF
0zzsjdmkHWkyrCsnyoN8aXfS4r8tdr4XJUMxlrhdcstW+CpM7sHU4gtdxlPhwxuE
gbzyB+xgLtAGmSIr/Uv0/alsHv2ASXamrF8hXpP1pF2Ib/s7X7Y9FpYhwWM8QEW1
VgcWNVc98IoidQq778aJGGFCgbP4bPb9xr1bJbubB00sSf/zRATheMPtsKVRQmuZ
jEnegfyZ0uuuHcjSIMantnf4NBguzi3PWg02NYRCRG+m/vwCG9He1FIfJ+1gX+iQ
UnuZb3N49YiF/dd1cSJ4OQISEskCklwZ+vhk0FBLAhaLI1UfWBxv43vyLyDhyo1g
duGbke3cv+XD9onfudDTxIZO4HtG3TUfzR00ri9EIRDnugbQugQfxKMIl+zXvmiv
4ZS6sgupay5aM7F2CGppC0uLDLdEJRgRnIfE3bTf3pdomNMEQO+XXdyreRkM3ZsS
/vnK7FLnb+yrdK7eh7E7FjWJqoH104lLnKJHuChtEdbieKGxpv9/iwVNI8mBjFuW
enV+Pa5anjS337BHVkwG4oG4cL1fDpXZBXHgt2meqehKNBMpqWJfGA70DNkzC3sM
u2VaRq0+k6gjx4LHkmuyIpF7siWc17a/qQIKpThnIYQ6GWD0EOL8vbR+fbv1AiIC
0quJYAZXW8+gB9j8IqvPIHja6zjgnSRY0ytRyMgpLXB5oHNvafKNyMBwFaY/JAgs
IAEDYWD/wpx4RSOIWi+7QAWYWZiwU8ODkW1+VE1HZBhnlPo9BsCVIaBwXumRoStu
TQuTmRA49bazvf9LUkgLeS9WPXd7dAAX47KsD9nT7sB6H9r18kRPRk688AxKfXjc
odmy3XT7AwOE54A+rMQ9JrTQwMG1+l0ynEggNJQK9dMCGd9YhBMUdBniU9g7evxX
xXQXW6SZ8bXsV1veskOM6tbWbE2gG+WEKksBamexed/JLSG4nnH3bxK5frDwQGqI
a2I0+ymFwG3+hg7qViKnczt9gZ1McYrMTaXAUunOeF5bua3m+vnQui6f3X9iju/n
PTBb5SmJuebDuRWUeJf5Z3Ww2EUH+lJrdkPwBsjrblmdYtW1mD/ceG/lW6dkrlN0
WvwRCLE7CU/vtBlexheXFhA5UEcooh2yvyGhEMDdcbnDrR6QIKmNPWbTqZNIw0Tb
bdRPsnjKh2aD1j4KJMD9NyQfRUqVCPxlcCgnip7V0lu6rJeRs28xT4R7lMW3dRjd
1StmDetTtgWD4ql0gcjt/XxGT18vxj7baBHcui7MOGmtaLP8AnKNrdyJtSQkJ6sh
pFJxgslN2+P3dUfjMpmKxEAx+r9FUobj2IY0jtKYk2drzEUh6S1j8VLVlF7vdal7
zc5KcnUmInt6i6hSTaIxufHTCsDHRGFXSqU7LNWKLbkFR0vhHaBKrLU2Ycd2Q3Q5
08A6xuF2DkGPcfXad1fhgst92XJ8nFZd1GKPeAh0w/XeZpcf0nwq3jxbMvjzFL1m
8+wxucjTcaDmalO8ID1r0BU+ksx/fyvsDbQFpF35IDigSg9Oo8fZYNO3LZ0R8oJu
QzealR9TZ2hTDE/olzXEipMvALgOoXajzu1++Y6X7JK0WKSY1XLGMhaOV7tJuodq
lMqylypIavG2uRTcicbgG58bqHgrrgZK+wz2CnBtO8pixzsD7AiDxBmDxx3uxcHj
QpOvNEGfto8mVGBRFiw0m4cNpCYJDtbmVklj/daqEL7iA2L4A8cdYIzc9ug1x9tB
W0qSLgcrVzmuWx1SSkKvw7vc92A237F+UAe8dZ3uTyNNLHtuPZ6hh9n1JDRajZ7Y
QrSXe5BINgbzeyxURfMCg7CFGku+ZRZLcENFzGsXuwQ32jEIMKZPNE/ddwxBAQp5
GB40XAyxEBV2F9bjoKiXAo58scC1yTFpN18Lplwchmpe+vouR8AGSZGSop/lW32R
LU+nombO+MhPsrdGKmGFw4OCO71VnDh2kyH+thDCcFxFx1cB+YoDGxc4oXTrKMdO
PSkj92E91O4A/bHsbzV2ZgyWZOOtlX9FRcRPLZ6Yck0L/RWjkpvx7NYPZJCwfVYF
gH3m5Z5NPkHZJPZctFP2ITFNssKIIbu2hJ9jVWJk8PZeeRDn8JESqc85HiTGE30M
RryNOAMUq3gXU3INI5tG93RL/pjuzUD7QXF4HxVCuwtbfjxD2+/5oUSVQ6zYP7+h
LfkUOUbxPsc49cbt7bO5yUGDN98oeuTpmMpwejxN2v79+DMPPR95hKDq1o+WaZCF
BZpIOGKKwTFXcSZz7qQjl44ugFI8v6Uc6xePSxXBMEBBmjWRhsDEAFLbYGzjNKWJ
bAoA0DKca70HS5AYOxgcnsBQqso5Xq3vBR8eLzCGkarEQwNmTr3wPgM1YFFSsKM8
qTnYXFHnkOAkG9t5x5H3Ftq/f/BvDLaziYmHl4AY5B0S6w3+cByIADDAb8YTKkMZ
sedpIoc1UbOh3bnZPwZSxvO0faQrhTGQZu1v1/GYy2IDNt6okjFDH0to4kuUP95Z
HjOj+VR0eH3KiEVaGCA4aZgR1K3EHzYXROmg0/vpjna4HqB948HaauTIxucK5GTx
DHf39qhjYIcVy9OQAk8HN0AVx+5XxEa8Saa2lwi3VxYrB58Je8fNx8QIBY0vWGCI
YbPkGLJwEoBPZmGJ03bvVga7xPrJt/QjhSzsjI2WC/StV4p5vCmYfW5SJWlHVki5
q+x4BcjvyfYZhYmgHX24eVmPjl1xmv1GYQWuSw5703w1vY3mVAKe+0/N8KWxIbF/
hLfXavuemqaBfBcHfY82VgdVcOxCTf+WKv07sEW4F4ZI3kf4OWT9XCGLGY54id+b
Ne+Btr0JYRPnlTsoOL8wr9tlV6uRg6f+k8Ks502/InYrondeSY3m9ulpeYr81dvF
wlg3zgdNamarr37/caj6EOhr0PHOYix29Lip/NqREIfe+6FP0SsDvnzYY/UDFURR
gyR2r6s8Nl7cOh4UwUn2UhnHsXT2rlATRI0SOb4Jo4P175exmgXHq/wbipWxHXRY
/p6k7BY5NZvK0btB55M2uNEUiFSsFn+k+opZSpdJXl1pqN2T71VHkFGHaFkZE8kN
1RY8A9AxB1dvNvCaVGdAeZ/bbuAn/A47WuJdzkPTX7FwvwxVIZ6GntjixcbCRwS7
80pAYmkbaQvF3W+0Ir5ETcRTluMaG/4euvqEHmPsSoaUxv/C/grYPf/4WdVVemo9
YWNFnkLNoT/QWvLpDPfdBB8Bcyn319DMAw0OfamkMeTyadINxu4hszoppTF4YvY4
MiKWO4GanI6srrwnQfF+mAemttJn3Su+SINUqdFKxzYgJwh5bCeZtt4/pcBPDoyr
0TNxOK7PnGUMLscXlPAR5hmQ9KF8BYgr5ML2KqFZNzBzMIrmdH73TL5qTY56VSob
iE7zKZNV1jrg6gkmYzoghFQXboBvx3ax/nPj6wJrxmCT5W2EgDn8oVKH6dOCRlG0
/ZjpXShBR+lxUZXNsCuCOc5tXnoYsB+prh0Ga+VuQAulu+kLEtRlBXuHRSW5Gixo
dy9drtiUG/LabwV4jsPbyqVVPyESVz4SSWOA5RJOZ+wAqCNkbYtUkXfRzaiD5joX
TE7DM8lgOWrG6YP8LGXcPuAiAfysBeazBFFeFxLB1Xq5Xvk33glphstH9UJK7Ptk
o002KWL9+zVTlr4PMMCYg+4vobO1KHQZJAz0cmGWzItdwf87yfelYq2+sBaTMktS
kaS2b48rUJuDUO7k3iL9960wlpiwCuvczW7QydKDUeRMsQpgsvNDA316x7hqPtyu
ntOlY9t6/jpfUVkgfdqCMvQNqowi2Ze73AQFnUkDiRzrTVq4bqrGaREMNvLPwy4F
Gdz6dH69mhZgXHsfWTGaiYxSV/27ooWsxPuHI7ayoKtnFcHnbBabKuRSmrU61iPq
XBdPgpegDsyFkzwkDyH4aGt/7RrIrhZu2HvcmmGnV/yaH6Uj3pn9qzyiszxi0JX6
hkf7VBmqkgveCgHnPj0Qht3qwFKopuBmy2qQMFl/So7CQgc1zpQ58EHG43XIJe4x
uDuqKjVcKSLkPz8WcLMtrNhLHkDklmZBFi+nWHYnnn7gp8WFYkye1OrOcSd7fNU+
7ZQiSg30wnMO+KYPzDIMs/oudWOlmEH4xTnF94b4i8Pyk2WmzMA5yA4yxaqikuUR
C6XeZ8DU32f3zi+0QXnxUZOf2NMJ+YTbzqMpHK2cKrIxzBYl6l3FNs/RKoQTdtFO
1klGvnC4mSgJwBGqIjrDfUpVSTGSvJl7AmMra+SmZVrAKCtiw6gEn+Dg20Q8o7NX
gNFllz83MwtgPaEOt8DwZpkCQ2MtC/LtqLyu8PBfOqVUEoV3J0vNy1jKle8/IeZA
O0Abquca6KEguq5ppUIqbvA7K4R7mtZk/DWRPBwUHR/9sIaS0f5zsSrXdifhFc9c
2SH8g+4KrAzRMGA7fURN+51/wGGzxqsCVxOImtD8J/8tld9aaN8yrp5kQ/1tZjTo
b+380qAaii4G8K6+5NOqWZna/cz3fp70eDsIaEbucArRVUNo1orI7oqy7qxGZsyy
DClN+MNcrbv/GoZabkOKGOBcouIv6ZRtcMLxCGJBAX7XS32QP/OKP5R0jKSMXo6U
nHF2IJ0TQk2wc8UIQrHYovIxUI3YjBF8btXIBK7Kuv02Z6f3KnOiByFDYc7Ji/Ra
8ywaJh2nd2HMDJH/ELsU1pZKAPQyHy1KVwxfmaecoHiFQPA/CMF86XpfoPEK486B
f42sWCVWjSDPSEZMC5fsFwU6BBKBjpMEmQMHHoA8gZqC7Fj9IlXsbYjT1zImPOm0
bYqXhVj6BK3Zy3jpGYH+85EYkZrLi/ojb1Gd2KNJaxVUOzO+6T7vo002XwPAm5sF
HjPk5gwV+jZuB8QeVRFK82JrTfHoWxoSyo+u6Z5wVVtPU4Y7dJYMbDU48B6pqRke
2Ows+rjS0i0JBARozlXNPtuXo85nx5n8c7PqdKfND+nyfpY0YfWTst7LOaWtX5eE
BGI1RdOrpskOXb8MLXXxeZMY+XH+Ov2n65IJ+gFjj34lumo8SYa9KEAkfKL1t1D8
pgJv4AoRAf0+tLdBX5wa3+S/ID5gUwzPGGjv02x0YnJfaoJ7qk4oHjGAqVE85tEI
HzM6ND0Ij/PctX4B6kPabNZEuN7miwkt7v+5zYaeo9Ko9r7rRimOedBvav69ER0W
rKZiv130raq7Y9KYDl17UpH8WLAGGvW8sPdBeJ1R/Z7KLiBJTVENesB74ofbritT
erDcqSgLZtqROVHdMa+hFyj0XnI1Do8o7BuSwkVk2fWIVqZVQSEm5wmsvakVKBo1
9v7PAfSerwoZp1gwNNAs1fXBbNQ280Vsz2LGYkkDgcdW0vqlaTb8IkWBXIlB3pwi
vg03lbzeBqf8u/gFFvZIVtlSYnOi/N/18l3WTTgYjdOcMrpxXYFVoyYi8iQKdum3
XHiIazOlcKY1cGTSV5h4ScpRtiWVvQ2+mOjqCfzO+6n4PfoDSmAXj4LAi3Ct9nxZ
zKtSWuONHiDpXI3HVeMNutB1CXy0+RdiZVBBOeVgODRt7H2rjYiqL3YWCxOF5rQh
Do9NJBjpkOI481l2X/wKzvoEtkPpP6QtDAUrTG71gP7HpNsl5d/MnUZlRrGIs0fD
Z+S048ECuWEUAiRKE2lBgisXgr5hNvc+V2Y0J3mHfgdQtTj/sc46di/T2l0FlEzp
UfAWET85EcSwDaGPj/KOy+h9t49cvp7uH+waqbgDYh35ohQsuWU3DZsU3FmBUz6O
TcY1e+m86YU1uzu+seRSX27tvZZjah9Ah4ZzbDYtD+9st2TBc8MjhcJlJTpEx68f
Cx2qJ3PLt1fkFC/EWzxcas0TAgwrQkHmhl0mQc7KnCGrSQEUAH+PCzENpBVITcsa
Wpgwel7PMdlt9vkflsIVJeBBHQy74ocOtpHqQPiyrENU5Csa0WUe5tdJh7d5PvwX
/I/rNNU0FGb9Pp6iIk6kd06pnzAVTy+XPKUmwpPC+PlutEVFED9jT0ts9AGdhLxi
I9yuDa7QTDcJwZU2oD1Iem6qd+axqmPBHEsSat6qdzQMeSnn0U0hm069tD9om1jd
W7GaklwIR0BsDoX7Kd9gH+fIMHzb3p/0tWqLWq1NrL7lTD6p3zy+CDCqVATF3vFs
7tCieIFuITcyAMwIwiPP0PKusIhocC/VNZNW9QNqeE9rZFS0zbxbDvhSNYaXZq/T
eYqf/9T7BFYlOY3K1oXS//YRmPAMBt8Wj1SpZJauZ4ZWfCSYi85P9NaBHUY0862Y
ul5cq5jwfqbJNdrQbCfs0PhqXr+4N4ew4aUN/6frrt/3zSeFmSwRLx/3hXASvYTW
uCVpsJ9o6MSIEKIPtM8UqlcfXWWgYX/I8zDj6z5iRnauhoW/FuBpWnuX3za15o19
9z2f/oBKUd2GaCKRUz8kRTEAKVCuTxwkamxImntHvUNpm7fWPMoamdfPtufzvCQK
CnKaMAnKxbdpm3+yRNEG5PzWvfDujuodBxXDo1dA403hGUZYdvoeQeRQ3T+hJtIY
KJ/tnBr0JvKnMFpDNBcOQeI9z+rRLb/4a5tkbYteJr9iBNMcrh6YqeAflASoqoAw
xlkw6/ZMXeKAFqTsU6c+gXrswjh/ZMrjNFYtPCvJhCz4FAB5nVE12SIpAHUF1l4D
jkn1P/QJlyv7C8nEbSS2qcDXSCZDsAJRlRP1f7UN5CyiyWWkcu85NqCDLgkVE+/2
Gl3GpW/FLsdHv59KisTuC2BDWd7haZ8th47n5aX0y3koWq7ayFI9ixzD7BSe7pAp
NeywyysUb7GTwQXqqe4OJEGqBAW+EhVFYighoTNghDQcWISWoZSWq1OyAdujFG/a
EVxlGisigcQzD779K1RxuRqkb/X9AGh0f44aTIx71jPyNvg1VWS4QU98tK8dSgh2
vup8VnBtm80RwXwOlcv5xSDIot88kkbEKIiTXS5v3HYYCRFgFCIAhw82/AJ0r8Sq
T3ziC46gVXrQPpDtXtNbDy5lnj79kWXlK3gXPQa5BK7IdhqIvU7kr1CfWXrtJXKb
qgmyACQLGRUtexfOWdyhsZj4UdRFIS2jlteVZr2HTJvr1ZeLBuByUQpvlaJAZ671
bXxcaMBF/bk6VcRSfhBztl8QxnIOhu6hxnTmXpd7dOGOp2zppp3TL/5K8DQyhfdu
0PbOdByLwMh6dkGZIvhhz3kB1g0OxtolgLKFofOFA7uNgIxYB48KVm91SkaPZwBk
CCA+ENG9sKRPtY5Vb4m3eiRiG4Ys9CFHdF2wqoW+oCQ1V0Se+w9jSQZbklbuqZzY
+jsz4e+OpmtM9UYCkWDwPK0wCfVe5pBKQU7sf1sFuaXpm4KvgFs+2gjUxeNgehHu
MQkq28XrFKH/JqU/UJk4IOY3DvGXMnvDq3N3veY1akY2k9N9jtB0RyIeZb9FtvQ6
MYBDJAgatTN4LaqHvCpyDtr/lE43VhI/d0P9iwzGuIUARbC3S42rxentHZ4ePXOa
Qgip7FTp+VLg1j76P9A7XKgM5UGn7tx/LtYEDHGrX+n78dKOiq7wFpXef2yDbSVM
6SRUj2yerX01f2fVw+Bbbrkd87vourG29/cHBGxUitD9MflVfPhILRtrA7Ydfjx8
g/Aj+O40ahvKvM99oXxyTkNiZHewx7h17CaEePWRTavO5FqIiIyaIDkaXfkMkvqE
zy/RIuVpSmByg/G/dTg/N5IM9Yd+UylE4CmYKwF43DNhzaS/yzkqQNQpc8U48KHu
QEpBi3sjnKxJmg6x4cTrnJfwXbsv1+jUTrbiEW94ixmXLBzAao2WP2JW9VONt4cm
Rb2Q1MKgSS/Jev1jsLgU+RyRJq3+cVQWf8keUoJnUbpOwiFKvlt373c9OVLEnDPN
v72ZISRuAfgk3O1HchhRxvkPErLeoexEDYwOn+UpEsTQPCSEQcPG8VAtE6Vhzn+K
JOlLDs1lAGKBYkSydduEcUqTcQvYzLEtX9Sak+2jL4zXHrf3d7gxMzKD/YE2b2Gb
Om7l1k9NPCetovqEUkCMyZZWEwNaq2FhUTBEg1GRuG3EcpLiqIDiFzIRK6QrTz73
7LyBmiLrasbC62mzqhBcM6abxitwsJFEeChm0/E9COFHVkmMHko5lLfGLJ7kfgjS
/sFLXczLazGLLwaEyAztiW2PSRIUGwAmBtnUk6er3jdXvyoAAqwPKRu5E7kVGFnC
I1mcd4pOrF67MT06po79jcKRB46qBCkmm8qbmrTnOo6fFI/H0ZeUfqW4xJ/PqP42
7OFw0U6nKQLYrjmvGvdckD1m/KnsCpBQPos6a1hkhcnW2znYeS3x3EoWC91Slku8
/Hpy0XYviCwPVHmItRQa2h71KAS6Ea33DOeHwgu0+rINGTCquT7CpXJ7NnfQ4D8A
qNW6gSJY3P9yuZSyebbSqjo+FVs4UMYuihQe4N473SVUbEEcbzvAGvm/goibJsbj
YZbcWI4h/9I9er+6xEuNsOKshy1rKy/MlhdI5gZfDwlR67WCf826NFQhmsESWLxa
2EG3Jzi6bEGGKks5auwhfcfsD+roJDvLwqAWzWkz/uvYogmpNHb8lr1rZKXfVsA/
Of0jm/PtHddnS+68lTofjpkDO5QkM7D24rEdTb+kp8EyCyWslW+OZ24cR20dyGBn
2BadlEml8M9r0OFQh8gePW/nf5KjJl/GCdf6Yi1hZcg=
`pragma protect end_protected
