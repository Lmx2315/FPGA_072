// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.0std
// ALTERA_TIMESTAMP:Wed Apr 26 13:33:37 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
hbFQcv1G4bYTuOKYymRSWCflsUsIs1tTxuMo9AQTUpaloPNFfufw7J+yx6oI1frA
JvYptiRus8W04Vodk3of3T5rVU+tpAId834wlYCRbIxSMHsZTiXx0ZsWraInL7i7
blqRN2MHBnbciHtrdWQ4Td98jem5Ac7zPnZWBQ6uLr4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 176784)
s2IA3B8UMvkXiXFmIsmG+Dul8eTKjtOZV8XZW54YjvnAfdP0Lk+tLREHznXgOmv3
oRAJ3w3FJdItF36z+fPYzFAWzxx7S+PGHWMpdE/EOOJ09PEE1sVHrxvtYrZxKk4p
oWN9IyMDlyQkTirR+iQUy48k7dj992yQhf1WTtG2QP7ki6Sqqv4wCZ4cUSjruHd/
1mp5oy8u2UdPlQxQcgPJM1f/UoLadXyoQM51SRmahHJMZk5m9vvjR+nS3zc9aWt8
TvsLk2WrnK+jRL+n4GvHqRMgulgx6y5Zv/utn3PU4PhqK49Ah+601sVPR6LJnkeK
gApgzirCa2zTACcqc6yPeFEzbSfYFWQruRDR34QVcVAhtuwlitsYCcMgjRPCoVjH
qJpcblXkja054jPLukwK25Vpv8ZNSt84AwAwxn1+xzWjYqbEafAzA/X4U5xF1KQX
1GPXUdbuFyZqz9sslquMI9ns9YHe/tyKQ6n1/lsQ7hOLkKvrbHcwQh3gi3L3a7gl
S22ymFJpkrLQ8S9WBxyOFbBap+djvkrtqpi9nDES4HxssuIAyQ/sVaaHVxbbwRWw
KHV93E8m3qAX8hD2riMst9zHBcVmI+/NZgY2iEMCCeJsZtS9nlU2awWaGMs/0nrq
RNWt84Rgvd3Pu+eFl6yRrKmVUyw3bn53AONl8gz/SenH+Jucu+ntRvPkUo2J/WJS
mccCsG3taSr6CQ4bcUVIcU8aTpTNNX9TFOmDbqs7MNshFZ8dJuV9xRO4MfK7MPus
hi0X0uUt7VrH71ZDBlusbvB0wMkkLHESzbwOhvKC6Sd1P2187TAmY1jqXxkSiwff
gcPMMh9R1OAaYXAdGHkT8cFMF4k2fMSFjfn8aQu6ZcJX4OyWTkFXnJH7hWZwB/Nf
7rZhyTOjVHHoY59BtVls/Js9R+lKgJJDW1v9yqsnY3F8EPqoEGJyqLTXhI0xMwmP
yF1U+vca9KHV5ZlWjokpPa7y2/LQtlBt+yiMj472wg43YzUMP3ufZnFiM8TIWl1e
jOQXOnasRyo1iIA3F/IdNK5IM5Gw97dwGsL5mR5Ih+DuLCRrSyy1gMeb6JqZaCuY
JPKAcnsAB/n0HiPTt8xZWOz7+F826k1fYwD0jQqotB61JF/7Ys+BBa+ByvisT0EF
0fqO0Emy8apkFF3crBjKQg9tlkkc9ki/IaYyQgLw03wTcWM8JEFbTwNPC9Lpi/GJ
kDb47BaqS3fkHfE2joHLAk+sSSwiYTVRlxo3k8eVbtfctiSMwwkAj+mG8tf67V6W
+vclXLVJTwKneORAXADnN6QqDbcWp/XkI4ERWKr5o+ETzH9A9fdlA9eSGf45QW0c
xitOt8uueyNHPnW/yFKnX2bWz6sXmiekMu+AxrjuKYQuS+OAgULpNnXxAI0foyXH
S/UJhNr00SjB2mcR7qTN0Lyf+dDaKvets3y0cI7M7g2WpfJJjfN+kRrS6CVxIGDf
DreSb9B+expV2Gc8mWZvtsmn8QoixLft+6qT2RWJFZtMqoqZfp2McfL0mp4wnVY+
sTNIeC7ckAnek3YPGMqSn1vCUn+6wXyCIhTIZnJ+2NneEHh2PVioirlkNUSL0t9k
KF7vjPKeyzfrNJugcsisJWQ9gj8ytIiFHJb2bWzrke81g2vbUCZAA+p47IqymxTK
73TevQzgRWtauxfq8ZTyKSk7cd6nF85xQ4MYyq9FIraW94+lCP0DxYU3w9UTcvvJ
N8N8nIHGh/0eRhbeJPc9CxTCnJ9fh29ysoxZLZtnGGEOzhGqOfUWPq/EOVvAdzgQ
tsmPAjHn62kCeiRB37uDlEU9NWdjcqxoHBiki9laWheER/kxjLd+K+BNHZ2e2Fkk
I9zlc0g2EU3tCqG20kJ6BXl0Pg1PbIZIT4X52Bc7PHOAXdNnAsKT44UeQtzA2EP6
RfAgBE3MJZm88TZWHWqKO6k/XVB9EUFZ1qK2E5U0otjqQQbteXG2hiXtLdg7GQDV
k+Q66MebWZ9Y73M8Mxs1C2K8fdt30iELvzc76W0H5J6yMEywtqtzipSF61tBzzqR
qjN62Juf18hdJWra0Ar/pj0eBOuwzE2mfaF785115PkswfhKN9Yr22yHEX3qGFnA
scCS6U5XbyxRQUdK3V+o4upgvemw/qWVXB34ch3yOX6Lpx+ggbLizAUMI0uvOxQw
ph1UWSHNAs7FABwgtO2Xi7igyfiMJbxjEC1yQAUCjXo0xiz19uS7V1t863U+9ncb
Cyfyw/jfQhRowpK2ixdE0LGRMNQjvwG8zOjN1qmMaEZgiLo5PgvUronDd3sN1v0V
lchSqsu/gPtIWEFg9KgDOOs1hUVrVTsL83tpUrAYtaI6RYaPSrBY3Xn7MNhXhuzL
+OjF/7fuVxnuf/M/BFuoCzUP2UD7L2DTBhaRB+z4GYuWAMD/H+GKCYERiUmky7P8
a8iddlisbffFB8f6xVSMSDJ3K+nZMJZUc3g6KKW92AGFuUYk2tBGi3ojJswcoFQU
sW00iiMT33NeHsiyYaVk8kgCX5Izmhcnyi+cQ+icIFLluFuMrCSDYXAQlJenYKiG
EgW/DXj0YJJo1geP28xTP73l6JmaosRMhqYzxcN4r+brpjvLeXiob/wjxxRWvysy
vNrYBiUlCzGWO7FJzqCkAIuvb26OtmpYCY+wkGJN/9wvWeJGWe3Qed1k6GPg9yKE
D1UR5UbXxD7vVnJDmrmyloyyxCTnpQNV2BM8Q8k3i9W1PzmbgWb3qUaBp3cngsGH
+uqxIkyJEdlXOo8GFlwhjGAH1wQwTMmb1SZSa+Bg4RsCUXvGE+szDRqo22mgaF4P
b1y9NM/c6i+yofPJp/glIq3Q4QqnQM8CXBN+293v8LDlC58BY2hryAvq2VtVoGuN
65pwv2i+8k0VGiHGhqk5aIGqyz5ApAV1F6D/UtbS+PnOgC+4+13jbIEki0u+ev4g
62aZolI6EUe3SelYfPmqaPIrd+TMg5jSU6UZC+IFN+3/jN8ogd9Uym0IcZjiZwfC
GR9HL2KZpXrJwilwsU1jm1+2wZ00t/zDNqcKOCzGekFhieT1CrUc4jm7r7LBNtv4
QBzYtPHXFTLMM0nSeDy6zegfD89cQrL3cZ+zkp6B7bryz0uI0FAPrxX0yH/Zh5Nz
yLTEhrR9v37+WznrpF78PneDlkfxhjYFwhszhJHU89+Ib6w8fVbq/QXduyI8BaEo
t26uJKAMLbqJsfjf1SPkZfYvmDbmjplWggbek0LwrEevltYNwvyzKwj9pRF9Pqmd
Z0IxFzsFiRN3UCOkrhNbhtO1InXuYRgplFH/mGJgv+qKYv6aYqnrmhxkTpVrG90C
MGCBQZBgbSIOBFklOuEKrrR1EiX2OdwQp6Yd51Lf9DiReUBHZQI0NF6ksUdc3EtK
BX01ysn2HhCaprKY+jAi36KI/gvWjY9lw2qYD6lMfwPRiMd2uSsSKSQyvx4W6OaU
iJwK5xXMZufrB9cnAb2n6fdfcMprY9reXVxV1GHrogKopjGEkNM2eBDkkHmxKGq9
C1rYUR4Eg+MVY4xadHhkDQoc3DF9ROXCG9sFMZ/AOOO8M4KxPjAKF1tTA+r/5WuY
DYwZTcGlghXIRO5YSJCi2sFAgw52RFNCWCiyHGXVNDiE8gIpr/WOudlT4OFpVBQi
Wq9W69ug3MtP2jaBP6Ocft2NoML3wTk++TldDQx8LtUkcMVQucqCALUbsYkxC4/D
0Hx0IR3JljmQR7CHOJRM1sZa8OKJK/UxwRS7OnHmLKtDGCtMWSr+lYBs+mgYzzyJ
J/jGr43bMgitjjzQkqPKQeP/RN6VwlGnPOzyWjGw4vgaBApRK44Lv901pr8+mEHU
tDw4WYNpLJ/MdkeVlneqBV01OaUPEQlnlvVVr27nePg9xj9tDIb7ZQFXQrxGssO1
4oOFURYRdmLJ76ZqQMCN4uVLMdpr5Yke8ySI1FRApnO0Sb5vmi6F3tmHj7IwB+AQ
Sbv4dy1hJf6yTdL2snTokw8T2jruf9PnLBM5LISRcLB6Nt/4h1PK3ESmlJJGqswA
EHMRXRa7KCeAhB4x03rq/h61NG2SAAhfnUH7BKhf+NBJEZDWiVCVpniPmIR4/7S4
TsqrMrnNrdzsQh4+gzyQ4GoY9tXpuC+rctOWUhVmQD+6y9y5hqXj91ShoCjjXVFm
Wq/q2eSl+8sKu/ypLQmIPcWgCltcvyT8rwPCWFnrseq/4pIc/PGTS2D/WuqtqKav
GAk2I2XcX1E4OKzFXvln4+DNvN4VHExq7eM0dnXEJkHrs6tbY8pt8h2p42YRovuM
/w8MATl94tGqErmxtEKQkQtQ440p4fCvsAcTVh4NRl0e1xJrgZ7HwXPkyAkS2e+N
/1Eb1RMLvhQyn/sROsNuqgF0f8nidnkAe8sFcLX5Tng7mXbl4OHxSQeWVcwNaac6
mzSd4l4LsIUX2KzgwzhR1VJJ29Sv9AC1c1Nu/mYjsXk1SmKKqCQRGN+239CQO6Ov
m8ZvPTOhSWvyLItLH/sjQ7VGWVZekJt+QUgi0lSG2Lzu7NSWo1BgRFIVu6Ur8gY7
7iIVTRi7HMXL5ue8P47rcTpXaNImu2W/hcUoBfhhAJQLsOJmiGJ5B7TD0UCIzqWO
Y60mGiq6FkgweZjxjBqAkuJFNzg/9Z0oHCQGLw6HLJShmugpTl14y+K5DbDimvN3
hTEMjCNsHm3YEZMxQLkqCEdl/kkYWFIeH4sVtQGKFPVGoBIErgIkEYLVWqpNEeOu
2sIK2BQ7sOlLEQZikRo2SAuUw0MpCJZCRJohQT5oxHPfXqvWTPSFcVbYD7/NBDje
hRNHDu5HBcvj7JAY+opPOcsCJd9HcU+iPFfwIc8LuZ41ymmCH8c+sfkhDhXXmYo2
HtwqGAX2YObW32GvWwflywJokasv1bykrLSq3NlFCcGluCmXW7Xa+dGqot8VspIf
fBUUkBMrAO9ZyckbZkfl2NrdpAX4Y6UTjgt3FztzlfMrHFAG+ARnQvXTxlrizbsR
E1oBA5WJWEte0nP7WjscwDxCZvAJkgiDpehHqUkgOOJqaBY8PDdsnm3S4CRxw/+V
1w7qUwVO8csV8BUlXOicVaF4LXXo+LJS0P5XOao+cPirqcb6EGFP+wdhyWqmesaO
oBuFoZjItWqxIpzSBuNE9xYHewgsEQDCGq2lpZ966fny905jOhOn+cb9qmgmUuiZ
EQkW4ZsGfM8z0Avt4f5oYXzxnz3n2HImNxJye+biHP4A5PsE5/Jp/qj0K0+PVuQr
k5jJO3YQphvzYcARE3uPAVb0c4mwiAEAw2eB5nIZ2GWbUyzFpSQHKgCeMIggyprE
KduN3CfyLIqDJICUBiDVEY3UhlAWbg27QqqNMucYdsaeDFBOXqQLvXiF+LLGVS9x
Ul77uDKK4Q2BqMpI8YlORTD8REWyp865XNQhxQB75gDKCkZAi1QNu/m9I3X2JJ4T
VTd/Smz/u2ZaEep6y49PMUGxIqCsrtnu2zZCkNbAQlIj7HhLU6+x4PvTylmffbHz
oywd5Zkg206WneMt5BmkUOHyVyehQ8kT2gGYGs7TNYKF7QmI6XhQ4jqX6FAM9bmS
aj1sNUIkxQuzALLWDgQ7JXafCPOZQ97C5U6SJcbNMPUx2ByauUWAcrIQkDmhjhiZ
cEbfInIivbgoJWey5m6PoxR8mea53S3vonVyg8JZmez59RhvuLgUQr8SZhMhl6co
I0pLzG66Ks0ye9dxlV2hraRjnzwBqv4+3ZSiAtW9suhuJvB83VNE82Ktr3mYPj1V
+oRy0R4EbG8gYaHz62ByTZpwpDNBdLqlB7GCYCd/l80lfJpHPiD4RAWss1AD8GYK
2QefKRazYp7GMLrUJmwNtX7REIwVnhtKf2ChMeUFugnvS1aPjI837lEPJXK8k6K0
EAZOZm8ktnDJieHpJa6WTWsus4TL5H6wq73tD0R+sZ0s44Uhq/2auwYMRDKr7QhB
cH0BO7nhH4hM+NRX4dpFhkS7610m4aSJ07mQsjWOYOW2V8/32dPfGtaSRM343TYB
kGf/Yf1o+YIJgCptidoFaIm/Lfw8aTaWBZwk53g2XKxqvDlYWwwYXoBM+fH+SBbe
BAeHGPemta7jrdGc/9asLrR2KAeinjbtp2WmZ+3bj9MqgWLcq366loX2tBEkZIwB
Hyq9aoBbq7vjZjPUuUwWgDwUSEwUYO4mdvUs0VQlkb30JvLa7jz0CGX3+aRDkbxY
JwxU7x1b7p6FHeQgYmZ7Qhnm2DN/IMM75NEZ81e3oa1vJNqUo99RObl6v370uRgp
m1Ab7aJWXT26QfkQF7CuMa4Q+QnCuDXaAC4UYF2aVxPJ/e3PwJGiuCxNUmMCjULx
ErxzkYjv+7lhO8oF6MZqHSmDRlqqfsC7GBJQHqUxVxMccLm5szQc55GgSxPa2a2n
RTuW8EtS7Rz14eh7s+re7wEHouvlYOL1qaFwJqhjgy1XUTMEdGInJVUxOerxva1Z
3cQMuA5oLc2Hab4f31pfLf7ZqU93yTZ6vr+saRzOZDaVy0E9+P3GIHPO/MVSQ72p
PO5pLkbK81Fm1Zz2PK2tExouqYdivEKB//1CNZ/WSDVP7Fitc+SiBdURN5lPFHIt
ffXNVVJkDOlzKjaM2le2NaS9Zw6o6KlM0CGusJso4jJ5BSYlNDH9o3sG0/t/QXUo
rXAeLcUDEukWJ+pld36P/wFtPXza0ZbRYalgF3r43occIH/Z+EkKZD86GIFTNHon
tgHZkhkyiCOj/DaZ3eP3WdPfThPHH5E3DjI9uVUgkB9kn5tOarzKiY2mVIJMKZS6
vDUpoWfKCZqXyL4ZgMLG0O+7S3KAnRGItJxDpRtA2pi0N+lFT2wsoE+APbm9EYKD
q1uIQtHlay6SkwMM31XssKp6iAt3Uy7ThY1YZtnoaxyBYDpqcI8W0XK3soSnm1WD
hKWFMnVpqAuI4WDlRmPW4BsClgLjEkh3YI9DVLb8EUZXhRelM3lfhh4QYi1zoRyf
rcjSzzQ9+TMzq0hoWgYrbG1zHYaZ7WXHkLqaZb+jB7re3h+KXvzYzluKzYOWhgap
e5ZuphpILAFdcKOAMth1TYBapoLIWeaZ1OMOKHZMnQ6o3EQqqfr/wc0YH7lFdGS7
LmRb4iHLerEfuMxlIMJtLnSg2tAl5eCzI7+FRrfw1RLEDU0ap2RPNYEQ2MTYQ3T3
DXjrqesf8D2e9eEm7EGa6vSxovy3wWk/olAD/WaJjzeOX+1iBV7jMCiIIqvfdUjl
vOA8UuQtZxNlmx9uBeFNkh3VBhyv4QZ7PyCXnC8sDFv2P6coJFd5M+E9k+uhdvdR
5kOgTv9TuowToq1gcxE+AqZIQ5yWnUTgRyicj0+wiCdRckHJ1ICnRU8emXXefiCa
nbuvNOlZ92wxTAcnyZYVtHdBJLydZ6EFGNTCO5epOv5njNbkwb1ZQGeKdS71Xy5I
yHW3Kidnrh25Mo1Gxf4uxEslD9+od78Gw8BB49adVSaiiHRokDPqrsz0FwWcK8zI
ZnfeZe3pPPowQNXv5V6qUTjYtw6YJrQVzf9R2VlWIen4t6663lQEpWzTw3RFcEnk
A012x2KL3WjLxfX1VqYKi5GdR0cRFER6unLQ8W6mUQPBClJy2Sii0SJ3H2YFvSd1
OLfwMiQR+ZyMRr1lWt+zbB5T7+7EuxrvVP13JFx359n/QXp7eGuNgNg80kfA5a+p
5P1R8eOztIK5wZK01gYoXgYYTkhVpkEOHhUU2qMWYWIFxtooPqkT9A6xTODtF/ym
/j+Hwukn7WTBecSOfI3tP0NyenF4xeAy9Je8kkyt+1PW9du5QN1eFazbtNafhOtw
LS9kW/F4COJ/DQ0aN1qYqOo/L9D+uMy8ZMURXTIrYKsJTzmFNHLlsQx51TyT/L4E
RZF3yV6Xf9Q20Y/rM7B6YQHHz916R3s5Sr+vx25vBgkYI9hoPvhFf1fnIhXzXhVd
4SHyL1CGtjcMytms5KFoAuwR1gt9hceZYUxGRssgLhxNUcD+7cLw91TojKxEppkr
EKk0IJQbYzhRkVMBHdXWREF5DhTo13ldwBmX/nmp7b6qj9QOq8l3y4/tNbCACcDM
ZiOz02hywaDOiotMFqzO7dA5RL/FuK0sPp9xa0N/9K31TzXv0jd1V8LVKgNfKJ77
LAyhoAWvKg6qoKtmmJ0gyaZ63J09pTc6ZKubPOhVlIk+uA7Y5bytrAngzbQgc64T
VK/MhmaWZ7gBbyuq0Va/ULG7aCIFamRuAsRh3Mq85OS0ofv/8twunPHbRbuPkoS3
fT0nc4rCaEH0Lp/ZWPhQ7ixS/bU9USN9ctpoXV9buzPbDjxYjy6bMXZcJaWa5QPK
mCEKAoU1+tKAcLsusel2iEGgsN/33KkEzZRD6knY/mdfAP2vXkRHNSg4McD7+VfN
KzCaVhQitzdX+UNz9SJJI1KV+lEyOmc0udXUXrZqyyylF6IHiPd4KWBk8IDAtXNo
osvLNrsARc05JLBtT97lTgAvTfdJvo/f9gjk6ccVFW7ar5I4Qp4sGq6Hc3m8vqUe
BFyiWcDY10/5gcBl10FqPyJNiqUNl6FYKPtiB1P+neFZkfIP68+P77NmI/r3I9mU
bLRURBj3Y5xX1w3AHOCdJnGE1oiv/jS0wDLIXKVL5byZOB8Ra5eYffZbjAWzkRfh
WjpCQ5GmfnV2umN+/j9RqslBm3I+FBiCreeY79kLWm64OCiplvQ3nVjnDkzIIxqB
s20Vi8o15rVZlgYaDLDZ17P722ltxv0r5tKEipx6CS5bYDwjwMe+T7Co8/Ls/KK1
FDgahe+mIUx8j/hqsaMNZa/pNwSjgwkuO/j3LcGjVFxIh/BLDTyN70rGIIkJWE/l
086+t24LC1OA+8neLeNAFdjeKQZiTpelZeqfqamGwdFGG30VbQvm/5hphx24z2aT
AVpHGGzEIMagiqWSNlfupZpxSlg1BYWMF+1TrRF6quOyUksSDeJ2PiLZ7cklnrWV
gXkWZNoiMy52fzfZffUAK8nxC7vyqjZRs6dxmUBYBQAfnOq2SbpnVG973QVEDub7
lGSokdyNS6QtsIVIeriMBqKE1wrS0agytqKh9ojN6q1r0l1RFnnqugksHdSFwl/I
CQGe+tWELhMEn21ox+0eD4RYwikAatyFK4GTD/P4hul6v0RZLJc13sQM8YrsK4UL
E2MfypwkrqgMFn6+u8ZKTlUrML1CwFrwHJ/dBjnyfdPwNboxdtwqvHpUQO3D17TL
hWeZTUnoPL8RwyAM0QGsbMM1BVqIuWdoMIuvBDjwAfIpmvqaxXoCoHt1oAxo4Cvt
9Ovx0uKJnTKFxsImmkwpRPnlMz57d/9GQtMVzJTVRpXE25FtrDD2zmXDi5KJZqsu
2MEM3zVAoEkxZeNBMGKHNbvGoz91GnwWXLrFn94adWLHBduBI/UDPLa5I4RGas1/
LIwHz+576NmPNI+kC42yC9qUu7f/heQ4bDWGu/qXm9OG9VuKK2H4fl7GYgBy4VeR
p4rxChf2ZgCAq/4dRg65VFVJ6azgx7/Y20TGWaEBeb2Qaoele/ui187kX2Q3V+Sj
Dynkb1dkPGNYwmPR/xKzUksfE25O1KZCQfWi7FKR0PDKFE/DbLUtQHdXIacvuoTj
bpMXhTMOXFPnePLmLMhpbH2BrV+WzX4YXwW6tRETGh9qkz8xKUZotCn3Mb4atQvI
2u+DdIaQRK/rIt+qyH/oV/EsE9uth6uFGmW4EBPju3KoTRWEStDTtEJ7bOEoXYxc
ardhbSqHHGX5MNm+T+IWsrDDyU/lkM0MNEr8Y2o1hWaKXdTXp8EjDcvqVXS4eSLs
IKwcAVrslrMaDaM0dUdYQ4LLtL5pLFtz57Psk6aW/DeOiv+ewga22qJruNzDq+EQ
768+QkC0CTGXuw6N+nZpR3y7f+ZmLKG4sKGBl6xr7+VeSDMHNLQYXHmKXeLQH3Vl
b+ZFyjvL8W9hCRYXkZAcahvav42pnrm2jesvQZZo6Kf3b+uiGZ2C0711WtF6rI0g
1VXxkfX7MnwUGdz5/4cVd1Od6FO2mGiyjYzi5pSVyzQixaqb8g5ToRA9ORTvJ+Wz
whhp68YBXtvc/Kwb3IiLcSOyop1vmq9MaNT64U5kwhDQLaaIS+9a6qmnE6oN52sE
or9d1ymNrEcUX4zhlawEFwfJ9ip0rO4aQSA2xFclYzzQG4rjYGc9Gcq7nhwWKI0t
9q8b8mPAwvE/rKsIisjFT8YN3yEgqsBYsuYjn0y6G5EYgPUxMsr9UlyZzwPU3Imv
dI599enqJYmwtQuPfemlWU2Kx6lyGINOa1xprnP993Q2UsT1yQC9L9rtpruDl8vS
Yy/YVcJ6V/dPT9QwxGjqUjbPVsK5FrfN8nwWQKo1jfB2OZPRavni2odzycmlmJIg
hGXjL6qBClARJZFG2QYayz9ir1I2ORYhTQbEOxRmhxhRrEyRr5G89qZsuS2cNSEo
nV+m87X0+UhWUS+/RXhnzgO/C7GhbpLWQtc6Yk2zMerTcm8wmhZRaYkoyof0YBtM
QkNyNbTRy+xhC6uKJckUiS9kKst7ga13QDRszjsY2wVKM7P9Gwbx8QqRF1P9QJ8P
GgfqSjV6E2Dvqf0Yj1IHYZEiM7yfy8MoVap71YDXdNRfmw4KyIVhz32Mg6W4nZJP
cL6CxOS3ohudL9vbONyrXZyckeXKGQ7wdEzuRFJRx5D3UHLc5GvWaXYX6EhlIqvk
nG2zQ/FtsNS4xwUI9Cy+bvo7ucDwak/iJQOr4RPzKwOQ9pYaYyVCfNITs5D0ESoI
z9DcaYQguqcQTU4KlbYkCNqX45eF/l7cCMeRe6y26KAQxDYVr30FYpirsZqfkSaX
Ig7fbd/e4zyvf6eNnaGpX4pBoLs9v4QAP+Y1gHUS6fxIzqX6Y3jrl4HhmkFkaUUJ
cNJzf+lqsQN0AfjniGcQOSfhIcaqQZhvoiJUNerxrZQ0ySddU1ORBe5jEWF75Otm
SghREZheeoNLKCqA0tnEHQ2hjUQJi3PMD7auP7rACmjcK/NMXhyDugm+5sDLAftH
Uda4xWaV89ywZtYsJBj15sXkyeZ/lNJnxhxRBFXfHxVc+bKzFmwxDQQ/9JpHLen8
RuaujtXhYCvMG5ABop+bMV/HTUHHoWH0qXxTaO1g5cMpNekPXBANDIjh340gqvc6
eC7J1fHFtyXNp7iUY7J7RwUjnMlj3hEb6IQnDGI8k9uSWmf5exhZYlh7yKT3gT8Q
/W+0Wl909Cgjd4Ejqiq1nhlj8fGZIp/uWYk0pypOw87D0obI4OOI6p1EliEk7OOZ
gVfSHmeqk7scRpT4WbEoaQE3mwNGW/k8a9VqDTzhrsciZWlUna1QZW3uefGziNpT
LLZXdIThoHIy8Zq0PDRO/YgHHQ1v5OkN8iR1dz37gIU3wN7m5cXeXLru+uKPQc9z
FOeOFZvaDYi+5uCqQuHnN3+CsqPgmaikHRmXqt+GqXzXdbfmC3no2Src6x0UpaqB
MzWlM5CHQIitcEnN5MYD7/b9r3V5vRlm9c4PzUbVklCIYPImAaMZV0N51cLMr9e2
2reKbmf82QwqpJLkFEPMnr2F+AdVoayCOlMf4NXJS77PzLC+WSSXkCy8lr0vEHCt
Te64oiM3HcPWWYcXDjtQeqdMplnP9v304OLmuEbkdx8pK7NXXeERKhdrNdVwnZlx
/29N6HeyyOABQQFuFkgQO35Razo0g0SiWP9yHbakltB1mvLh8hUhxCO23c4sr98d
I/auhJ0TcaUv3IPhvB1GgCWWaKEm8udIFAYzWng6Dn65t6RB6CztAVLBveWqDrDX
q3hJIfnn8bW2oE99l0utJYUiTOPEpF2fkWmt4p4ph99Qet98ljBqxn++fe8Wfnhj
QU9w5FERVGbBQ35PKebapa3ME07EFMLZ+IjTejhZBeAfFHuRAk7/l8B585agsnpb
P7mF664gxBBpg88+EXXhLxyYB8vtiX1zrDdSK1QcwBPKCTqRivfKzW60OzR05J63
ej2bT3mg7OOzChitJc0sFFlus3EKVWyyZs4vfgs1suQke7+F4cUYr7sdTqoKbKET
YS1CZOwebv9XvWCG4NM+h+oNJPZQSBoSuW0/ajJXv0yA1Pox9HGKIXHLZhHfjK+m
sK9vJ1Ub0cqzGoSjWzoZnD0qyKv0ZzASDVlDF0teieT4MIiqvzcCVBUDkruN+Zqd
Rk6R8bA4Xv26e93fwiTLsi3jU0BX6TFUwmJ0opu+yx+Hz5m5PYkKZx1b4y/k7N5o
oe4xYCrRgWXVA2O07ZwILRL0CVLAmIVSsIEgPdlJqlPh0XcwVDd69LIZSaVZ3RTE
uVwmibhaZURwi2qXAUupopaH7au5umgNF5sgogq6veZrCW9VSnLRgOVkLI8NpMCj
FrJ8fBxHQhnx/Gh8o0wRLviANKPYhAUWwRt7wOiypRcCyItPTpYDw0iBhD6fdcgA
xYfgBuNHzQmI+qFt9sRGSRxfWMaGVVj46nM8tdd7F8PmtxPnI+29P0N3aha17D5P
z9eO1v/JYv49CZQRG4ezKwF8NOmGL9x0B/r/iPkCCgYdUy+AhkKvumj1UxcF09aZ
mmkiIn1584R7FzUGaHMpkmVhCoIjKCqcDn35oV1tzWkpeuRr+vmLkbKjc2gvlgR4
S4UfGay54JhKz6nwAI8C4G/xJ/6GCjaTx/xKVCTf/SGqEzwYXv1vAVjOLAs57W8G
fa/wf4l9dLCljLMOnDOBVGmLv6xbOGOkGU0Iu5gYjIlwbFrYaLqz14uQEJCvWmIg
niptesAJYNhRp5yLMdkuvd2qoxirdC4v4alThY3c2aczdRSPsWov2pm1+9/QWyxc
Gz7D/HRlysDgg6bAvzAdpzH3JX2oYvQlwQJNZIfSrdeBfBWf2hQyTTcS8/oZ72za
m3rMFWsNbqEfzaauHLrjZWyLydW8jjDIPRbLVcLmWMMM5NBxeWKlFKbQmU9pZ1vK
BhO8p+Wj9w0KYQNJNUA2tUib+pP01Cey1bAOQzDRizaoVHrrmdEBYCCzcHXZVnIj
RZiVPDwf8HLize3Rm3pn36hpzSzWq0F0xT0GeJxzoWYp2B+2FQ9/WHrvQQxFprgZ
CjxVUyaZ1OIZ9M4yylfPepJoRWwwcEa95RfQEiQrwOzCHcaGNEdGWDlmxQf8UvKu
LNeTFpyHvJYgy2w2WMDEY6gIcIvfBPUDv8nJCUOi4OHUsxgdcGrjM9w00SpNoUx8
ZExmSuJs+I0O1fPHap0oynRJpY/Rka0B6UcBDM5Mrlc3AweCdoMFnP/oDUuKCz24
b5izYPxKRsk1gTGC4oybOZWi+AtWK+xecp1jt6xo3svqP4BgdheSAx7Q5sx9H5sC
k6gJJTe8fzFSQ7uhjC9IWsuLd3iaTPty+8ZZe9iEVOHqk/grlMDRGy4o3p3/11Ag
Fcr+APDFXaqzhr7tx8LtNZnMa28uyOWVjhneHlKG9d5kZFQJX9e8aMwVF4nsXOu7
f4KmuxsMt/dNPJDZ7zT8PYLdWDNb3G5AzSzhP3onQ7s4Ex/qBwEgviG9kTkiEia7
fwAhi1X8lDbrY/Yi4brpJPt+BWW/2dI/tdBAdduf9WMqrLAfYTsRNvsAj+UBzJy1
c4N7fln2OWA1C6MaXhwHViQ2rBiN9NECFOJOVabcv+lTeNeSzmPObNaU0TZh9fKW
iDJDTL6pCV9f1HhKdyazkkRoCMEBt9SVbnMMvfPfLWpy1fsDehHxP72bxmxGStWg
BlNXXsNROEAnbwMKgYPUfLcMPNhYxIagNnscX1qQS2W7xUVcA3QXAH6tHHGCYPVJ
0J8FtL6aZfTLbh9oXiClc98zg4EtGUct8gpCcJvzWxy5G01uvDGHXHGvtHDqtJND
QH6Hov0v3LdeRNOuQu9kbkQO2LWAcdQuZhWo76S/FaOwAE4DaCkF33/byuTu3jaS
i6bPrAdRbWWfUq1UP4X3WcSJO4vlpic/x95aNGXRHVfL0ibnI+5R4LA1tvgMXxB+
hnhBaOpu4c8b3m/OCwvaotJwC9ICGgi/VJUjCBYab9SdUpCWc6YskntyCIz2P4yx
M8mngqW7SBPpqW0LCNvGTl3Kf3+5C9SNwBlG2XfH5Ym0JD/EfwAp5Aq7RhDuJATL
x7RFZa6aDOcHfuL7E8P5lNWxIO1i0onplro68kKWlDTSDf20Mbaj+bisyPIDYy1D
0664VqCn5IfDuJI5ZcRH9v9fMDFhTOWIaksBaz7B4wGTgQmR+boIY4ti7Vc2dyXH
j1qJhGJpn+DrIeVJP67WOll/4f2Ib6Youxp8xeDA2VW+GLvFyOZtPpj0ejj2H3cP
LrrArc1ghON9fzpZZwEt6VaZ/HODBjH/QwEUpmYel7NQT9nCdMKa+iEptyYH29s2
ixa5d8/KtrAYIPWevuKcPKJt8kbfTxVBh4ohYVSNzP0EtTR9mGH13AbfuJuGLq7t
UbdCeHmRkrBOvjm1xiNAKGeJwOxQ6/CbLVBfJz967emDqlLmHBzTRbJnOexmh7kK
x1TFzWW4KlAtXzdUvUUwU2JlYWRLpmo/n+UEQBprxzM3BT73xmbgea6qsUaLEAas
wYXW+8oRJOD9FsvZEsArsFneqmu2RyE4Tkn291182ojFYymJkjx7PQsTjZEdfSTC
iKHfJiPPko06jZo4FUtiV+d3+RbJZn/Nqu6OvzFzitJCjsSpgw4foW/aagw10pEn
j8daDj2FFiixj2iaWk361tFySl1+KjBOM4KI0CgTbqluELFieOO/ECBfpInMev35
mCHJN4Pc+xlFhpaAG0IlfpOGkAbLQsRuWpwIuxc10TuD327lZscV4xTB+oyB7+d4
BWdNn20YYBWXoBS6dkyCAhMzSZqW4onc806QcBTSwFrDEWHkjn0gRC4JFDzxEnJO
4i9ysPackvbYJd9fORLDXn2BqD0wlxmo8B/lIBll5AQEvS7Hvm7OtWy6oatuVuFG
TO0KEZQ0zQxGqpuPqH2OBDRss/e4WHl10hWTm0JY46bsHMLy/rtZkru59/nRIXZN
aBkLH8PVGLtn5AbCymSglQw75BGjo9G1aQLTmihnevoNp78qZRMZ2oeAW4HGreQi
tEDoNLDCsaitjj7vRcX1lK+FOVh9V5T576XIDnGvWQMDLO7I4koEZ40pta5b7nTl
ZtZnhwj4YGuXYTOx5C3zSdN+AfE9fFXseuDx0NyKwsDF/vMzn0fzfuZ3CFeK8X3h
7VOimHXuCykbG75MX2i49mB1w4yQNRY/uQwrC9juWh70Zz16D5gRB2Mi8WrvL6nP
ldhtkfkdWiTju3nGp7/8dMW1KSYXMrGXB24O/jHcwHwUdze+jdcXN6AyjIUrzTUu
ssipWOPzMlVIA1qv+yyJd/0hnqOg2eJ6t6JlUhIbdPI8DXW919txxljKu4LoxcIB
m3wi3vpB3skSK4+/2xZibcWK4SjS44UIZY/A2kA3aM2SiAme9wZ+BFLN2RM0BCK0
NMh8dCq3O0g803Yr7VGw8DcttndQg5E2LxbC9aYyO88z52RayIUp/uG5VGL9zCG+
tya+MR8oTMnu3ZReQXlhA77Wm/HFj6HkhN5+/6FDgExEcQK8a5pTz+xVeKE1ikxS
vrT096qGn44ctL5Nhh1+bGt3llBI5WAx80tCTIm0kYteYiUkQ8F8jHrws+/aDi6P
AfQsPQeRySqbUl/26qKQBA34rd05dfFCISubbkWyfiVs+26TqRSxDJDcU63gxfQZ
BVCCikflfNjPDNOCnQxf71lmYR/4Zj0ezLQTN/9g9zbvFiOzz6V0KUTfYUQGh5lC
3/bhYI1cbzkZg6Ey59NuXRPLVPE/v8Arbvn8o5u5jDYqR6pdh/6n27RCjJjMwJWl
/QuNP2wupib9BoU9WSU096vrvK109EPpBJVEOSBe6FiDcMGqGcAIW+hdqwWbzn9r
So3VPtdA2LLEmCKp8W3bOhQ2Elk3fLUZ/8A1SRBsGu1fgeri7+5Q6aOct8pns9X/
gkZhUVhQpyU9cSs4pH4rIfip88N0G9pZEecgNgwDs9L8ZnG01K0YuE8qFxICsWN1
sJjrqMZCXNwxazFlyyDcHeLErFddaP5vl4XmAekwmvRJsWKxoQz3epxCN8Tz4ir9
GGKqvTLrJix9vcrxKe5H7y5L5QGVRMw9gMlfeQcAQL4PVX3BrczrezZoWfOvFWD1
tPrK0+RkqVTeteT37eCc4G/EhHb/839TQJCoeGgst6FcG5941JnbCz8S+BAOJAoM
LXQ5kjX3UOZl0wQs8Nyd7GCBT1Fu05hV0QWYUUC9KYPmo42meVo4ZfFSj2joA6TJ
75ERV15YpvoNKqb5BKQLCJ1ePezVUuq3NeM1yeFYMULeSAyQTl5wb/OpWVyRfW03
AYZSWd1/REFMCo+v8C8R7SvERknSjMCbm073ztCoJ7Gyb/McYEo6JjrMAJbV5+3M
ddOLFeKQ4PfN2zLncoLR9QOi0q4PtEYZaFTcgxjiwN5GqSBGeQXFQ+kADhjADgQ/
vZvc/NER4TMDPFXEde0L8s4jHJkIEGHlEiflRarlfv0yEbDaHJtYO4sqxSBpwMaO
oXddvnL7n5d5ZR4HNIr8lwkzaCfhf/4Fc+nFhl7GCYAz7odHzYxlz7Wd0cF9v/i/
/SdezuCO9TVtIFgk7fCe213116zhKyH9kSOalpPKsq2udrF+YzvT9a31EmGmA7DT
EY15sr6yDT/vZg0sK61qlvoCn7GE59mnUOW2Ficoj8YGSozuwcxNEkTsqMHcVgK0
7ivY5yod1cJstWVAwfSCjk2buafliVv0CnM1HqNwgJPxiHeGjlo4NpOKxQfMQdcm
g94ym0GF7M29ga/bs0fLs4cT3/x/l9oYTRZrq1y/t0K4pizgqA0jdMdAcuSsnlsK
4bXHfvrb9SCpx4MApADDZiyu7jBFNZ87o5b0KHw493bwka1lCTytfZaHzCjvBm92
3YdALLXSbxfCzcUNQu4a3QRUcP49j+Fj+g83ihcMxS6FDg8NnaYE2Z6l8EQu7j4P
1YHE4Nv8DRnWYI+RuUxlB5V3fx/xNnSw21sj+nQnrp7GtWc/4gggdIb9tLmEc+Q0
yJCHS4NvKV5XpKJsmyOUfx3VKHc/apjKqYaXVaa1nKv/ymXnslD99+8cs2HRj7OE
rG9wWTYqWx1axdOLIWytdYn3xFO10urMvhzcBKq4LuLy4hZiWIwbqzsMXmCRRtez
u75guiuDMFE8LHC/yeua0BGnv7fQGwigwXP7a+TVe0FPZnNq+j/avJZMt616FmAy
beEueqwlliQ5THX/hhbzvs8N9XXExIB8DMjqThqO2EKEDybSCzTpj4jw4lY/HpGs
UKGZjZtxifAO/0fJvDBzzkb4YPAuu3BEEhGk70Ssc/jiAIdKdFo/7FLYxfCKrDuG
U3Dk9bC2irF86NtLCrnvOXu76sZThmavJdE9VLbQtfGk0gmteB2FlU01q+kCKEAw
DwBK+3ST8z51LtMqxXqS2VchtExMPtqDMFSreUVI+AqTeIjzihMYkb1pwoNHtVO3
f35StjSFN7WLctGDx/FMua9w++kfCHz8ButP0PukL5MRl9oQ59D2KDOHoLgjy5wk
c+ZgJM9VRqLaSBIDywW50TNQOtQyokuPmtKXh1VsTCufhLKd3cyGC7bIfyAYB0Sp
6BH6Yy3SUiu+6lGn6Vn3xL+L23JHVdOt3oL9FVCGKmDrE4et72XM+pITrD/Y382X
hh/UXAMnVr9wMS0qYkk6evyECJ8NpGtiwbLSusrjZTT8TDtJiptp6tMz2Hx3pACL
0eoFUNgCibST7lq5VYREzQJCanZErZjnnEJEQ3uBZQKI9GnK/n0p9fu/+ceOSXQw
uWA6zzT/4S6HsZn9RLGBAuGKRr869fA9C3/RLhjpfWrG1aMc9UwtGwYsKrwVmo5H
Zs1Us3HPO3uO+5YHO31wGhnddnj2XdNBh+c9rcICnSagrD2wh4cyGZeDEyXLo4mC
yL5KgRfsjRkgKwlUQc3N78XclVuo+LdKEXZ5h0lJ+tYyp/nVosO62NGet5B1t6sH
5vXI/CRUdSoltVt88N60xe6Uzn/TKrEprDAAg5NFGx5CcnY09ON+rc2zU3kFaYSr
kO5OSwuIFV0ZyYGfC2fbnWJ6V2ZXsFnRH2sKVMqY7VqfwO2hrMZ/k/I9wxfj9MaB
VHGG1VDbb4sylCrUknN4QgkKNnGn7y95Z8gjXI+aola9SJ+qpgaS7RWscV+9sC4l
WdF+IgXsCI2uXTD7ovld1Xoy4oeAUTdPPKWTxWQB+1ofgMLSSDtZoYKZd2QQy+ob
AxrAiBqDQl85i7QwbwN5i5VW/fncZGGhZQf1g2Dz0aPG93jyME2RsQSsXYhK+7PX
ps3YuEI+QcvtbrODnq4mob94UN/gayNHNsPZldgPKbPWjgxpBOLbEzCVCjpyNuKg
cNa4Fb7vVwct0S2kfHbV5avucTjcvCZMGow9v8heb4tua4K5v6pvfo60NTcz02Tv
1lMuoiQc/JR8ag3+9vHsMA8bfw3rT6k1LVQPr7coMXACsqFm4Zu04aeWn58SuLNp
J+ZobeJUuxeBhV4EG7DWUn3GK+ViDocnehBDlCkM/Tvv8GXM35q44z/vbw0jjcYw
HnczFJVxqvEdAeItlLcjR5TPtfHFI+l1tiKkZsoRUcVTecMZS2efFpRwVk3Rf3fh
d2zvYe6dbOD0eO1KyBTvpFs8EtcoYUrQVHPJM33UJgmSj+jWZSA1NHEYQBkJpNOl
fY5LeNh8mV4s7fCEirgp7HwPN9F1x3T8oj7mYkirWe6762wg2BPUSGypmhC9PXdJ
iex5wu08pMmUVkR5cOPPqyDs+K5UE6Uij/X7HS+8rJqG13dxk/KlZ0vDxUfVR1pt
pV/jzVROqDyaB0N2PdVWxJ3zewNkEF2Mvx1apwCiyK6jGc9MKHXMrsSAXiT3qkrd
oofemuiuuqZW5ZZJSPytSjXocvQh+hP3mCM+vLe7HlcTDfwR0G/WKPn+sQkwRvV0
7ox41ZaEgXcOZ5dZmxYFH5SK5jCtKjQS/zTG8Yyix+ouXqTN1A9K8Uora4DfjaAY
7+NzWgC4FPk2XoLirkfDrXnVlU2Q3dTIcLfFfpI/LFmvtsQyiovjxbIYFHbK9SQn
QA34VI/0Qib2t3JYRECagPL4Wb0Sog5/1VDswVbsAvKikNI88yReUBEu2zcCFrx/
oWAKYuHnaVrC+s4T80MwTgUa3c0uqX4qlC+CJhz0AWa8OdklFHLPPeJoihkbbpGL
LKnkNtV9AJO5uV/+I8ffuTfDs3tg5njtBpvgSHFOYBG0xvJGpTICPjhvHZegEZBX
07dZ8pDoKHcVy0IdwYIRH56cYLMYRckpap/PzvG8vHvt4uZRzPBPldDAG3PBcBce
AOpmsTDEBotwRqdGyetkiSAjLjVX8y8q+ybUyG8hcjGcZ7BRQhuDA+kZfo+l9507
4ErqsPV4XQgyl3Ob8R0ThvN4pmG1hbn4VLIH1yfBeWcseXmJrnPO5PdrtB0DS/P7
U3f3+UzQ+1kcv7hUGbb5yqKwvPNYhv4BW/y2MZCIYT4JSanT4t9Gk4nhgVd/QHTN
kVneMaEPgdmieYu71rYiXyCwGWL54Tu/ta48yoUrx/z/c6Y7q/sjpwo5WtUyoVdD
zwOuDYVM+4LVCBATTYpP7Zs5AJW4zfm88p9X9DukWh9i7aceiBNApwOcmt7HTXhi
HUhFKOMYbyQPNVz02h9eQ7LmDHcqSolkdTinzf0/zXU6rQKnOd7F+xItD6T/U/1V
p6xKliATPcxKy9MV7YyrDt2k0BihSmydyKytX7HW/Nw92+YF38EW4spkozv6UyHH
DVsX/vufaAw9MPiBXWhKDVl79lvNBAUr88FuXVbjYnW3hMbMpFb5kddf73eW1NFr
o+XQcf1ynabhHlnUMAbBzwnV2jRgWQPJfR9KxewLEHmunutucHGgH+WPK5skRgmU
6IwyfgPoizkl/vOs3ieGGMvjWXsStMeVWkF9Dn400bXITtOa/MJRheTLgfLTyNNu
XWKTCg3FDchUQGnw/Bl1GmrSiZWfM7agM7mHTKvLLyp6IdKQbQnZS8LOEYPWjTgY
tqu3bLpOCD+IhQyNb5sopqOJXYTJkxwsMJXN3W5RsEnxEoiLVkix+pajRRi6kOoq
rfbDPbO0qudFwh0W7fkFOi7r0ny798YAAJHcBbhaNNJkHWDg7X4vcCJvd5FxPUD6
wHzCHTNNCqlgfPZUO0fQFykCZ4nQ8U1O40KM32sMh5uYhOv1/j4dPKC77aG+9Mlh
t9Z94cFoJ1pFV9F7Co1pTXFGdBCJkmNVE1nWXjQPs5Kpl2TpQPVajmAQVT4ttvul
DwhuHQ5fMgDSlfg17r/8kveMf6wkobw7mQ/e+nSqp1dO8gWrJG73Ktc/dilTAfiJ
DUfHfuu6JS8Y0067RLGKSK4Hnds4BFQs/7oHpB2MUSZKW3fXfrxgjcgfm9SyVRRL
19XobRMKtqTrqiIlCvJuCVMGHMfqIkw9faoqv8fdK/z5b32HpkQMpaQAws0wpwVR
9wTVA0iWjMMMfEX7LpyNET8iDnMD6HQtQXqmIsoiTb95mjSGXB0H4hmhqrs99L9i
NMAhCLkU1PXGs+9Tqv88eRC1fABFycmGqa3ld67icvCCpvLYq2BnMRlsQnegmxRh
g0BpA/JsDDlPC/GTQkSqLBgu9hXH3YwCvlNBuTsLDutHzox64XU2Ap5fWit66nsh
8Udx1rNWAAJAIzJABdE8ZWTyYYq6jYi/0w3p9hXnsv/xmFgrZbmZIK0oFNsmRZ1t
8lWcVGv4aWc3w51bvE5b2TS4o1DpSEHuZuARDyx78M2Nll8Vj3CqTeqRfK3xBrcG
kXgfXbIkPd0pNtT9LKXVPkaZZqdXRSNfYK36Ucoww815MkFSEhfLqTBDCVs9+ZQy
H6O81N+79mTByYTnAzw75wf/S3vT/JtUKY2se4TrcG8RJJfBAKeP+WzjsyvOUvVb
opsKI6Loe3ZMBr2RU6maFcDcSy5edHSuIVgrsoHz/tWdFVwdqOsZgz4WP4VxGSmv
iGz5BQSJ+jASKBvtrKAq+UzBw9o1bWUe2csaFRux2R/TTBrTElBazjXx0FoJCZCM
NcOgRC1aEhBqvkLyyE9svpdFoYXPnOtAmLipXkKyY4n+tHI2LQOhn1BzEK78/v9i
s0y5sLUZmsrHfw/wXV3ZPgcx/IHLVxmHlhhmbZpVPaj33WLXoVcGsz6kpDblvE3p
c7RQjkYQA6iynnW/p8gc66itxoGkcQncaZp/+rzkazXprhG6nUnRQXCuZa9yCyU7
wuPaYzstFjIFD1nqmQor95bR0WtMkkRkF6gu/7e+mn9PIXkCJMBEpTo5pB78aJtq
QZ7728HvCti9pZpZ/FrN0M3R4G8zkkr4E05gt7w9v58bBsoOasRi9SU6ZeAPxS73
TihllnXrR/0hf8awkUaWzsUJuNOYnfwNQ27iVSKODc+kLkQCAiffRQHoqqimSdHU
MXdkvlZoxhPe3+g6QQNeHtyjn4nvCK0xKR2xPAGoZaH5JeViM2XyXC47ET1ExZ/a
+e8vN/q4wMMyCHZIFapPInfUW/4GQo8azvGR/bwbQ6hVB2VBHYZW1aWMD7YpQugr
4yPM5tSZpbfMrBr6ymYbG8jfQpROfGBaxv0VmknuPkx//cneWRxV4E7If6WfUJoK
KrjUyfaG7z1JNlra7Pd/r+28Hw4mLi56/hyZ7WHqYKr7UPYQF/T2bFsGkk6nn9fP
Aj/NYVxZtbMtOGnmq9FVPQ60LbDztQdjemVPZ2NpzWDmHSw4owmf/AVuXyN37xIs
Lb/NQdVUn2ImsUy1tlDI4AIYIfhfZCeAZREVkmyJIbEY7ueUISh+KACBhFnB19yV
zvEnIfcSA/EP3wea4VabkjNyLwveo67Uhn1yzmt7ip0C7rEYiVSu3kov6j+pLVDx
2UgRSv3WMq4FcXNsNwHkgLpyG/AiKl8eBcQOdzLFXT5cTEcfMfhlcz83q98jSWSN
0p5YYEVUGTBJbmDFCCHZphbnS0YFE2UdWRE+bRSL9h9DVqraN6vymF07OM387dO0
4SmZxrSgY1OA7XIItJufL8J2Fpo7pQxIquYa0N9oMIoBzFic5sJXWRVxXQ3+HKb4
38Ev+iscYyZmK8n2Ef05nUa9qMGRhTuSFtCze2iJZ6YAM/zDfmMX9gopYErZ9mCP
n7PmBaQrxE6Rn7aGZIsvdm8sWUtGYy2v/rqpGVdA95se6lvRnlf4A2lMcjHo6Q67
tT5yy5yBaewnOp8oJzFndHzeczIAv4fxBkovb90N2zxbOrA9ApTtCr38ovPLYb4E
8WraCmCV3kbECRfoBvV9GZLCPXxZbVWbICg0AZwuEtGQc/ILeAu8H/qJ7ITk6iSl
Vh6uS9FCVYQIQ+EE5dyAp8wlCHImfen8R97rr0sVz0PqQMk56Z+Vb6NWgkPVL0TU
hN7+ygRvCu5/DUVfHjmQBmiUVytA8xXGWLnbwau2EInytTo7Llz+8Gp7RzcC93eX
dS809zxtBA2UgkoUGJ/YmIbCFN3h7OhG7dghHnMhWrGqhQW/VwmhFbkdcyOrM+wV
yfMnMnNsuw2gwREqcZK4PUG3wWuvNYTIwsXOLgjk+b2/PX2KlEFeGj6Q+GGRIRB8
TTg6pqn53lN6Gn56bk8W1hEByvP6PSDb5mokE1ZospjeVXzew6gZKDO3f/3wDvaA
4VW+5t2pDepPc2H6bMRuab7V6B7/3GrQqNHeJK2Q5asM7fGiV33Ld1r/Sd9gkTdb
5LCS71URWe6M61pk9k7o4r8gMPMPXcM3Y2a7sZWBns5VKhnr49n4ek5XdHhY0Iy9
Vt4iFHVwIaWgRZTisifcwS+K7NldW8JoOTZE/t6bVJcstOnx8DL1brpLKKG6SEM2
hLagGuncPhZmxWmZrpadD4L72hvfPkmmKfN6K5HZc4E4npFnyR7Sxnrnjy4ZzZXd
QstLSo02EV24jI+l8U+6nglBLY8l77Nd6eT8jtjrkeI4xJBss4epmWIPhFayQU01
86FLOO255j2z8hIrkrRCBhubF5G43lINiLknx2gqEf9EEqU51ldlT7T0/3I4N6P3
L2HwkWjwi702UgTEsVuqz4IpiIkr691bhB6YMri1UOQmaKvNfAbVSmyWBY599wv6
P8b16ImzK3tYa8Sh0U67fINY71Rb0J2+/dcS6DPYHDuL5TV+wuqPsX9le4ysurHk
PQMNJ0gBl9MUuGF/Xm27gmkAAfaR/7C9QQE1gv5I7BzBzTYlbnRKVqwuKD9dsck0
FHF8J/zwur0Ytdn5iWieoqeVfZ8LdudjW7oWl6V0Tv1MFF+vHS/N7Mhar+dpEJ5P
T+u4PmENBjmaih6CgpP3IVdZXUOg4GzhTPQea4b7iiUzYBx6wfKDqNfnLFUtnkDU
cEQ/2Q32E1+ZQ68HgtBf3RozTZG+j5dK7rudrkLGMPi3kGUVI11A6gKCuUrvSmAJ
IKLjlJfLzsH0yzkU+REgOiEAQy5FM7vuggUJMeQ9LUsCruoQZUy97+lQurWq5IIb
IP8gp+1UUtyERnwgtEZwJwTud7PHQT4xLSoCMVOuFr5EiyeXzHpot7ZdxIoN7Svw
NFtzTfNKEGNSEdy/DQidCpXTH/sudFXneBK85ZS8J5kEtdAyg21xOlgvrrPtHcis
ofXJxJAjZN4TwClE5ODt9A9UfszLl+zArlowwlU17iCmA89pRBfpPXhHUPhtgSNu
ZZXsKZqkssGPkCQtg0KgpqKJi3UIa4vs76fDJFJnPljlw/oLCZWZmYkkEddNJz6F
3fY6ZZgIFX4Xa8Zvjck0LBfQHD4Dq3gI0QLEDqGE4vZcK+Pz5nhdIaYQF5KTIYon
DfPmgPuEgHsWIBhSuWGAug2GjIGKBXaSYna54kxPvGeoCLQItY60bYP4Ssolo65C
u+6DV9NQBkSv6/NmhrptYNdcQGl0mGDo05PLqIEFp8H3n5HKgJkpyXPSxXVFLTe/
tqXPQ83+eFSrerAlrfKZSNnwAPafH0fxLDJNC+Rh+Zlv/yq3oqUZR1ku7xW0zHrd
t4dippdSZmzJ2eRZNEFt/Vugsj6nsLOqzsyxrn7j+hVocIIDcpbmUx7heOt1P6/p
sBmZv25Ol0MMPagYsL5fTuiQqii4rWY2Zwk0FwQ6fegK+c9H/RRVNhH0hXTNGVTW
lIErRbPci4J18qtu2c+9JeE8BmFYEhgV6PfcyeOtnkCwFG3cywSRKDsN3Eaxqh38
CXkRx78tIAuYE/AUo0N7+jlC4Cg+7PPej/m+LTq2uR555gIC10qBn5IoQUICJF65
HQ/PSnHcO8l2lru4EC/Ov522kVmub6JWpcRpEtu17bWyvX4uRr5SPMD7hUj/2MIc
DKQBY345CUokGqd1loKf0M8ygHZMMQ0hMWWePEkLe2Qm2PdrwNdt+M/oEhPqDuro
5MdqPcJBVl9oaky1FFcM1QlTuCoPFbwlTQFRzU0WHIp9LOa5o42NLdwBYU4YjNav
q06JR93LfiWDur+TPk7TfUNIt8cF0sHeAEwN4U1XQ5jEMYBzm9KZUrK5w+66I6li
En1rhZkgaZG4/Dah1FAwH62VaYA2Pn4WD+lDCDg4/uBD1oXEW8MbPSBP4koQFw56
51O5xSKTexbxe9W/ctP9DuH5ZVoVpsmtiClgbOOXPHMa2kFIak+OjErpS+xQxJm4
eS9N3gCrqTAg+zgwoBaZXaqmv8C9lYfMdzRzls9q4ll5L7TNNfzFBeuM7DzsqBbi
M3cow03Ro7hY4ESO+0hqUE0uk9knNtsuhGo0fNzAes1IzqQ64h5tOBWO4sn7zbxT
jiR8jMBggZbyYWQWkJXHiDZxLrhBaElQ2NMU8I5kq73w7Xk573p81CXnWg1dn6OR
He3FSV3EYkZNgxDAP7D/C8mqbgdkScZIJ1YzPtehyBS+BzW/dCWvS9niJp3LJqfH
nuFwRLb5HNtwNlMfMWNpyZaO+vetIPXCUofMDwLogaIsQpDL6Ct7BeZa2ks9+N8Z
WWrS6KSx1qg+8ZtRfur7ZWWvj05MkErGkmUUCcxRupQGpdeEWuxid0tyc379F23m
xJp2JM/zI545FzsXlMfYkUHym9j5728+R24Ug2CmC3u+Sem8TzK9r/ZN7hD7gkw9
HJs0LuoMu7zgIvRDQJlMIY2KJ90aMpqm16qSG7ohVZkW7sNZCGagdYH3QTTaW/ws
q58JGTbr5g46GaNN4iMm+1WN2LNPVea1zxdiRoIfe0L/9pTH7C6tz5+1HZy6Vnkv
OGFDTf2jIP8u2Oj6xIvxUEMr/RA/Ce8c5bMwcK7tTPmavOXX6d0zKESQS2G7gzeF
bz+kjfJIdGgX/oPYzR9Y+XMrMBEflDDn977RYTuo7+FK4LA8R0muRloAuacwII5n
44LiQfy/G/GIC8SFm2lYSwjbvdLhYtKQ5uVWreSoJ5i4onLfpDoecpmEhrf/vFHK
qwtxM/hPoMBLaJYvO6a1OQvdtcRYz/WJvyRMLuMY9Aytbao8Pxd6JNUALCPrYoku
z4EXlqZCBFoervExASduRselEECMcaIRKQjdMq25KhMbiilUnsqT8LphZQooiOzg
SiRryN7FmajCHpGvUyM5yqYfGNhjU2TWI9LdHBampFHh2QzU8yi07NSZM/LktpTm
T0Q7x/a/lm14imO6DIL5Tgrr9lW7kZIeN1Bwyc6yW3zz9ilEDeZNE2l59QT/N5Fr
Ycq/sOJLS7aiUnkHsM1N6GptjFHh+W+fZB2JHkyG0EBaS2euwDSm1+3bYLefqJ+f
GfInq2MjSvyUOBdqAmBTJYKrESTfc5yCJSTL6cuUMqEfpMNJRphCKhO4k1obXn6F
NDT+4GGVcWOpkwsU/dL8Vnj8QfLzHSCnOnBM8mo50EAv2vSIjcb0oEi8zBhYnvGE
/7Ht2U7I32u+wOPSqKC57AZ7PTifoOP0S8V8EXFLlUva474z2OrG08s2lZp2vzIL
p8UDG4BtSHWkk97bFtHqBCEfBLXwCS01NO/Iau3uoD1/88QxL6z7XTa1s3pyTAGZ
SpeOEfYACLo0G9CdXl3SdUasrsM24ymCfUapUUXcJlYj0PKc7FPq/shQONEg2JYK
ehVEDIY0sQm3KjcUB8vpayvxGWxosyfayJ9do9i3aVh0O/YOf8uw0KqyjR3hnnwd
QJBzBLDPyEdlpXlH2vj2ga58i3c+Bmh+lBBnpjJrvb0QPoMZRHDv1Ugmbs2MELk8
R9Fk4RMKJ+p80e/2ytHYrEfM/ZUipXtDuM+i/n5zvIDz2uqFdaCVEsZRvEDbgkPl
TpCFB0Fm5UHLowEBZphPH6mWh9s+O5MOjsAIIA8vJBq8VGrkia37h8y4ImYf7wBG
SBcqp+x+EP6H4XRBlGzasxjKSzXIqypaap+DvHr+BhFWTIm5TGmhl3Hc/njlNeIm
qwvkc1D/VEJ3mx/hswv+ZBYYYFE2a0LHajnsEaNrkLlFBd/5qu3hrPfOCd8LdSqD
zIRvuNf+UaCCZWQQzTW2YD65viynLA0K8QUKExB95Dlfg7f9E2upd1bYMI4ZAHIO
g4zE1H/yJGzVUXzlAaG1vPcTsya6VpGiIyf6X+8fE135MuKqeQ6OWSYPZkKXZTFq
I85p1crbVaJqag2Yx+QYhVbC6GhfOlRuXtjudS+SiV4RI5QPnRAe96CHZfekaqxD
zglUzenkSzn0CUgm5ouv/nGJ8GTbA9QLbV1/5Ya2Bxbr6doA794KsW5NoWlAMslX
ntAhAOMxyegiztAf/rp27tQAtBFc4WUqHoF4v7zMJVp9YIbCRXSX7V2mjZs9QArq
J0DzBIUUDDWGIRFG0hPV1ybP2nOIqwfHnCEhedtAMzm2G24iWrnsfq4o46SPX4oj
j7ehUzL/7lQ/xxJDqjgBge2aj70Gxi2HdpwIqauzuz1AxF1wjJXQDJ/hrjnNdosX
mBjftJmZFph0+xZNwB9bvXUNwl5FDIFmFSFRM3QuWdaERPyTCiG7NWwYAZcETahG
v4qoIThEno5XxwkMDq8l/KhUIXKVyucbcCQBpYhO40SaSvYlJ4+caJe6a3dAajl7
RZGwB9l/MWDXPRgy3+GPZb6OVkYnZcOPxdcK+nkLzLsfWuze8ybwfLsIK02pqD+3
6Z1wxXcL17rXAb9ShGPfXnd7lDZ8fk1fOAIyerd3Z1kKo6DnoH0L9Y5+6aU515gt
hbXpR+cus5tojwzdkZeaIXQb7zhEag64evsTp4CdlmaKy1bM1OpkCT9vm3TDKvTj
oyJZC45GB7FsE16JjWOVULVkKQPP1+WVIO+jFoT6tQHdr0EalV8Vx3S6NX37Nhj8
NjnOZ31VSkh2xVvW2dAOvoz8GSh898wAKs8RcXala18NN4dsBqHv89XPBh1S7HKu
fWJ10TBUAPGrC07gTdyu3aSy5FI9apUSli/V0PGdeRQFuUhP35nkLYbJuip62kNS
krMLa4s5UWLnCm/2KTBTDs9zlpVunVY9F0YZiA6bTM9/LQi6Z6A+7HIuUvfcELef
UIvayvEUQI2td4SDyfuQdB+b1bk/VE6qKroJWt7zSKojo+PdSPs0y0wiwiz06bzO
vpaO9ctXLwV2bQb5qnH1QdJTgZcV335px/Pkuj794nNmfesaSwBug8vT0l5O/K63
jB8hLizWWXLdtdQuHWKHcVZUbpAEcHohJ5boG1asqxP5H/6+B5oW2Rvv150OCFQ+
hxgooByS92KTm5LnL4anHc4FyJDnqfN+x9z8sEY8gqbkY75OWjoacUMUa9zvCNV6
7J8WEuaN78Zo7nP62Sh8hPfxd2g3OizgmaQYSFt/RglZojMAz9Go3CNvEZ8AAlny
LYK2ID5KjvU0L8xqhkgXCVHbRikrUWAJGPQ4QZ+9pe4T2R6ixrO20nA/NzUzfxJO
SoW7s1ol6g6ZSi4OAYdUw02lTxv2UKLSMZke71Os2+Ljpc9qILdhNRG7j2sNvBJO
/gx614TFfwo+srp1s4AtySYRjrlKK2VmcO2tjW7FJ6pHYJpv32J6C0g+WTGzmoVX
k1ygbn/CL1MY+6eQK4yIDAfaNa9IiwTPQc9nRvFmsJla8iJXnhHGa3v2OeUjEjgf
4L9mSOoEiOB3GwTDAlyFW0uA7vqZnGj7UAadj6u3/1gshObZmiMwbLwY2GhO82in
jxsw4I2GuERU6rDp2jkyZQAhengt7lQpKBG7R12ZJvrilJJ9a7VbhG1qfD3z42xE
WzrMZc6NvvCPyDxb12KNHS1L1q8J+ckgI9qDWJAzF8W1u8Z5PoM8AzuzKBQs4Bpn
BpHFGT6Xx92nAjCoQ4ePq6cqiPk42mf4suYT41pnk2Q1eW7xTjnPD3NHTHtfUR12
+QAxKUlmQBydzyVWiYrkPk4hjjKCnzodfjW+ZBCZXYzyEGnDxERV3Cm+uRQEivnl
6VqcCc18b1IFxLv7EvBIRbiK8rbHuxu2Wj/zHtizs9+GlcKDmutbl3s3GdfuEOKY
kpWi3tmWnyaMZOa1s1P0Bp/F36zHNG6TKr6sIWlgEFo9cC6wvRDV0K/cygtku0jx
wcHaSkhB+uvhlmvSdtQHQSZRK8Z5UUp6OdgaZRGP2wMIVtYLVpIbQ+1eCfN6xyfo
bWZWZjCMSJvHvtgg38f/jX6jmrinGl5bWRUQbX8jmAY/d+yFZSISwLs3KRIYYt71
wXBFnExVPbT5Z7MlLgGWc1+6qpt9gujq+f0iIeSaMNo8p5yk/ItKMDS5RUMRVVZk
/atixtlKfhZLYsrVyIoLs4LB9lSg7sSiM69cuCIRFWHAndFXz2wMy44Uw8PS0d01
WqrPKtbI8KuxkuM4zEL9lugcym4YYt5M2LYi2VH8RZiiWwrne5RX68/CSSZZgo2T
fuJgq/skm+D8qPpWCP3FVX6eJxSFHaBcvDWgmZioTFrmMQxyFYXRm03URk8lS1cj
ftRB/uhb0p20iKdN0UfE74q+/TidnToGnwrIGuIZt+9BX18cvcnDgjo8EIPJObVJ
BDhsapc5bG2sulogFP8zQGZsejro9J3UbffDD62hkjOsvvl50pz6yjFoelmhuHb3
UGgIcxaOqHjyn6SyggQ/H/z/HnLvWM6jUm+CaWaMc0dtThr7vttptprnos++f05u
z2I0WE/IawVhvH1WmwMIkyDdOUVuN9OXWY2GlnixGl1max9V9A70PAYBDcZxpfvZ
Q6a5vFXMd+Y5mWcjfDqAMnPn4MnAzFGrA4oUMO1/Mv1mct/uu4h7HG5/sOt1Y/ex
D3MdfoA8Eg//ysCaXLD5U3kDU9PhOfDB5AQFHWuAKqtZcXfXrLrtZQ7xw0wmddlI
SJu5BiSpyBsUaP7WL0IydXs8Y/LfN9KRLaQcUQnUOFPaGmMPYuwIsZBhJFzN4STj
mylodV1PlOo9MPfKMgpWKnSsV/ieK+4FI2FK8PVwr8wljAFC9l3Neo4Wpp/ygmSJ
N4EIkzYyVXKVWowo7+asRX+rnNfeyrWmwlMrfEdbvhRYXhDDlscJcgxvk3+LklQn
CBPZMwZTI8kjtFK9GMs6wLIh43aO4yaLLQBuEkarem7p47SQ5harPp3gheFEz/GW
AnTXbtIaIeCLol91akDbwNCF4xUGxdYWYlLdVJNO550me3/z01ZhUjUm6EVHG3NK
02DaLaA9haL2zDX0uFALsAltvnsmkCQLviGjfxn27RhJ2XaZUHkZAoaWYVGsWXso
OuenlxwIGN1Z8k9omk65ZcLlYQvR1yDF2tVvXqXNwe/iqmJ4ZDL7zT+YUyGWxMCf
P5XproAeCvKAqAsXpdmE727obLRFJIdhzu1DFowrvyIovbScPm8hRKRsdUbjCYwp
KAf6XqkbGf6O4ZBNGl+ishxhWqzjhKVIOaMj0IxcffGoFUAk4pxYJI4B0OBR5zrT
Ys2R0HZUo36DY/V1JBaMDs4PXG4QZTS/BlWzYa2A1isA5Vt5gM42ESPcBOQcTSPA
ZBItRW+YultaaXXZ0NQeb725QwhPRYuWgoBjbbZ0FvuwoWK60ZBV1/IThZhx0+1W
ErDAkytln20Af2KP9nbpz3F4xPXetzTHrlk48uNMeSpcljEavJI7CzbfRKqDq7FK
izVJIACO+cAaoY9TJuHGs7u9FXRvy2lhZZHYnuI/vMJ4AT880r34HXWgB5+E2xPC
lRThJvP2NVwBnyaTlUGE4cokRLcXd8eeX6BB+K9H/jeEN1jUPiQ/W2o1OZyssXsC
c9zxAF9CyaQObQIdGODPL8Z8fAprUVrV0Ch/DL+N+Dsax89xDckN7RmThJCNdXKX
ofpsn2NQDmZj1CHyfp1j+ZEASVZR9QGm8jiY93iOHC8pine19+hkSvEQ499xbtED
UEhNtJjhZPaayuoUo8uEw7YTP99dPGtGTeukciwaEUJOxuoEFGNd2lyO6TqPXonZ
rv4/x78OCukQLyeVJ7HjGw0EbY+7DXK+5iPLp2HsU9CeAwj9DK5vHWtZ1DBV89jy
iRhbAYCnOyVotw1Fet0o7jlnqrPbxbrJVRoUoCZCOMiYkrKetd91eKhg9Mmqo572
Av3s2Hbsllj8S3EVS39DbkORRGgxjb13pKM6Mm2Vpn9zFot1sl6N+dXEhH6gdz1t
bRpadvA3qsDXT1IhHGW7Eok4tG87sTCZHWmjxhv7RmB93mIuppdkOEvXX0iXITsK
V5dh9JdEEbC6NymTDMG+V+oWcH8K/iy75K2KL8fYNWxOIEryanwvR681q/6CQtmL
6b0mcND1gwvY9XLrF2eENS4gme+ewhiol81DiMUs4LJGPWMmIBGZlcACU98VmJGc
ByVJkFe5wSQPT6DFeK0011fvLuJuqa/gw5QBB36Q/ppObjk/L8xPrB0M26NcmTq/
qu5EBZLjsZ3/nvmqYLEggtVJU4SFj2qA1DJfU2MPx3VjrVH2rjW5+5qrFInV+aoh
h7SCakFlmR/YX+hCK3JmDITwdMEEbCOuKrxkXs8vgw7cexYcaI5j796NiLK6tFdK
2MACRJNeI3SHpFgFyHJiTHL6oHulDLhwsN6/fHtM5Y2ly8rOscsLsvEe3dZRLHt8
HWhDnxxRA5Ily03H1lQ8Ob9lYgX1I7jSHIyY/Hs0Vj1eVelx7g0qxQHePurtYV8u
RRGtSvOZGBijMkAsGZ1CeQ4/xl+yUeR7RVx00dFN3FcERtuZJZgdTJRtmFIkSF1f
0x1nmeoFWs4/SQ2QgX/DnobpnuiqOkGIh+Ef8ENyRPC7XNPWpMm39lzVGO4wyQNc
mDD2VL+v7Wrd6LPCMe/esSeVwgbWbXs2XWLj5xsOtQP9kTnP+sVqci5k1gBUV4ye
CNEdUc3E0RXMnIk3ygpmeIdpxX+3Zm9gMqC40Dw9eOBkcf0UMUYJV7s4pdk14+pM
bb+vxuaR5KnFnEtqBdQKswNdtGEkc2iVjvBXq2rpRkcBeA9G4w6q/LjCB/r2a0tG
w70fqVfxQfxD9+G63zGTNrKxY78n0+syT8TU6NZ+jyL+r8cFlTrRuZ1EawqKs5H0
f8ZVcCy9zTL9FYuB6GjYtWTCRI7TnFy+TO7qfACg9TC6y9LlgbrMdzftggvoSCTQ
X1GAk+nCezuIgvC1fcPnMJFu/JlkizGMTOcKGY7EUHY+S6qb3+QoSYsvgYGlfAEF
iyykMm+LJx0qnhExI/gQCssg0rFN0YHPELQPqoJcMC8kDvGyQCMqn6Ivau8rjvGp
BcnpBgmLvTfv0Nc97SC39JeT81FtC2/bOYELWcjYK8YyTOJOdbDOu45tuFhY6UOX
Hv1ZF1VGmZEVB++hYYGIoO6eLuGq5JlmEsFxqg9nOIogpaG9emkwHrVRMHqNM/oO
SiT+hsM4a52m4UmrWgVlU6/V+u070AHWOAzZPSf8qy7tor8A6EtqI1W0hUUXcSu+
SBZGRn1wAfjnomzT/sjCvGnrTi06WMKFBgWOz2te6G/w9iSJAdNbfO+NcwQYMuTm
wxv2tJz02TEpY/YN8/Kim3i0wEj9ihwGijtO7IfVNHrTuEPDpUaeVAAGbBBVpzTL
G/6n1xGnzwk60c5veQRUSot21EHcQUROak11Sd2jAm2vHIM1cGGuCLomKFouDEjM
kre+vmpyJKzItSVhDbfqLR5FYqIy4PG7gcIm0tfBJ+6Q2odEO1N5VmKp7DoM1vwj
6ucnOelWVuyp5qo1Y8ZpOb481X+wR7po2n4pLfEJYQDiBAWxWR6ZA8prH4U/OFli
g4V2+QBkX9xKec03Zxj5eI9A6Xqd8iiJPbNpezGk+/t0/x0tw+1RX/ZliXFXnEUN
TC8uPRDLY9q2NzMfDuZVfOid8aH8MyrILwBb/FigowcRj6K7+PZRMbio4yCyByku
or76XtsRmMJKsRL/eN1oh20izO2C5cPnJ677dXO/9i0vIreAopHYryW/FkE1BATc
6sn/pvGd3u5OJVgIZdpA31afrZ89dVt2eeDjfRRguzmf5p+6c8sPsnmRFM4kf2QS
l9tKa7zQLrfW52Gbcj/z382YEKAQhG+LHv5s3xnsalBOA89fHy0emIUc1TVtkfiK
8OG8lhpjrTQhAosO66dMMynLaKv3VTphgqDlwHuumW8co8Sj0i1ZiG9cbBILX8o9
5Q0aSK4xbx5A5qwqePanE2smiWZo3GXqLK9ZowRlciXRx9uTHD/FUyyrUhGIYSd2
3ETbMSarX2CeV+iqfIgkbMsIk56EHslQ1o995ewXSTq19SZz2QDIJESp+RHiQusm
Dc+bOYEtupCtytQB6xNVpdpObq5f0HYffkOfuNETrVnCSWeCfd0FE1a0p2r4HuE7
lyc1tZc6yQqsWv8fAu7cBUGSeLpOIHmwKoFzYH/xX4hBJjTy4qQod22TP09JgOVl
ObM1rqVy5hABNE5GXJmQnKAR9nCpAz5U5E/aC3zJZhLChK7mga2iHHFe2bGbxulg
DLNw5Gs88o8Q/dS+qOecfUuQIL08DNrTGXbutfngiACXQYb+jw4gzQRukdNRlGgj
4qw2tyPA/3IRpC2UYkjDIroC0hYNyuH/gJRNYKDGjnkaDeSedLrg9z3FvwlbU6Xq
GS+rtEtP08pwj1qhlLGMN1T3ZclBSw17jIb0qZ7P6fFZdxsvaiuoPY7OC55TKGX3
o12PSwMxzpXp9dYeH1TYd2DzBxecvBwDah049b3DhlUyPqykt5jAO6YuXZCSTanE
djWTtPVkLp/zkOJwj7/Pz9WDsUbbKWjWdVRHMSou+NcfSBpFCj0HFCBFYvzjNPLj
oWUWMiknNpvAAVEKgmBLfSf4bnv+v+ZbFAxhUlMB/Itw9vT3QQk5uRjxfYZxhV2s
P4QV4oV5RoxuG4CpIECGXsA2nXC0pVua3HaBcoCP0nkUOe7T0923t720AO/fXks8
orU7P3CkxLj1agXeAfhO0uT3QEWlG8md2PXKmMLlxiByQ2UL/Fgk7BoAfmjubfdE
I99dum156JszX0OGBS/CVSoAkzj895UJaekTdib9T0nDjEHI8VrYlnFPyhU0M2Pn
JQZSKfJTbx/s51In1mmByTfzojMxGZfkkHgHV1dMhnVW38KYtxprs/N7r9fG5AIg
iwqhqdhUPO4RRbRjr/RHfV1Z6ijD8IIytqvOarcPnP6f/D2D1rqgp/CFeHk/d/XT
a/IcFrAIh5o9QaE+V5x8rplKasJlGqMpcjhuhP01AOFl2OpT0Vmn/v6GQkNvWEmT
I81z+9pnUFmNnz8D2Y5PpemOAxkAqM5CGDTzIluJ82DI0PdfZeFqWpHBUjaWb9by
NXa1HqH64QYPJIOfJoFR2n3fzcEGzgSDP1NHS2UrwiCXlb0hrhTe3iLmRRWGMHKg
5iu/qkVOfiJt+ew+M0f+xYTSlVGMGI6J1OsPcuP5hTLbVQFZCc4c/5prgStE3y0r
rEvKa571g8KLxR9vSMyF3q+uJJ1V5I8Yv1Bi0Ng+48PhQxBlIaWL82zFMtmVh8MT
RJQwkDFWGoHnM/uuGwH0NrGYhL54ZX6+4VECXUspEYTdh7UkcWfXGCFfxQDEt5qr
+iZgY3BROSuPRO/H+p0xTDxzqFVRyT++0o0DD7MC+cGGZIcaSAmi+ldCdOnY1F/7
SpYZCfg2Vb8zV3GJ03qkGJXBGIC5R6qxzZWglAx799olXRDfjhO8BaGzy0C0P9O1
H2VBrk0GKvuM7Q1DRuN1JtNr1B7g8Nz4QZlIZuEstSKbAcGbEUB5sDquS8voTYth
qAseClDbaCoD8toIs/iqLO7XiCxTfFJBLVE/Zvfn6dwfZMz4SiC18GGqBS/lMiUN
i7bQx+J+2JXZQm5heTvIOY61jBNroOZYKQbjvFtI7PULf8dDG7V/RGxfY64ZEMF/
3UBP6W8FyOsJHtWtRqODvy4jxzhzuBAPMevW+kJ4s3hWjDtedjz8yc8EMV/uFBQt
DTdNYYrFgxqKFHqaax/kbmrUhQJw/PeX2K5JlcJtS2PXCQUyho/BLwJFOlwrQ4vm
JpDKY8Q3/7kRIxSaZaBvD8bCBJCyzpq15EeZEAWM2hTW15Pk6PmxQFf2HZFC8VCB
lHEchZ4YPhL365F5woKO0BA+QCNjMTJqKM1a8fcwkDNm/dIGtvIhSyoesSYqz9va
FcuHhC40xAu8D+6m82XmyoVOuENCGPHwPFZoZf8GWgApGHug/O897327fj3IN4Rk
Du8LFCxzCyAZCeeGEoNRbNKCyPlOshhEgb0sO5QJsvsLuX4nJdpAjddDvKXy+UiG
3FtZAbwxJ0Rpif87OtTZ9ZLnqAyPy+hv+sxPP+anZJQ3w6ccPJA3UPc8eAQ7WtfZ
OVcb8G3YeLMUeHACnLV6asKDlYKN4QOz9jf+Eg1PrjGpSJ4nLVlRjGzKaK8o48eq
cDSv35fMqFY+zUJiZrl7Tup2CpgJLZibnVZG8s43sOqBmb6xqwffLFvI32GCDVhC
kUkRGDLxgL3GN4fgpTI+h493eZUivdKJ0N6EPCSwSgxBxxD0RsyU8Zjj8Albk7yo
LESr+JJvTsIpbgu1Rk3hCd+88QyKe4qcPQKRVQPa742N4DQdOHSZoFtP0ocQezaX
MWof8h4HszCANN3gJqv/GLHYsPpqueHbBLn5jmWmSmIyTpTW2h0NNtFYcgjlv6Kg
e8Ec0opTkhWNTbZqifRx6KrwO8PL2yBauSD+YeA29hxMHd8+18BwQe/DpXfUsv/7
52itn+GMaPomPs2RX8ukcObF8FSBW+9PckXNOhiglSrByS5Je2HJYREv5JnUBdD7
J/HATdx77hTzyLwSDhrALZJQRY3h+vASAR6K7U/TC3dDkaiXkFesDU4sxwvPwne3
MEheb30/ys/wNCFoz1pk6Mzn9POMfsZtXpovsBNsbeT8khJlHbsTLDxYPsZQJUlh
steldEWTs2Qss5WumhzVwVDWkm50Mx8s//+PMjOsS5RZhNsrOm6rpIy7JU4wA7Xe
fwcplnA6KM72zMEBM/IJJBZ7doTeAnrjF69AEFuTAy7sBxoz1zU9YIne6JY3VT/O
wNJNSYZCnjkQt69g8JWdPoBafP/Gj1ZmalPRjzwqVbHduU1lEN9U0o/sMV9FTVQa
VXWXkmN/F78q3bzXbF1yTGLomRP71rA8IE6iEwSHOvS3zLsZYpeGdCKD0J2jdGuv
mUFKJPCVAccL9muU9y07cmWxtRugSu7ssgSlyTZfbW4x/DjmVddLQsSRm8Slswox
6i1PjLIpSZPo4j03cr7fdH7f24+Q1nNQYcUUC8LZy/IuqWBdX3FRnEVPLH84gdoW
7nN/0ft1aoCVUkEp7KK+BWBcz1NE32MljJww4tK+XD/O9spzgsjqwSgf4zA/SxOl
HOLTJU0Z/6FPGM57vkOKd2z9NLHTNy+AzOdaTJAHI9ha/s33yGSMoR6ONwiWdPN3
fXtt5GkxmEg68vRqh9p7CIUu3ra0GBCTcTJ0SfBRcjnJHZtMyMXZY2iMd0gNzFmg
uktdJTRxPg3wFRChCBYf2CXXiwmeXt43k1bH2joM80puWmGE7rhMY8RTvuEhLTU1
zlp/01+vZV9rqpgUOu+Z2zhWD3jZflf06w/nOTHhQ6oHcZA6dAkn/U0yHL9aiEOk
Vx4/KZjfYQoOzki2DHvl1m9CIVs5TctMiltmje+25oU3I49erin+kJ8akQ19BnRT
IAmElIbk3l1ICYyLLbg1bvkX3xx7Jjt8GMUflATmFcJg5VlYEAmVtj+/U2VZZR2A
aiDwBNhQvy5SutVq2lji3uEpC3OI28BxYA592YHl4qzNmq6TIHU1NFx9vuDgaRnU
u8dvpDbCZOD/DPaH0C8w7Y1HWuNRHZVmx2lYWOEXUV19UR5RVc3X0/G9sVQFU+g6
KyTh5LyXNu4y+dLtaKcqMhUOCf+V+4IQdFmHKjskoQGYXwfZ74lEs8AIXY7D1IGt
4belUcaYe+a/I08OhmZ6rl3oKSHutyZxxtbZu2Mc/aEkasrYjrMK9XDaePSKUhee
Flgm3Sgr5Vk/0+6Gj3oroMrOXA3gNPLkPjV3FgOSvqsEEGP/jINLkhcMtJ0/JWot
AffhaZcEgVuakncjvZVBK3aRV7geL0EwytCoYXIh3rEvvihI8REnBN68FzRHSzuq
OLwwlWQdMmYY4pE4Tq6JZrVgKHWx9dNBDteOuWqyKWNWnYNJtjGuw25JwCtRRnmU
uOjNciXBKUfVs0oYf7/MNM9cez5Pvcxb9tDkGR8hnnIG7Y/LYSGM6vr9k88P2Ret
dGt7MnUx/pD8ER4SiNRF61PmvpufR18Qn+pRxcbzgvLs4rK1GA/Z/emicFF0SlHB
nsh4SdxvoRDxt80TAIh5pEd3XUT3WsCrgh3nw6pcQRaYM6D1e8QB+HQD4QJIhPkw
L/pov5x/bg5ZIMruhj6ajJzwkc/Wmq5PTGigs+Zcr/hgPglCtEBaHXuMFzfQckG1
gvc81itwpMrKzwDtiqsH2Lx5PSTS+JVGnI6sP4+fXb4+YwD8lCocbUPWXoRlRVrH
U6qsq8mGn9FXSADxcN10l/TlhikSzPC+3YUlVhB12izxESlZTUjqUCRhVFiuyYuM
t3y6YIMGLtnsuYNDYO5SvCDs6kTZgJ/mmuHo74rwx4G5pqtQnPiyfOwl9PpD9Bgf
YuEq9yORP10QpriYU5M7d2JbhTNVqCWFefHaQU8MXuuZrr247qr+uNQVxDo+V+JR
rjPMC4F1Uh0x7PI7DAi33nk236md3F1gK+oE02j6JEKPQMFqZxErSlSAMqs/IV9F
KlNBrANfTcPLBboqJeYtd81bycYstSbVT7UzfU7qiq/kSTrzUU0ivu8hwSQFUSo6
bNYtkIMVHNkYokAI1EsrXjsOM9Ga6pfhdsoWem2GZ/q5sQGKNw5w4G/POVGKgf4r
d0m75+GWBqQfKJVXvbHWbV/rhOPXoaD6uqWGgBYakaUkT5j61bqXKaDM17wevUVc
R3SzFmv2ROihuBzLxVsjrr7f54y0uQaD4u5daWXsUaWLOviPxlSgnsdMegWX7WTq
mscYHKfoJRHQn8hsxAXyrFE7RGx95GuZK9YV9E8fYh9OFh6gwuznWps6r6C5gSNZ
z+SqElZ+bX2cAhq/9bIPtgymcldUSrI6lsBjVK/ly1p0iNIpk9IkQUYutrdcIlOv
f44bbxy5usi+AptoNzJ8941dUGT8MR+sDAA2ol2XzBR7m2VwLfvNlhV3ICDvMDFw
1zZwz5Mznp14islbV93+aCD6w75Q7bIMB86secYmF7ZKLzg+yFfPbWCteASGF1xI
KlaeRSSQs+nngdPPW9W8y0SRK7Zll0k5bRyD2jNqimpanJ4B75O944BF/XdTKeyq
1KxR8o4em1vpdzoxCGzN5Gyqu4fxSoSczyqcvF1K1O3Kq1O3dPmGzdla9VuMnYOB
qxAyl+J+VrM91VI4Du+ClGSHG0RUeE6ukFJmMRnfvQlF6ESTF4fQ8VPA6Q532bsZ
3BYZGbTtpu2g/7rP2NcKYN1zMNmxiqF3Erprf/oOsvDoY8WEyF7jRjoXlMRnfQzw
zSLUpRkaxyMUC28CQ8c4h/AXlPoTuCYZThGCtmHnj5kC27xBDF7gFgF86fF6XQVQ
8pKLcweXqedbfs2FVrooVUEpc88sE7bEtc0TWtaXSujAjaS4NytY2lJY9CuaYDnQ
XdlFBkEQ6aS/UAlP8UVl0rukaLuLSz+7eIDVTko3VrCdHC1AuDOaYkJ/n3rdifFD
ocsMqUImdx1hJXMQ6Hm2ffnMUQXQkmd7cI5hXAmuUMMbxA6iiCyxRRE3TR36yG9y
n2cDdbbmkuGLrT4Lkm8Ret0KGJI7RqXOYtnV0IziPpBqOwl/joF6hYuJHVz3VmKP
IpDSjz34mVHqIVkasCno3bub1DMYgpVdkNLjVQ+7ikWdsXamfK8V1LrgXjTsk0oq
cm2hvUWnWmeFlCXsksZiE4qx/vSZm2vSxtTk2fz//aHzIvjODkiGyxlkIWL+UJzq
kGWa5wsok0udbykf/WUJPp2Y4+H5RW71S9k6aMIHpaREgwYdaZt8BQsBXq1ulzmR
CQxuLU4x9KyMDb+5AlbW5GOwXrDJx52MXpSquTrJrgUKho4Rie69tMtA391fK/rU
bpahnvB6ep70yOxfUM2sO6tlMYE3CDiYk1cuLIw8hdSXdQWt8zQnP3DbTh/ZdeuN
2cCm9n32LER/P3QPz9UFG0IjD9haE/z/MqieiwFcdzWnKO4quiRd7rjgf+34pPmL
+h3XUe1frQCODV3jYJFRDqbPnNDMy8vz9bEPSQSnA/HNu/W6jd6TxzeWwst2vN0C
Jqyvrokx77YENZgvhqJN3HC7bkdHt/Y5y4djb56GTpgJ6h/Xcoh+skC4I1AhApM4
uBqcQxaek35UzaqJU1DQRjF9q0+Kllq3UXTMFhKG3H/XvV+hEj/DGm9gfiZkRWpk
AGdrFl58IoMONKJUha768dfZvb6rDVNJus36AIJpM45PCsNBBMNqucYObbPY6ct+
wfZnvW88wQyq48WZ0ozlKDlXzAqOHF0clbAXFNI7+U6SRJuF1b83+fTxB4uk3eVJ
8aMX3n4nUN7EJj8igtxypzTX6nIg8+vh4MaK7wxaHYX7UYSOF/wFkXFQTtvSaNaQ
X+mx29RA+MF99ln4eiWr2yZjWG0+5IO8bJL3n2DevirYxY0Piy2GUxyTOc3gdVg/
xEbMeNt3JdTRXSorqdqkTsDsLFOIc7Xqc0noDWQwsy7+IjWw0BT1BZ5VWZMiGJCD
ku2I5+/1Np9g27bVBqzmAAsKSnDnwlePyF64WmO7uOBdTOqyhNIxGUtOOLqeyag0
LTmenEvyyQ4e8zeY3ExRw47oRA8jrcX31DPBeMQEDehODmO+cN2IzAGITllWkqVS
N2Vr+au18wma/mIdjKg/ht7kdFGWS4pD3rR410DTT9SaeYBzQzoUILCnVWPwGBVC
U8u5bDhcppAvL1BcqCobJ5D/TJbmVwUdjmM1z0lV9H8ym/9ckMprh+9b0Tq88JQP
vJO4Zjuiif9kGWzbulqS0sjhnXa0F/EE8V52OE+Jgpm9s8OG5FevYqusQrARYp9n
BwN7RIAKzP4YpFyhcSWiVti53Boro3lk1uLfrWZa8kKroSdSX0NaWg5hdQdyYSVh
P0LZ6/Gozdx5hypYXEOxVQUOLVN1NaMXQlRV6Kppzq7FD0Q6kksJXR/B2wjQwhgX
KATbdv1pl7xkL7gApRU8C6xrm/tz/F7xv6EbhLv6oqJv+i2OLJ9A113laepmGoZ2
8Nm7DqgKdMYhl9aAc+q4Au4rUdC71BnSJeOIjHbRlsWrZmUoQFrGhG+Dp5uabPua
DFQgihcaYrAW1c6qlj3amSqoMXly42Oq3FUMTWc0GcvmVNyZCjc5491CljcIhyfK
PBoiAN8x7fJjoColpJ6x2u5U/XAYHoW6FhnB4qfsqG4s4G7+r7JesctnQfd1xZB7
hydCcBy1BhJ+rE9enPHQS4ceDRG6JM4v3j4e+qkzdVXFyoLVvi48gCyrrEOtndxV
Eew4JHAHo8+EUlNtQTW/OGI+FryzqmQaaTBuTgMxZUXaBKKAzU35DoVTjrP/fREk
91Eo0NWwko2DfHrG8Wh8LuD2Cu0J42XUi4ioUOzBlC1kT6MxA6Svz6epSbMN0xEW
L65j3U7XNWakQJGzJSVlVN+sCOdIgYi2EAi8+xDl8QRUI3IjVcqBVXbgYBTbrZsK
C9j5K6JJ/mlT36hzjP5BQPMkfddPMyPhetw0z4hsAbFMZFOsEEp/R5+mFy9u+8iW
1wFWlGan0uLzxfbsQyqS8IlPZ0VW4gyLfcs5Gz4TX71nu2pfNPh6DO0DMJafsiC2
Dfgx+XHMeoJEoPbp71znuGbBb+pXmdwM2qyC4kxAnRApELSqUKO+UC80pqzNlPjC
F+s1ejJrZZF0b3f9ZNwkeuxEr0i5QxwezSV16PLb1d+4rFT9gVd+yy5yQ+WBwyO0
hUSvzKkmtJa9JQwHUM00tycenbkWkNORe6MSEZyioemNJro7paTSrhVo9HCGvV9P
oH7Rc+1fAUXJ3HXpcrQ9TPSd1+c/X2Il9qC7XImAQHdKPxYszjr7yGJopsxjqTdJ
GgUvU0CysRsgbV6oWVhfeV6VMuBTsuImft4YqD4hrXMSyIVcMvyfKU+2icU+ZGHk
tdplro6ZIipicMK2O0v3AOOkaCUsY6P1bCEcmSEbK7BAH4Gj5G07XBVdNxYudIxi
cpcyXQ38m7Oqk0CS8fklfj/an6NzJnHTlcv/p2VUgdDunI5Z4Nf1tFVOUBguveVP
Iwolsn+Vkz+f4FKX8U46j9ziKSDBO18Dn69MU1VeIS20VZ1PkOR4TdMKJ/UoJk6+
DwtK/BVDPVPlOIHMt213DdeW+pDj2X7dYw97RaUeCBcod1U1c/eT4+i5kgeq8Kfd
T5krM/W0wvCyl+lptfwV8/QhcyvPHdcS91rpd1n5/C/4o+3CMqPezK8yFWsW4CG4
6ZOWjw5GqQYL4+4Vl6oLgsY8S327zXhzguJXFvMcAyCatRVzXnv2eNHMZkNmqLmA
Hp51kZu5cci6lqNUTUuvkOXPnrFfn1d/PdqrDXv9wFmBCaPXBDUNlUxwgYaqPYRK
3WpLcvdo+oDaD+m+NxFQ2jxa0WX3U6imNCdk+qkbhbcNc63Lu7N4o1FvVCjZy2U0
kHSg+AawYIVbHmypScE39xdm5AcW4NOZ2MHcoOP7XeTBUq4vWOZRg7Vz1Ht2kt4u
h8/+hx3m6ZuFhwneqauPsurMD46It+g+Uy7q4hz6wloebGsHdzrsIZdzxGE6/hAh
O7+npg2fR5JZUUrclCW01ghGY26FiQ8nKzu0fKsCGd07tpRJsgXKnZysKMH+SAvu
PRlrppTUA5MsbsqrmChROTa52MBGtpTNwwtRpjS8HN4sKVY9y4YghP+o0rGmyLme
E81BYihVXShNv3LbXZCcVGu1dhsUjcf0ZhgvkkAh1FMAa6lR7xPzgk1HZ6Tn+ly6
P/4wkXEqCdM3894BBszU20g/b4aoy3O8CBd5IUd9cRXdlxyarWY5O+mVZs180s+x
vMDoMazsPK60b2mzHNAo9BJIX49jG186aP5xSS5GjIywOlkpPkNASP0ysTu++v1W
rYaCa0Pc2LziRtkwv6aPgCOE8FTxs9GIrqCSrT/uwm7C55TA4g9lv60KSmJjfagR
72MeQindYDGfVCuabYO0HAcaopHzj81ujz3mXSs5Y1sk9Lo3aCpupONqNIwRRQhC
OSOvJ//RCRGm3aGojMBLvgTmoHgZPjvHI9xD6gKpIRNygZbs9BLvuVS8rRTikZno
RU+G6c3znwC5WcaOhDUOyi0A2puQJJyEyPxy9O9gE6euUoud+x8fFyjtrf2nMiEm
sy5zBND4luiYb0ijKNbGmktrwAx6lKcR7PC86bNsiq38hk8rGiPZJ+LBKtyDUns/
qKv2haAWahVcKNJY2HlwfLZoRQ1n9klZeTGKPF8g98tK+cURcj6nqbfPyFyTQ3kH
4nba0kP3FWViwc0vxyldeNaSajAtv8xAHx79arIwt2o1nJN4m4G5RVNxWHwx6xHh
YTc+cA/73qc225iGZZqEVFPj0uuYvwvDePhq11VbvTh4imBvSzctYCCZGnZMUBSY
LQjPgmJlbECK9qJqs4ADm6BqOLUGkCzgSBf3npTweWtleUYSkTieoUJAPf6svYdX
mdb4NYf2SaGcLsNHFL+AAtXThVzq0VkkBQgL5vQpZSQ6hfweliX4w4ks0yGTgLPg
/8VBQvS822XXyJuprw88EwW72GbZOLYhUcqVcE9FLycOVqLT72IBHCSowLkg25hU
qy/3t51fWxGjm123Q/o7AK0gulwICEx1zt8eNM6FC35o/aIy9S3ceaSvZ8Klag1w
NrOzM5lX64h09x9M4RJPPpZXt7nvaNsz0pM6M09TGh6vXxTSizBb+FBWO49Eit4p
RoZDbSdX8T3H8Nbg1OEbhXxh8tCZLTj0pZv6BYzE2Syf817pZCLQi498+TFdeKz9
I3q67R60Vi1e6TIZd8qddWH2gqzkrwXN1vJVnlG7f5XGiRM1bxKbGxcHKzt3jAhh
r++Eq3pRdptCtr+tJx6YE0WDfL/A14cwctmhG7aDlCq9Fo+q4Y9+EeeGf3zhhXWK
EpO54L0JqomfnAjH7x++QRpUPLMTIp5Q5qWgmcVJdgalZUi8b8Cf2JTBcXss1Qgt
MlVVwNGkq3+Z1sQe+AFXPa0i6r+c+tYLCzs8viskONAhQfAVwfytP/5wmUNhYqCR
Yng8w1oFI18MhIPaPP19vqfbUISbT/UjMInIQniRbB9j+MGE5LDnIbff/YXotiFW
CyDOVG8kPo+HJW9E23H/nzbjgsnDO5YER2QNJ+oD7IgGm5kCL0fcG/HANeG9aMRF
tBf9mgwNjg6sF1UEZKhi7OV8jmqEIisSqnPSXfSk2YCZqnrQne5M/ggxUNGwlHFk
RRdaXuzArAK3VmAv++H77nErEso5cJ9uAGE/Yl1VrjxFXM7/54mYhz8fS1MOGMkd
rHfVD5ClNFMIHi+Fdo0I8BQxBqYtYLEhMpkvMHAw5Zh/Kyl4FdRH+QRO3NeiwVmg
2CRPzAhQnTvPhlK3SbeXw7Czu56ZdNDxMQcwmHvn02pDuauRVn4pPTbHEOcRXuML
y9+58woX5bclly3Syxtyq5D1N9oOtpPP26EhtDbQ484KvGL6OH3RhdRiN01wKwAM
Rq3sDjLKtGk+hmXRpUPgpluoFHDTkDvWQFJ6GvatvdZ4GUzQmmaFWgvSEQVmtZW8
uiM8sveaUeeuZDFvNT9U31hwt/DK0wTel8KSnXfQWIEgtBbGq2Jkfm1gwCa28/zk
Faf8/5sCh8P/0ylmlNLLW807eBYHja38qr/YqZRqX7l6ce62ADKKKmryv/xZ3t+E
mAsvJ8OsjSUml4nPb8N7JzOApRYOZrPjAeEuqjhuGePtaTGWbYlsFQ+oA+zKEB2j
GQSaeEWpyjfZHsOsDO1ldepAPKeVbLrGn5GMNpfpJEnL80vN9gVFkJKVIOL8xiab
oUTVbztP6xLasD3zCpXykbBGlvrog3SfxZmbPnocXuat12a+/VvOhaQxeY2trvvO
G+wwOHV9NZcgEcPUT1dMX0h9sRFYQL89pmtoylFHIo5OnY5XRSchNLyqG4+Ljgla
J/v5k8L1clqodJ0omSWvnJKjYKZcawamuHvFxdusvzyMkPx/1mn+4YAMWMM9GURj
R1wUz2DJmFflDZAtN4NJwsCw0P4PGFvV3tu8tZ1V20sr/FCuqlXGeM0/qEpfuJ1s
zFbfMupPwpMeH1kOirP6jO9W20Sn+SIHDtnJuPaidXCqgoiZGP6JGHjB0PJb2tSe
lENinPSY7/Dl4kfJdIiA8dKa+zuib7xC7Upl2A0BGgSxDzUng0j3S3nPKA3Ytkyh
wLcYqSIdrAAVdyyz6hBlIAqLF/wA0mykqGHOIQqplBlhDVlAa4PtD+Ddd8xvQs45
zL89SnsqENb+PROu5dK5OWka4Tf2lrGKMrZVhzcqZ3nfEQXr4UqzCKSoquQFb0it
LUfdsNVrsKS0LhVSOH0ou4tHLbhgKqMOu1SX9/taSd1UCgZBMh7BEfSCnlguzxdT
m36LHVgrDLFmfLOVhWBhoQMb1YejYJJjPsZNosA+IN5gvpUHmZPFkrQVNahL/PNH
g+1kgEXkRQ8UbYipGIq6TvaoKZYBvEwvH6bwQgn0WTLDRo5so2mj9yK/1wzmTZKD
LY22qynOiD/e4LFwzGu7Mno5B1fOMkONtJAVfYtotv+bFdq/sQQNI1JUxtcTApBm
Ce+PxqpWl/3RQ0WbIoJGigTUVaOSvpZ7sskjAXshTKIM1guRGP5+jabde2EkjN4x
OssWql7ySJ2Sw8JZ1tvcQ+UpMbrfGrQfDfpzqA0d1Te5wjSgvvgBcUb4NVWTEXOY
2RhBkvme9JwPVM75NEGoXFie37PzJWo36VVfRHp+0Gb2MZUsjsoDolbtnhaO+EUY
dM4kO9HZlUh9nAUFnjJZwThipBnZA61dS/GFEQFrHI8fL4cuL8ArFIY+5vCC1+d0
7gTmL7zBeNRI9yNuYdbVOXCIbZlesGrfO96XfVpFNNWBMDD9Nyr6G0Cw8kXGPW7d
Z+LcmZV6SSHfS5PqPB0qgPiZAqSmIQjR8Ydgh1GQkdmEDeY5pDUTUrLQhlnL6HIO
kgwy3Hk/lVyUd4Es/rhQ+D1jWmCJxM/4+81f86yRrtHdcc2/rMdrvrQmU+QWFxWS
uPZle0aTq96tbLoavlKf9wPxlZ9nDP+14QrM7BsYbgxt3f+PM3rsPA2yIQYrUU5t
/n4PUayT94LsPT8DK9dsrLjTdJ0GEbtVdwj9ODY2Gc4wATzAaS0TEIZTgN+EJotE
jTi6+QnKdLcSnN4Ft5IO536Z/ZS5CPrA5ruy+ybEVWpc0uci1+fzoT7wq9JcKRyE
KuHnf+/RH49btWeB8fnqCSviXN6ppWFrY4+FGyuk+NkMJvL4Zp7fMoAp+Z8EBTRp
8GlBJ1Py5eIkZ432g18mYW8mVlDjvo1ZIRjGLnEw/WjIG/NtNQ32eiNaCxcdggav
nICyI9qSxaBubgssmgTwOsqyVGG9NrSloRSclCoupJ6qJfcTP5vZdZJAEy2x0fiH
VjM8uvcK7PaG4W063xnjh4z0j6HQCtYmaM+8ieG6fbzIqdAi/JUHepUrw5NsKW1T
FaQQtCG9sNYdjWsZZRyNDGCEdm5MPREWYXNyVUWOOxYFouCu3cRQH473jnPL97Fo
XRN7tkU4lG68KKP1NlGTAoEosWrsh1O5AL+Y7SEcmePd7bVdLpxzAMc3RN8asx0G
oRoLdUXzIbllH4sOE1H4C5Agj1Y/c2kPqh1q0I0pkpqI+Ppx/noS0uF4g2s3i2JB
RXjX8fA8P55BUNN6mwtSSr3U7i/Gj1xL7o71dcZLJRNU6va55gHOxWZcceCvyyRm
L6z79wZHYwziTknBY5yv6s+zZJQU8JtHeQJW53Rl31FDJlBJgy8J0IUTsXuBfrga
f3ir8BFaC+4iUFhh5napGPaapy8Zknj6tpAMajkGLI8oJA5dbsBGAjtxM7iHEf+6
cb09FMN1JHdoDbAYA3zHhqmkP5uWMOsUXs1wygWEdKt/K35KvyIXIbqyzDS7CaAF
iQPm50QmJ0XHIHKOv4kwFIdpil1LtVdi6Hx1OBk0PRArSyvfb0C/HaysW+XY3QI5
0F3c0wom9ge58JkrrGu8JMHYCtyuBAVN+oGRez6PAaz4Af2F73NEnoOERw47WA7q
QhxqHwocX72dK9SybRNRQ3NEC0akccRKevfPPpYEdsPrYcJrCk0IYCZzWmIxC6ax
c2K1Z4FqpLZSQ9DACkImaz+hWQRNG+UBuWVDQbCbOSOKAEpXr+I3aKNEjmh6WBXH
X3kN03qDLp+t/7yfpu5R0lApHxgbdSWDxrt6nEJIt6krKKdOlb/8Ot9ZC3P9plhV
mT2UEzLxf8d+wlwDTZavvjlC8diLKqqXlM90bpEj1EikJzshrfxbyVEm8DBmiIfD
n2oJE/saY56BvgPd9jAdPQOBfvo/fGgTmz53eNqkxPSmMZYt+3hz6sXL+e4vmodZ
GcyuGyv04u1vcezmC729iJ3G0F3GfJ3XyvQHIhcc2DM90XCwnYyt0RUNmy9N1blO
nM3ye2yg+VM+/eLjA+lNdIv/GMnARMbJX38LshiGlpQji+RJN7KbPiRlNqK5NTAd
LMcJXYdssMji2anBF8H3klo80memVecegfWWiCZhqa0AvRulE4Bsg5WepVAH3ebS
VrQMWzPXJR1f0Vit76NK33FZtfinXxOYyA/FDvn9TledF4X2EQmVrrMr/qw6q2fT
Y6L0elQfJyQ/ebTu38SXr0cv6hcSlV+nhW3dJldTpk1WCAoBHD+UW5fprKiMkukX
GwVWUDX+71o/M1LucfRUZ4DcBZHiconsrfVfv126YMql26KD0pbqmLiryPNSJECy
NTgbrQcVBSGJQlsNvzu6BwMpqyWYqFA8/p3P8VM5M+oMINcdoYvB92SfHlIOgIuB
kimeQvaJhOhzJbPBdsYnHcnRi5pde4r+YXk/e3HSeDABEPKPHyqldYSpiEAH09RY
JwbPcFPEcnCR4Z9rOUMZa2dW8csMOfCG7NqLahqccr7dICOUMkDkulQQ3pMNTNTm
jFLotbLXAwAx5rp+7CtnEc6ultwFETt0yKWg83DcSBBTBkYVaGgPc7/j0BWexUJp
95YsF12nU1MeRELbykYX7lbxoJqppwghjOSmjbyYpdu7wEG9+RCx27aRGTLRQAjO
MwKriP74xb/WWjzSH4LwoFDrGhPj7rq+mOaltxuhBmNnXOuYRT8DkRdWNki2pxMe
bMI21s6rCCusnUL0v8EZdNURfI0oKjayE3avzUKcbHULtaaaUiMrWAmenl+nR/WM
RISqd1RTCBFj7bIrUmjwufxQQQiYilLDrJgvPREzGW0Xl1rw2Y3Oj3H/bY5AsEgs
YC79Kpfu5uKNdQ1r5lc8Y37ZLcxwr2sozqW+cdiSFQDw7wSUXEeXJfoVKjvzj48W
9q+eaEgiod96twjRvIf5Ek0WwIm9U/Uw+EjOjasaZJiG5hqo52RlxvV4n0xuOSpL
6C4vR/PaOsBdXWtWm9eEKftd5/hjHKNRCcRdNP3v1fSGxpp24JosWFYPnNl46Y7a
3aiU7EJUJE6jjLSgWqXskQ/D4M8c3QUwu5o1IisS/+iHXxsyfY/XGqoX+PrnaFr8
5yjjsfqkpgm8A5Lae8EPg04FQq217y6pWG//0W2ju3CR/4fQAZF3zaTWJ8a6XFNj
/umff9nCGXY4wvQAuNrWW5EJXNMoPEwCktdz4BMNL+wHYDNzoD7wX6C1XO0ew+g7
qvV+9JxVaREBdymA4n3pMK8urEnZqgDIuNH1WBoTq4eECzslqcYcnhVS5tu5mKOC
mUv4Cue8/NN9spDafDfM6GD0oiaGfOpxpc1TFI1PEdxPYZF+wzFAYYi7jLXRcJDj
XdO/6HhQ8VCaO7VMexok4sjuXoE197KKDaJokwhuoOPdSkvo90zvQ8bTulnGqN3I
8Wc+Q80Rf344tmaUyhawTv6Yn7AEEVKDNMoZhLqoDuNwQ/XBm4uUZRhL11OuUuew
L3rv7d7rMXE8NIPWEUhvKtLHYGHZbT5Y+yRMgs1DUfDUp/VUTzCYH4VdqO9aaCMg
L/08D282Vc0vTdwyVbVfgt8uE95qzTNm0NNyR1pLK+5Nr0Prfr6BMWZ+SViWkTqA
w59c1zG1JWnAZtLmYqT+tYnF7TG1sPq1BuLdOnuEAvB4f0BTB0UZItN0gG1TdjGx
W3BNJbQr74B8hD9N62U+69tHMwtzLOVfsGr62g0dP2c2h6yr8qzv8azBbmWrfDqe
pvratei0tc71VgDmkmZVJlkv3WwuXqoEY2DGaf8XygN0gcd1hXT88b4NWKS8cK4m
x3pVPS/P4/8pE34RsWkr7XsrRhJCKdimXCr6/daHaV4uNZnfN3b+Hn3STHget8Av
DbAJXl9kgimngJomOytEYwS+88ewMJ8E1Q7p1S1pHIlHrwPdM7odEE7XzCQLFpze
I3ohJW1V13fxTtBT2LnTx3CCl3Nj2m+hlJXjMVJjqoD0z3ShLjP6Fbqon56HZmJU
W+hcp0UIOLBUibrc6d0DXTxAIbU5lbNR40cgXRlx0RQf+KqjLdjLbvbNDSFMD8WN
pWHDiLVcLUbo23rYcbOz/d3WErvf63UUl2hygE1m24KquOVZG30KLN0MwVeAKuzC
avFLHJm4cglyL2FosNJlPxPsvevvbqJcIhs0aykjinCo+agP78JzIvavlLeCMzOJ
8lGubCWNwZz9p1YjmgL5NjPU1g5NGenU8wve1HabB04Ar+exEYD2JXGYX5CWERKy
46le5TmMvMtvxqdJWY/WxqPZ8BkQ+fUXwhWUeP3BI7OzW54Qe+qDK7IRoyWj6rUz
Y8gddGsRFIqYYYayU0body2Uz1TF3x6n/j8T1jCaJQ4Jk9PrDDNIcjyi4QZDfdpB
ifaj/s1ZJP9fY0IJ/uHoyJAuSiGfoSz56W3NUSx2EQ2ALtqRHI7ff1SxwpoeiUkg
1Xz4l1uIctnGPFBntDme+F043vMndONZmvmZmG8jgFE30SzJgmCPSdTjHC2PYzkQ
fXVMmWyInCNiwCZ5sM51URDHkIqLlFwsPZ9zSRpGQmZdKBX/nkNM5ywC5Muruaua
I8Z2+fYyRIpMMEjxTHLeCqiTUAVDJX3kMzvf5+ZgL8lvmBCf/W/dM3wlPGhlDl58
LALCANfzodgxoBueDgB6euy5+4aBWuiOPuMlzsz4ZykvcAkUp+eXEi3dHJ0KuZ6I
XfWtUBY8hCj77euyU4eNIvAkGb4re0mKl0Htmit+qVmI8FCdWP6JJRk+qDAy3D9R
QKTBZ+tivm4lB77ZgWXm0NfuBX+LA0oXx1TVwa/hdXrKYw9ne9oyAdyVR7MUnZvv
L6oHZZ2Bg53z42JmzJ9oVhm4FWRp2Y8vRCo5JgTRvSIR0NyPoEgkDFWvFKwvq6Y8
9L2SLU6VY0pIS64BlOlXuQJD9DgX4SeIXERQyUianePDdXbHtqaXg906K1AZTyVw
ZKi/oIBY0ZWkeZVtuf7thoBqSq61h9tTK97f1BIm21cRUJpBpwmPePRFutvQC4C+
USU7y5ve4jLpbEG/yG6RRdQaBXSZ00A1+ZyavClJQZde10v/RpxevgzJs6h9P16S
fU1fzJ05I8kH8WgahDKbgqUzhg02ES/wqk88UbSJwE6h1v2ctHdaQjDpmrNRaShg
3yzmFAziBgoehrniaKIYvl16U4qvXnPBPdrFh2p54Ntm/k45eQpX8UCxGWbZS7K+
77k89Quk1Bdwb2C5ooCeOAcj/QWXCuav5bjo5aNu1OSukGchmghG5okbUVcBrAua
1tur7YFfKM4z/KnMwu526rfX2RA3O1+GRzCcdgDxXsZaXXYVCc3zBnbt9MI3jdzO
Uhl0A3aXDXIFGjJbP8aG17Ic0YYnlXzbCNWI7cy4d48LEuknKUARAgd5OIczpj+r
MZHi4DoqM6OwFGMaknu4DcTh5dLzOTjZsF8L4uwBSH4f6doAgONYU6BxrLGZgJjX
bExYM6Aaw3i/qGJY5rR43oEyn/Rpt8ZW1obmVBvqKIQNdx/wqz1AQP8I4KtpXa8c
lNapEteQPIA2GtoCuepERF/IEwU5ZJGGHqjga0uWx4YI7rRbVlMxJhi9a+De5f/B
Z6bFZ4yWUdToSIyRBu6OfNeuc7Mw1Zqv7yuxZrMEJoNlmEMIZuklJb51G0mpXJof
QK4CmkoW2C8DfewVjCFz61LUgma15uAwH2ZxfloWKuIeEiFA0sSGDeDzyb/nq8kV
Ye7f49RTpVJGSg2BACt57HgjUBA1+uYIfvGa7jRDGBdxEsb2DK25uA20xdv1NCaP
YxMI4qR7p3IY9AejKh8YfJF1myktzAF5fMp522AxT7Ra0h9pE1h4YtNG4mfvuqKx
MWAU3kYRXt/FMmzL3oU9dXc/ZpeLI/NSZ1LPN0yfSObJPLJg/aVrR3uSloLLVrlv
fDDJ4Vi2p0ts4LeA7VPkE8xq8//533w9ibki90kZDiojx4Nw+QSa5xc6ixPOsPW4
ZzQ1giRXpIh2duIeXdKwMP+OtAOMQ4j92NyIoRgH7vtCaEKOpWk71NC6GqsFZa1T
qJ6KobrU/gKp0BW1BvUyMEdVrEcAPGXIImKGMpOBNDciTTdG4EQRrgmBN6wc/nIr
SqiqTrrIST+ssvB+fZaXjPmBWmPLgE/J3Arpb8j2cZZIoMS4uD+wKGlaGWEEekh8
Mnra7ggMuLPpqdCvOaBPtBph47PuHWHmCjRC2Ztq4ii8AiIuIIk3M+3lESi/AR1/
zcMtfeDHfyoMYxTmOLLGATMKkCu4BOpkv6BlRndtjQvzbpU8swmEo66CQvAG4ira
3+s4pOOpPRwVlWKNwDMbbu4XaAa5ETomVx+7IkL+qkYhHxsq0X+qLsRim5KALaWm
WBU6FXKi8HYVXXIaz97OfSgWFWrIvCV5QBR+KUk7YCaISfC9skgfBWAcYb0ul2jZ
Z29UaqOtIsJexnDJ2W9B3m61pCsM3fzIutPyWTE1d4BUg5IjtPqs6ekr49BIb3Bj
gW7ut5JMbgyA+5rPb6TH/dcFZNGcey5P/LsfH2t7Hx3s19dl/TZg+YtxKT4zycY1
YnRxlgknAqVQaJSQbYvtYSlKrWobqqBdvUxLPrzVlWjVr3uKR0rcOPIeH7775fiu
NrVoc/SRSB1I2RoifQoGfafm6mT6zNfVsiE5/AFRqKM0FDXKK54pIAsh6CmWVDp2
EmLpoI2JH3i6D/678X9lNd6HDnRKB0qZhox7m/CteOMn4JJ298lt/R0HPrcqChKV
SQR41QClEVhx/ZBqYXRGS+bvLyXwuQ2bjmoiOxp3aXVO8GFH/Z5Ex7jgjVrPeken
kvnHQG/wI+ZvzLnrWjnubdSKZ0habLlAKuJKLzMkQBMhmqBL3cuGJOIUGLU2FaCz
OVYARCdESeukZWsO7G7PsFFmweomjlmRZZaTFJb62CI4AcxgFKzESyW9j/Krvurn
btT1xFUJkZwYkRqw2z3VPXMh03f5I1qYtDRKzOLDWf366qQQ0oDUIWFtQ2noBpvs
NgEK8pZ7N5AoQPk0aA6MUHTkDmhuMods2Dzm7zItZCrhx2nOCC9O+h9Biei5tjxv
q/zw77UUDYCnSlXTo033/jLvjlgCqYWbW14zYRr6+4sVBgwwd5/mFeBC5o7wtA1q
sbWO9SxHDRYaSEau+8Lh23fiTd3Sbt9oZlsQm+cfm2oG+2tjhwuXSXTiQyqgxuol
PV9o0cQFdLfWWGkrtpQGQyX40r94F8ZYvZZY9EyoC/dHr5FlW+fMpjen64nu/REs
6msRDjghxIWZfC95RjTCEwr9rjdYZgHs+3ZfoCCdrL7lB6bM0Qh2WfpkEcQClj8g
crjBZG4zARAABugT3CSVzdpSoGAq7g4JG8JaNAnBXg2SP4yjRazBM+uNbMYY/CP/
BRylYYYitPD+8eqcABKpnF5C4o2M282nJhjkPaRd1Zyv2X1UWDKPd5RUq6ikp76X
HEPR0FJd8RJZe38odomcW/aRJsNlIlOTV5/f5+rHrdE33zQ7rgFnGETRnEj0gEgP
6y2z0cCMeif2p2Lz36oGmwQkNiBGHdUcsonWhJvn47P3XyFlWl4ybHDmBU2jDpzS
i/0WMbfcme9446gcO3KVnsDAAWEZxBzdc+X4Is6YGMf92V/4nnQcx686UmqLBxYV
gZT8dlhRQ3X3Q+PhlQWUHoGYTWFdPSbb2KDquynTj558NJHGW0R2dBnTRDZlMDoy
B7R96ZJkPihks5lmVd91vfNW3skG4baZ4QFqov/AhnfGNTpzUgu5TFM86CPdz25s
JZLoL8GN3/LwEbU5hmpwD/jowpNJ/yh3ZFvqhjHDDpcxYUPosnG/VEgA5OzQCIpO
dXZYYNWKpylmZcdh3OODvG2Ram1K5ub12/vlUqDUMK9B58NayLtczlzEnTForrGR
4C6VKr0p8W2sse0EOFm8pbG6KZYgrqIF61wb/3o3enxYwUAyk2B0faSO+vMmv1cb
mLcntAiGIvNoBkNFFjfjIRKfnHagLGoMpa77K4EnO5+CkNdbrZP86uciTGJqRXiT
89vlg0j8ItsfXu5vhC8A3OdczsKb6vOTG1VTaYG/PMGEDahPlWp1aZJtioYiALiG
tKCLkWDKa3QWwr1REo8DmJ4XATxEf6flUXttTfu6eVPrCxefHXWgLs9QonxxLFm+
fHDLORl/1fjQVx6f+T+7MNjd1lHCDV91OUpWYLALyshvZHNluNrW3Ht2sIWwqrhl
SX8+oNyRmzT8P8NSfc42sbVXva2jboswexzFHNM1yFAnIEesluacPJNuUnUOG5DP
7gqBQXqTMvgp4eAmLA9ahWWHn5fEh61uu9Sr+qNABjjnj+OichP5OoSfWQXnO7iw
pMq04k4OU31JMIDcCc4AdE4WIfnqAG3zbeCjZiHqBeR6wpohrCAYuJC7degcz3t5
V4K9CAOc5dZjCkFxjtDRALdXGxnljAcgEd03oB+Uq+HEqgoL0Z+SKyXELX1XoFLC
TMi6YHn3Jx+Mb5uwRHGs8WT8oKu4iQoobLGCf6bPSQ1zvzDUgA97AukOt4Bzi/oR
x2YgCJgtGTqUpQ8yoC3zJLv97SwmpvoJbl4dFa9WiQh+jOOCkwtONJ1StYl5hNYH
vPUzK6HEPk8zzLLTCbEVixsLb7gg3I8HGjxQEZCZ3Di1c86D0GQaDWkj3JtVRipC
wEzcEJgfMoTM1l1iSRTT1BdDqXxL+jzm2lMNkWdLdE9E7ZiN9BhGOYCo1pxrE1nd
MtP9FMpdFsSpn0aVfEXBM5S2bXzBFOsnBxCNML5lMdoCx9eMmwRD36hFY+QVMQUe
YvlU1iRgfXwzAb4xIVfS2m8BpsJpL0tgoU8t8R1UKRcHD9IXdkJ6DIGKnwF4wFGj
WapPT+LhxvNkPqicOnwA2oNLYOBs3BdKE8DiMxG7ZlPWVoKID7gKN+LqDrMbwLmN
3IA3JoCM90iwSqEcU+7lI9Pe1WCa7xKtcoNC4LQpU2Nrve7pAl1RYzzfSz2bLI0z
IJEo5Sle/zWSCKrcBx1ffh630F0qOQUFcP/I2j1n+g8brSO3ZcOpTb3UfUyKUEHU
ExL1RqSJLuiRuOxNXKe5B3VZQM25fjyPOy08DBYjF6oQ7cQdp2Vr6ZntUN0PnuQl
YpY7p07g5WSvk6K7jzE6nY7SHICjX2yfdH6gYUWyJgqES3jTizfjHds4J8IYRYBL
e2fVSBdoscrD0mm9xYt8jxiJ+4op3+coSL8ITv1afvv/uQsqWIOdIS1niK6mio1L
NM/cV0tEpmcS6VfNpJYFzHXoDquBB21G0dTXuuW6ZOtIEEXaAVR3+Xlq8NBRUKxO
x2h+FEsRC3xWGWZ5YkGJ5gS4WorsfQ2DRLYnVE/hne5VDFfeWw0k4rFzdiWKviaZ
mj7r4x+TwCOzYe/b3K6d7B1+9rDnYju1QdbEOdbAUMdvRqTEjGs+1bq66R2gtGrg
iPqppaN1OVA0lD7hmrK7ASce03fE64qMUOBKxyw1mDv2rx0ZUh/ZcZVgutW77UwO
4JwfscmnXFJxEH9eWvhraMNeMtT9wEiR/aoF8kB45KhbW5e3jsWZm8uvskFJnCuy
WD2FVdN7JOEi7cwNjC6b4Nb6ESz/Qs28CZfoSpdBogSMqtZkc9qCSQ5e906v39cs
NDpuXZ2oN2djJTLv/Zq9lhtPncsTde0Nva8jpS4hE74c1zSZetBdCcdOppGQhU5T
UORyf5BdGnmsKE9svQD2N38DqOF9B1+Ktn40KYJiY90JXFRiypAo4XcFy5FyL0Er
/xqgfXItDIfTgLhCS+b086SXJb8gYre5tsmJYI7RBIxtLh6WeR125i27lJPurgNN
x+SHkvUn+if+Mq3liHT35pW2qOHJzzw21BpqXjAJ0SSihPdnRrsH0fZng6b2gsJq
1T7vdGxF85uJqRMVTffBRabBwHYn5QfK3NVAW+99xmKrjmdk1dICYq69q6Aq2cgk
bpGLVRdWLVt1Y7MMPwZ8uVwj10mOGta6G4OBY4XkZx2OlLQPwKOmLYLZXkyc+I1d
+RwtxjH7cqNx5xh4W0n4VpFyUfo8xIrE5NDHF+6AR+bgUHpl3x7Jz4492vtUK+o7
5E1tJwb3/Ys1tpl/8wz5hOid2eY+K1hGnsQm80YlveTZIT5WzHBRX04L/j1hBkyF
PFmFSPuNEN1wE3gmEz42K0ImqfXXPWFzy2QaNQynuu4MWICAFJdiLWRgbkExuJvx
n+fFl9iO2KKZYJNVICKGxIgyjgPx1Sa5OfTL5zTT054aIDHQyzHkVcldemJtDihg
iTjCnsMGHI2PhWv6tmAcnra48kX1/tzo4XRekmmbdZpzfYzA7/8Ao2bdghiN14I6
zuWD0szmjlRSHVlq0GDae7NmyI3eLakg2GCt8rjZ5gvM4wM0fEM4zYaJSob0XBYS
RYrz+VNlI6iIurdb/R+KA1onvtFnVDP40+A+hAjK+AoRcuFsJSHOjqgZvOzoBPdf
kc55bbWZ/ZSUW2eQukzhakbcHfDgQIqdEwF11915Rkzs1viHCYqOYiuPDxM9w6gG
bKjD2XNvUaRi1+8RSiI4Zb+t/mZ4F3ILfWQpYal0irzvnlJGJ6EeLMC7Oco78Biw
z1YuSV0kS+kVT+FGv9jT9z19f6pRV9ocNy/rRTh0/+5VYw4yEitF3CAFIMUArlzE
qYCtoTZrjWDTuae80YziVHx8v6P6720MArNRCro4jyEGG9srF/dkRKxjtScmDzzp
OcPBrgvR/4hKLTmIC0qBb9K6TtMACRR1UGsemypOzuRs+/06peSZabyiMZZsJjA7
AYWNkMaieUead0x+dnWjGvTcoKS/U3tEfOnf91V2+CrEhJK4NPeAL4ot+KKLwjTV
A460PdqfmRfWmJw/5FsmUkUqPqObQI0MLYyujlmdi7j0u8+t5AzbOl55hVlzIWvR
HD5g9iQm7wUvYJ23sPo1YwQfa3DyJSd+Kcm0qnDLnqouQ4uuSI8ZP+YzDn8hyPRz
y9ZdxQQlgRqGjXBjqKWrI5OLK22D2DzQRhjiq74qmm/F/CZKgQ+PNC4zw2YqLyRg
wDEbWrUgglODUbXIAH++Kfi8a5q5MDSRT/4bZgWW6JNGgVf0VpYgBiMeBeWN8QDs
34WSgch/bvYS7LV1nwjxW8TpC7bh0WJnvpGEVVnhFJjqrgWlxELNxzVDUPBwWIpr
BENTy3QxObqd1I4LEob61vn7KLB72NpjHLStxS3brHTQxZrrGfjZrnHp0+o+jckl
7pM66lS5l3Urhy1w3JxDAvYNCu3EZHq8VyQpe8CDDFL1DWwpC0j78k0Dqyz+WpvH
K59INZOyF0RhNS8Vj0eSzS71wJE00qv/SiK9gJ18+g/eA3R7Z1ZDJRpSGLhbiMOB
rZu0eO7B3LkOAJgzfeqPYBwMvt+LII6pSjOeLhlvAXj+abXmyfHAKWNnoE0bIR2V
fJ6elNPqq8xfpiE1oWvrPYFsjLu89bgA+6ZMytvZXuNzAVsdaVeMKbFTQaqR2GNT
mrg9vNrPZXkqXuCO1X/BihLRftBU+IUK/bqk66vlNG0IDSqMReaSdgYFuXGC+Cee
m11BnRT/Z0SqZeKs1M586M8LpTwek4sk1Y5jcbjKsO48kweX4BpKs3tB0KMdIKrj
onXCs7zBa1JXBt0oy+Xq+8tXMUqQfPuYd56k04awHKF7XiR3Bhy7SM/Rbxd/TmUE
JzaQNEzpr+jh7XFTrCwTFEW5y31wnklEMolvVOStXVJ5Y3BNy62/ABzulh/Xsc7t
KeVA7IMXWlIm0gaeH2rpkECJuJ0WsTYrL1Y3YdKBSDGVZa2qpLAlLfmr5sxQ+9Ax
KGwwT7Q+J+hlwifAlh/eSxANu3P0ot1yNuvtVG0SxMFaAaWKJ3BdZExr50ZppIfr
VjGtthqBRqMUX/af/lpox+A+t5g1Cul5QxNlFaa1Lv73OWvZ1yfgcKpSNZ2N9TeX
8Hzk5LkfjIi2hoCYXOarJfy+HEzU+yYCgOJm5R4lzajKad0hqDrFXoFFOD3nHWIj
erCgikItVSjzzwWR/kdGvClKgv2Izi+IDzNx7nchRoR+IpKLf8muLWPRAnE6Jh6y
nsP6RCf7E2N3jfuaIRJxQhtEHtJXEH0mbnpL0fU42joK1OfXgPxFHc0n32lJUuCz
d+XIizGxOtsev2t3BBzmHuHnrxISmv87eU2hH3oQpZWDNBQXpcXGVb0n9iS2nLpk
W0T15bUcHSFoA/Fc5k+AAhQNaF8B6Fg/NdjTK74BZ9uZaJWUty0lVM5iliFoyR7h
rK6q1taLBDRKampSc+9e6ZVKgf9Z5qoNTOaNmMNC9kPTzh2G2AmwMAiA1Lehi5b5
Tf2kZDmmWbpuuRA+P9eUt1CYD1GxmC/j//GdEiFlC9VWTf05iw0wrrB/k+bRiiCh
73oHXLd21rcN5jSXVRNcgDXUQXi25B8cSyHE0Q6vB9Ux4Hrcu9kj+/NH4Ly2ZcTS
Ex8Fj6tH7dPzcZXX3eXbCBAdnCzqb2u7pZd/WHqB3NNV5fb/1qTV2QhajtEGimlo
JBalimmpSfpanEs9TIHyoIrRsOepFwHL49ZKtgI4DeJA6NRzMpAGxYYl4/bye54j
L9TycVj07DgeWMbis7muU3oRmLPkwBCfRUW+QCWEuVvBivx2XvzCpOrWhVHkM+Ui
Dk62MYDtpSHIUFFX4/Dbh75njaAOs0PfQebH+lm6Bm27UF7Dr1suIPqD5tZSpdln
z/hNsgxDBXJVv7RXtx/OPXdc/whY+ywCmNSnaEvsylsjzFVmOWccG4T8aRxgzSKD
Y9RVwrkLOEhBV0y4D2+8+3Sd1ND3ONxkijk4+sJB+4YkGgo/ok61BpXx3C9y2hwW
tjjchAffVVMUNFluyj7JTn89x2OKR68OHVOr3UBikGFaLh927Q4owBKw/CLKcTiP
sg1VjQrhedmyYwGVKRXOxDKV9yVT4uKfmLFWmf9dDsO86TzT8vJZCMHKFJKa4qYw
P/eLyrvXSr38EC43rPtTM4E/Lvdr4V67RIq72mD54L4JWmP03IE/FdL9niTitrhk
CbL647x+0No/fF175BssrzTbaf22Y5VRCNr+AAvuB3yk2H/QH0imAsY7jghfDZ5m
hpdGqeokyFBB1cH+o1A+2CPiyzEe//iyBplpcC1Y+wLG499TXmoF3CiFgFhrtTU5
YM2AMMJA+aeHYuLuaRJ247McU+S0GJOo1+0O7UYV8Uo0I3JCIj7AR9ZQz9UBkZRv
hyZuF3GdP5IKkq+dUDlyXBB9GTIULR7OOWsMDizHThyUjr+4al+JEVKZeely3BgD
ypk56e21h2l1FZ5BARud83MMRflYh88yGYsbjItOLZ6rPg0VQi07DgJtcDdzdcCW
v1e/Mfzj09sfU0iBiEE8W1937qqX0LpDUR0+5eefb6R4U2XbDThyu0wmUpLLr/+U
yYNqkeEWurovYzJdCQ53HjVsYZXo+FCLYqtr0g+F4aU65Xf7oB8Q+s4ur2afC+Cm
goa6z+jVe+EVuiF967JBb3PNMnJ/9T2blI+qoSDQDJon6ggwEhL/foUYRb/0Hr4h
w4txr+D5cRE0EQDgPdneQQiMDhPbVXsSVy6J5VRELVT/xDm2Lhe9FkN+9zwbblUT
chG4avkXt9CiYFZtjb0drreC7J3KChKd0c7NgZJCk12QIgOEi+Fv4QCNh8NXJ/0r
O2byuskjQXwTx/aw0Z6o5ZQ4R4jl572A3ag7G4JeqTHqXOKfgbRO5gu757iKtWZH
VveepcBWA1Aeo8d22EOxYdQ/ZRPLmxXGvao7nb6DmZBxkH9h5DbWsUWTaQbHRTih
cnp+SbXfznQUUl3c8p9BGhyks/wpEGQVuiaGGcBQDE1IK6ZeTb2t5emFAOl65llq
nBAxWaId/jp2ysFDNrHwHwxIhorCJ/mpbZ3mVeE+lIM8dhlUngbdL3t5Dq/Q1s8U
Xo0D5ygT1exMyEZa6vxvyv4TnLSicO1sVR4zyFUAt/tgFddviNCR+QRJq6d+k0nu
iGMCVL/KSN6AKv8nQB8cmo80oU2oJVFQlp0oDnANAuqXE9Y9XHvxm/W7WARgNKVc
VGMW37gNfNvReHq8sIejpZXUoGCwC6h+Ea48b4oqXKg6ezd0jzVfZsWql1BEzotp
z8+StKLXiCJRIEzrhb4hhRWygksldpnuaTSWR7lIleYyjgRZPhqljCu2tonuVko6
38HgHEDZhfebwKZ5D0hX/q8zoYomwPR/o/KUQlt4+IIJLIV3aVWxYXGavKl8Biph
CSrOzQYzpoY3zo+6KroKB+WjszHOGS96k1x+ZBM910j/F0QSs0w3yaPT75THye/C
2EgbCklkuetBiW6IOrWXQPRIGR8guT6qtrHEJBVX+suzfibcrfjZ/GjdtgASeOjo
GAkqo2esE3YZCH7t4Hkyc2kC1afXRkHup4k0j1PMzzKLetxPNJ04jxwwA152BWXJ
1QD5pNWhxz4bkL/mipDDljgZ7e7qlANJzds41eNXwKX8WTZUgEIGYl+kAYLLq2CY
MiewxIajbq02uAYE7/RsbbLTvQUqnD9WaK5f5Cl7QPv0YZSh5SW3zzm/Ws1NOKm6
7X5c5ITw8jRE0b4wocqMeEj9yMQ3TDhzsOitWeONQt+/Vmf37uLkUmKID1sSrbvj
25Tf0cwV+y8l6SpHcDWt67KlEOXneb6GqoRjITzvMs+wPq2s/FSzfbgNWVkSXD4T
79Z5U7a5LVHFaMgAwd+Z6i7qSRUlZ6K1Pilw8Krdg6AxKcvTVoAK7s3Xgt1KHQUO
c8SSvvAeYcVmvm7CWQr1aA29on/GoaecqComspiYCGIGXVv9uTlRj4Xupdu9kQ+8
shI9mLRTFX7jhgVD972g1fKwlSowLUXaqR9cYo3JhyUZOcE1Q/u5bV9QrIhcJ/rL
1ICeIFUDxGQ9kg8blHIhZlOYCMf70dzDbPfdGTpiby12PSN6EBgtyQwFZjbHDVei
9aQhUgUeettDQM+MB1qyCRksF5XMO7cYfvIMa4/GpZi+DmZqUeAZi2YbtxrrzsJI
7WKGJFx28mQgFvQd2qdUycRvsM8K1WzTFB1z+SjBC45iRHsEMtf+kIwXMOi+VCV5
1yolNrZ3f+Xz8JLdsp1OR2b3SRx9FUqTfm/In2dmpSwYRwe9U7/mydxQyHG4jW9l
U7iLFrmcWB5Sz6WKybOgsPSc4SH0zqZAYCwrHmjL5pp3OpYFT1xSw7TDi/1Ga0P5
X06jgbFsOIl+naHTKaYhfY5nHTOcpAlLCdUuEmQDRggfVdyjOBOTPK+gP5/0Kukk
3YFp0YM3HG4PrVUXEWjxAhEEABdzie7LMV9dkzQzNf607Rf46xcphKdQT0Tqi5wE
zd9PQR5ALL7aPd7KvxSVv5ZEfyCc3E5/8zQbYFwvMAt3X2Ytwbz1u+gaZfhILjR0
0tb8tvZdF0YiL/33KhKqAjuFXOdK3fbxFeCu/KsXsBdTv0DJ1hIoBk2+8vzaDGgj
0NNSbK9XKuWGZ0CeG9Bf529U3RO9aFOkk6g962Et3g3ZA0jEYGX4cab5XhriUn/t
AJ85PdyXwB9pR9Dm5Qt/LQBTkxqjP1lxKfgtQy5gVyugOgW3RaTfLuO9OSeqQzi5
CP0omdWEThGBtP44vESS7+lntaBIqNi8uwJI51cS4r2HPo5Tf3Zgs3WULL5zWaJd
iKdzLOIH7D1QEg4iAMb/+qIEEEXC2JdeO05n84WYIvb4XaELixKnPx3+uG5Vpp9x
8f8VPWzeI6rKGp6yqY4uCkJJlBvzb08KfSGl353gxbHLFy2Ex8sE0IQ7frca32PO
yOHLJbA3Ww3pcnZCTdKwQU624+Qm6vk2cTk3pSWkgPGZxkiw4FlQRqpTOYtiUGn8
fR/Ie+zkTDZtuK9u5F2uKVgM2Y0n6ZJA1wIFShArHJfJZBRxIOUpfRBSn98pPKeX
NdSHSxJ1tgC+ICMJaAJv58hGnD+8RPuWsTTEPEHk9DiKsUSqNPlM8QpW257xhtR6
89pcBiZ4ftlnfd5VZK8719sC9/r8aR9mAJ/2tn1GlKYNm1N4wqnVClW+cU3IOGW6
gS95u2hcUYMcNPTN4m0AsDoOBYJP2StBUTcajZRim3UddQaT4QqodGIAE8SZLLVY
UKrJ2tJX32BRhV2T9ctUEjTAJwczLQ1vs7vsGreRVkgG7dlSa2wHrf5MTY/PXayQ
cm/JXPZcKFVuRjnvwXHYCK5U+TdcDxMewwGNXwtNWOoQxTA5ZzmWe56t/8yOBbMc
2htJVOqTHXmlTlVCs0rvRe0ORuUOCqVSm+d4yPX/ay/foasF9T1FQDKmhSDkQUWX
MRq+4qDgrv83eAWzjBsSr6SK2QBt5AVVsz3RuLLOk8eKz73a1ZyAuZZ7gc6UbWQV
SrOScIbf4uex0p+pDFzxQ1EPha0b7l89OLJjSeRuJcLjMiP9rbIakit3IIlWKIPo
5sY3v88Nt5kUZzNO3FxdGc3bBl7JrxfLxrkyvX1wCaryS2GPhb0LFHazGxqRbTfv
VH4SGEgZ9yDEaizmJtPkT6neYzhVenntQ6X69P2LVJWw5SXzlckjUhbWOsVqCsRf
LdjdW9Z9N+Q2IADeUHcj2XgmIXcb2uBUy+uFxqgVoac2OJfnuF1YbXM0Ku+YsAiY
av2fHKJHOhRVREm1cYhxE5HRX9bSQ38mnZ2Z9ObImKSAuj9Ze4ZeY8l6m8YeEhBP
GBYwJlmQaaRI1mbhx+MsZFZ7UkpWPK5zQRanC59WmLmmqXcGmfIdJevaOiye+rG2
Hz/rY6DO/QkaCFNAWPkRnF6oG+WavoD2oqwriztX9YUkjlpIfNTxRzbmTAk/4Bkf
44KWMZJinOSQfEsC7of83FgqtSLXsw0gXDCkWD813oRuk42uGlBbhJPztNAY2qMy
iPYNvj6zciiUiorO5fE6xxevS8voDUM/jzkycQAFaTF+2rOnvb647mbrKeZtognE
Y+xLMS51LCPlCAMVjkZx+zeo10+4k/6hFS4o0H/tt7QhZWd1pDzYpgyCC3m2B8bC
tbHtRKgyRifouCjvtLndlqkXsN8GCjfepCqaGECBm4ZetOQG4DouLkh/OhAKxTOg
NuY25QzC25w43ZA1alNWYaWZc+0hSJlkKdC0fThs0UeURxZ6rfwlDlY2DIqaBHjH
jaqKhER7Uqt+452mEwQHu0ZaKW7OdYODGfMLe/5qMQ1AMihLKK55kk3WhQ4QpSlE
WcZOSjEuSDaUXeEbZJM6EaAPkc2LDgpBT+jqp1CrNzUZiDRurEmOP8uJVL4DuHdF
g5zL0m7AD1ntUo1Ma7cv1JbFbfU7ctFDgEj76gufQVrt1Quz6cwG7ol5MhjsqNca
19vXbAKgjxj1OPWFFEPYcYmt0TSHnyskTgHEROIIaDZJvtDKQLNyf8pMyzyqER8c
dgs2Rm6c8r9Fa9DYfnm3WM5K75VUWLv6b3m7fh+2c2htF6uYrhVaA/hrjpThtg3v
o8ZbkqOXrF1/oXAc+iiDLfDGyvl6KkOitWi46rPZCRGJjkiS0SkhcNn2HKZXuY+M
sYcrCWZkYWM3Vr0AR/MFbj0i1NlYWh2NsNrgtToy7Dl18xg3KD3Hgf5WsYpZbtZu
uO2YnJhCe9eqEjDxuJsdS0Xt3GGIuFurpprfjY+3tJxNehSbmLvS8CwNjy3p3FWB
ySSquVyDg1NdgYY2s9ZUQ9SwW1vxtARJuX+PSaXeQ5GolJsxb8/UEhbnPPwQdLjh
sdLK2mxJPUJIMp51NnOrBMLprLXUr6AiKsWktOU30KcWZwfOYmIAiJE5eUK0DKdg
VDV5SZaR/oMg66CebWNNKH1PBRSeZPwDwfhLVdTVe6jEaIxI6+HH1Mg9Brb/Jsy8
d+qUcpDXaZGU5Kfkns9BngRbIdw2u8GgdBEmf2R69ExLvivWqrQ2qz7GZrW1AvQT
xENMXXvjOXL0kQlpiSi1dnWIW5AX4Vji52EdrgoQb4D84XLyBwq7hJn6zO0O/M3i
43BwMd+YIPhHinM0/YtShq6d79pYD9uNPyfg17nxPCdZGhyBRwAIhQlgVo+VktG0
OKPBqLRV3bq/LNRsZGdmCMmnL2IVh4/k/2rZngBaZ/t3N+hMtbAzBiee4sTetaTx
FIiV7V0RiESHrlUmP+seNFXTa7m9xm2OpV3k0icPU5YPwfF0MIWQPTNQB0WAkfwk
V2IzuwoIvpyX2hLxABe5GMW2+8BPHUsmdAUplM+L/n9R2pbfrWP+fX2+czI+xvgL
1ycAw6tYo3EzrCmWqLRxemw/sDKL9IxOEkNhLNNeK+Kj5OZAjOCEAhb+udp8WrFD
PQm8EcsFXHWmGYVURHFUUCX9ezTpOO7cOylAxlle4bCZDv09GaZtQh2Bw4lVCqll
P62P+Mh3mMID7yEu0XWqpAmKvr17LjMdDLjuX1vFWxrLFleBAY+3bQB2Z4I33ElZ
ikonYYZV3PVz+Rlsz6H4StUwIGAJ7XlBqosewgE2B1ZT58O7iUdYdcMKkFOJXq1r
KE2H2Cltu4xLlF/5JTkCTJpTdmKrTbEwN1J/0DPtHtcN6ezxzL2ON2JtdzEPxpYP
bu5NKye0+ly95IiMludddmm58FMZ4tf8Bs35SSZFiKuJnJgq+QRy/hkjxcoiHYli
MihfLDPWzYjor4jKjyJIX8fbqOA7F6Y6fGLpjiQfqhEKdx1oKlJHJ18NpuxFFCGz
cm8k4SfD+OVevRxkexPzlqf79W0Ns7bm2nzSa9aO3nJHjh+gbnL2eXx8ZVAioZw/
6HANl7Xu0Cb0V6y/yQ5WQ7dRex97CP1SAmeYcssl7AL/462kMoDGj8/lEHGpJ3dU
uAVFB+9VvW+KUi96lO8q6IqcsApGqY3GqiuEIk46m3XbOCj1secI13CM+rTRfUvM
UAOfMyGYqrZyyMBIB+cA7B1MePFam2AKms03hyNOCLcEwbn7til2QRnW39nVfZBz
dLShPh3f4kvXmU/fjLmvV0yRGdGckA95MDHjtq1XFo7kAgcNr3mrAOLQHQ4H+5nt
84v3BLWN8EaFyTiWrYg3ZklQyI+9JHEVrivp2z134Dn2yx8gHQzOBmCQNl300T5d
XHOdnEJJYbX0j//FFzfnZy/GU63F4G3BuELIKfELVGarTJyYSKuvFfZU159Lmyck
rfdfxWyt3gd7RKzR5VHUv4taOLMrrVpAT8iv2PNncMqxC0EKIIOKpr6/u9eIqjRB
sUia20lc82UyxLuyTkWDOmUkcuiuJGDskPAVZKbUYD+HLbl6d+fMSkkXI9T1rVo4
nPF8Ee4MybztWa2A2K+UIMkE1YDcmOjWHjf/GTHjiKX46jTMiKSrJZy38X8magdc
0hrAbJrit7vhK1w5iPB0YYQHvmE3ezMkSbpvpPBhDtiyHVkiJsqtn+z5aEAQk0ZQ
vE6kQpZ43C8gD/dno39+9CLkay5cWG7qfd9s0SyJ0krrHlpC86kkLvowTFjXXMRY
+Mm8tSu4Mvj4dzAwGxGksUR4oQqIf+K7fDEIOYCsPweypAb2ghUYvaoKTClycmIn
KIpj0iK0glmlAWKLE/tXu5vXn6L4px3wVCRiKb8FIQmPVXyL0lvlddl3e7bjjgqn
7Ve5dbwADuTr9Yre7a7EiT1GMNwmClfsJ2+Ghi09GT8j5D/dVqSUXbbTq/k1Iz/m
SmJC2VsGqDGKYD9MqAviwq4W4cMw7ZJKoYonbc8+opSFltZEFkNkIVWkB3zPNjBV
CySjZKDlKm/Tv9gzX6VtymEEHFYQDlSUUaqRulf7azrINX8GmfdmNC8WMkjXfR/r
zEv2OmFgcireDbYWcxvH1aRkqGbswTAp5C+e4CODWWOeOdM0QS6hKPt2I/4DQdKu
NoOl1kVuAZ2BWLjYUWxf3XXBm3cvnLQviDlCuCwXLZF/7ZhrhBerikhHU6gcTdrR
rQeauHNxBTjkn+9ivmHoHHTcIV8YM6Fz/5842sF1aQiOnrBQQPcyPIkmr9cANoSX
Xwh/VAEPZwYNRIdSzNU87V7oqMrHPdDjheewoU8CqOb1Y6f4rNb3JSZVrEekxRBA
wf1k8efyzT2CA7Bf3s/BcRFYe077r99ZPyxcJ78zK5IBT1PBXj3BG7HHOs5F5gvF
P1Txaf6a6xOVKgmv9TQpthKMUuemr/bDNrM86MZBALjgRSxQIABwXPJWczR6C20y
toZeTmM6sVDffZSVkPNXkopM1wj6z5n6v++EnYOkW+UmyCfCN/k6OH5IWuQjqSgg
A3K2DjqatUvQjTFrJFg4xYpD29DIvsrYsmWWGZDcLFYEpNKpIn2NZ/jYbsVhCH4M
Btxt1PXTIRqcUIUZTQQP5gcNxsbNrhF0p8Gb0v2PEjIK10K+vwGq2hNrv/VwHgk1
lh4pBg/AJDPVEO7pmpH4ZZEp5jsnV1wiUgvOgtFRHgCRsr2+YPRuTF2s5KAQHWd2
+OZMUVbgzRfl+9bbeGdFVyQwOqzsZ+tehnuOu7AP4buSgvF/QUd7asLN/VQ08gut
fugRSQFc3ANjO31h4svGdekR+RaMs43ylixmmxcWOtyUez3Y8TtGLPl7ML1TDib+
0Z1ecC1atdCK4z2ZsA9erMoVTOttuk7twMhTXoMpRBvYbBf9Zdci1oJLiJKBDiL+
o/UtebF5KDCBQ8ZuoxMjSeuF0fhF2FewBi7wqztPW27jRiUr8mx7UIV45fYFDPO5
tQhyedN3qii8brtS74LvMFLWRcWcpBw9lXjislwE6TeDIe4epVg1ITfHaAKhNWSI
4iEIPRUV5hcsWE1UKdnSJ6yRuflu6tqrYdEcxT5gwlA+wvrSEKeCWgsivdUkiDuf
fk+DCq7dV/y4YQK0g+0NGhugRvXWkX/bVwF0PLQnK0UNkC5/O/7VvdfbmP1bH4/T
Swa2y19j1/h5Ys9zmyj9CNly8kf0s90uVmxlfc1KHYudkrIgoGFS/XGCxKJBRSo+
L9uxBcx8ZTaghbXhgpb/mn8P3fbIwQ8sDhTIlg5+L0lE0eqTnnEg77c0iz3fq7Pj
vVFGSai3HsW5D4/cjDp8znN2UvJKc9P3cIOhzBSPmdHF98G0/pRUI3aBqorLy5Cd
o/5hYD0a64sqRihWBA2nqRfCvw5bt+6YXE5mVFCevlPykpMIdMFtNcVVyg8pexAO
mktVakPTAFOalUGnI+FEEDPHbp9UZ3Kd1qZ8BYGXmxZLf4R9sdqVHKADd8i1T+pR
oaod9rTGRvR9UfGfUFnu796V2VzHND6Op3MwLQ58J1Sdj6PKbf1dm36uByDUeXO+
74RY3nP6ntitGiHJSw8XirLTesp0Yfwidr8BFFXl8toNUu1YHbiAPD2PBtXKv4HZ
4oG864MWv0//1e1KJQFWqnZH1kmxMkCT2eKgQbzAjbGyU0/X/LObKgYMnu58sumM
Z2nI7zTYcG+SgYGJ/uFe/E4f3dzgNS1jjN8SaJfzJK4lR9h4ib06ZDZHJUbnB8zr
xsPCAv9USH9bRDd5bRl852cH2+5yh/J19XeNo+DIVVsL3Kzy8pdNzaFjW7VC81an
uZOH6lnsOVwpuRuVnFtd1Lq1BP+bVEliZPcJ4JYBNSpIK7fKNr+GBkz82cROk/O7
msqQroPIxWLsMt22I1tk299vQYLu/2l0MI6Dm8fF0vG0V2UUqXrgwgOKEgrvqdum
+X5lcyDOCbLdbTsFL7Ct4QCRLwL+o6JRqRNWlnrsYDO3KuAxX/UMyHkERT7I8SAQ
JM0+YrmIi4nCHhw+ke2MdnLoJpjQFx8gXDQYPVmNDdMiW5CgIlyM++/2+RzPPqy0
8tr5K5+CaiG9688fgeOQ2IJBq3EwT4zV44byOF1o7ZqgYf8dBY+DdQksxUGTgU2R
7O2hyP4R2qOV54XRfvReE8UsxuOpR/0MSeGqpcCH7NrKIF8d9ObjvyHdYgjbtrec
Lip6Y6KlC+J+g7phad51mPHDI3rdk/V/Bnc/VmZ/axj30gDW7yhHv3R4PP9bc+WI
acVFHDZ1GlY2I317fsdn/Eod5pGykExZIuMxWM5IHFg3mW7K3i2KdrvpPRVLuD51
FwVlq81c712htFBQFDeuohrN5Yxzta5wDC0gJ9LIptapXW84qExNyJbVfF98CKDD
v1c6YU9J4YCEO98i92ws8+eU+ZeBZDCip/GwAfQtzdLUjpUJuF3MMNymRzfcqljH
uAiGEHTnKWObKjYff5aGH3Y2ix9idHwxiRYlr3Vr0FW+vxJHE4ojMpz0nlBRcpXj
LqA45J1VnOI0TZw5lD0LG8PRHkhZqX31zMNQN0A8f5+JDd/k6e/yw7gU1fbjr9/b
EfQG2fuzAPoPDZYKKQ384hqnAJmjkQXIpucQwxXB6dbmY2YwFxEI4oL7OxtRlSh3
xDc/A/FhE+djhLj1yl9v80aIfU4tcSe6AxI0Sgu/nemRloHOJJeJL/SX4/eplVRW
au+PO6VP5t9nJASuvJ28hl4ovoFyDDLSudIkGfEtsRfR2CbQ14HKJmQGGdiK9iMG
n/Y43KM8+feD2cr6ztp3qiUlO5rKIhLS+QWWTNXmZDMHEyutl239mcOkdX+YgWNk
PKTrIJsy+223JwOjzHcv+R3wgAz1DjLqgS7XSPLpdzqr+Xutz8ZRlsP0gTkfHk6W
SyVnvwp/LHIKLfiVfzhA7c7a9WpakqKTb3y0KNGjHBwyNhDmkPNCI+vw+LFYj5uy
jpUVqkO9QyqCVOBYRtnDIHIQdTH4p1AUZCfWeD7GhUaJSlputNWfPzegP1A4QXXL
U0I8AumtS9sczF4hJ9fdoUK/dwjSXz/DlS/Vp/oCBRxb9llPphdplxGhtGmT/QPg
UVjwGNadLtuGAabC1qX6Go4xm0JYL52lZSea12228TsHslf4mC+aG1RhB7sC2jX5
D4SpMjxIiimzcGi9XxQmUVkleGOS2tqmoZR4UqSRNwYDyVMpCJJDg7umRpKJHvuM
upAlEJdlJuw3h+OyMFF0004EFT2fYtRXAWn8/8Ltg2XKl+XzUR0JEo2Zp8A47eaA
hYuSp+1ToJvH26rZgD4SO8335I+P6oqHR6lT71KofMlcIpr1LqXpITT84Y0ChuK1
OKccaYrVY+d29oJ3NZ52MBeUexHLrVbC1MesR3Z72KQ8fN4Cqgv483nIAZ/JZK8z
uLr2rG6zZcrqUnIqDWDvLFeWwEOdrDmoKMAeOgpfOvLu+UpdLPGCtWJLFDcpAT0F
b6osf2QeO6Sabazd+GH4wCAXAN8rP+U4mYixtL+hy1jiJC4O81lIQ8zf/7FUPft9
jK588OYsOpe0w8/71ytxb8NH+H8KOVgTfuGyq2gchwwzK64eEcdaA7P+PeGte07f
UiZ3cw0zpKifvAaio/yKphLOqCcFJovdJsAhdVE3EYdBBM9fFC8A4TuE8+dXEmc0
gUBR7XSVWbdelnA4+1ClVsaJPzcGJmgcRuoot5uSchtUTtw8uqM3gRuIgKlRWmf3
+ML7zxQPLDJqCbzCpTh3jdQypwTf2zbB0xoQMlu3JMm4MSpCSPwiiHbNxtRiuutp
OOKCwUlZStyQ1hAC3uH2uVVoezHXYq0j8WLGrtP8CHsevXonB77c2juYbcrPqE3m
YVNUv0LwhFxPpdXTqIsKvgwGojNSrLUxoezjy2i6zSf999y9VNjyn2MCsI5lyM4M
5Dz8kSnMwELtpgLy87IJj/Z7+VQAgBe2nfQU8qiWk4vqbP+UVoU52l7kl2vyBVMF
xOGEWv+hWSQTT1Vie/gt4a3z9fii7dl3WOmOgWOjAZ+g6qpTJPrisXZnYcQgliHy
fg7uGjgX8Tqt4MSH+rlgDlU+yzClgIWilwzfACuwD42K/XUra5CRCqVK9rgCN+5z
2hz3YYPGHNL9u98d4mZngR8B/7fzu0C9HiBV/BTG1a9ZwodzxTykxHCGUElZqnf9
M31J3UFc63ep1Nj1v6B64ZVBBj21P49O2BF8kc2BckNm4GYkH2NOZj7Y8db9s12t
fsAnab/lZRboC2YwrYG2fcYgIY+MBylcqC+fNRJzTl4wOjnBCRpgxqKQGzqFtxw8
tD0BrM1jKKg7D04cQSPz5EBK1j3VCQ+qg8qRcJA2k+rIVEI9IorHJfSNjgInds71
D37vtaKe0obbyoCT0pEjJ7MiNuPFZ+3IWS7LJGoXJLvldcrYFBs69dbdRxxbUeFD
rna9Pg13LvXB6qy830JCqLw4ZLD1bWF01mQPdhFB9EZ4lCJrh+VBTP/nzfPpMtjH
D/6opFCy9QAesLMbYFCJrHFgH9V5RsoR56/NzWd6lRilok8xH4v/ieZr9l5OLiIt
jef8RmhQFBd2R7f34zbvhHaSv9Bz7KdTS4cKdm3aqh4nnjpOymUaWcv3m/ZlzNR4
eqSPSXdxzBpbNYc5b4L2t9d6HYCpNITahq117I8dLk+bFNt9iVXWu8IXJC9xetEC
AGwBtAp1VSQ/X3qphumXUlmDK57VxX7TR5KgzgoI1lgwWl3aKkdiyW65pU8/4Zmw
3PNR17Te7nJt2rhqGzEiQQiAgCvaFeHM/2Y76YpRTHcc+x6YzjLDBa+cU/IFIvVO
BvI9ivdaKQrLUmdcxU1FNGrXfhjyof+/9TdYjrDgP4XBPd7Zjfq6N7TyerDMy+iU
9NKK1uv3ykoMIvpBeXEC2l50Qa3OhqC3m2KR25yslpIxky9TYBH8FbVauZI0faQ9
I+5MEDVmNhP5t6qZKaeXURFPL07m2mCK0I38T+X/ST+SU5CO23YUn1JevSaiJn5h
iOKQbTP23esf9uMZIVeNcgfJB8LQpddGHSysWRx0oSz0Nf/TvUYSVDi+MDwDqujZ
RzwZKalFardI1uZXBO9hR1YtYZO+yRpl3+a8V0BagO2MyBnjtL6KukFNGMJmqWVw
SbeXGJ4GeePMLejWtI71x+IB5TrGyfVAj7wVI9NH8i+hfstctdNZ5nFAkFqYTMgS
lXUqwqw37X/PzzBnp01db1JTI3WhOkvTUTBy3CTowkySiU3X5LJfGMxPmiD0+8Rn
2naDBgOBRhpafTebxgorZvuH92PZsMvB8BYdoJo2kPxzTisquq6s4nxW57aOdC3w
JmnqSAGm915B9mj2kOxeQ25tG3chzQiAtj3Qf5ryyoJ1Vke0fkfSxH+/ZJJz1nXG
e/ULBSJLYNJT76ejRbfB6vUpiVbIz9gK9nspltdtq+adty3aa2u72hlmahtUZnHs
xLGUXSn8s3SBQEqWcpH+wY+qSXheHgkQr28dCyn0K/U0pg0oE7FhLDDxE39V5+vs
ALzXLUBYS/yCD5tJUQ4603yTRkkuteGM3G5zCCGR/4N/XB7nR2Wew6XQ91FS8cNp
ZMw253tL6ykC+Rvqk+6Mguy5+PqXAdByDwTlTB7jj1DA5z0QUKzXUni9N06/MaDp
3l0Ls1S/d17g4+2DpTtwAkaBF5DR2B0DwS85gFv32odicoPsybHhYvriB9aAccws
oqDSFY+amUdDfPBFfZWvqiBrH4kzDEWQvSudd+nYngqIl4Xqu5dxzFM7mxjzqbXy
zm45xAvBOwFEvXnPihK3qSzmg4Oc6eDHXuv7Ua31/V1HzVq/4PQrLoALes7LbSkV
qSZpiWqSRHxlyb4hYF93dFZtp3ap5Y2crC54yfFwda7QzkgK3mQSLsJFD2q0h/k0
oPCs4aJQd3qIrZy2I7/aIpaHpMyHRDPacl57ys4NGLgBsJvq/ibM56g5CEWAMPc8
Jzg2JqMokMXbEziqBUnzdIODu3cH/5B9SpS/X3UaaTdhQgI1RxQhLpkkcrliR/zX
hn7/+uoL8JffBdzg5i6s2yXGvsorbVnKQagHVp6qWFYcS5KKA2VnSd0bbX0fgTOW
d/Teutj/H+Ono0zbJwxuPv0JkSRvWyeYueFxkBSwnmOoKtn9/aDzi8V1Io5OLaGY
d11OeCiT34T8N5ByLR4LnjoOjND5sV+2m/wo2cbH4C6iJmaSxvXaDbS8u/oj0Qoq
wmsJxyXjKPjJ4X/1ZfGh3NLEl0A0PFfhIWhT/Ho/QmqkeYTIZSlxrXeZZJrV35bR
HYE2FCj7KTAy0XWIuDGPSnr3FOg9J/fnDDyqoz831OuJkomE+K3gLXnij/IGMdz4
gmlCSXPA0f9O/jsiN7Iq7NGb0R80MgyMT2nPL8zxC2ruD9NFRnPwRoWbV7GRUQRS
oxZj/QTE1K35C+Go3YSU/3dCL2gYHCqxWuh7KuHWXRQpk0lu+bf6yTiO1coyIYPA
Ea/1s0/ALVfDRcQ+x2pK/Ln1rKZoxKq4W+26U6W+ZmnfER2PjMpuhfo+46zLpSvU
Ub+Z0QBKrlOR7zxljGpFSkJsV5tftPVqP6JeoWtwXVb1gJGjQEFCQuHtkot2IKTC
en6UPKs/+VNet4UHfpS++2E1INnImEQYsuD6kTybVpJ4UYKWqtRasT7fu4JNfpwY
M4Xcwkn3L7GK3uDswRwrRMJG6ClIQrtnIj06Lwk4Va9picvHt7/441AxOHFymHDS
rK13qVfY2H9FUb00oZMKe7q+RFySyLfMaABtgHi3hOZobBJ2ht8RzPZnVCE5H6ID
P2UOwJ9B5sPM+SsRakg+VBf8z9I61CmKNY+mvHeZ/OvOQ4XgbZGEFdHsLr/uYZ5W
p72ergf6DGh4gwAodfvEF6arPky8qgYjIx1TIvuz7D0tk32txejCdn7sO0ijXcr5
yvAdnTBZDSouQJPDrEfRpcInXrbcXgtwlXut7SnK4oGEXzUvnTrXwqvBezEX/uFY
V2Ma1mlZNWNPD8CSV+RT5/dI4f3mnT+Dfg5oFhdl0N1wAZdQam6p9sZ3KqSaFw1/
s3vjFu5TjrcIMCnfz7286r+pbhnJ2fdfa1YVM6YxsSTdgt5j4Dc6A8H0l21f0uRW
3wHRO+YiC8Ou+meVGtGYQyNFk9kGNy0FEbHVe0OVTNOBL0bvUbqJGf5LllAlkGNs
2y1oinqrP1H9auAq6d153iOZzGjQu7HOzAueZEmqKJ6JvhG0hs14r0M5cNMcyixK
DrDTLhch5/SGo2MPSJ0I3wJEIJ1hdl/+xx5LAphCcymSA59dMdTpVjfANu5SgXoa
Uuzk/6D/KMOdU7vc/cgo7VDKUjs/Qy5FmakBLm3VbzWj4hRaMjPQU8aEjKqFE1yH
xuEmhoXBvDKabcx1MW22ODbT0OjsuvYMskwwDeAWK9gDRNnqQhtCZelrmnt/gTM0
9+z976FuQI+i4ekaFA8C41bv0VzoOGO2UuFdk1rNvoc99DKI8jzjDEYvKH9c3GiD
g8r8CMGeHWhDPfosaTbr1SHfjan4P9VC0nAQZRi4FaQrFgY6FtOCXp+Q6xUsdmEb
WQ+Gf9cj2MNHfoda/+11Di8bjYrjZAxPd2H77qPNI6vdC8aPpVB+oFnH4IyE05cY
Ag1QPKPzcVp84TzDSDvVEyaui3j98XY3+RquMEYDX8PenC6wEHGPP9322KTJEmnX
ITKGjJsGoPLgfvA3+VYRt4SO5W7BAxyQNQpNUgr5m3HfnKg+7yriOrtbl0qR6JuP
8MpB+O1hYATPe3eTEQ0hTh2kRk9EYycBrb9vuX7FvNFwgGSrfF3lXo5hUesSdOAU
RCISTqghobdUdFXtrShT8xnf08lNf+UrC9duMg1NQr9P69qyGCkyUTKzlR7xZqQ+
A9Ij5S0KtKH1Rjlg74l5qfUFou4l5fc63thl6UFgkU3GgobtgCE9q5/NtDJ9NyeG
MrjcDSyqgL8p9upCxzXCXHG6VeaW09yfX6P0NzWnzRuXD6xI0YEzQKL+DTLVmxxe
m9HOt6cD/M0cCGt8KfamZiZEF9X9kvFqR4JYYYSJVtcJ2WklFQ44jfYZaoSJlnNX
MZtMx++ef5n+QSxzsM3flXzjmf5grfeSGlIx4zeVmv/LwvUgv+ti5lv89hNYW+VC
rK9PLRvRwa30FCAiOzaCTIhd7hBkiwIR857DxDhY61U4zMnSqMBNuS0qGRt2thtp
PI3ws/r0GrQgOjnXBKht3OxoS1NEDHEAghfLRFPO/8mTyZIiJVqqSQBCFktZnKLI
JlwF39o0ZJRLtMVq3X7W0jyRlaSqkL4S/zsZMeaydVBebP5qd57HZd1oijgovLKZ
uOBwi1R35VVKacB3wxPknelK6PZYEplqSKyj/pSl2EtQniINIJBw0b0txdixHFvK
sz0hLNUQwziz/dTM+FRq5w9+ygMxAKUKWLeCePA4l4ZUL1HaO521ZAYAS24UuBdX
XegBxlR3NqyAUHNn+LQv6Gf6kU1EZeDAJe0I5ipHQVvU4CRVO+CaNuInF6GHxZdn
Z5QVaLQSV7yvidZI11Bi3sf9grg/OGMEx+fdkXdMKllN3gVeceCP277P61P4hm6A
+MuudI5/FO5nU+G0kT4k5DKutP2kDOCLyn2k89lGIijVYJrYukVyC2cT8tk6/Yke
r4A9MJxwo+/2zsoxFtm+ybVNO65aErJdP4OfuOFxP4XRj5b0D8rYiK/NpzAkR1be
LgrN44ZsuDNk4f1tPR/BsEfN6VGqt6paw5Be+hjxcv9Ce7kQfbidj8k2t8jip4Lx
OFn7KEfujm9ZmJEzlNJii87BXa2rVa989qhSY29NfhHLpKQvWYkst6LKraMj0Msj
tMWsWZr7dgCtSHI1iucX5WlF5x1a7UVSm58dpx6FvtoPiykqng9GSblP3mz8h+z4
pRUrcGxM6zFDtfih7YFAJlcEJB8pdEsauOpFbd7Wq7v4eXkPnSIjM39GyhqCjVQP
TtfKcSDK1NMhytcE2EocNCabDJF3dLsJ4NlGRJ20uT8ArSnLs/SttB767Z3OAJG8
NZturaX42ToQiAqD17zc03qgzyRtWr6mUQikR+BuiRpCEquX18u7MWs0MCLxk4Sf
W3x7t5DOeS2ULt/5+4Qenmind90fH8YYtkF/X4U9LiscO6yfMIU681Xzxul3uYlO
4+qUoLaVBhcY3SpHTrXBcnAYR+dVj3ts5edb5XFpgdUw98NhYIUA7ATN9LZ7ScdD
bpEgkW6IlTbfUqGJzStK8RJuvPZl35NnB1aFlwPQ0yPtE6DUi8B1dKCLaZ96wwb6
qqMkgt8nAdZCANIbhCU9uzqJaEewyLoFaNCKuZ+eWPaVZ0Hmd49JC2yoXrcHhHWD
WThrUUqsTkgZP2Ilvxa/pBVMWhrp4lYHubh+KcdL7O0SkRFO9NxJnZoBZxYP2cyk
VwXvrWYJHfXrTnEcJ4XKmJIWlTjcRQ5XLW6tXD0T9vG+t63lWoE+uYcXzom5zNxe
qJ2P2pDL43Ndwb+UMQ5b+l6uGIcaXQazrVJXCcdodR3UHcBrPCer75btmjk91sKU
B+otgvdg572i/lvLQQhLPFFVlrREgxtdXB0q9/Hb6Rd8xsvYp+wnO9mcuHUtxLmk
u70KSQfjo3k+2gXyEtmkluPtzi141WUhNEDr5fnMy1M5gDaWbTvzjofKv6NFDOCV
VZiXdqGDLqbgb4MbHirxnndLwWG8krKNaoXOEUAoLt2p6mKnRsqULHPQFyBepq43
tbboc2PUJzcVSNQg0qgM3w8mkSO4eUkk2VuFFsv5ghkCyLfZE1AYJuNagBKDJrwa
yf2EEOhcuaUGMMc/km4mlbrwuMPtrJAsh2KmzYxZ7bF2jpngTI4gMZkIu/tA21OB
twcSCZYAIHM1XK2jQfTjxcqxwrPA8ZSN/3RStV3Jjwmeon76rbSrJgI5RC8+sWIC
/w890MiC7189g+aLWk1uFZP9oR8Gv2QK7rRQCTvLziT7rKKhABO/RWCp3FgdYZoW
gWwH7anm26ymtA10ITaZther5Dgibmkj89yqEeq/PWOR/8Ez56USy5pA9W55vIZf
S5QistQYI/JeEBY1K2oXjVWlwy1obTs9yMGj27fvKLv/LRo3tQ9z+lMaqm0tyUCK
hrodyS7h0tqIhvFHuaTwrj576pgtANlAUbF6GVkfWxUBrZ4+lotBTCiWXCKmplya
oZenoGMZ1TJ14zUlnxV7amlrAUG/WpMEyRCKg8ONoxhBE0PHht95qp/EScOgY4fY
bcdVjxkADjFLLlp2h6OhXi2wz0SA2AEfLvlpJCgwPpiD2h5CZcv0M4DvTTM2/qzu
zYSwp28qVAf0xGJmyrdmjP/kBqkcRFKtCHWOn5Y5axE365+Ces02YW+qMfmM+PBe
ODjWcRsot4BmTXUg47gSzznXUDQWcUjDGNmcftcWcRqXVFBiqaZrtwHsEWLXbdTx
AxzcszI4/PLDRj+sSVza1fVxqTb9+ndb6e00v0edqn47aPYzxzYN5CHR/Fb/8PfA
zKkWV80zSta5vTyqJ3SwvDtD5Cgw1vnxkgH/7V5+tjPqkx9zdlnDEXlQXOy3QuEL
1zGr5RfDrkCC3t8kTDGxfKgKd0EbW2VXOHzHOsxw+zA10QsZ++PfO8eAlCXN0vq3
3gsh2A0/D9AY/uWQb6q6+dbUrfaWIGYf/maJqP1vtZ22WfytggOIcyqjZ3AApvKL
+FvAAgGdxG/V7jaBOlI4a4fLbGuHG47uj/+GFoZNtAB+dsCjAht0Od5a0zrumkju
ZOV2wqYxo5akmTx+PbzMCY2xkQ0euGOcdsolw3IrBu+MUSPkkNRAV5+4E7tW1oHz
twne6pOVVVUlPDcjigebExkJB/cGYS05ZMe8OqjYpYtCLBI5n67ZJPxlplQGAmyO
+MpBaHswb9ps3rAhQTw8xHhSpxGdBpB0bQyp0Qum4iE8ywaPHNc5ZyQJlH5+PUBK
/JfuBOne4mSawn4KKtNrO3qQahBAB7F0/PIMKaCF+qxUo25LTpRocur8tDatrprs
Az2j5u2VSFm0NmNs7tmPBrsSt7ga4IIAeUOQWDUCHZ/GVnCN4ihfAodNm8Us+LZu
/KHMY739XSfwj9b2TsaCDa1xo+OcGzAh7etJqX1ETuqh4KB76Ui+noSWrjrAGyAH
tCcEm71BUmqUrWGXHXO6Dupmh2LyTGPnppEHC3ibFy7sHzRpKsogNJnO380qUEZe
R3Ea1b/mKA4o5Pn6PeAWwoEIs1PD5LdlkuuvCMhA19agSyqMjCmcgoCOEqcgSQCQ
qPQC4i0IzganKnD3ZHjpOcVvS3uPNDR9BO5wBy0d6xrX6THmMf6P9VnyW9HbZJ1b
IXXQKkUAT2ZdbL6OtICVCIWa8JOwFPjg/T0Gv8eVIkWJIuvvxR+LXu5mQrwy5X8M
YXWz5MvGIevc86U3Ve6xRh1YitwtQQ4WEOItgftE15eyFp4Al//56RzNVHqjMBhg
pTLnx/35htabdb7PtL5jAotvpblJb4Lx7RwbupOaPMAxMzX8hYJj3EDL7vuEtmKH
UDiBN3phrGK32rJfO3k+AdwH3/NR+mFnoSA8/tQ2sNFvYIwjZ48D2vS79MCaLOa/
RTCJF/mSrdpWr17hEKwg+uUxNU4wf6ZYyu+iOWGNnthatL2EDNx+61ia35t/9qBV
xOSLLzbDOjX9b4PsRI/IgKN1Z8JNjS2Ke6n5+9rk22GdXjiMztZVZCtAWJGt6P26
wJUx3Ol8ZLcUmpoRMAVTB6N16li82q0eQFBlrSkL1ggrOwybN/BLZGVbFm/nPu5C
7AHlMNrwxyhkBRtiFtFcH4afEbjDFyI9lQ7G5G6clCUYrQIQT5MImK+ToCSn08ow
UxjQop4vWAuEJsjYaB275O9Q0qi90vQ8vCL9bxXITYItKzsQzAQDfuA0aV+oTOkw
qi7pJGi+AiMMSqJTjgJ4mvmRUZsVuyDf63AjfLEcrwMx3ed1jK+tyc9sI/S7TfIb
Vyhka8ZuPJFtwmRhuREYoCOGbpXym/4XGzWzJaKADoG40W8gzvI/ujTudN00fLwL
JrasxyqRfldcHYcM3xrs1nrwQ5hJAFALgf1t7KpokIUnSm9vsIZlaEiD2XbsIg8N
rZh+AM2206+objcoCuhJrZfjyoZMEy7pTqgQOHEhF6Y3/BiVChYWpsVZvUl32DQC
kDIsn5mNroKzs2QhRjtPLih1FQwdoGJe+GW+d+1cxDzYg0PcZFDmNyqDvvN93CJX
/QCGCsZ/TcHrUye/ONGSGsuYGikqZsVqd6JyQeTyZIPGFGRGrmqYa+Zw3A6bZ6b2
Pw8JakVnZxdVZ2hGJfA4TVZm1xYf53aEiOy/a7anpZK+c2QFtQBL+ZScjpBEcjWT
4jTKQM9mX/P4PQumaqLNSnBgRuzUVKto7AdnPxzdArLgn1njsgTg3vq91Syls8N5
bABc82n9wOgPspPJt4dnSqGMZLXjB8YvgP4FXyEH2I5lttD/tlKHSMKBMWCKow7Z
YqrGXR/0Kj2PCJta8D/4ktc4HanV0kK66WxOXJqB+F0LmWZOLz6FJyq+l8TlIifQ
pT3OO5Hf2V2D4iXlXvIsPXnp5HMvpBAI8NGS3/z37AZREVW+Xy90hkdYL9r6d+NE
UO3PWrfDHXTHY7HHliWuR0WTxpgYoHQOHF0PrYDGjJ8FhxS6XKa7pBjGKOkVXLzW
stuNnt0iCv8LQdkSCuVG3P0H1AYa4cRxfg6maRLy0p8L+n6d54R4I2RzskLr6rsH
8bLs7SE5Z5vF1ARQLT4A+lz79ezGzwq9yc8LFUL8+iT2W8X4UpnmD/uJOIXOWMVq
mlpbmyYQEqz9jxsSaRZW4e4skFuNh7/2Wl2tGx/vmjGP7/39Nq3wbOWWsBigKGuP
sga9/gksn1WuI6wTBL6QzFPQoJh1NNoCTrBv2KfdWNeQkskBkMpkhlCXlUFlUtYr
Qic9qPvFFHwvCeonflf/CPRSKdpdi5ZMUG7kbdhEI7Mk3oXoJKSNEnPk1F8pszg4
5xrz6z46h9OqsJSE/6f+dwR9nPaOUAiQNKf9iTlqgr/Bg2AsFEaWdpgk1CU7V6y3
/ritJICj7Bq164tuN5k1CjVcDyWrn2G3xG7+JI/L2dM+/e6ZuPyqaR7fszuFKIzw
Zy2eJ/9YkeTzB7FinD6zIs81fo5GTjZ+nulg+UzEH6iOskUaMDanYFBl2T+ScWpm
AekHG4UYcfk+HXWqX10cqRlILXbj0XlzcxGIvvwJfHHvvhA9bGH6jKgpgIrszCla
k3YJYjzAcKAHkEUBfQ1pJTiHDWn8eq3VTGKdriScszNfWDK8d6P7ByF4AfcZEKG3
7HqAlHNT1Yhgy4RonYCAW6xVYZLG9hUscCCIQzBT9MZ3jeu0alfa5CLEFEUAdOLC
tuxqFlcvn139msBWVWwViv6ven5bk/4tH10i0KWAFX03gZ51K34dokrDEU+TkAQS
MPjVm7NAbH/X8iDgXqgWHY6b7uev6cHJ+46Q6jSlb7nzBP4QO2cQCIwEzWt3/BHE
/6pzHiFD/rb0aXtos55Auwm16zhZQYs1e3/VUNf2G7J0xtzMvjxQIJIiw1LpBIt4
WkTzkvA83bo4U9ArMOpTTvOYMsISigKz7Q52cwzRp9L/i01eB0pvQBH+t2BQnRsw
qmJg1Zmu53OZuJOQd8z7mPGUtIm3mWwV0dYCH8TidF0LZfRuuPrIpVJxkws9++3d
1WoTcxpAgGEfQ4ce4fZuDnLHhuqKhl+JwS3zQ9m4cnXQbDiQ4DIFwUIA+IHqMq4M
nlkdXOspqFAUuwsEoHaPqgjWMO7HAdkO0lglN//VD8JjtKQbRU/NcQe8cMrzlXBx
TnkIb81t8Lhtw9DFmu4XpgKpE/AJVu5qAPxRO9gyZ9V8jUlHGuqhbhgqR6Wxsx7o
ehWY7P5ccQ3HeyV9Dhszp0E5+ountKW+Hycii6QaPz/nC59cIIr8weVFLkG2xn0/
s9adNUY8eIyMHUFuTPbUZqNoA8Mmyjr9emWNPNs25O9AAzOwsgQt9pgSqJnAx4YP
KVMKRxp4KspNNG2eMdT5WYhVBSYW+buBvgGQ7ytPQLSn4aC+EklWbTlQpZaAGZ7p
EQP8bHCNmlzqcjrbrtSuECp4CgysENVgwFWc4/OebhswXDL/Ez5HOmeLWKURNJXs
3XY6iE4N7HF7mN7wEL9zbCoRWf6yWivAog2PnxyB7TW9Q/xqNJ2TZBvTFSe0+Szo
sHHc71aytE0Ia0++F8rw42SoZ+tsIILamJHddS7baMDzaewD8HRrUuRGa3wcyAHT
EIYlY7zneBNzP0s/Z4gpKgubWdIPXhScecEWxmENzyTKYXoX0ffrsKz9XJm3Prmz
8WgGbhJrLk03DQTZ9pRdJbuoyq/uHC7BmNe0JH3iTLNj+sdUuVaHWwh0ac2SeoBF
1vDZXHjKZGdvtT1vpIADNgZ5tfai3gYg/iJUuxITvHqFjC80sZAFFxKnenz/w0n8
rGkBF+0MhYOiggWZB34FnXuCUFFUqwQqRPmyQY/zpR2OaFVUBZzA35NWU2znKzeq
3oRaRJC4HytPl9+YwB1SopzvIzvRSKw/RWQ637VZG6MZbylNpt7ROYw69AiT/+3B
KGK4f3s+O3jwpMCjxtj94y23xkMErafEp+GZWlQVo/2POlylXHXc5ztZb8Ctmne5
9+PCtEeHfwm9GBzVeB/a8QgWtCdOYtSZCeQDDC+fYp1Um6+K6TlpwpxbZ+XOSAay
vbU5Hf0FW5nOe0sc95bVEtpRW66Oz7HpQpibK+RnY6VZbDk6sl+H80M1rm3RKO6z
2oJsmgXVglyOGZsr5sUUFWN1AgbXPXw8GaVVwqjI6ICCkpN7ff5akEhob+z1XxIq
KlA+OLblHk1juCSzvr8anDaUf00o6yQLWvdYp9jzryUofiL5en30g4iiBvXQfCZv
7RyWp+i23tJfyg/V3ol6KDFVDg1RGwVIFGOUhrIXBJBd0t+1/XccynkwvN6/u5sN
smgKZLIbvoNkpwnBKueCgMcrq7Buf1WSWvjaNNnSzRRZadcvGRXyp4VFfx8IOyd1
OvL+pgP6ddSFoI8MFTDpnYzHMFE6e89lokp/yuDlgCJB/mW1sOzQsT9AG5OJLZ3U
iuZsNs9yx9pKaSuGtsSacTiQAd68LxUHDMVpUi+jdc75eli6n6TIfbw2JKnK1/dz
XBvl4sDSaR8HcnmNSOnsnWhRZR/vMnO9u9lWOR88jI0VPtasPjPVEO6yUnX3VVq9
Z7Rt970qg4lxwG8fSHc4aGn5fl/m5ZjS0pC6nZZc5uPlhl3OJrtPy9UsS3scwftg
+Ew1GTZGotvAvdbvaHJuMiJWxE76AsFFYoQtj42YIWl1RMdBLSQ2ycpsjUO7smTc
scJYOGB/f/zejaIelfQkIEvyyuNlZROYSjx73YdxelFKtWFpzl9NsEvs3v5tVCSN
vSnLMqC2qdaB7fx32GdPepx+J0MjRw4MBl/AxaY+LEcDJcMPOvKBnu11vDucyORR
KL+/2E5UlKlT3i8T3MY1Kf7ZDrQJqCZzhF/oVoz9E0FhY5ITXo2cQwEzi4ZeEpcA
p9eHnHBV4EKssF5/7jWpEM3ifeLgabUHfotAqHafNqrerCr4Sro92TAVLoNRcJSA
OFd2s9VLcoSdKtIXbFog6uvg5wpVu2Kxpp4lq5IwuuvoCJObZixdyc67TzLl5KSt
3htJMOZpUU3yJf3KbetqD16FNC7aKI5UokhproczlGuT4X/WxDP/+U+x0nj0ToTe
zbtt/Zt5iuiE4CrvM2Xdz49Zx2haJiCs9Eg4Kd6z4qMmrzV9rcxbwHmCnzNefRu+
jBN+hcvD28XtwsXLZBo/mj4HPaddT+rAMgO4bmF158uamX2TfYADEEIbehQ4UfhG
N3qBiSSel0j/0alIFGClyKhM6h9M5zPBhFoxitoG8LOfGQPe41MOK636G1E+3YQJ
B374qSEaj5rV5H5RQMGdtnnBUi5HAsoC75esTIJu4eeCAXtX4zV3w5x6jY0vWGpN
pCyaFWCX/O5MGf4/wHwwTHRkef+auaApI+gBwg6g+8V/hhhS8gS8PDX9fXs3Ap/e
1UgSJQAj7dewiZl24LuZT7iRdWpRGR1IjcmWOZxGK51vAiW7Tucx1Fxg6crUqIgH
mOMPQu8vXj3Fh1RKNs5x0EMVlsCmQ3aMQ8jvA6m0B6nUdcWFXB8OC8lGRlT4xp2u
96XBs3xroOSEypaeRYWtASEIZlaUn91e1LOpxsrUar6Jd/3d0NS7y/unC6OGaNww
ge2an2NIZMGPfYJ26TKI8QXstZZW7h7Xmi/XLtqFYXh28i5cGWCutBVzuEXWsPMl
rbWXM8OC1UU9GpfxK++/b50Uijrg1OoSv8nkx4YvsLUeN+Fljqegcq3efSDmWIo6
sRcXlYADaWubQbMhG+AiyJR/0yFwRoCASotwK5JA1HGpxdrYM6CH2iSJ9f1hXYH6
A6g7TR26SqJyq4tQDg91mPQNG3g5QUBlDLSnzHV+bssK700Sg0cBje8dlRjqZ10o
IfRmVu7p9ZArPkG3b2MuJ6nCimUtzGetJeIflOmB+pNcoHD01DSYvB/qL5EaZeZn
6UV4qcOhL5IhYKav9YQsRLp/HrZivY4J7tDeuzxJIoiX3wqSoa5VT4ODrw1Y4+Nh
IwNPZZdU7nWXYObEiQkWCQLw1+A8CsBNBscB46GYCSjqXWLBNP+edpQ75TV6x16t
k9/5f1SXgHDyIR9G53OQDVja4hROJkn/unCLxihz5cgOhZ4OqMpoUrrmlVqv21TT
tQbv8sOO0NzN0WOWQAqD+a/nBonDso7qHvvhuNL8jo5PT4DbghLowFYWYPLb7n82
OTRRfjXa+7/rP30qKKZeKmtJYzoPydSI6B1VAudgjQPvpjVjT4dj4GGamIgFZKcc
yrXt6g0c+50DD41bsNE8B0mvcysmMRL1OTkGWOfYMisGDEBK7/dvjFVTzQO6LW1h
lmYt9xHHCcACtdVvkvvftkwnaXU5lRLQXYhllJlWEaDu2CpDZ2ZPbIBW73sorDXs
VlroCwGtQB+Xgum8wOXC5kvLkwt+nFktGZQIuLzL4GWRejH8p1fGvj1hNghS/JPd
vUuVTO+rzb45ZY4e6KI2jSF3VGpd6yZ9br/iEeMCo64Ta9SeDYA4mTrOZ78PtBTJ
cT4EJnkyJz8MsLZNQoM9tglTkOG33kN8iOnn3aqHyryKM7ivg+E4sWMP+KVVTQWI
lDsR2jAxlqCbdHif5ycT6aWwWVAKth1kr9C7EkwO/6CKS/7MNy+pRfaKviUpDX2R
cqbuptIYPSi2i04qCjBSdnZRNpjDc2IvXw++t5yIYahRqcDcLzc3HGqlzZQcGRQg
fYZmGiw4EMxsKj6HE1tCCDBTR+BCOeV7sxWfw0pAYSAhFZXD5Bf1DG5XdKKgYF4c
qmlMzMQfrb8qoDH27j16fEFYmm7JbD4ZyM49ediFGPBx3bzGKxbT+kArR6AGqzGd
XJqtp9dQBHbX727FqEYKGNL/tk/nwA6erXGjoE3A5h7g9YJ7rUyxbMk5b4gocbcJ
SZXKLdtwfsC5KoOpyDVT0zQA/xYIs3W7vqJIv4vkaG/jdRnVHQdHpt8nrXznuotT
J5eICIv/4s8mz9fJXCTKyJ3qg7Npt43najm5d6maiEZ2J11bRXkKoA/L6IkVYisV
Ny4zdcaQm9XExW6/8ePpSKYJgcV/vUJIVqFRJZzPb5euyxVtYuUqpr7tkv5Srt3s
o5MphArAcGfMB0zjPt7AagSl0wxaz936Jfxm2UWgHqTtZzHzJT3gvEXLbaH6CgRE
abGvJAVli+ZLOkScGnvAuPk0uZUB25lhWNZ+un5EfingOwCxGa7FVvBmZfKbzOwN
t0U2LlYhBhxJHHamhghqtD1Nz2hJtPASskBNE0vJnuOtJ8i8wHMuym7Zw6jcdBsr
wva8Me3Fd5sjJ9luTRDGixUz1dEtF6DKFJrb8HUeDYjwg28hcG1PoN1hcSou3nq/
OQpvycHYzyENfwlpKe8MXYamYwGic+7YGXWJOPsSBITREgKA9Q57MQqto6blkgQE
Ufcs9txt1y8BvI2rLbObKtW236C8J3SIvW3JrD9G9xVDHKq8wq2axS3MrM0hfIzM
y7ohtNtL5d8AlRjThKv6dIZdYmZT7S61IboAmK42DnekOEihq3QB8Hz95ra4Npq5
OrNOMAhqAyDUyn1OCGpbty5HSFZVYAZHdeNbeFDSr2GP3CUPtWS9RWgGhrFDEfE3
+OxEhjDNug9o38Xk+tso4/UGoFsVJQSra1VFZxJbQVPg5HZJfhKxjob6CutWfly7
TWD/sojNk/6LqjD2L6M2XgyzQYB+iuEhDBpq2HL1On6hKoo5GsTpSZZTEJ7ips9o
hH4AKk5FnueLaGlWRNEJv8oKeS67uF8P8wIS2Ax9G5YAnkoyhPEpB4G2jr+efS9f
6kl5ziZIxysQNlQJ+dyji42MQPGwTbfsQ8FAMv6HiD4bHhPJeh+f5nMS1fiRf5fO
cyLg3lV6cCyatoYkm/m2cMqe46uB9R5Hh627RCCaLLoIUJdNKCUANeGU4W7PKk1Y
vnYTzsx8WVYPw6ix/tekScDyJNB8zjUNiTNK5uI4rFvzv6UJY88t/0l1+FgVIMzn
EXG5dgg3SMLAxgIo3gF7xAENKC130iFNSFtyGsOkZ/OZG7XbSB6BDPlMweg4p1D+
Po5QT/32K0B6JxG80aLsKmoEFM/We84VhyVkOoRrzFsdeKLAO1aQb59MMmJWGPXh
MIrAQd7RQQOkqBEhqyesvea3seqQyuuZmM3FdUExlj2hJk6bqBjIyzPApn6fbX6a
iaAtt1tUbv/Su0uo/6HdfS+0izNuyMi9IBt3zJo1ddqt32wu6AC6WNmzs7SImn0/
HmGdElzJd0GMhWA2MCpt6HNhFp/0gcLw/2lewEjZrGqSeMoC8FeN7K4p5fPRvAW8
GsXOaCZDhVJF16n6o67alZ7bTqxpUz7e39e2pPk8ZeWqlWNE2pNjphw6rOXYadWW
kmpFnYQsnBbps13RCv3/lKdEePpoN3ynsSZpJO64huNqVXLMUvPpWehNL8LSiKCk
WGoQaUcg2/0BFk07xe8btqoyeT+kGs2b8Fq+VU8WVSQ0kTykXMcr96qrqZEPtaBB
w6hZ/zza7eHoQAcXp/74sJqMiW8STy+w20Aikd1uxHejWaAC2fEfAQXDi2GV8vhH
ojgaFQatzeL3IDqJIcHTqxj1n7E5JpIhjBl0t6IxYCPbSOuGkyAkGLeZjUTJ5WOa
6LzQWJm1ruwPWz591lb+2w6XpMwwBQDrkV3E2raTrPkOqeiD5gRGNV1QE4wXMHHX
RXhLPFQlNyyh6XNwdeizeqrz7fxwYQxNFcdFLv8rJ49AhGMQbMEwD9oVHT2efM2h
bBYlmByE//geVuNRl7jKFVlrmB2nTINyqIWwSC8tI08Z41bhvWL9KjDiS6wGPv08
XurrK3uStdRho7jjJBurF33bDM/tAuMYsbUYzRNkXtxmKBNiDUcNINEbrQep2nWN
6QkR9JminAsX1STmHXkgfnEUuAF4qo95wHkGcJaa0kBO+TLxBUqy9ydPnCeIEgSf
MuEaBKk/QwTeHbftOzcbLCu808HDhiGtKGcV4qJAkvnrmN8kVOHitoYF/lUDclZJ
JwiPi+abpZqTb9S+2fP423NSOsX/s8O/YkagrnDXG/CwZG7MmWPLSmGGFIuvrUhj
vYVAz0rh9je8YHsLYpQ3dXaBZNaR3LeBvEs3zSbdfmLjizf47NWKxj3n0vss6FBc
YGeONt+IjNi9vzeXHhwjuQR8CPZw2/W4CX4L5D2gt/NHWfR97mqggeftdtZ4fKBr
9woPsZS3LTsYnOzRj97tIiGruHLpsHpC0r0kELfQUAzWa39QdJBSVAh+MConthcW
jMffYgARC7wpGYVohtUtF+D9vextaDjGnMvbg3gnIlzjFo3B264LgpbP/JbjGXjD
9qVxycHLKB37VqdYC3PED1/wBEtVF7YY7lis/R/Vjd/TkZdBoi28kRAXGddGP3Qo
CRPGWYmzhy5anlOfI237pZqYW3x/igplJplmyEhTqrNf7kY2PT51rtX/I7wCZMPO
L0bz5+tY02YGsdunYpHIxzKV5M45T1wPEWhuMWrZLKhgPVkWOTQfqsge4gj51cLs
AUvoF0FDes6bK8tDrPaWRT/neaG/uZzbOzW2n+ljKEsR65tqnWghwa7Go3FcRv7X
7+Ar0krH3/OZNWMp+tqyd4ag7WTEQK2lpfW7BRcaU+YAS4RTd101Z7vTHC8N5J5C
O8o9FaAdbLIu25QxJg3IYsTwazP8uohDmfx0ZcQFWoz912tAmpmlorRF4Cm3XvOX
oLvtl8hJNjwwl4mTLLi6vAbf1brrpf4fh4vI+E7hPoALqbP8zhwbW0E6nEnWCRV1
5tbqXgQnUM2eRWM8uqubGTc4wDSkVsToMY9U4S+A+08efaggqsl5ouu8EPp+uYr7
4i4gwkB7t2I79fRY6AyUcTGqlv8x4APUV+SsA6qtxCm6OcoYSXRC7Ba9CYSyLSur
jxz7GqwGdk3A5SFHCjfHAD/96g3Dq+URpD5VoBolvGOc/bDRtakhvKXrpLBBJ5Cc
vj4rPZBvMEIQG8K88IWjL+QCA71C0Ui53+2Xl4r8h0WNa7ks1smkSHbVh6QMKj2V
EeYojVpKSMFd6b9aefbgC4xVMR35mijMV+6bu89S3u+LtsbUyXbfGg8b4qs/xQCe
ZKTaV9Y/Zr2YMWpht9ZBRmA+kXDBoxuFI1kG9e5fYI79PgMwMCxPTNz9LEODIz/a
cIvpiNJ4sCnNunUBzRGDreHBrd2jxIJ4f+eLHC7Opyc4cCRGSSKqiTITr/wpvb1u
ZI7yt8sW9rTZP09Hm3XD5dWbpPqQbPcW7yopWdIDGy5jSiaUAKk/77dg5NjrCYQ6
O/fkFkypK38z7RMzUykfwqon+RttMl9uPOnC2nE32Q/iA0q1Fovu5ap/DTQcZzWU
3fAW8Q+Jq/GKmNT9qHiWjP3ksY1tAgrClBlMn3QCrSElwhPacdkZgAxY74H9zaEs
hc2C5DzKuXbWo3JPveJjijmoS/4az+OyVRuLMh2OgDC+4yZbYkqGySLkHnFN2Fd2
fqXHnq6W61f+1JnIus38ZG7yEenOAHAtzxZMTpiTWO+s5O74xuqzIqZDFRkp2OXw
plYMVEJnpi8QD0poI/2XTafXdd+6S8OlPIc4TOejKE0aCDus1q1FmCL/FbWKg0Le
ty7ZwvfeSJstzOQzcPBOQOXWoOTxksOhI8Hs/Y3kBIN6nd4FMUtzejINHrBCJhvj
0B1nU0wN9iRi5zpdRro4fm1E1HnvHUBKnWMIxwlH5rkik8SmTjMEy/j+hHez8T8C
HTQXoH5gh23WgcE50t94OKVkhImetteTCbzFh1/l6oErMAYajL9HyfRrOomupWQA
br2oWlLCrg2l0a7oz9RFDPTv5WtMfYx3II1q6yPo8i3ul7yLyaKCZ/ubO0Ljq2Uk
KG17kKWHa7XS4IpiRKanIKR8amCrRNRShzZEengXrrWHoDSks2y3ZP8blUCRX5f4
hnu3Sf/FSe/kigT8+WOYWdGi1nfQccPl9HEVhDmOv0ellYq4G0v8cOqfu+1lrzsy
97W+eRV/nkMlKIyCC5AsJ0MceKCPpIiIusdFzv5vAoK9igpe9084wSY1Chgglp1X
qhUKSbMESos2Gk15AayMOuJC9BcivyGay7VNuOnPl2z1lzp1NLL2MwPfVW+9XcRR
Yt3La6ez9gPkrqPQKNm3/IAXzgGcEcbHTsutyQdgR+FTJf3KwBaC7ecy4vZAGR6+
RLbjvk1q3+b71OEF5oI9RTHYSqAhM3Em8+YuzL3xtuudvounT1MbAZVOI7ukLIMd
dCsjc4zhpp+mtVA8EQfBhS8RrpgU/xqAMbQ+L0q/I19ExBGh5oJsIgaXHT3pviAi
8GjHi9cH2Y3Gs5LqHQFaiD7Ne4TzSNQJL23tvLXyJ/je4QsU0qcFUC/uaPlJXT3s
Poc4iqlr8fGWzzUcyIkBmimYEjoUgJNwcjNLjUA/gBkNNgtt4L+GIXTcTP9uqQC1
sF3SvfnywuR43nvfJwVWLWshBsIb6UcigPj0ivqQ5ktb3NcVm3J5whfUAd0gAoRB
sf4gomUUl3V5QmnDm+c/vLZl7urDih/eaCba+NtxMrV/TFzuS+qUf0JqSseMsq0y
SosUdAlG4XTfTWgu0MppJ3IZz+7ss9uHtsSBujGDPQzzW49VP+RGZL5zJ2s81AdU
xLV+Yz6n77GgptMYkgjd2uJAVZRdqnlQiHhMI04skpwEskeRK9SGJj6u3MM7/x0i
zKjrA764pvzYZFqBfMb6OAPA921kYc+6kJCq1cBkSnvhHLXkFDJ+scoNONLoNhuk
8vHlfbwDR0O5ebaBd/Ja4oZGkeSSI7JWxTY9CC1bk3oC40TDQa3K5iWcobOfO5pB
1n0PubtHC4WNrsUIkQDvzAChBm7eQyBugL5pNt5HkXcDFV1v93RAjB6d7+9dAOQg
1XjY1BmCSWGiLYOWmx6peNKisjdDLvJZg0puEk/KIElv0jnHVjWx48/uN7fSgiKy
dz0iL2v5X4m9WjL7eVQH9z9Otd34DP0cTR23Gue4aIe/Y5s3ZwOTLOb5eszuPb16
fwaus2Z8+B7aF5EBI6oRXy6fT09ru8/E/Kot1iIk+ZQ7J8xJFjKYguMBQAaDh/Oa
7pL9/PXU0igREP8J1/XlNgTBvZoO53h7ff2hj3V38oS0GS6I3/CtWMK9BME9VCXu
/4QHXF6nxBNJ64pfKH14oAA0HuXz2EjunOB7c+VO7DhPm3g6B1fJfByICl09W0nX
VeDHUyZ0aBokrxdFbjvUh4WdqJlKsu9W4on/vhABSmGqholFIgqksVJYxJ6O+RQC
ATgeeXTB7zvPA4LddgPx5/QpMMq+XTIf3g1s75wpXnF5dwAXz6tT4k8gXKTQ4d4r
XaVqOW1bbyVImRV03r6gk/OG0sxFGilicDx0xPhcliEovws5ErqZi3YIfvEGgGQ+
/FrWC7SGa9N2cZPsY30BC8g0KkYefRT69PFMYMB5S6ZcEcu+ZlzYWcjKkoOwIiYV
Dn8Weq/RwosPN4aviCJjqt+V8oAja8iLA+9lV9uhIOUeGn88ptWUjjnwtX4d23DH
ti0tpGewINWzHN1xpygsvpQSB+JO2Ss7FyR+ZooXoIsQvSGeADEG2RLMWE6fAnF+
dPpmuygN1bJydPIcU2L+97mDaIRmJsh2oGKReYDSXROYVglyZJdrY65pE1v2udvl
68/fops0YKdPCizTuYsNA9lazMcIIyx/U5Cacam9cAC+rHhG62ZViSYR3Tx60zo+
4FZgqfIfHOvcp5dsa/7CkNzCWkT6YmOvGhg6VOrJtCOjR8dZWEW+2C+kntE4B7gt
MidEFGhY3wnED/GXmnFnoDzzAXqWJiPzoUM71K9shNMK851TpyKb1iAaWBP37H1v
w1AdiB6t6IKuHV3pW+0AY+bhBH/lpCEQZeLTZuBv05QTDYwnqxl4VTqVsdA3zAdQ
NwHemUrFzs8CKrMSlouZkdDQgxKuCEWFkN8KYhY8yNKNcN90Z+JXiW2y2BQpb9BM
d0u3H31CL8+0XnfiriW936eDA8BP8045ESMXuA4h97+mGDBm6mGnl23HlP6KHsvR
CmQyN0AeKo/2NkRCxiEON30Ja3cMrNeDQmwARYao1L+ri1QVySK/q2dcdZnyona4
Q+EBXtp/MFa3PaVuzeXenIxmVlF3knwQ0ZqBgTxIeH9YOlbYV0t1j0OxNml6Tw5U
HQbvwwfRGdCapRzrJwCwBt5WtGyLmdRTEWKy9mMUa6d/M2Y9GAgQPN4dum3UOWkT
IPNBH7aFqcjZOGlLPYjmuizCQwWdsJ7lyypONI9uPnHIi2Pus7cwhiybz9gnswfK
Qc4esrZTiU9+9DKr76zu5gifTLyzZGiTNiSyYZXhcuwuL6tQNTyhy3kWe3SpmFOW
gqVl1+V0+1TNNLonugNIwPrxWT1SQpe6Cc/Peu0kG4m9V308yraKet2UtCpDUQkV
N7Q2HAT2/g0qa52nQhvAxNK0ZxB+F2oiCTyyu2rW6D9O9LrZcAE4an8QGQVWtwNu
n5djBU7VTMIITRGI8L7zoxDIVxSp5Xlphp5TQgaJF7bc74Qox3YjeLnMClcIFp4d
Y2kTbEAIvEsCIw2XeUBau2Eph1MaIiuikVI0DQDjKsKjf4B3kl11YRDHt8b+fyzr
IV/ni+fqhEkjmmVb5Kc2dhEu/teSaqfMCHtAKsa2mXDYvvCsov2GTmXjnVDVp1Ws
1NUlBnzVCcpCYtpJ9zDdyIKRxHF8THKoB+eIZ73uEdqLfhoKVA/PoJZ8t+Uvo2+W
hj91lIZawIud95jMGGKqWo5zi8F7odySiulQO5I3hPqwH5FFuzm1uO2gv98FOjK8
xW88in4fsw3qYHrNFnUganxBVC56JpGCV6LZBj5r468lsLiU4QipIOY7zvlUUZfo
Yn5oc9Hbw3ynG+kyVQI8FEd31b7zGucs2EolE0W91sFgp6uPEYktqvPy2ee1uIKA
4AcVWmem3oyZ2w2SFmdH1EQpcoWEbLdNu4z/3LXqjYi7IayHmtSk6bJAct4uuViS
YLY8ZMENFS5BsjbMSV6byOPTt9pZ5QbUQjXYCGlwoRrT/qj+0XlZ/nt8YSLdRIzO
T6rkk6FretjgSF7FMWroQcY3YQgKycZPmJDrs7QxotPFjgs5jknxP4robeP1+5Fr
7PN0kwzPpCdeIbw1XS3Vq3gI1DCSjNQl+hahuxghyCJqF92huW7jp926QP955mBI
lGRwcBWhFz6IjJ26SMQViV86L81BAHXT1Ai7VxMIMZXHeWZowET4pruKUBOxCgE7
cHIhfOk3Y+gNupYjRRKnvKft8py7MHC56MyWqVxNYlz0Mkt5SxWuLpRDi5eSq3a2
EJxuMxgO8y1pY03KlSsjZR7V1QhU7Pzpd6kO+Vx1LRebVnoVnyl4dzfdibg7S7ii
LSmgd47Hnc/9xJ9yQLzCyTtnS0UCHN/XQY8xS5K3/X133pMwhwBTuCXim84dak9D
lnljTz2+2RpR7F77+eH+V2k7DHd454Et3Uu8mhkAlNr9OzXGcHakUyxJM2x5b1m1
FxZBYJ5+Hb6w6ddikg12oeqYCIAVrmsUUAlAI2gxfdZuLpuGGvMbk2L8chkl3ZQZ
R7zw2nQJVgUhaIgTaX5BMTTGErghF/yZuYjbZXTywLQiihaCN6aKKpFCxxuBiVIo
qy4xGAUEcU/lDuq2bLONZZ1AAQev5+5eNFa6q7tNkzBgKjayK5tfNLXutBM5PiZf
8+QLUjJiiyoYuKGncLIQioBE6hKramtuof0O9mtqcEOXB31gWjqyhYFiQM7vrvA8
2Du0l2bgSuA3vC0Debm0QIJB25FhEcvMKx78plqMYwIE9HHyh6aNwlse5jt3p8uu
uGy3taGjj+u8/BbO7zovFRnHT4JjRJPA3LyOngRA4YBT/7UHfzG5Pr/gl7WwHTSv
eAPCoosm2AUj10vEEkrLWxEkfgrwVVkhwpW6RMdFWGV+8i6lAQrjfoQRz5CFaS95
Ir8k0cez8t9als9wDT4fah1uDX7ovzCfOH0byxCs8MTkcUyI2fMNyjFiMuMlLgUW
RkwfBJRreOcvrq3FVhZ74agGt1O4gBVol4pcmL6l857z8whtpoCNjn6+/ioLNngd
yEHMjA+ERhIbDZcqCZXyp4sysjjNtnGh368Nu1rWlj3gZSS29My53I2Saq9V3Yem
8tqfGnli7uKsQFvJxnBPkKoZivzob4sTrHQM8mvLHQ9cNa4UIEfhojt0SpZEldX/
IA/7yVxVkSKjNGqdTB7Fo/wEwv4jRMXhDb7ESu/BL0gnaI5dO6KQMKwDVvp0bfOw
QxTXJIaM/NvV9MHJJ/I1GVTLCSRndDRU7XxQqzj8UkOUh6Hjjimhg7R8wYVTHcKW
IvnIJa17rM9R/Myn6Y4ozyOIsFJ1tIXO0NRKcE0bmU6WBEPhlEzpH+sY8f7KSUt5
HzlxUUylZiIRiubG+bIunDFaNS0coJBjXw407JgROACwYrIsLYWtJ5G4uOc7bqqY
cYxPUjcy2o7MHC9GE7ecFKS7pTJ3n5O0wVeRlkNV91wD/5GF9KjW7qop2bxplaDz
WgFXsdHyn87q5BrfdYrenC+iDQ5LAXp0uF5qWbkrjIyttXuk8prmKcg7g2EAY0HV
QMBgIdZxdGppEiStbTye3tT0geuU5qovXXseIPb/UBWj9k3MAF8JwnJS9Y958veU
9t0gd0zW8+QUyawwEqO+LC/VvfiSzLyf1LdltMTp/uMDB2iqgOuKhXdRwtUAU/k4
QZJiwlIECE3s4wQWQr6Tqr3iH0lbPcQwUf5pObrtzbyOqwakIX1ESuiucZEFbIrG
E7ZzzNaPpbKn+Meu7S+FySWV+HQVSsVj9rnBS3ZJBGB0c4KctNxFoQbKa2M7eVba
lIKqnKP7/5xrkUjpbZxLDlB7GGnjNQpvnn1DxcL2XXcpBlEwO7yqG0IQ6yfR1pAv
HV4ozxgWzn7PRvWi+IjZxr9qQzt81yScPdaBWLSQ29YmXtH2B5sJKw7pgRLqEK2t
OavfNLfYcT59Wq6Ll9GEvoNILej5bdDOI/LJX8UbMICI6RoxHU7Wn4icHsJM5ZQ6
gi6PupY9e2tPUwxyA6Wap9FASUdCeYudShQfkzaYv4WjmQrggye1tUUNKE6G+62a
NnfnmSBdh1tZYqVVV4kXDtzzrrEtXIYPxmf2E25mLfVu1SzlceBzPdUs0VSSrEj2
IXuUIpx501VY05UFnZT6YpDCQp8R3uMQUMvbdUYHC2kBNZ4fXgdoM2yzFVsshxiN
gq3fhApzAaPtwKWk8MvoNe9evia56D6b/D7+qsjfe6ZZ6A9XnfTa8W2+rmy+2jZC
eRfMo+SYO8CqCctfjLcI2qXvDBc4RB2AElT8PCrHrwFmrOKAqXN2tcQTPA2nbxC+
VuBJnsLANJd3OweJlRBl1H3ve93vHFiXYH6X6HOO2F6HWx4Epr0Sv4u98phHUns0
qSjTsbLeZKECJWPh0CdMStj38ow19JIU4rGUFN1o5DMoCb98IVDx7oyVBPEWDCLQ
9/syMN+4laGxitApF7F7Lir7KAdSMpdfpyU/ld7ok5KpPo5peQLRXo8oANarbgRB
+ZZBImotMvckGwwxTUORjrcV8BKt0M7e47UCYZUMypDCs8y+Ltg7tPZAMKSiRTAU
LkkdbrouXopKZZvYYEFISGe3mZ7a+/Yzohs+lnjJzt/YrdC+++GRTAQc8tgWwxQd
/s2Zl6EEAfaJrRCd1N/BvC2tzBfAgEa7JKUmR6WjEfqAu8h8k4Zhx4w69DcNRp5P
rLMJAQDN5TcKa83mGQ8a/XXzavkTd1UlVlhVoXOVwN2OABb6aKwjLRNyS8vCScY0
VsGKnGckQ2+YyQaQB34OUQFMVhJzJFJGI3Bx9FiSb3iQxLovX2XQ8OGl6VdPvP0y
az4d97R7F7UqN8VgQloivxQIIPPwyggP2KPJQWVMsJp2ktW6J/8/oDL/U7dndaFJ
zHq6Bi/oUXf0RFqpuOJnNptSQ7JYNn0jDpQUdkj9Nu7Jxge9k7RE2b4ueGIquSNQ
LLVTcaTMVVDz0Q8bpTqCsPd85CLp9rbr0ZlezuMFUQyBsdYTRVKMwV2eHd3bkM9I
54vZeqe2v3fqZWLn5cjHGZZLVq6GLv6Kh2jyv1PZxHk+9bzR6/wFkZ9w2mrW4JZO
xfl4Sech7nInm9kty/AFhrsIFuCC+GR/EM52jzACzgLsdpitZYgp7yernPt+QwXZ
hQy2n3VtMfh9VouaZt6GC1mDKy8ZUHDzb6f61YaeX+aVYu8ksfL1Qz2jfU1CJyi+
nLf4jcsIPYs0Si9kM91C4r+Nx4abstytFBeFRaD6OrkjlyjxYZy8YkDM9I5BAGaG
+LJwcgxNjHEj3JxLdGhkyegmi2WmPyyLzt87P2zsNoR7kOUW6ilBO5IvmWeUy1Mc
7ag8KiHq8LEVtoBif0xgSc0jCf9DFZweIYNyLilXobVwfnUM9IsrfmYdyE2PjQIc
0KDZpWDbc/tIEwZLigPWlr++NivwTu0T76fVs5nTF+lw2YfP5MdGa/DlkmygSI10
t95fVVj4b4N2CVkFYaDD7ADrfYNt+Hko136qdUjitzffkB5L7mArlxDHxdqJvrev
4Nq++ptEDXfeP/EMDMpkZIyx0+QyVNcIzBc0fGAKVnOkTsO5kn5GinC2MPbp1idj
VnymNvYd4ifjeb6MXwTHKpHfFo0pd3Uj3whwkDIRxe5c/FbZ4b9QU7AJoI34N/he
xNZQjaWZLcyVElcwVjomYk1V2yMpa+PGMX5Io+ytzlLUytUnxHFTpYiP+bbjBEFg
eTI8UHooAYK14Tq5/luWzMsYzkc7t+CBgCGsCwTpJh48/ZjcLTLOpieSUKvqXYDm
fzA2LymaLS9rSpSSvyapR962kWzj/dwtaLDW9N/ZQ/JrrhxZU2dnRHPd2a46ghrq
cL8McWffvWdVP3CvkdMEauCOdE14SyPOHo2CAuDstqpwdgD/4FuxOj52Gqet2uSy
9ebDcCl4x7CcFVitrlIO8nxqbV2xeZv8Wlmjp8jzxuCYabq4Tm71bAzkJ8qejZFU
jRYplgf8BcGDoPUn2SPDVuTvvMk4yuq/FxOzUQKv9oPtArco+ZmuttVUXz7H/RGG
TlUk2AYvqh3C8PJhAJ0z4TbypTs1tjJFh8fQT1tdmPb96F+GGKv225il744njpQg
kAdk8lOCqDMZUAMlOpOhM+ty6HYp4tc+TW3e45hgXtqv7D2bRnevev/iA+U3UbZm
fH8fQxRy7w8owtYkq9NSLDz9aRpqpG2oLFsiFvghsT9tVRQ4pHPcKSi7ZjrVBdwK
4slXfAd83eKtpj60tVmV6uLJkRn8FuVbJuhL4aI4DJOywpVKyobZKrSi8Gy/4HMV
qUG72lsg5Zvb1RDGNjkZQOe+QP8ubb1R6+W9OdtAy2Yt9NXGE3U9EQUEYDcBin3p
95yJQJEMfxHyvfJ6n0Kid7xqfwVkYntZm1R+KbKbeAHmS1Bu5PW6LAwplvsgPanQ
1ruMKBctakeLqiqNwuvxFOb0yWScjEp8pP9mtOx08nLiPlHnG7QDABMSFAkcQqvt
kYYgA1eiJtZ0Ep6R1CTAtzA38lN6/drEDXMJ/qCs829U++I5K9WDDLKLOQ+LZx7B
dxe0qDNcBPGloEfQ+w0vNTlKxBe1ZuEpzwLs8yCNkKcv6xxUo9v0ZQT81UTcUb2v
ttRTQaW1rWa0F965xRpEzcxhkZ650nWfSmJfQV6ADOL+EycGGQXJpiMImZ49A2bj
9VgJR0w2kuJa3/1nnd7rKZ19NCL9IoDP11g9HOYNNxjvIMaU+xqriQAT0vDLLFKH
/tQW6sh1UUq2JCGEe49mpYY/nvgPz2GfCnIs5ZmS753MPiZRdAi8+QsvzrbpMP13
JWTKx2/IntjcsqyOgk3OCz3uM0G206t0pXrkNkLJJGJumPkOs3/WAeJVWCEIrg0a
VTEJpM7JFoPUVWJbAojAPew6zyODbdjE2Vfi9AdfHvep+r5tNLzSfE+kVKaRzkWy
FWR9xgvrT73EQiL+5XuZIc0gVAszq1LQLCOl6RK2k9RGZ82edKWlpKaC7B+I36VU
/hzter1jYd94rXcqJLWgRj2qr0ch6zdfRk6uI8+Ecm+vIz2zGf1YQrsOQD5X9ed3
kuo+87W3hiYbJEPWI9OFwWDVPzhvP28ujDvj2ZjCj2uBTdh2qRkA/KeVxGcaKKXn
Q+UBwctSkWz4EmCx8LoTmw2uNMeZcSQyRw8YFCPCpjEGZ2AJjG2srqlK3hw+17mA
53r6XD/xx3rqFpOE6bUuHRx3qy8V/zAe2QOcBe9Tz+zCR9dLBjt1mfOhTTNKUUK4
9AvXYBrTfdscnL17H9skOm0SzqFgSBMDXT1befrxU4Y+4+zYioYLejLZYidnj+Me
LMn6nmW5ENJJKU3T3ewXXexdEkPhccOqe3+A91zqzzRcupri7KWYNLlgmfPCaOpY
W9DuJwAmdrzFpo1ay+BkhgDEjH7f9D7DC/jB+Lc8xD61FhpNL8292JYzAQq65oIy
soUYNs0S1NtCRbxBTZ//LJEKSQ/LCi7dgC1CDm9npz2mrM9J+EGOzcA4aqFpV6Io
xq76wjZRERMc3VzBouoDiO7iRE73ULeIag0F19C5X1DMW9qJ1lIxikjfNDKVcRZG
mrwVhydqauDEcgcf/Gy0yvdyTrkEM/LUMgdOqyEqx2N3BqSMQ+n9GFDAp0aKN2jj
C5nXxBtru29kBBN9c5vwMqcr41z95O83L6YtvJPnoRJ8LeCmeG4OGb+/GvdWP5nn
C2qq6Ys2nNWU3YV2Z/YjbpAn6ho1TXiHfEHy0MLsyQveKLp6NQRO68gEbtKtEGLb
6WL7k/HcfCoDxq1LICOEMaUx7sXg+zVLAM0/E/U418+eDEtFO2Z8JsFRxhZ61cQ5
ZzdvXGIJAUz5KqrlL6Xf3rCr50X2PSdBncqqk6s8y0DEf9D4PYEfdE3s7ILbuaNp
LltCh8tAWtR9g1qo/ETo8/dl8V9ZEZjIcuoYMurXnKHOQpU/qHZxzEvB+V5zb3BQ
4MrmpnTqaGGCFPTfX1pvkarVyivPJZV1ydgBWVQSd9lkdI05zw5a8t1hqTAnJez/
q8PX7LNVHFHC60s9+jE6wvUPA33SkHmit5+Ql4Kd+ry3DnINPZBf0oVlMFnqfmaZ
Tsf7Z26l2NReftTEWX4PQp8gpPrTET2gH3Hl+FpNSgQwWyg9oSfhp7GY1EC4cSYo
xWZAfG55RObWIx+eaHghUgxl+FS1BM/x4L6YAnB3YCDYtGgJnx7yPLeh24w91m+4
dGzIF9Laz3OhCk2q+ZdsattjEXOcMlBgAaxZMTmdjrFMF56vC+7zeu4Isl+e6AtY
cGBrYqL5dA+JWIqvf/ZansfUiXrHFclw6/g0eXl8FqlmTWN7Op/BygsXwnQfhmag
vNDocaCMJrdi1igp5SXvH9AR77xRmeaAHt8po01P8bE6yevSq4p2ZFXrjbElbskP
CW77zi4ozncRV4kpoVrSRUl1oYfhIA5C7l+YHIB8NjQV+1K4qG9JOlMCAnf57v/0
pnVIFmBasvvXLSj9/+W/Obxpy3udJigEV3oc6aX7q9DCIdAGCyu2qqRMC+pcl9LY
kxRKOS2ah+vgjfsqDayQKI6yzJ92ZaaDukp70WdktY6ajQ6EmJj7brzhJPtQunEC
k85jtFQoFujJRwylzlni3sf4O6H+45StxdoWnpDT3wyMHKnXwjtLtzpxtCJQ1XKw
jo0A3TfSdiGCpvO7V9f38arakf9fsTsWv6nvlCA6I8bUPCWe9XVPIMdiJdKyN2FM
35GO+hztwWjxDWn46TEp10fhsaWFuV53kTXSIzHVtL4cOKG8SeRb26EK0DH6Fi9S
hhZC/QAnA8P+yEf3tj4+Ck3vHt3DJfrZ3KEOPDi3Zq7hj40mdjagzZ4T9qYt25+b
K0sSOlF1SX3GdF6YJHvNCq2LtsfMRy2IsXLXN6NyquRhTyaeKTA5sUuqpsrwh/fb
/sqpPTS2/BF72f18fsq+nXHU2RgGs4ZZCAXJRKtZmd4RtSStAm4ods7sLVqFIHiN
dAyGnJ8D7GIE7IZkXM65BpzzpNb+OhzbhdNLMQZ2HOXYhUezTteXlFPC7gJrQV3a
HAtRpNchFhBStTNd5440z5LsenKoTAtnlGnNvuAmY6knxEMvSZBK32Alb8sLUD3w
yU/k89XUBGtdK1UrKzMdtqpbmKxCsaPmQfeYFLXxzpmekBMtzjQMXLqc1k8JSOnM
FqAO3L8qneAtsghJIAVihTtac90BfelO6Y06GUECIAYibSual+wFY+5YTWpKXW6p
lDidU7ge11V8gx0WZ1v7bRfJVab+Ze0qYpYDu6CEFthbqjt81kPn10oEXRE6oGsJ
fQj4AUHpZbsfiMBtLiZUYNeFdoWVa1fDS2XiWnFV3zziA+oObwXEIMwrx9COJCX6
YoybfNj5rXNN4p+1Y/YTLyyLq1EiRPmtoF/MJ1rszxfNBaGy20/6gmXbGBcLiXru
Q8l72vOt46viu8cuWwe1NWHIbH5ev3FYR3SF/RhB9SbdPXHbwLm0pVv1kmu8aa60
LoOCrbqHSdQwb2vUJPSvXqKxgoE7P8iD7Depa2So5ibuVJdANjAizlswX/oDsz8Y
kCQh1XpFda8isNN3O7gw9NI5JI6vq8Zaadb0jZiO72THb7vvneKr6UkMj2BYDtUn
/TFM1lM97fZTnCMJpnkERfzLJM9C0LfQhd1YkT3I/zPhkrpWW5hZ0yEUYdRwmAkE
Ax4XFopqowzFlc2XcHC3h2uCN4094IeFHHTslFUMSf0xyVa0szGYgS70lywFMgXw
uQ+KLfBZTs/GGqTc6KKxlSYbOnT4jCLWxexP7V6rCH1Z5gddKGd7gDZb08tbf6ac
SsQsSkZQ24wmP2EttvKrOeRbCqQ9zVvW70Ez6CCwG5q/fsAyEZDcpLbuuTGKzn63
9jp7oXepywI5zDl2jutZJtWrM+rBGc5k+KZi0CZxofVGeCVWgu0I3aOm34qXFu2C
eH19TAMD98E8s2NVpIjaz+yrQWYPi7v0SzwsN5/hftJc3kfaFKaw41ctCOD+n3XD
BRcaf5M4Quwzt3ULoJzpOtypm6+sHt9hyEG0ZUIvnDAfRveDThQf+UC/mrVhjBG9
hugzVMWb9b56620wXF1aBof6NGFPbK66e3UuRgZb91w0z7zSF+4T/DiNmkVVvKDt
5Q64m1n7JXBItrQt7P0pl3clcv0Saq9otNuw2NRPFCPPkVBTHxlGTOGnT2914JMO
5rgLVAPL9PsrBfZEIHYk3dSCN2/Quwa34Ph9OXxNYJC4DthtxewbFHZ1CjaBSENS
OwFnG19rEmT5SazSKVZg5vcWBy+aZInYDUO4W+IW4pRkK0PJ/ldSBw5Lf2Hicggf
4lKmJXE/ZZCdD1qgmbjGDQoebqT3WrfuFg9o7P9J0HHuq2pA6374NytEJPxeuuu4
AWz0aX7Lub9I03xhrTPSjZTSxj/+153ujisLFtsrjbp7+zXIKKV96NGAPQoUU+Bi
prChOSWkAf9oyCEip53Idw2Zg0WfmRn1OfpEHQ0hZFeozkFaRYotXU87C8zfiTzc
28hS34dGSL8273/JhGvKIei+0QKE8tOQ+G+mWsXiUUKB4UT/GymE0tbg68wsn80g
2PEWwLUmZ0YzNHjM6rILRT5sCXDIPE0dZrt/kAufxLvNUWgKq+G+42Vdqxr8IZBK
d38yrrS6ZEC+sDjMFA7JEsW4cVwF0Bai2eEd2+fbbZUMxzZ0GiQvV/WZUIPU1MG0
IIIvuLzLI9GuzMp8Lb7W/DKL+nLdN4UUQ/QsltOfUFqLwYLkZLv8hf0yJMqhvJ4G
CHVrl7/4fyBgerkaMBG5Z8hi7eTJ8tSp0TMCeZ931j2glmJRA6YccYv7hVIXGis3
lzJKlgDgySIZS9ddEcJKrvAHJLX5rRUrxDWK/vr56ds0dzhtTp/WVJIEdiAzIKBx
dR6Ir04SGDPAhhFSuotE/Ow9OcO3zAa4fz8MTzy1bV2+QGtrJHPUGSarYLJ/9reT
7OMW67xpoqC9hzAiJWhshHUe9bdHV3xZcOH7CfMGcpmEZK4uRA1Ex2zyR1JJrynr
DnH5WmKziHfsS5Gv8BgTXZkw+uwwZ3j/zSjjYt3lMQABPTjPcnMef5CUVytExXmL
4nXbG3pXg4DiUez6SU7Fg/Gr4Tz+G9E24wBJ1sbhrWwS+mp9McObvAwb6vMfYFe9
A8zWsz3uCfNwo9Q+6s3Rnh+/2sSi+pL/kzYGb+On3j15YMVhlj6TzDyxsGd9EMv/
2DfE5iWZCd9oBda8NzrdlPz0zRLjIIrq8/uYkhwmuaESrolsrSTgN8NBoyjtKEeC
uXxo10DRaK1wEJx1nO6tT/P6LaQqVXcm7KE0DXlbtBaAeZthLInJmxJuundcgUd4
IBV+mjVo69T4Y5YjjWx+CTGMLvPgzWwMqleU5xIghkyz2LTcQJ+f1MLCQbO/lpfR
FKOoi0PKn0EZ/fNL0ljg+nvNY0G8uk3Fr+uIsm4AtjvT2qM8HIHof6jGlC77Qbvp
09M/ednrhBtJD1bw6qYL6NqKUOnLC7pKtqamxVx2j7gzRaljpafY825KTVdFXePy
bMV9K//4Ez/bYNt/uWSh3weTcpY4OonVGQHXUrFos2QzxUHz4oH4DwYbUY8eejdt
jyyFEIEfdUBU6i/TVZLPYMIkJBS3CmC4aM5OM6AnijdgmTs2vK6e+FgI3ByOaWCe
PmlJXMpJNZATarN2cDqf56Z11DPmh2H6cPyBZzrfclzWXDMYifgSYpSIzT8IGGRO
gfT0zSh+e3JUAru5jLmRuAmccYbJ1I2NMfJqoxUp5YeCev3xH8yfZIeSnilW0rN5
TdhgHcipCTTAveUBLJa9OLa866jylOWVGqoGueov4ePM4cMmPFl/XDy+xp0jYoqr
vlJGrLUQEf+eK47FlvmmeVC3TIS2w/W+93jAXln74X5xKp4UQlNQ0y1Af1fMzlyJ
I8/7ZMTAJjZ96Mfgrk1ii/h0XHmqNz3fTeX217RdLesEwoe8JD8Off80n/JBihwB
/lUGtEl5eq54HC9dvnZT7ZqISwtz2qEwmI8V5WqWK4nqcCpOoEEzZcuKh/UHY43A
9mIzsGhXR5J+oRhAHnVd/wdkcF727hZS1T40ethj15VXiFbC75gFHEGMMogi85y6
Dra0AtjblMbcWozQyxVCT6j0D36rS/TRxOMHjGM1InrB8MR9mA/j4rLs4hMyao4g
iOgOhy86vjWVDhF+rEMrDLEZbCsTSaspYMDgRJk8ycme2j3uoWEzyJhfCvygBhFk
xTu1jnlPGQo3SrLMk9mnQa/YwP9hN0IL6Vs28y3VHFslFDubS3cC8BmweQA1034O
v2qeO2zdrXpYDSWQZKUY5FzL91cGNnby6258gLvpxmSAvNnkbql0vLiEfjni84zb
QtOdErY4NTssI3heMSZn/OQ2/lCjGuv9spsMpjDErQ9IvkEgwijpIFMafPqYdb4V
4G8ooFM02XIYCgHA+YzTycUXqDy3EpwgwKQDvpAqUG9LmBnXl+heFFXh7Vc9UGFf
ziwZBsAjXbkK8ughsYz75nmUfP826GNAsn3PGuXhLMU4+ELwfdN5ScgwbeJ+G0Kc
zznXO/Wka5huajfi+7Kg/2QWXGhqz4LZMa/1lA/eXJDOMWTanila4jb0fLA2bWFv
FTnTjeYaVh7vZhd65lJ2fk4A9QwZK6VLi3dHVaOhCRGAR0/trnBCE4uGizTlhywV
StgbOWOH3mH/bbqYr4VBVWr4TGgqc3syoXth1V+nlorxh5d5Qx2V9bpegat65wep
0PS9mkpDQFSv4GolRtDUK5ddetPolIPh67Fdv0TEdcK8PXs0drSxiZBeUS3Fx53s
XqdEYqbR7biBsZaF6re4oaXuk1bi++h0Kts/9tsO+yjWH/yjQDS7qAM2rup/MV9X
W2S5RRlJt68PqYqkj1eGCMyIKAwyKG2ajUgA7eJAnZJWj6GED2yFzBCSiS8nqR6Y
fJiU4qP9ALe5x/7ElQoWGpNLb/9HfGfYi3/jztJR6eniUkp9GWnr1wUU635RcEMp
vFASf7zqpCOp6cXkud5LsPtx9HQxd2/eQuCPbfK1dUCJudqsY5LOAcLL7JL1gfTc
JWC/aB1mr9Yk7vrWPdNxS+2rFA/oYjdkYGl9Si7UAw39uK9MmAl+ZMYloLTBzz5h
c0Z+prj+zBfrgk5gb5/G0UMIdzdOARndN/xB7f1Bpt00Ia1HiblyLK//oCcQBVtO
XRfTFfI86+u2PoGJt5QtAe1rgkmn4hfTk0a+K7F9QSinHzBYcRUVuvHPEDAcARjy
On3S2Ke7ch5iTRb/z1Oaf7zsr+7BSuYJv4GBn56UaSL+PRtPcaG9tCKvD2L+NH3E
0trNqZOVf2ICOmeTTykzUzMKYsbJhD+RHlwALXRoEmpJMRC60w+GXaFJtOwUg80A
Q1E0arwyQ4oKE8l4Ue6SaffjVrza5x4DkYNaSOKrBXVP/0n/ojnvyXMgmyryaulx
7gqlpPxohO4dAlAYqsgUUJe7+REll6ie/+hF7+kuKx1aZfpWFea4hgOI1pqsC89i
PhteiGtGewKzyQeNP6YddnRNGBvB2YPaNl+LhZwdI7loebj4/6gbQSVUI3cIqpel
CL/iXiGXdL4oweLdkX3jsNKYqs4ygUZEXRX9pAlX3lw/2Sd8q4g9HmQnSCcSHmG6
8Q3U9vMmzX2hLtkXG7Dqnbpic2jh5vNgLe6a69xPl/Cny8DRAwHlXQ4+C2KDARW9
pmwU0/TrITsZ4u8lSieV9Dntq6Y0sQBvkr86L8KIRXlFfsXBeuYG1GHsbm6uPjWV
BXR1l+wYsxRTff4tV8a0JwIZVcNK1NXe4ZvqIUiaBnr2K3QGH0xLmVy0vlv3oK75
fNz+YLaOX8CPyETJVZ4i0G5iKTS0PUbFF5rNW2YnKKVhE/HbSUG09uKbCw57Wwjz
Sl8KEaCkDg+KntRuap/wPrslUb/2QmwSYm1JbZf2lMquV8bZ7HUDb9zx+xTYqe0U
XFP6ke3o3xJbvb5+lGPvJXcjDgPf+X+Frit2lJ/XRBlFmtPmbGbV0YS4XglpdbiZ
NkjXw2AENH5OLWGeki08dYanvd82IQL9ITLrZGug9DpjgazaFWchihOy7PMgRGAw
2Bv/kGyRzH9U8b1jJfxpKdxB+AuwymB4K9/kKqT3ifpRUwl0ACadEkzWJ95/SlDJ
J9QwCvgrOoInQGj23U6h6eNWwCwQtpbDFCu/9DGPdThvXUD4JqcvEK6/LFYQ/EUI
A8ycBOisNcsWJ7PGmLKcNTNyozqQHM/ZlflhS1RNHDPpRCuHcrK+94NnB2UmqdTN
rAsjhNNUw8xFXSHByUJDY7nlDkZ222OcfG65yIs8da3KlLih0SO5FRUh+FZumT0G
4A1bYEeAJO/NWeVrcqd+UykImEEFEZTqqgFrYIlK0QHANNNgnoTlx0is7DDxQ3Xg
PXhFjgWyuKJVFvq1y1R2R8Nk7qT5QVjio4GxoC9R90v4ctPNJy5q8CIiJTwrVuxC
VHVmzS7QnuoH4rG/xJMdbCcSmncqL+emC7SVYKCB5fsdLVBC/t6ch/9RhjCG935a
SknCvXZZ3a0X3OxDtspBz5z5ip1an/N21D+lhi61Pc7vkPEusEEmsVpS7yD7v+XR
zRMFvY6nJFJQ7wC+J9bSCnDxcfMsBRenGrljKdQ489sgPTx+MeshfrGheQqKFtUo
uIR5AzxvWGdyVNvTKikq46Nue9ESHnHywxAEzAXcSeo5CGBURJYw6jL0w2t87Nv5
N7UIFsSc/pY/ADtsUOz7Xv7xjU3QrniH2QY+DLdPIAhzA4XW3TGZtNaq9dB1LKJX
vg34Cx80hRaRHz7aC4cCM5xa3vyAqrvBNqgfH6k3eAy3CvV3nCQrTtV9q5DrfmPC
a3fFBDZHe2GjTkM/ffl95lcg2zuPH+PiCe3AiAubYJ4OZvY5Lqy5o9X45L3EE5cU
Ut3YMy4MUEo2uLCw5hl9CAsFr7BsIYildAJEzdwUCJvsjbpaam0xQtLl62638eEV
XrmKHk6mdqZIAk/kAFaTfSihAZu/LnvfXTKHicDfIZPaZdHnXjpDbdod3FIVHbjM
Fh/DKd+ST4LZwdNAif8YxQ95f2KrZR80SPW5gi6y2P/54+8KounLR4wzLyxqaoOH
p+tmVHOvzWB43wPJ3o80ceuhVyTVKH1GnMzK2iHkiCuvQ2RZ8WD0Nx86nCYgrkxR
aTTWLXXyJg0UeTx/EHG7aN2kEdQE7K4vgxjpGype0FXC7bawMioaebfQ9i+N4sCJ
rk81HUXTztKMMZL7cYhAKyqa8fIkd7DbEngwM7uli/g4+Lm+ryTSHgnAkb31YO+z
y2S3dMqT0cNRO0FYMRc3nLa/pKOttZj3nNWzoxuoTaNYjFjynP5rOY0zE8cnuFh+
KGvNkHFfoBUil+FXTckARwqN7BuDyG90O8WB51OglJUrruPsl0sgMCUv+Yu008J7
GHqEEPFUgd2tUHB7T1yUuSxg5t6dxUSNXhfbNzPg5fZ5w69B4a+J1NaHjBLtLzh3
TFC+0KEJgrI12pLF4+fCW+5VH2yqWBQCfQQt51xik8SUxIlWOiwqW6uAkE41z7Bx
WndYKqPA7/J2S5aOHi7FYtAy05SB5xcVrtoMgQ15xaVgS6sxnZIB/572GxfD2aB8
ay906oFu/GgpU3AZyCpLvtrTCx60SVPFXDSHw16mLU06qbmOyt3Q0Z1R+srM7TxJ
VHUEw3WqsNFoLw69CXDEJB2gEVCj3+yum0tnaRDrCfKOO7QFAiljg52LOkMFbRt5
4XO08NAss7qQVmAsOGNM/rKtvCjZrfKoDYnuH7rYLqiH6lhaSW2BBYlfYfDw3Joy
CaDsJmK7FyQuG8JWmuZXfg1AvqO2pBknC5NuLFemFkLCy2YHz57yDp+fL48+nVJG
3V/nMQcCi6Q5G6gtQcemlWIcyDW78cYOABvqHdpQmj9TgSQY768Bxvru82gmuD2g
AWvuATBaYbUFqvIDobA9lKlVhA9n5TzizM4oywtj+leq+Dg0VmYh3PBPMAGUpMRR
ikUNXG87z/qfk7qJCmE4nP2xkhstuiPoWrCLyg4CoWwL2X+DYLxSKRWzAPrYTER8
zoA+6eyNntTMoZUwip38OasdIIHud4Q3gbKxH1iS+btab4oX86GG6GCkeOeacyqr
UPl0B6s1KL+8hs0WAHhHyZ5T49Gdib4SLrC6YrjK6nFv0u3PVE2z7yZaB+fvTMH/
HD4CAHs7X7PSDq+/QCz0QOyvCZvOVPn8fsUAzGzTIzMNnxJvMw3vhHOjd7ODr6zW
4FV9P7O6mXOJAteBxzUCUUYzX3msZSergqWMh9OAXbYtfryQ8aeqZEbo0Pr0s3QO
pEkaODKeXPlY31/A4f5SglhLd75HNdNqFFg5y02D8+jZ8NSapqZirSF8HW1SsCYp
AVgpRrp01lKVriMX/xTvboXRbuwIQH8HbNySyhbCH0PODAdV5JAfBtZpMektXsgM
7aQLbGwsFihQoGGiPt+MMQ3YnK3qdUQmhXLs3KKtPT2T5TKGQcztXSQW6wWwMJu7
CkOA9bkEqpY/+1UipDJLdYRk6CpXUKAmrn62uhZaG0ezBWUfeF+pklB3OFUt8MCu
iXhAc2XFjSS//4MkZhquAqfG7WZF8yglyIsDO7gmIpM+pqjhtBmKGG6YmO8wKxPL
dElAn2NM02Zu9srdhmmOzszqRckk2NYOkgK4fcF7EFsjG621w9TjJiyHSDVoENm5
dkg8tm3ZDSIrmvOXlAhnOs/LHPUFKFuwBOC825rk3ClCJBtu8gltcJUxcjJJZF7m
KOS01H/Mom4V4SgbjMIwI8bQNaSJ/aCzl1yBUjN6wY4i5eE2YTlukYPHfF1NQDLU
ize1XsU3jGhlKnhgfoILIZp1Ucwifqj37zaLFqzEuXVUbj8B0JoKb3jYHM17LFgc
m1tW6AUfArsBO95km3qb7ats8zW2Hp9pN9ox/CzB21dqFIXQPE9zpLN4iHp+G/R5
86YVI8riB85lwJRz/Gxu89M3dNe84cSwc1ynGExmvJA7o/HVMF1FpIVbiy3OzxRE
mzzwWG+EhP94qcXiQxd7D3lPJ+6hi9XnVrVGYeMLtlAuZXrM7bMqT0oEzoHi1SY5
JKcnI0kF0A3+aPjK9ZgDbO8l0/d3msv7gAqd5UWeWoJqEcI+GNkyJpbBrQwRAm70
bZjAU1AXMSwT5IMxBZ8vDEeM0j9kkfJKDyl+3nUheOJVa8YCi8xd9fmTGLj6js1C
j/G1JcfvIbcYk7lHHVRdtf307jx/ldzVxk8sBF+Ow+t0BAnN+uJ+MA+NSqHoX95k
6riXcxOflObJOApZjppQ6RoeeJhZbXv7tBVmE0rSLgRPgwRSNELp+JuDhN7z/Dp9
tpmV8M+2Pw3+Ce+9IQcqwhT+Wifsxy3rPh7diiYKink6z97EXVcI8b/Ch9Pb9KrX
vDqQy+vXuFEG5a6Ehdb6Hc57++3WEBs0Kw0dqMCpbHNIqXaSdfePh3H4OTQmvFkR
es1VwAXGWTVq1W4oceXWdBv7ni/78kjClsuCqbA8fiSEMqH+qEmTP06MUUKH3nJO
uxdbbfWbx6ylF4JCnt2sxnY+77pO6JFm0ir9CgRRSCAZfPqD2JGtdIL0bYavfxKi
MsHztSA0UCf/8QRAtEayMwX8X6qVc6GmdgNWk7GXS/PDYCh68JporGjQq4xds9UA
ZnLjGKwenpJd21UA4jvgmf5xWX0Y9eLnKFOvbmQipB8L63wtfJgxTWfFmlryxkxm
JQdq+TCeTgdIWxN7MJmlmoH5Lw2Kei2Yq/qK4zMF+9AcIjKEl3e3OjIpBcKm55z0
bH5tDj4iyxWd2VasAHO/Q71GsK7k447g3nr3NdSj+BLmoOJ5IWPoowuScmaVgRo9
7ru+ox1Aba3M2dfrOsVDGzgKhiqGDu50U6HKMijXRpgvIgnGHT9O9buQN4+MV9Rr
p4eih1+BkaJM4yRLT/jW6LF+qCLva2zsL/E7Y22b3Df9V4RTs1XMHsyn/QMh9dFE
ifZ6vUv4KIJkfqnO8ej+ueNJPQtSFe844FAvy/QQkdnjY9QSq0yZ1izOw+IE81dG
4S5UZdw4ZsHrcYt7T+Yrx2lphexkP6uwvGcNgnG8PSm3SJg4+FB8vAfYbES/ZQO/
k+tqm14XPHcE7PA5ZoNfLnqAmcUQyBq1Y/mFC24RDi059JTXAup0hutHtqY+WQkJ
UWckD+UhXXjnAIem0M/O1tnoUdYccByzvTW3M8XM5rbKOO1LlARa5aVsRW1al/xB
E5m85hIUmou7UQoRYysv2b8sT6rgZTIwalHNJBUy1PeSFRwOp+1nUXuGSJPW5KXJ
reZ+MFNmRf7LNHnwT+Gn1Ch76WDbaRO20sZOxVDPubFdfqiWihonXT4qSiscXLbh
ir/1My4fCoSS4Bm4uNeZsk1s3v20hjxiEKBWBXWGC3ESuOBNgWU01HnbmtxHGZ0A
/tyESjl3+86sG8cx0dKWymjWY4xqvKoXqMNLc+0HBkdUbL56E86Jkh6iVfnV6WTD
ubjCOB+V06Oei8g1NeqbPM7rV/RObvXcV6IHZ3ZBTo0RJbwKgSt9ReZ6iI0/PMi1
Xrjpb9rHP0YC/faRWvLtXLu4x422WPGJHmSIdaeeefe3OqC/qwwnD8MiZ8ieC7AT
vDzUWdDmreC7hyEbsIuIYnFMAejnjLlsnwGs6xmCVjGXGoZUhikrb9jfqu1ml0BX
v0O226nOVNy61dexxHHKmZ8QKa3eiatOSSzgM2e2Vvj1IE7N5HAf7m1gzyC/NyuV
aTx96gmQkOte8nwmN96mu253zhuhqhvBGxKl01flu6kthgq39euuQdCYkEkHZI/j
2E0ZoXXjCPjLtYtfuNfkI/IWUgVh4vL5ShwBzrh8s8u2H1JUmnTFUq6qcwWhj3uM
1wuk08aoC+AEaVCBc3MyS7xWZ+WUZ0ZmO2EQ4SYoVCEli2jmu8yU8KlORwkGXz9b
H7zVkjXA0Yg5LNTt9iIM5ueKn+2ANmog2rbC1Xm9Xz8OdWFIviXv0cfokifp1nI/
8eWq6j4b1l8oo8+A7x3bIwq+v4jGSquF40mCMlF6uR4uTBL1fO32nLiIj/asQBF4
wwvfhatMRJwK73fzB++qsvk0RxYtrkp3T/A9VeZJpFZXCgdWYeU6JU5xas4+lvFX
VUOyBwzi1vle+uSCEJEiPO2JcPikvFsEkMXLZczmdqAd+cpyJC4GwCCwhfOx8L61
L2S6hJdrTQdgmKabwB5N1PRwFwfvP9RW0O3ojHxLZZt2kYgWYNfZfyWm4RXB7+71
BoY7pMwt1Xj0QNw4bmJQTINZVfiPqtBgIFfpfbuH1+YKxviIzlspi3I2cM53C3pO
ZJc1SUfk39M7YR55DlX3/tEJpfOsfXb/2A6AOPRZO5WhbKKRJkz07z6Vofr95Irm
UuBNN+NTRxfVrUBzw8R+2Kp5xDAQB8MSNqBbRYWN/ueTCru+YtKG2vnHzG6CXCRo
lxYNP7qHqI+07redZihKc3BnrsS3xcyE+Mddk8+4VnwKZOIw6Fsu2k8//JrCEnOG
Wv7bBsG68X5rth36dq0fmoeLK+FqRBWctgzSHGtnttCYiMq0ZDMhgBRsu7xWjSRa
M22qSszjaN3a0+0UC3FAtXOzDJr4lnE4Qk/vUUHJKfy2XadJQN9scTny4rLDpeOp
DMojqY7nruceOkYyC+Yc/BThSxVf2DBVex1VQyAXRWn0BBS8e39NNUjzjCT5twFX
w3GNLpA219v5R6f2rVDpUEI2O/h6w376xvpRoDKHHrRyhCwBfZn8CPh1NjRvF/PB
yBDBiD7hSzYHGLP9oMCGFQgTNvhOxXKpe5886yppjzEpfOqpbv+QXky5/jMdWPSL
Nw8+Czpw3CV2Ti6pvMNnhndBFLMu2r2ghJ/B9uhrfIFbNUe2AivkaqOISEDF0AwS
YSLhXYWU5kUM9PlgZ4IrcYZH+78kVHiIgycmD513fXwyDSm5rQK4ESsXQigfy40e
6iEQ/gk5tM1qAOb83ostjWprtIoEDuHp2z3NRSaYeOCHNs0GwYKwQzDTe43hYCkU
ir7rrZzKAKfLsYADICV15XkkgnzVW5hvZRCCp4Dx61w3NAhH4JaSAQdmKvix/v1j
zJa/6MM/Eg8HKhgm7w/0QLZNjIxfv/1Cjr6+EqWIOAf19AQU2eP2cpZ5QayiSBlj
CCw4khWn5OutlMlATlRelDFixKgSp+0uMEFe0j9CHhxadXt2BpyY106lZRKNN8pF
bJ8L5WXDGrZw6kDu73yA7dIMZVl/w+MWaYJALdzodOZC2wynBTCfEbcnD4U0e5+q
JzI4iFr4pKvtw9+b3lsf9aQ7AjvhDxfHG2yQqt8wrNK3yX8gHQkh6ZIEPgWu4GnG
lqMl6ar+C3ttEeitv9ALFw7ih7obJvvAi/TtlDPgmvKQGExq0AXyXIgdS0ooVOtK
FYCeL7fuBTXSD4ePc468o9yqprDaQnK1mhAOlVOIoeu2WLQ8sILtGTiFA9EqIG1V
146I/JLyqA4rojkSoOGGVUl0AK5Ynb4meh1ynO+jQWPT7B4vLIERAG5WI6TQl+FR
D1TPUHmZuJIz6zAVwwQrFmDWlAfIcQctPfNvV3+EAVbVGK/WK9cD5Qfncx9ZLHEa
w/UAXQHq6xR0yi1/2GrYvd7vhgoYlfv6j7+riz6REQnbBuY7BoradGEaEMfzdxBz
pKDN8j1aqvz8EgdWpcUZcBZQ7/qSLYb1MnMetVHgGVLnzwJdF013wI097FuapmlA
4RUtPS7IPL/s/svWFLDKGvYTsivqBZ5UfoaZ6sUrMu9C9eq/z/uNx/cx5aYbPk7l
8oGxQAkEe8JRWfdzfGSFCYHDb5BicT1M6xxmjYDbUC7sOjmbWicKtxR/dkMDyb0d
rm7BND4oskv8cdNsrD+QwxVWHGG7rCJVcQWRDA66FsLG6XyzsYXAS9l//16Al3NC
eSyu9vP09lYYRoINh/86JBcWVR0mZv536KYKb/uQbDFdFr6vYXCwHJZzpxQZ3YXY
BupJhv76l3EZnadbuELmWL1kYwgats2dbqGTRjl6wEx1mHJNYHuK33fBfeTIZmH0
gwHVIRUsF7C2sMR4YtCNBk6GKmCa5YwoQ9VAVqZipO5hBa3Gc6q9M8QsGQwwI8XN
XOItd1RC5QrcYs/ufvu7mkno/xDs/2P8Qwof3ENBBemFRNrG//gMOQKffIoYBRvS
OtSr+L31cQvB6LcUnehC2BdnAdQyAgCwV9hPbCNIKp3F3kMajFcuv91FvBt81JRG
4aXlW4I3ZYHCiHvX8dNswMDSxFwGQMeWm+p542XY8wZAQ+lg4Fh7EppKzX7J8RLl
Q4DEfnVSrV0VPYZHstUE7UvNjgDeqNxc2S/7ez1vqhRLZfL1PF8+F80+zMNVpads
WcpQGLgReL4CkDi+m3+YtaLO5/Ji3Fa/7ujQgFeSGwad6IYHSMOfjCvqXr/ytIe/
jeFPvODWUM2LOzYAv5aWO7jId9PXEdVFKdJ2qspE3FNdvDf/ExvddSJd6UG38D5m
qgjjE3Xas8bhbYPpSwED0YfIQfiPfCrH56n09cKfXarF0Oaxx3ZHkNuykpgEwZP4
g1fsjwMj//EM+nnPHMgH324Wah1t7y7ag/G7YWTdDfMGui+xxTdQuAMuzYTKHz2A
F39KBl1oukSBPJK/JL1Mq8G5wvoEkxfqu5pMorItWTtDM+IoNIrGvnmEv4ZiXXd4
enNBxRHC+5zscZZLtjfd0nE+zXJ9+O5HVC9U/M29kbV2XmmLBmlcxHvofLh7lBWU
0qV/gMXg4ZaVdnfqerKb7Ny29VEeiqWQZkyj8cxINmNUYivPEp39iLQR5b0ltIJC
850W+zaaBkAGn+1dTJj3GZ1gcSQLAIsoRU70xHDBqlfznCf8BhQJfuXRzCba87pk
ojH/8S//rNmbAGV2+Wzy48VHysBz63Zmoe6fRkkb/Jt/PNhd6kjwmVx1bbQ1djcU
SsT1CTjMNM1GTjaxIma1Erw6cHy0liUujSDhfWHl2tIt33AW6pMCi7DSaRAAE64U
Z+Bj7yWIX8lGtAftbW4xtVUAuG2d/C4LoTX8GuOIKWQoskJnzgqHcK369q6tq5+r
RWCUKb1kdV7+QGnvny/wIV1nzJQbbXj/01W4uc+Mqa7CV2SkecRZJTct9e+tY/Kj
gBvIK4Jk+fRxcH0YUVoiPxwD7NGAvAszfSGwExAdsF02LhK3wcV1o2zu56UB1KzZ
X9/pMINq7C5K2/WjssbvSh1UeFiGsqnh/IqBv2oIKQX9GcH58ST4Qt/4WNgmuSpQ
gC3XOsLomtz+Zd//rSbaWXRib11QkovWegNusQaCgLctz+0/Sk3rtVqRB1WDZrX/
Lx2RmmwrVBthoSXKVpg0X64qS8DQKZ/LP9JyhTyBNR6h8krtl+XeE0fboCazSjt3
lkLxjVVLk0t3Y+SFbq/2Neexo71nUMLIusixtBNJVROovaADE2+kC0u8o5Usetq7
iZKBDntsDjO/nknN9bzYUnyfKw9vvrceeAa48GY72tYu1R9fLnMge89izHsEGBBo
e52EtvZE4y7twUCm63ZlqoPdTfDYkUh5mvqgH9F+w99NYK1PqvArNPeeEO4aPVS2
21KA7eqPiQFq+70jdI/j285AMon1uYXM4FEXCWvrb66Ie7OOC7KPMmp8H0KIDugl
KxG5m049sS4ZG79AIKO7RUmTWQL3b0uA+cdKXKwjrwD9wOIg0aefpoRU/gfHzuFt
75TrbyGviR/cYCfezMtSLDcGvowALgpejcgtXWXZ5o4J4be3VoOuWQPif466aIB9
Vtfrrg5FuTz4bWH6mkPfgwTJVhWeGznP0HPJdZ7wx3vDM19HD2Hd5gTS58iWDOgN
WB8aMgXM3MAIXRtQ+HVKL4951ZyIEwlUP5MyZd+xZYyFnYbEwL5MiV52cBDcgGW6
gArJfJVznQTdSWm8SWm9GkcMW9jO51Q6rN9J6tyEjnFn2jyxqfhLJAzpoGZsVU1/
p/uHLWM45fMab4R9zT6y4tTAZunFKbfa9VkZkC+3usEafhhBxgSy1JxMu+wHQfw/
imUhGJUavYPUZEqA0q4GXP/lbQOJOnrMLGV4FZ1sZ/EujZRW/O2YfxL9sbDewKqc
lVumtWDD7PGi7l69cc4EAsRq8mNfC2NvKdvRmqX1lUlqG6dzha1CvfMn/dsg0gse
BduT3TKxJH5AnDSWWoGCkpoDuoBxGIpe1OazkSS2IyEiCffkJgTRcnJAnGVwKncR
4D32F//0dxbVaI2cf1FJoe6Md+wz+K6QuY5GMu412wtpH7V1gNQ4xkH1uwXKEs8n
FJd/PyygZpE4QtW5VS8DCLq48OLEurrc1y6tL+txH3eYktV3ydYohuXAM132PsBi
pDHf0F1Ftqq5kOB2RA5nx6Aj5X0CbcVLp7rj7MOcTGiSzIsZtznK+ERrttbcuzxG
CNblJ8FLPYB8vSzR5n1ESp5XHVFyEepVfHZkuFNixeDgpQyRi8YMilZeTUrAQxPY
0Z8WM3iAFbZVZkoJRu8estXPLYPebPJA5F8pm1QuZlzXpDFkLcmoOec28++rE60t
HVgx8WvPKfZ2AhB5cjtG0I4Mc5JfIFy/jrHGvhZeW/LgqXObN2QLkxfb5tMI0pxG
zO+VIjU6JsLrvrfO3bJ6XBDajzS21fCZDtIruVtX/bR73qawYxBi227QPs02KRxK
16FwIvy2ioiXPtBXld4TFYpm6VETXk1/Yo7wqieFjvc2/HUAhOILxwsPAuATjUZ6
lmbg/KCTtOdhAUewX1YFugxX7e5xwCCIAJNRVFajbk3LDT5W5U++HljG6S9P5WkY
NDvABePM2xdrzH8Li8SxHlBJvqPeomvj/8tOIg6uQBzoHFgoFZ7MXz+Op99hyLa1
BSLSfVzV7mE+0rxwqHd7Dow8UP1SyoAgjsbk/hwhE/dCOM8rb+ufEn5pVrDVo+Ml
ZE6ENF8Xh7aXifEusgIWsMEr75mSt6Yhs6Epx1sYZDi1eJYcK2pi3hZlAv2rJ6lR
xpk0PTYMNJxDRkVjiZ3jf3LBPIzZqtzd5uLXT43Jngbb28J176aXxPMP5cC5CRq5
Fa55/IgkNhrvtwXSJlRJZg1VQYZIZapwsUzTidRT+BuC9DxGbduzUiptjwEhiPra
SiFolk8nQLQREd/1Ee2rb7qsRrdRLAm8k1ElqTT3bWqUDrfv8Ush0bI8SLXIUUpJ
b/Z+nMzpHxGnrqBrdBDV9cq07CJrf0N6LBB7plf9X//aCcU9Zz6I6JbZiVIAJI/O
IXv73ZEdIQz22VkRPqvo3R+NmQmQIB6tEXgfCOmGgCyQWwCiwkmpuWyOQXc4uPa8
oppKT3yqEMgV/FeOgkYzp0NdLGVyByvxLh9sCdigcMHOBVJONujMxZ/RBsiF0Qeq
eSoQN2O07up/oTcl8aYpWODWdANYOKhI2FHWjhpqo61K8McXsx6UfnyjMNoGAtg2
UqLr4Wajg90+au3G1+vuBQttyFvI03qKICdunW5EssqZYlPHJOZBsYYXIWtg+f/T
Xff78bgcKik/G9ZPnZ2noFiq3FqrkPST292kl1uBrYcfU8B55ao7LmuGHiHOC9Ty
sv9rcPxqd/S6a5h7R8ZGNmDOLHDUfEYnLdnbpHeNZRpTEmWNAMCQv1hFMLeli2k9
Au/Ciy1BK+5Xezqe3n0Myj+trALM+iRE6Foko1x7U4YhiYRb3db0opWhZ3haEcPu
d5GBnFsFDQWNYsLgBqlXW1Tw60xGiPejSkgeM0pVIYhjWEKWdeQaBEpqg0GSESKW
BATsdwyeRa2naIhokGBo7X5avW1ythKb59JD1Vwm/4x0kmSBXCWn6cYFl9fN8P+j
y0lIeNx+g+dnpDoEEz5KGtPmLu6zjDJ/Go5wEs/dMGZNLxuT/J2B84VetB+s7Z3/
FekOAWdO/kggdnx3AFikrr+MAxu7ng6bRHZmKDNZjDKeCIlNjl76Atv8mL0TYOF+
j4AGeOEJ9cKmfLpqC3LY1rbFE4he6ncAHmnrqFGaTyzq/7fUfQY1b4DZ0tWXZ6wN
CoZIZfUKd1a2PIKIjSH/n5Tr5Tj4B+we/YNd6FXaeAZzHGOU9Czw/Cfbp6Ti4Q2W
lSGTv4h0VBLkNhH0Qk7FiKpPg6Lm+jhfrdjkzp3+ZK+Fl6SawUIgtKKJOaFX+P42
JEKv6Zmy2Vm4/YLMel2WRB2wwa/6awhWZ3RTaSKeYU+ZGnIIRj1pcoMudEOorqf5
PXZShTXkAJkd4ts/aZIIGThPwkDgtZFBK2wQO5br7DOwJ063MF2ZXz5fMolpBEr5
DplZpY/XK39wtibsW6lkSCHR5QBKeYZxNDXYr3zTyvDA867kN1TsMmCxQqoZnPT3
ZBmUvwDVFnfmenEJwCTMRXh5bw0OFS0hOiYU0aDqStior/Eupu4DLrXTgPZldD+c
DdOMUrmEu+tqGB7vhfJQFMyz1RYi+wXbn3OCtERS1mKGpLzV47pRh9tLr2lvhVde
GV+FDL+tnSBe5bK6/IeSI4H4C40vQ0jzrJ2LdDqbr11RzIEvmpwzRH1xNe2VFYNE
jQ/slxRTr9x2Mfl0dbn124r55Dzs/mfiG/AEaFFS91S5wWt23dqtjhZKDiwU7Po0
alHZYrHO+FPbX14StV+ovc8klz55DmXmcCtSztDI6FW9tl81e6FWDK3kbFv51nwG
L6hVPq6E1ERT1kCPHbXI/9pzIEPywtgroYoCCl2XAy7rFO3QzdZlsC1kvnm7/MMf
4HqPvTckKSCz79tCXalbUP1b9cG4uUe/UEyZciBGnaPuLFLx90CuxXv2aG2j+xt1
Mc3Nak2VJdqMfil8n5wfTljhfXqIdbtI8nT0r4C9KNpPnLYgSPuGhdYgTrDq4aYm
VIUo4m89NKNucY/s9p6N0pCfO401uEWOyKQTWgE6yOBF96l8/aFQL6yGvpsZb0FS
rNl8/waENXIAbguFD29afuLZD6MdJqGruLUyff2N7jVxqdWPXXV6C4sIv1796FWB
cpHrUkhzPP852gUO4bS1GnVmRa+O84wjSsc6xfOBf9WHQJYjyEAAg8oIXPPTgKqn
fzbCbA5KvreyIi10FG21VCQUacrJx8EFnCfMeMh9Ljm9O72WC2SfjMmiaOJkoWKe
mnjrxDKSXOflyDDSTGfukKApyRgB5M5N3hubI3wfd5hYzAyu//r7n7X1B0EG/Ljt
zfQWEPcEV3kaY0VbK8joN2hp7n8/2cV86RY0LFYVjhqYa42LZzkUL6OYeyAhfu07
YpZ6YKNLOrvptJCMaxZTA3p3UiWK+kXqDWC4BBZbG4STgChkDVYUXTt0j4EwB+pQ
nWH8ATu1Rc93ByUTMFVpKURBdWyJHR1lO7kUb5MN+pvk7kk3dhtgu7gGcbvvw4Pi
MwetL1bTTBogC1KcGW4f3n4AplHbxAYHbIKOdLdc2OllqLXO7x9pEErlpX5K15We
AZuW/XE5t3NVtuIk99NuR7yJp42S/izh47OeNC7GRqJxb+JFco1uGkpHx7653Hqi
IsHnT0OnB+PwZAEbdwyhBTB38F8PDm6bZRI4Nzn2fpgTyczhQsToP97uX+dVtUQe
Sc5/qSwhpQ9IjR9novtXsbyYdmktBNQPBKJxZ/cEYyfygm/sGs/jVT6FIr7uyjen
v/zxiAPbpXBGxzXvSB9+9IJP6YsbH2ZM4rVYKyNH8A276Hv1fKQTlOVn1t+AbwyS
8gKFGQMaobq1waFrwI0COGPQVxg7mZ/3QZ0FfWrmG+KrTY92ARQ+/is0o9k78lvw
Zz4d1RMBxLSTw8s0rUQzWqOAx4SPv3VJyBVG89ips4/EXStvK6Mm/whj6PW9GbmF
TSHjSnJ/wWI/HQudtAZtAO2lrnHbcneWkDKx+HV9COEitYkhPLCtRljrWcjX7FCc
Xap7WFbV00emBJ7Ktc+ILzUCQARrDTgBZfx7tMlJylL+Od1XxkbKdcTqf5LmJZgm
eGSv8yB17vhrsBTy+maEEUyEGQRytckzatHCzXovzu048I7KOAXVTYpM3YT2MRCz
LUwZj5AWv1s10VqxzmZtYJ7jk8nuicX9suyh5ulQ1jxOJGU3pzYIlrfwseAufxju
P3Efvqp1QIpKIRyhRa+P1rFX7yzPPEvi7mOUE0itf+LhGsAAAauQu7Q7qwqoHcnH
r3SvCKlZ8A1CioSOqcN9zAnHXigSyP9qkPWEnK/ygTtULw42ALngSxbCVkPxxDG3
l9stVisSFXW9gr2sJNfnt3cdYcRJLF4vG+sedj+ChHgYwNe0QyR95iWmf9dQ2WnA
Nrt7WDq98zjRLyC0tcjpAEb3yhV7quzj0Y75T6jNu3pSmAo+uOw5f2uNXUDYOGZZ
gQOF9gqpu8zaDQGTESKdKGowpkfg72rVyKUSlIl1V29iL5j6bKaYnPfr2FIBL9on
ypVsoW2UN2wkTmQcvLjMqzSiX3qoI80nvXrpzE44d/PYeffe5SWZNXc7XgU1OpRS
TJSNIoOEHNB6ZIkVDejPsHR6YcffDL4nCrJzquPL3OYdMYo2Mfdm86r/GBKB/f+2
l/EQzbhWdWiGAkEL3RcO7EAuhcY+4y8JrKoWkrXP60cEFKatPGNOMuA4TUZMFTg8
bUUYOmScCm+fAnD8pprZfPvGJv5KuDz77PU6m9HQV31cuB9LFn1H5TDwO/+aihXU
Xy62J7KtU5ZRbOvn/JOn8zocVX4tnWM+INFYIp1eqQXx4e6Nl85lcHVcK5vclTjT
vsC+m507/mPoWhZdr0CXwlpgtLAzrERSYX1bT9U/HWEoNx/rRLzL88Q74bZzyDlJ
11hcJ73yRsdml5u5yQxTNeiaYzJnz1wV54vzmJd4rL24q9emRxS1U+UtI2ktcDFk
a3Jx9NlUx68LjylgdAeOXXRUT/cy+DwrAtTsrh+m6OSWbDHQvK6n6wiuAZxssNcD
06AJlgT7bNb6iNybfqXV+OaL97zg2C5szfO5oyBgBBj+KlOtIgpCVaYvcUIdJan7
8twKyVBxzEU5gbHpYKfUg1vQCeILIBBgnV6jQrK7VoAos7UGYFf8lZtnm0hidYcV
6uR0zjSMgwzIpkSxjAIgkhjSYcDA8TNQvw8FMpO1mvVPCsd3MRRf+FExV9qhVL5a
BGe9rKVXiWHp0MZ9aW9c26+Q5YyxNC5dUVo7OIG21dq9TcrWk9tclLG9xi1JzIFu
HJCi13Qmq+m9fsXauWc7Er2AvYwTwIJKvXLCHdl5epyBxgCN8+dK/4E6S6cSMHfB
jKo3TRVBHVhghOGMH3yMKJhubQYSvSNUvftHSFpYYooNLAkqvQat0Csp/dzbhRSs
bvibKlIoT+dG9FPlbFfVdWQqc97G2BpxWqfkKe/djeT8sBDBNdPeppE+G2qplJ4v
F0W2Cem9BLxa0oLH1OnOM7BFQs4JfqXEifxyJU40SuAecD3MdBv3/NXvWEYhGKIB
VDE0GTXVsroLK1nNHP+mRSaWl69HI5oq0M59t+4HoDzl8bg/6ZTk+AMopXg3iOMg
XI/OhBMFLeHEXRVXEuqya6HmiDcjXvVy9jvJKvnwqI8TK88Sb8LhWTcqgauF3VDp
NBkUJw/rEx7Uz+CNe1suy4oXMmER3qZcylWJjaE3SxFkQVE0sd9NtwLT4iTKoRcH
6E80XfnkXvNntmzt8YzppuIf+eEGlrWasalHbsHUgbOZ92OZWdRZX1tWcSBwTBNr
Vt0AtgnhMPfQLdBdAQAucbZAkq9gcX5xE1w1J3auWUimk1oghRwsb8jDQjXYO4aD
xM3ep6DLHCa6W7kYaPC5dxz/CKt7E/F15JNdQk90XRBi/Jc7+FPeC/5dVVYC2+gY
EMsSKKuJpq1x2hTSUhn5+eAGYoOpECkQEPdWKDgvg0wHrwhcPmVdKhrO6M+10M2w
6Io/7jdxKh2T7GQJ5/gOB319D5G/pwf2jA5YItyu8AvyhorAbBXCS8Vl8Bb1fQah
4QOqLBgaOQN6PTayDr98WM+iJHwS+BpdaynjG3ZwSO5YJuBL7cRVALISVvNM1TlT
wRAz7MWDjdjm5T1wXopTuEgAlfEoO7j0pLEaDoKVIOrUpRZA0d7knS8JP4q99YNh
hnZKToUZnaP8WwJEYtSMHJqIA03Ae9VR0wuT3yWLk4ubOPjAyGyvG5H+QtVk26aV
FU64iqLnjMHnYP4KP+DIokbGd7QGY59J650JeTqRpdWHvLDmbHwm57nWNDKYWboI
9Kz8g5qf47PdDY1hjaniPfeBuEgs5g6USrsOlrnpX6XMZ+2zY/CZQD8UDMsVfpXA
skgAckigojjddkDf+ERV8AzycwtqpUV4pJtWn3vLj+KXuLmbAQ12c1cJ/Iml9VfF
tIWFreGtWvOEPnyMinVQJML4tUlmxhWmnuXQZFhUXk7HXTrDR3YOVvMVPSKhpw0K
TgGypfyP6gtklB+2BGIoDE1A1dJzoQOlsZ/vB1I+OAOlXYRYbjObXTJOc9uTfMJa
VSYfCHx6tcBTp9qgO+gIoyDyVne89V6l3Cvcce8tiOWt9b49ePQ3XJEaB34kfa2J
E8lgETfA3+S1uNuJhgfPaJQgdo7NBlGtBdUVO9O4yC1J+iUClxTODqbJ19bH/qOL
47KK4NVYZpv4c82De2Nk/1YOBGI8CDXhG76lC1CsPqACXsbDPFR+TrC44OPX2YqK
aJ+c5n9o964RZbnCPROnLpzLo+jW2jaiJznVcb9qZ6i4awSZXPOFIqvs6nrwRUDa
/BHTqY73w3Tzaod9dIwM6S974+H05cIDgoR77lyDkTveUQmGWPmu2oK6TwMwQ6F7
T+paZRuiUW0sOFL4aP8HITignWzQtCvo3+uIlwo1/gb2fL++shDlDK9Lki9CVjQV
VD4JzPg9AedGlod/bEx+dO36JuwBowfCgfVo98m+fn+ur49LSIFyd7sRbl9qSp0Q
ZcV4i5x0tsapHIQBVily2/XlsAxQ9FN+0DobtCIRRRGbv4VI9kSKoHGLhPpAR3Jp
RypWStj6K208VlSu8QPHKcIHBrfdgMAS5KeC7pCnDpjFyaEatV4ZjvNy+Mgi2ate
5KwPXVoUC3vACkm6TpmLB8Cq+MAkU5taBkvlxbFgL0qHZ2FulC9KUCvZUQpL/MiO
3j48Ep7Gy9so7mFhBS7JOHRnrdsc7cDhuqLffYF3k4KY8e4+pOYmAWRnpfqKycoT
rK4c20/Ia0Ws1Z/pLG5Z1SLqzUrQrRq3msEBNa0Qv+PjXWeWb19A9E16Vwyd8H8m
VVrVKoN0M49By48/jhxSs8WW9wzuksYj7QzhgRHBW60jiRk1AE7WGQDwGesV+ap/
OEeNY8S44j3JjsNu21jF/uKZgY+Qbkl3kXmY0nG/m5KrPnVwcf2/QmzS/5WploKJ
k7/r3orARviAHH08xovvRscc4fHG6w4Agg2sNajIEz3SuCYwKdka/M8ncCwVAMti
+rvHOf1pRGma5hLjFEATXqxyZpBtKWQQu4e+JAIekUMgAjH9zPKebiHKr6DLIsJn
B5QmwqUvjxHrgAL/RojHdhNrIMv6SF54ylqMeJNrm1qs3V4yy1ojZ9yoElVtbB4Z
c2jKkFI1bCjD1MTlujPsSgEzTLbJ3yt1VGKJw3M2xq04qqrWQ4jfFbFu8knDKNNc
M57XHPCnZ8B9/KnbBtQElRxrQ008M3Y0djED4P/7GNaZOeF8e0pip2QmiVCiwmZE
q/BOQ1fbiSaVATO0NgqfKFcH90pQvCApFYyzNgOdTSMb3tn6JpQSTJSIiR5dQTye
ybMtiEj00EkRMzI8iRKPUHHa3rwvkeOYNkSjBKAxQrih7QR2RaQ3G705lqraHtFw
cLk8DROZkrYHb+chfLegf9Thc+3Z9tq+o7OneAgmaKEYSIOJMVfxPSyqq3ayTdtY
ruh59Yys/1aHjgli+yMsPsq7zfYNwCpCHQPbgivetgSjJqJ5WENateax+YwOqqdR
WMhs1+pKLG4P2hORrkAxcMFZs/EcqIGCmIXVL28fiZx+A7SNOJrtUkXAqayxaIa3
GgPPVrfADC+2VNmaAXGpNkFRh28CbYC1KFCRQXQYL14pEPAKYUSlSijrZ3Cc0+Fo
wONUyH5p/+2RY/SQoq7AmCUeEUnALZBtFfggE/CwNUcOG39DSyvxGijgIfQnsvbT
ebYnkNvXKTkDOY744qKaqwQF3hzm/UdpRs6BMKCVbFlwCmyJNGEKZ3eNyvgAdaRA
dL62SPdJLO2L7+0LBgU5auCWpdunt09CWgoNT6Srap42pLQ8T3NnhwfkGx0ErFMZ
1MeLbuEyp6N5Y7IRrKE1s5qpxgzpd5L8gtvTK0G/a7GNRb0tNqLQAEUDI4V/qqHQ
9ae4+yyvMdLI+ZUcp4HAnPTmfASswjINhtT02u7rgUf7gAmusd4acIvXXd0ycuR2
Vq5LwYTK3f1Z9x6N/qjBiejEIv9B0T88FSJn2c9SGwTBTSGnt3Q4cLAJ+TBF4Zh+
aeLfDtnfJ6PRVSMpP953u8iVgTXtnq/Q7zZxuZLrMBU7EIOoSxAYalxtdiyiMOPV
75yumyMSPz2IxwSHyPF7xTNRy05gpCGQ6sDhBtRzfOzfIsXnJbTSzBQz5aon5c+n
NKeiYpE68JiqsPGT1SjtDm2fpGJ+aVh4xeRxu5Tsl00YE69TndQaON+2N42BGXhK
tSrLXg0tUyzOa8/JUgZ7oWE8J1c1I1A53s3kpPawB3BfykCWhkktLayss92cAXYN
h66xfjinNHS6I7lfgN4rK4akROuJJWh4bJkElBWoquf21d7Iv5Qwon9iLnIsBIcn
dqwEAQl+qsx7VdgCqDJKB7LRAHPDjiOnOr3czAOBuluuaoyw/GTnu+jD5yMzrntE
5rfUzJEh78p9QZhQE+7y7cMGVPeBm3ogSshCiRrpr3hB4BJx1AXHdHqER6OVtAjb
DFA7AbWSdYY5kGMUm1x1QYYitJHf2X6s7V9Y98Bpsy2RHqApnwZXRMW16Hs/1Qd2
IIYhz8o/0MGu/7/tWUTMiKgthP6uORGeBk9YVP7JOWJ+h/DoerKdc9BFwQE5+cyB
OLHc9p2AaALS5Q3LmmZNm2utND+PdcuFsHF9hSn3GvG2fC3FqYB1pKzGeX0mq9S4
7JhEoAefGForSpKXIHa6aG7aFr0Kq9R3U35Ai/+61CD8vzimjV1vEGFW3oK2j+qU
f9j/JEF0J1OUNqL8fljdVmGB1PVDmRSGxQt9fUZFLv5LqMsHob+o7e8+dgev/J8y
99AXfYlEEAKZ1sQKey1IOh0Pb/Y/aZYZwNOzE8h2hBV3KnpFsq7GVkmbuIilu4is
S6wZ9XGnz5m/+9jJU3Ab31RtrhsOQFvfHt4hU9hEfULgXBMeM8cU6Rs+ZuX9xqbc
LmvGKa1HPv61ZkpOkaEgtdJ0ghQh3BLBOZm0hdGBclt3URPZQUoXm1BBDj9TCY0f
6w4No/MDvqS+Lyiv+/6JDNVBO40WsYjlkvadSTxXQrd8kS/zf+CH6P4unYqa0rLU
4GrLBrUkvzpdE2xQXdbxwQ1AM9gxivLIwzdf0SrdwJaJsGB+vipH97LAR1TEA1kM
4k5pPu5+i2boBOazMSyoCzI/bHM9naznn0KyhPN0ja0GwJu1uTGOJMHmzVY8alui
6oQzkh1I6xNejyCybOkoHHhsiGeBdMqRxfz69HURLd2la5UZ8T04KURUAzajB4j3
sjtE89UsLtnfbH4mpoR3e1/ryoIBSyeIs4JTxkXaeEfOlTxF5ISi6XpPIjtdA6CE
KxRLeqMXuv1gCzgjRaNxoCyfvCHftH1sAIQRq9ooPe+zv4RigVCl8TXsLAMaC3d1
7nM0Cw3ilkC8xGADRVuq09Wwk8kLZFl/3KHQYCKYwvebXrq/T9BvtB8OKmtOIXKJ
4IEFYZaXVJN1xobA2S/sAJTf+DTcfiV8FN+uV6DpwSZcrO8e3IV7xAOO0NJkoz7n
ir5y1m0o3BpwAYZS+DYt3+sbvK55btnsJU5Uc8+N1xZZ1UOZH4DTj9KjZ3nU54Fx
soD/cDu3f98eVn0NBDuTZ6pbURmYI4iIlFTQpj43KTL73LFfUvbx1CIaIwDtqcX+
SXRJsSxhIyLBR2WTSQwbglYkMj0XL4sc1soR3ajEHtD5VAGuUSznj1YZeARrSyZ5
VlENpNFTuSvHbK7wLmQzQqjgZBC1+E/uJ+dCIzo/Qm9GZecBzxEBYXksAd0k0Peg
bIkh/oe5WdiLwbyi0WsWRevV2Xnj5zw+Ny3mOIElHKowyYlwknbizB3BlDN1ciD3
UkpNfg5aoyeJZNV/i+584Tpxs4A7invJCnRhw3xDw1pePHiAQRMey/77Lfdyc0/U
jnLVCNzIpK2IcBsPsgsehYz+uLc+LvqE1odCkIB+LUMJehN0YzeKWLoxPHbrYDzW
EX9LCCVCEYd4aqHiHfvr4Uxk+P5U/zR4GXmpORnp/YVLvYEoR+0kaPzLUNzWOSWr
9s1EzRG++UK+Cgw/p8JUcjuqDkDrx2eu5oI04FUhRcR6jMfc75kaOQ8IkdxeMVmT
bE+trPgV9u0+eHCEbx+QRiESOk/+tWY7Lwpy4TYMlYBN+NIJrX6n5BlaVMZCU59T
D6JTQGbPVjKCDwgorlWNlS1vaPh/U2PQWEeZrky4BF6JASdLq13Uzxk8b0d6Zmr7
Jw9qQA9H8VgiLYt4zdhe5EWpDh/SN71eaq1IGjgE+j5/1aV/MHr4sv/ErMgVaS0U
1RG36+GHzWhKDsCw73a7ZLh7NO5dLpC81P2oahjityTdIn4biVXaEK2q/JOklwsF
ziCGzap3INxUW06vTZAEaPmAlxETdhSU6Xpxv/TevjFaFODaBNko01Ay9eeMsDDe
KUHl6aX0qtB5Q7spc63cOwI7FLZea2RCvuuwXAdiJfQDVkLRqjW9MAn9YmxuLt/b
BzfXWqZar2U/sTFbGI7pvX6lBXpvJRRx5Mn3TQIEQvw6K0jHVKQ5TIe1Xr/ed3s/
T+OwHfHSS+Ybmbp3m+GxtG98nhdagzudnrk6ojLV4g/j4b6BcEGAWkc0xW9IP/+s
18lAFRx4RxnMX/sM5QqmYJxxrAfrY8muHNZHfzyOV5GOcXwK1fITS6jHMmLG3lv1
qrS4yf5Er4P6QJx9IbW31P+HQZC735guSE0YSvcfyXFPcKRVF65JS9dUSjX0kpe6
mSKfXvFRPZYsCnhf92KHPqMkimJcWe/0MSCw2rGZmKKGMkdxXXSipN9fy87/JuFO
BneW5mLjjjLRPvOpcOtSo1j/uwxFPR7TjeBQYbaM2KFHuPC6DqEFBbxz431JnXLz
/z27tpHUgc9vmv3PV05GDGOzLRFE/pBvt6qAgObmMnVaoMqS5ZC/iwMKMhTXEBO+
37W70a1twtLMpy5YSmoK1K1OTCVENITBxZz6iGim0hp+sKnZnjZiRDHS+eFx2NJd
7LIJgxhqKKxo6zSZelQx2oUtzuhFvHHqHGYtFxjCRWSSLjbBVdjZiC+BGokpiFEb
mz/YQeU9dNxxH5H/bBlJJtv3X7/XFAcu0Zh+aNIRN7+HJ9OoML4A4zSnisLYEK8b
3b5wp5Y4CQ3XeEW3Is7n1JJPsC1oDAPJ7g4c6vEogONpuUChAIBtNVyGqnTmxbF1
uoVaY/uthnoW7y8SLmPsRDAOnKQ5lDiWToqJZ5cEdOcKAdKSnU+sz0i+iXKHxFC0
bH/3+zF5pchD1x+WV8cimL4LZmatylOLALU/o2gN8ZY2rn4ADwxX94O8ISLFyyT0
/gwoDh0XYmmZ3ES4BmCvezUK4z82+sMFn8RvVVRrXPG0G6fLbVW4HvRaQXzy8W+u
2kCwh0j6LcPg1Glc52o4Gl7VdQ40LFsCN+08baUwxZ6Hg6warO6GFeo7yeqqsuKQ
mQx6Ib1+R6VMxOI+zEpRQOX5RWcYahW1Uo0m/LVhPne0mRsNKPpdEZkrQpEf31Ao
hYjXqJGgE7K6B6OpCOx/t61XREzvUhVqcYlL/eXG5F/egI+LYvxRywBrlCwr6haR
pL7K1akaL/WvCqMRSSEzEe3lp9uXPG81TkaObNGpVD1mP63whhcSiWETscwa2ucw
R/dprtrC+XQwjOHoeV6p4k/BIB4P4zo0WqhdR61z9Dw3JtuMcQcFm9rEZcfDBOUd
zMRZo3HJCGHSMjU501tAbNxLdEZ707oSislbG7b++GmsspfcUwNr/N9CXS9n1e7j
dVvcb+GoFiypRONBbUBobJCHhtQtAo8jcStXxNsxigHHYYahp+UX+rFfFHYVuHP+
0711hZM65SCgL6mJkiFK2oSwaHTK8zTbdb8RjS9Tj7HRQF31vrv5Jyh+wmO3fdSF
6YkodPxXAI9xt9OzaKWjk8GpOh6edWwZNhpEi2UYteBcdW15I+DJ9Ol1WcdhGTmI
kNbh31tLZwN/GKH8Xx4nq3DyZ08FBA1M3DkaXuQ0unWoxqHp4pGmwtjb8Wa3VT8Z
1FOjVloP+N3H5jRNsXMdbM2mOhR5ZfmqZTkpUySl4qeqycMrf240+BXnFD7OXyW/
6ItBKBuNSIBGWr6dFyDBlQdRhwWJA7K2XXq8IjaOZjSGKDp3mUPV2Ylae9e8E55e
eW1HyCUAtC+LVwKAi78UPqpGDVSw2/ESCMQcFXDrX7IPMVYAxbFuPw4HcGuZTP14
OvGpqD1O7xLpIZE0FRJrZoDNzP4hTG3LKWRegWMIeRMdE8tu9Dnk7lTKu4W83hio
Dstfp7PtKZ0PrLauOdkc9TQkR8cRo/g2EPeiEyJ4cLzNAEf0UlzIoLvwikyAuok9
yB8HH9TWjDyem9rr3ua2X/Y93T3l9adX9hlumfypLgRSch0zUpcULsKpfWxl5Wqy
tpi/hIUECorhqfCCRBbqsUiSLh9O5uD09xQ0S2qziuX6uqhPD36GNml6+ivot14q
9D1BMUiqMIvU0+mqxC4w5YAATEmA2od/7Mlt+gOwcQ0OJJPMeMmoqXXiLerT+5gy
QJ1n+N2t+KMiiO6xFvG9O2ArfipShdQv/lAXra35ZM3S1nfdmonvUFBlrlRSzNjR
sPEWBWPUjCMMawOcQvEGm/yxVl4WS4q4BPPzJa2N2su7kfFgMsfjJbYFAqesBpdu
OxsGnEIhse2MEk0vTgtW+RzGCGwEA518XldgixlvmCliE7iebsjqAb8ltiZuICgn
hxICIQHFMRXN2Cu3VwLhISz/IQsY1Dlq95VNWaqqWllMwW2vlxluC/SRyXKm48VH
DUy+D6enZ+ijtewA58VAfXlWl5xwOrN40GX8WYzeSUh00ZUn0eoYe4Z6r1C8tIEN
QolY9KseOkFqm3emYsvpNliBsWZivf57iFbomJxjXlqRJ0gQ0B++mjie4ZAlT0cp
6azHHuTDwmadzp2h/Z8NUYAzznQES3ghLa+zXfpNtLUiouGE0GorPtouvVDWQ8q2
0So+ZtUmAv3OG5OLogwOuaaSG/vhvx1g35LQJN0EyzStdMaQLkHQVuGwteemCtRj
v4IwR1C6fvN8gDs8peQ6/nnqnlDq1Gy9xEcZhSaWouizqXfT47SUyC/iRGcrJWmX
9GOFSsvyaYzoTPVrb4lslxyBYB+eUxX63Cgmgs5VX5v9AgLoWk2/RW5S3fd4WFZC
PEBDMq4wenlSv9ocCzR+q6MGxUdNjQm2BdgXFvk63PHfYQoF/H151Wxfl8gUvGJR
wnAuy3t3VHAyRQt12emb7j5pnlw7nwiIN0xEXLaOCdKlBytVydt2b/Gz/xw8LcGO
ypjnv2RKR06ENaE/CzHxVCGbQiSq/0CxXrQ/lZFYqnHqyIIa7KO25LYahMpCGWlD
fo7Qt/xw3UmTB6EQcDrNJXBnoFVwmA6yLQSc2A5PJ1g4k74C+iHruxXRW7ZCcQ9R
x3A9hx+NGBzavn7uSHDo/yAElNzvWWa7yea7ayqHsP7DTHtXrlxBZjxvbonxlSG0
txNq4kkTffqXhEeBXEqr2xYVpMe+jMvLOwgvOMOL7g0a+svWRua0E3nqiqAadqn6
6ljc+aXSL+9OCtzQkd2staxy4d8/WMaPsvva9ABhLgY+0PrgG3HOJBYH2CeA43yy
UghifGgR4klBE0w5ukEW0kLXzlebqlHQkUwPvXocO3aVAq8cxKQfPNohO2qb6wyN
+fGltgH0BUvxxrB2Oj0QwmXo2inK9nvhVKiH1aSbvONghg4crPyFz+QvMfAEFj7a
VITLPI3VAobra3nxvVM7G0MZQxRqPV4BjktyxaefSpZVehXzTN+i7DFUcajWEd0j
YUaAnhzT2Z6Wy9XNx5BUv6cev0u2lm8qknUOGgj3qqPbuDF6W24IULBYzjS+lIOn
wZoPmjvOuKkDFE7iZhEmJ0TwpwULa6c0wjy8tuHogyAgaIpkDgW0k4dFeWMoD6dS
TjdGlp0fuIPI9waOf3uicW3nd7u9j1fp6uzbtFHSol6m1leruen3M2RrkOOxcn8E
GnEbT3ikt+R3xWJoAbnxNI4E43UxaAqonIbd/xENmykFLSvhReLCC4kgvi70Zikw
1Hk7oszQyctdIvRFzegg4A2VRQFBfmCSu00gfBN/VEV2csQZlJB++jTetdUXg5Na
i9S8EonaFDkmadfCslEvqlxJzGNMuTRsvsluQgV32llMTNaMp8jiJCAxUxx4fsSt
PafgIHpfrhQvcnXRtn8a0Kdw5vr56Dw7yFe0p6WtlAgbLq9AL2KHGreCXz6qgvI+
12zxTFb/N+iG4wtmXrjAv/WRx6vipc+ZoLxiqiVjxhoaA8DvD2ZfmjVj8MqnKO/A
N2enWqynMal20IyQ3GB/xgxfaFuNBpmej1YJR2vkFK68lHnBB4bpV1BZ16hh7zPf
sPdEPaWoUOKBKY7xoueb24mVF6q3RynaikaSkQfFCW/yyUHCXDuOrPZTvPmvExhm
kvAdglQxm5pMNJ0VVEDdo9oY0mnpIXSO6NuaRVvC+zKq6Pa12sedsiTmKh9uquHp
BzdLkoM1LBYkCYJ9FmTAJ4ge2IbQwgNbNJY79+DPoiiG++NCBVM0cQvQpos6m02S
c8htZO0V6jC2kTap7nLDc4hSc2I7KWtBNanhLCky7S0nqnWl6dV4wemJq+OmyoEW
bG9fw4Cq6WUCXoRwuE7eZIP+LZfmQc+v+U13MdHgBWUvHaXMXvVslY8euI8UqaN6
ENoioJ38nPwlyqYBitPNacHsrwn9E7bgk5ZUR43N2xXQ9zjeIbZOzp0WHJMV1USC
w5jyblS4B8GlgZVco9mb7kOX68vDhKKsQd5oPhDKXoBcUeRVGfUvp/dnQgV0X88N
KjiGE+dPcAVxCXws/wpn8Ov1WUGFKglW9T354QWFmwlwy0a9vz+1tk6nZE3/TZ76
YzNzlB4uCLu0QGUdaSQFAUYfjBfF1VMciOwj+LGwW2jgZ0GQ+/EKXxNMOm7iG0Ts
BP9xmC9Jl/Uv+7DEDpW9FjJ/1A+O4sk7yVKxLuhD2jCYglTaKPETjoWqBj+Ldb/N
8rfAg61jOKi/F/xJepNAnbpRkrZMLP/JEZsycsnt3qEhONm0rJJ1CW1YQiS8hkqb
Cb4+ZRCzKATZOlkMXTG1frMjUrKfOCBkXl1M2w79+b2jDeATJ9E0EtdZF2bYhBHh
ssoAPMWTbQ3halNMp/CXVWrEE46xmvGJbZjQARIhNk4Fd13Sh3mbB9G/QU4vYffl
PMtACgVH0+LlFFpGqv3pOT0aYJz1X08UJ2Sc03oluXYHgLgVaMo1+2Bl4emT0tpL
8mHIw0NAdzK3UFIxurSylfp4L/bN5Lpj9yhVr8yyONTosjpMJYMZdFjNfxVglSly
vWoMmt/ckrZr0rNUx82cphLGnH4wjiG0XJQfymhqfkn0oB1QN5VwirVi/WAKuKRP
pKIiCmASV4yPRMaeOG+mL1CkcBq5MrM782Z+xsy00T7q03kRMl5a2kJek5xugwrb
o5Z63FQUTqTmP2gjVaoIDKG/lnPAfbBy5TBJrH/md8jDLQv0mE9NCXD5rfz9POaM
BhflmVCiJEwh4a5OHXtgrlm8PJQolqrKVNE2als3KRiUW4xwVX5QmeBNlr+mwwaT
5S6Mdwo4vw4kkYpGDtRfZUDxGAbeulK+EUwnW73GpQuxmEh+tW3BfNNd1TFMF0yj
fDE2KFxWNUpTD3GeDK3EVxprPUz0LYHOE9/f4FVMbCHNqVOJPHoRoXKRQGTpP+ON
1IOJAOqGe7bKnP1473Y1J4T5Nb46+CijVnkEC35l6OaDz+piFrPHs9ssPdGl/9VW
KDQNPKWxd+ZyaR8ipNzKaHQRUHfkBqguZ9R/jguS8DxPTSOIeMmBY1h5tvRoYTbu
SoISYIAIA4fVVNNX/jWCQ5H45lPcepZTBs37xFSaq4Gtrh5wG6ED9sPmWI9Kx/z7
1JfJU8BtRRfXu7puAaOR/vBADPdyaPUtrqa+WZvC3RFrOQgYgssRLQOavzLZyV+B
oOeiSYG4JIJyDilwShYplnzaHnhC8SnaLD6Ub8njCEVyuz3PxVSxQp7SwE940IY0
HlPozwh/paI4qtveJ2MQEMtdSsIaYLGPU1RmY19vKpCsjNzoGkH+V8VXmhELD5As
bPDcI+Lws7LwcQse3WUtn95n7ZJVsw02mexZwZK/l+pXYKGSbbk7T9V4FlO0wF7i
BJh9sqqHyMfMVKXPrOkySpjK8oaAED+hlMtOP6G0/wyZRZ64AT2h67GRFhkl4Tkq
6bLeunSNRmsOSngW0vp8V2pKYuZiXZJwA1N4vOf63k36aVvV0EffsF6ysUd0XcKa
MCTxCO14nX1Yvq0DTobNQ0CZJlDP/E0Gslep4X+gcS/x2o7P6swcLmQIbWO8+ym7
7TWXwCL7q7JfkDKoxL7BAhk251xYOv8/86p3wUsBapVU+w/s6Uk9hkfXRviFRlmS
zTcyZV3HkGT5MWEocSljVqgyBtUc1unX2QxSeZPgkBBiRs1xZpWsRkzPhHdr2pnr
SWXYuiumgelsRzvI83ZWaAkqqTYWzgPl4owXJDCgi/p0p/XEegq4aXH8N0kv3liD
5lCUubCxA2ieo/lO8fw/Y2vAa4t+RQcBYFoFmDDv/8UPQkXHeBU8wRgc7kfkNUA1
EU96u0R3YwtYccQ7LXdVCgEJi44neaNqVrY8P4Fuc34ZhOFFLf1L0ZoBE4rko5d+
hPcCDgopPEpe0HtKnDNdz2PzSaDQzYmCXY996Q1oFYWohjeOLtOU4iSXWOlEkcb7
vi4Ma1ywOdlEsCefc2PcxvkB9cSItJneZI9KClyOM0HRhvRJaoxGnaXCN5/gr5sc
KLJsuQmgOiiRb8rmDiZhuXcTXQk8KC4pFMfUgfShuxRkSZZBLecjmPd4ORgBOiVj
5K06a/a7zhLYHfqyIFlFSkJ1qR4Z5zTm6Jciv4xMDCa/peKx+28trsadoSwIwDI/
/14JgMNHZKCgtT0mb11lDtkTVw6uGi14NT2rY5B/BFkPtaYPu8VD1ZRHD6EQQ9ed
g76pqOnrMAdxH9EYK4B53JjOykg3GQ4mebSjgIP7HC75jztOgajDV9WeMarvVOtd
swh5LO0IpQ4JIPCCy4PfrV8Hk6oKsgmH3YjCJLkzB5IEiQnk3IfB2gAH5kh3iChK
RL9VqBkFcHP058W852sV4sANpVjDZ4V4PeNsfs7qZHBRGt2J6Aq9MrubEhwl3/lW
8ybFydqGPG4VvnimUoWCcQKVr0sGCV2R2F1AzMi97jUIPtz1JIXmI0ETbTjIdPA0
psWC2/8ewzknstPX8bhHyLEfSeL5ziI0et1LfhTHqn7WLKc5E0+5mDqeoEkTHiKZ
GMB0GhlB8m5cLs3x7zyvcvjFNPbo0d3UmXTYuF7C+iw2F+DZ80elPNPHhdU54d7Q
LXI0p/tvNwK0T32hpIDIulvFtfjc2Gs3+gsl9iNUjbSFDfUcsOY1c9A+J0Tsdiue
8/d6G+cAGkmkVDUT232XCrAAZDbaJiDrTe1VieIW1YfUAOtNE84VzpLHorUmACCf
fa4TEK8RqC2f8GVNu08MV+XQ1wFzmlZRBute5vtEVbRNCeWm1TEU6r+JcA4XYV6c
bkke5eOjdF0rRDI1Sw3J4EgCckgjoNV3fMb+Tsf3aRQIc2ziHdO28/joTjr4/54+
NTSlMB6/RYPAWKhNNenPV7f8XD3QjP3y1haYE+a2dMLrzJtrtL3Bg/UD6p7KMP4s
0a9WTazhCe9C980lGXf/ZPE8F+YUUPKRr3lNPbsU7odin7qmWwl8LoavNpNcJzas
XM2G8bMg8jlfklhRQpHfG0zff0Yw3axnHEWrogbKOoy3k/Qiw/DspbfRr2jLnhzW
1EixII9BV+2SgHDoz3a3KybXMOH/3gCE60zpo6m8MLGsZcb7J7lPSiVRABJMxmHT
SxuMSUOTIGAEZmZ7lJDxRuIJSlx2EToepEyY/cLkqoKhNiFg0jqiWGdygP72mQjo
s1Thf4rvW5+uOqcaH8Ui9mwPnRRKf8HiXsziUv5+bV0+lWsAO2KHWjW01Q6d5t0l
V38z2isSET5qmsl0f8VQgcJcAjiwzZgTMBvazloXtFLP7dg29B/q9ACdI6cHxPsz
n/Vnh0WX40WikVTHhkyfhn+WaIYC+BY7F7SQDXV2zMUPWG8s7KozaNTf3pB1r1fE
0WAImiheiPXUFtJl8HYgQJmq0m/c4ljw8uen78xGThKzCANVAw91K3C2XAa91g4y
rVYmrrB40yswuOYjL7bmWY+/6XOxjvvvFva5qbH5n0YEhJ4gky5fd+7xotJtflYQ
ekhSbaktWcYPf9IUCygjEt4C2ObnRIRsE2GZLZNRi9kEUN1kJdcf0dawWggyXTZw
13GpUwTgxedLvkLk0LIXESiU57z+5nV1Acw7NCT2Qq/b61iDYzFxdGXGop18DVT4
BGabzJ6G6+qMdx13OrZ8ZNMoT/ytBnhZEd/C/QGQhZVRW75hHwZekpbBja+y2Utz
zswd0hTPcILMfKCq42Nii68kWg9iJS5sre+h0WadgpxgCmSGdeB1puNtvvoxmF36
9CZFXw1K5qlu1r/z2PCzS6SZPrKIxz2E7W0FIJMBwT3F5kdgSNDsPgJL2WwzHQQ7
f442/zBbQd/KQbEu9KrNZLjdB5fy8xWrRnOvCEqz1wN9B1iCU8Yn23hlGNqrCyyW
2e3QL50/3Qj0EMX42gJfwhfn/d7mrmKBXymknS9ZPfCAaX7ZUQz2O8leILnrOh88
IERXP08KZOmutpwU42aXOEfNHbmUNpsUdXCK4MD5ZccEb0uN4Wzmu4ltXcGlEzDL
r1C6FcfZehYF6tJjmlCbuys/3lj09vWvC/VkLEX9eQb0mNtt1u1RieLjr/pnqVve
ORC2HQeKa7ycbAGORMOxkCVNzUnFqPvczeEmjSON7jbF0QgDw+ND2y294kBmNi/m
uPmuVuQQEjamPUAfJAkYAAnx2BluCM1jTAReXu7Ay0NQt1L+Ecdmw4UERC/IXM0r
OvstXkVEkcc+BSro1nXlZwXGkZYINmdXpdhRKfO2l7DAg8z3hNOiz2lQ2ZUZu99C
kHf4LCrgmE/E2mSqXQU9qrSeq/AiYdMB88/z0VhraBcC5/Gb3pzZpSkMAlAZN7k4
eK4OXDaqNhL2fwoxgVP/1e3tY3i9+7I2BYmwMVDG9XetXvLA8oZPeH85Gzs7+ASD
K8GzOE2zOZOUDVPqPITV1RXm4+4ffBtB6wdjM5akvb2wj5Vv/kYcS6wHrq8VcBT4
Fx+cS96gfpZgliNDhfFnVkDk9xaUE2uUTt+r57MdFCuJ0NIDkucFolG5m/AhzR+u
tgZt6XWmtjdJxkMbXQ7bH8k/ztME2kF4HVSr8mglbGMNAUs05/++RpzZeEhXWBZf
CQhzuP3n0kzuEPulmPMO/MtzSsaU/wuBv39VvbSgDTeKoFa6bPxBu2avT8R62sqX
Xx00w//2Wrb+wywU3zGP/VB4E68yJdc4HCzfFa4SEH3mUNc9p2PqLP/tLXKBr/NT
bRQAtHWfcB+bnaTRqrSIDCR/64zJFIQUFegqznLAPSuEVhD1ufa470+nyBRfmSqq
GeROilulCx5tVk8MsR8i2Ie+h0MBSOvWy4boIK0vSBpwuNFC4QXu67hw61PMKUuC
IOxkkc2p5wCp2ge1YlABTJiRtv9i1lwhuVjvpZw+GlGjVuMbL0glZ5CiC5hJqniV
92Cp2fHRy24Znr5c+qu3WgaLjULAwvxxOO8snQheOytR4so85HF8BoWF5PL8f375
S3pjATpSWs3ZiZXDmXpu/FLV4EkcWxIDoaCZI+sPmA5k+sPnW0z+/otlVENhPZhl
pyqMwTDNIt3PknuhI9NfIdb3ptmMCCBWsYwlrZNXMTLFzHF6v7krpgigbF7t3HoB
RyeMIwsWPaOAfVD0dIcKFy10adxFD5CLSlpgYUxYGdwP0dp+UXQiyQld+AKD5yEN
lLmwP6pZAIIrj1wxAwu51hmd7ViuC1Rr+mZ1sACEmUty4fwwASBv9T7Iw3LTQZAZ
z00laCbXJHUT+s6q7x0CaOxeum2n3s7951GefcquUdlXZwzjaw2XbkNOyYWYB4HR
geclcAYb2Kv9VX8Bdc4He1+5Zejm3qazSGsIe4EUPxoA6H1IGf2L0/mZ7sD41eZP
iq6viHWOj7YLmAQKPXUCuP9KjWg9q2LQyV2HI0Z0FKZ077pzF9eE4cvsBxs39yJA
Ns19w4orkSR8Lw1Mqt2L6u6AxRuxh+UCWR0ZNck0i+yIvtHd1dSdaoumDs86pCAO
+kfNvxChIvTWqBg2rUGT7cAz/KrqjrTGzaR2ZfcxPUe7Vl8Rblohp6CMZZ4b0IJB
wi/4GZd60ZDpjh8Og0EnRladrn4CIPLyKZl1CloUW9V4sYP+UR51EwuRv/qMqzud
MHlJJG09MDBA3UdH8DEE/av18Hq7AzAihsNuRj9Q/ygg0yjHWI3uxiC7fMbnIpa8
PugzFQCWB1I/DA93rZIwdakuwJwjHrpj5Q/aVjOcPEm6DTOsr80ukTfURqCxi6mr
oRK3yWJnwcurOV0eutWPiVVme957jfP1YWc8dkvnTeLlhrlDAXJA+906xTMQjxoy
UEWjvu4qgw1t3nNI9t2M9Ak5hGVV+5axuZ65YKO/dSHuJeL+M1UU4QXOlyJ35DCh
olKD0h8YR0kwYlHe41gO7AslJkbS2GEvICaK0GUd0XvxxagVHwRxwI7mfnBWe9oa
jz5T7x9tBg53ALIoxHiH0FDTMAd1QY6Trwz8aXu5dpaIMbjMMDIxYafNgrpZx7Os
M2oLlS89tytOvPO2H2Th1wcyR9oru/Q+Q7ygVBE+TCqt5EXJVCSVcxOBG7n7l0qY
HJJN8iRspxbuNPI29CJTYoomn5BJ0CqEihtd2Ftxs7gxHrURJMVRcHMqt9rAfEcN
yrAvozNQRqebwmGyxaIAuN/+DDb1aP3WHd1JNfJp7zokigud7uZ7Ee4L14TxoV2P
Xa/Jeh/7OH0dCxXyG/eANEODIBA8p1yZUluqCiq48PCGfqQ1qE4+BBdYFuudFRkw
7SJXuDkin5FZputPWbKjbvNeXdPS3ODEjwbJZsqfb5UcgQ8LndYB8GN7t57sql0J
0WMIQjf1unDEGnRieIs1AeYBeePPwgXVROktq80hgBdyaIHVe7m0A0rJFd7sBTjg
OF4qw694mvz/iqospaAjBjJ2sPsbIfqlfzxbJSIA8HA6J/sQm1zreRXbIC9qxMmN
n79gPjhHHC1Qsw27WOejPxziePwGkD1bUAJR1FrGGXx6/Ys/EXpz9J8fXgMOY8oD
ofB8GHTMjrDa/fKgZpPODrSzl5NqIeoa+ePXRCxASIXahTUurXnCatvnLbxJ4VJZ
BMdTh5h0hNwnDCcO6/kwWoUmljWdWWB2DkHwzDMWkGEKTNxcZD2I6TniAg/I1emQ
aA256rT4hasf8Si1djtqjroOz8fdn/354jj5ZothCkbwr+Gc7ttpAXZUFHOpFZaB
oNAUXW8IDMm4Kap9YPzhy6Qgw63cBI6vjBbDx4AlBNvgH1+5vZ4tBx3edWzwnoKh
mLb4PQ4K/WEu97+QT77QfBJsccfCihcISk5qwscB63DE0q18NmBNI2lr0vNHVj1m
+9zLR6qSpdyKX10j/EakYU9LWiT/2vGNw/4grJ0FzmG+iFXt3Nbjtk0l+PjhpbId
LxTGo1yjMeD7t5u9i94jZY7619hdunptXvljBQjfPIvFBMpMsoBc1WAbEG7WHIBG
INz8I8TbQzW62T/yYZzgs8uTW6tYCVXz+ysPh7MFvd229I3CpmkMv1Z364uAsDXM
ETg+jNZq0AbmiHp4HKonmE73Kq6rMas9hVjPbVvn6MKaeq7QE0Ie8pAtiRUApBz1
sXx80++gAYeCV0uBmTMO/IiFEusBoeUz72nVK07//JUvSTucab2Ua0UZpbWiZQpI
b24g+Sv5+92i1ya/dPf5er2dglZA50dF8PcIZFk5RcgV/weadixDYgwab6J6Jap3
Hrig6BOcfislox/mEwfYX/3gFHnloFCjcub9G3/elWQWNbjpxWH56gVPcoQuwYta
z31IroEBb44JJEpneVOr0C4xCBcLJNDqsc6KkbMY+1daanoSWNzPlZO14wfcp/fn
7kflLT+1ZBHOEpiQhHe/ktgKsL2nt+cemXTkzFFnrHPBj+CuRZ1jJWd8rhWFECLY
CqI+F0DryORelAvL/v4sxZIks4jaMIaQ3ngDqHBTJq9PRsZxuSSbN1rnOjcrPFMH
N1K/j2xJ4J34gf0+ZqoNykZkK4GAfjzQtogxUeXtvjjzLfnhd4j/PrPvlLZjKy8u
2MnmscQzpvqZ9Lwo/9p4RE7vNAEBqFI2Rg5YlFJ7aG+ar89mekuTFex+ifVU4kSK
sJwFxamcvnCwmFAPWP7eovT4AO+PfhTkQ57Y4gfzD7TnNhgJbsrkLvEPt0c8sv7r
+3wzOeHhiHvoKxAR2BwrPWJ2nWcp3EqUSuwpftJsUYiI8hJ6wZXB2p6n8Q8SANES
OR7kfDBFVfVFxO5rJiZf2ytBI8TMRT8KPT70LGN4z0wKMlwTUBbP3+3qaPtKO/L6
yAwnEKXCMZqZV8R/9ynQRDjusC3kOCs6i/AULtRY2WU+eHqeLGDYOVLRy8GqDzjf
P9HLgSo+8bIZhU3B8euu1JR/yzWkXIV3V0TScPWx7z9PTbKSUgB6jc1hcCMtOIqE
OHS15PdIpfG376q6FdOmwKTfKsqHivwXXWod6KogqFv9xDFVMSu6izTlAsVwwVUb
Dw6LarJOel7kfUswdj4sOrBMrtoMrsNWGvooxwaLmgvVdMxUJjERJjHenhJ6/nnO
wtfA4zrDqXyJWOxrFBZRPTYuBprve8YuLirzjK005cIkFYGVA1FS++I7ZfFTqFTB
LU1KKq1DmYZWbuDxe55MR9eOyH4xy7Sbg/JSe8aaGD5zeLmqCGmV9PlkZw1wD7Q6
/WZ38K96k52D63z65hD+grJpCUhoW7RMAQtkKpbzrXNfx1NQpa7v1l43HqLBmMir
gilU9uxQAfJr7a5Cc3T6CaynemPRsLzRAmw8RacVXaFzPB7C1wu1+GaILyyexM4X
0uOw7akOd55W10FJOWxhP1wOMBFqxoMUEiCukzhOHP3lHkBmO4C5Gq5pGwk68yvz
9419zRhgAaOgGYGdoBstFn/Nc36BSzv7hQkgpbd/J1Ve/AmGEbW9PA6cbtPQZYjf
895CY34D0UstXMXnA8aAbGL6gB8lgluku2o3tWa5w5WoXEq581ej2/vjgK4xmf7i
/7/qJH+/iFb6t1LTZM3vv7iv5K2QL+vc2Vgv/+S2F84E3jU/xk/b23vQDhlMCh/l
Io3zzc0qYOKvZK3oSPoUjbfLAN1GbenKQ6D6Vs25akhLp4uEPwMywlyzYHUTKMEc
Pi9Zmegr9c2fM8tHlyG46iHw7YF65ENRqr4b1nkXenlhFv4fH6P8p7VVYoBNkPgQ
PbxyWkH+byB8zpFOIyAMcqJyDJ+f5yjVvTXDpD57WYk/vabHiPDU/9Sqt0x5SMnC
plxPvJI2GW3jnaxjOKmM9kT3Lnf3oIOypCwIENP8MJpiwLeL5cLFDSuptkQaTHqc
OpBJNs6bfoXGha4ozUzGdJGQQxR/4QXg7sVRu+CrRAhO8uPfP5qzOjsXNtdaDAA+
sg/kJWse1QcvfDdljerAGFLrfo+bzcZW4+IZJpZuo6y9jK5L82JuCFVCC+QVFbPR
P7Z8wHgU5JlsIUwOYpUpDqk/Kq0bc5muxcDoUiy/cOc3t0Q5kx9BsQYVgT+vHoA3
6lev2SI/P75d4XuIzX4B22gsAUMfozg9qMn68UcNej2AgrjgNUieL0mbGGIeWu/3
SVeSK77BUGIFYtIZkJEXYUwqNXuEMFKMf3EGokLcCT7nfh2Mqf2TMtapstd1XwHv
+9OSn5AzzxY+pP1/NwzmqFUkIEfouwczg+QNcVYQVMWtKlA3DJnQoRRqEsxdj64J
LK6oH+ObkUSsISontaYo+I9G7i3KwiLIcZv9lpP3+8XnIhntoCBlPl+5K0czOebq
IbwjVnzgRQ81rjS+6HkGYjMNmWyCJfbxd9A9+CgWgLa22k5hlcMIDmLQvo9EVe/v
4elVb8453n5LMUtr+MFOltScDteuoFhRmSzsh/Ol+cIRXBH9xwEQfNSgn/RxZoqh
UGrSfK70YiV9oX0m0uZ1AxVXqACGkm5DrGYxzRvyI1GOQ6g/O168nKjnamWDi7N/
IWy3Y4eyOa21lflvGQ3iVth2j2tDaehSJ6iB971uwfQ5NDLcx/gfzHYZOXj9qYA0
BZ+bJW2cJErJ133Mw/9I5to6alx3SRkNEfkRrkw9/8/CElsHXxylZzbl81kZJe+o
3mzJBLGUbNhpxlgPvtVdGdiD+UOzYgaZHXutwa7zHQpLdYkNVCFSspF00Df+VBU5
hPs04Lo/NZ7rsQ3XmWizr5X6wElE5fqD3L35Zf/uwD1JcztcqnQBEem/k1byDF6Z
46OuvwBQxGIkCt4olKYVFksypIR0gxcDse9gnmZReGNXy5P/xOtQ5qThHvlB765V
ae3bNvS74ir/Ymq3uruAgbvU0+E2PAZYqNu/CqrRRmdnlqx1Pw7WAGCMuMxbQV+r
dCnW5qco+I/uxWBNbJYjGEiKhr52OPIBOpEP4yiLFqhjKIPA+Rhs7+o8SopZvJqC
ibi+nkN2dP+bVPREUiSVr+84pSsrAli55CHGtiA9FdGLTu7cT5g7yAKy0MIJkX18
bkj8mP9u0DoYX6GAggd4o3LqP9hHicsTi5ENGnCALjBBXmeQ0sK39Nk1cM/3avVH
mMeKgn85r0n6bqNzUTtVDRQvNNYZD6HHpxiEO9zTsLEV97KBNn8NpdxivLPTTMMo
eMsy2/3sGN1YBSi/5Z+fAPTijQOO2TMEnMXgXlg61Xz92wOkrgcwdFPPtSUGTgwu
1qDNupYKW8BKMIuzfLZ3oLIcz4hJsN1RiClqXXdaZWy7LoR+bqGpWP8EcOV/fzGa
1ZxTHbOKg7NmOf3Tud0sZLZdJtz1+w9+c2d1QkwEmujXMYc3c/ZFbS+9JhZKOYsG
qIAO6Fp/PDW2eLXIY9xfXsV7EBC2ssivMRhqNjlZuGIaAU3D59jVFjXREJXi6dHm
RxBCnt8b81pXpS7DVYT0xMlxKZ73W4TPhX1yw0oBoaxuY3yS3XAgzNkTvjYSSOJ6
5sePu5woSd7DYpP04y4c8D6l84mtQ5a/LG8GhXs2FzaQTUBDy5sNrLECPxcUsiHo
5ugkQNIHgbJ/TX20HYd4+S94NJviz5VGfcXX2BmDXJrRzn7QSHNIq47vAsRdy6Rl
Em8ph/wR3rDI3X4tiXcdJO9/si34JZIn/yKA9rAgE6JMx60AHIa5lxOVarqaWmo4
I0kyN8oQm1Nd1J/QasRQoG6I0veT36abDbwrJACRgLym9VWST8zN7Ol32auzFpTR
ppe2EjIaGiF/0+QbgI/aw52S3JMa5bUDqyrykW8Xf0Et4WWJXe/07GpVYTg6lCOE
T1c6ZNHKGVVrsLBHCyM03Gtzq9OuX6HMa9HQrvqC+qdszClrhllaK+ZV9t4nCkas
u6B4VRxMReQlgYh6s1uUq/Nzus1cdcr2dA6PhcpCcHNuUwvriRLf2sDPYB5pwoRP
ybZb1P4cTLXifxjL4afOZU6p7QhBo0as6iVFzqK7cepDJ40oiMd/mBHeIbqBNzFj
DYkQc4FyAtWUhDjdRz/HnNjx1z3XAx/R5/cNYFobiTB02BzQ2vbc6OF7FiDl0NaS
48r4MvyH9wrtO4kgJN7L1NVS76Z9kew6+N45bhywfByA1lknAXFZVL51LbyD5i+p
ZvJTPnHgQS3GUtOTnfNXTivvvfMbYxxjppoc2PMGVh9sT3CX7oUaAMnhOg5j+RWK
GxsV1Uv4pQCK1iil1sigi+keSL4l2oaMT/Gph5hyA26XmwMGsfINdHpSrGfYSi0X
XmeZwu7iE1903604wDghGAS7dbjE9CEt8FL9+b53eS0tVUxLHQtzBQ3KBrIs8Thl
Q0XjhR8FkSPIdTQD+dy/0q6xDpGUgwkkHEHgcmpucmvaq20TbNs7m/zSEO+i3mdE
cXRMYhNX+jj4bKIfMdh6gIu9aaABHlK3wMODz9mgakcU4ZXYgPFT9wKxnYvAxnxQ
Ge2LZHsWqhgO9an0gj+SMuyq94TIJFVRV4+xVYLAR67GkuOCdei1EKA5zuaQG2+9
TLg17nrBnpT6iJcDo7T7Avkk2wXRGUmL5SPng1rlxQtU/3M+inYa01qbYI0pOcUP
egS4pBJt/ZeDsNx+cKn5yd71uRS1nYVnnfXiYP/Qd0VWlXkGYKKyOeN/hJyB9ciF
zTFS4IsE06aEsfDjevpXiIA53vvVWDSnHBGDYTd6rI25vo0dRdxzncozcC74WAQZ
LAesC+c3LFRNEddxTWW8S0XbKMjAE00aCFF4icVeUQc9pAKhQD8AGlvzwDvHVzsf
IxS96AOfxyxUP2wXsr1LZ6cvv5aQPMdlv0udW2FrUJzEW0j4XtfZoL0botcORort
SsETOk0Uvxf8HR4Y2mOudKT2GWX3YEpFA1KqPof8cnt1DPrQJ9DMRGMy3WinHMFq
V32+cb7I2TsKXDCrYggG44crKSTWgGQnRE+fHggW2RFeoX1Zsjlxr72hHJPkWej9
YbX+uQe5DxilCoSNeGNi5OcPlDyEb3zeWUc3BPiQB92mt8M056QxRaYrXIcyZjR9
eT7t/OLHvExqbPj34mokectPKhLeQo/VlhtL8bLR5H5PXnuIXYyR8z7wvY5zQ5jQ
Ohyr4Lo+Mv1ttaiWimVDWqZQ7/M3JyyXzhso15JEC4cBaKFhZFml559ESFduUVFJ
muMv6HwSWwNhRwDwfhiBfgzRRr2QhNelIbW3SV30xiMZUFzvtAnVud7+L1VxQMno
4e68Gct4Q2n+yn6DnNwklTYE193MkY+Y7dRfNqxqCQt2GoPe0rOe6Zxo6PhPCYIk
38TEIRfUtaitxhLe2fG0c1dKvATCezzVQzJYPHi6392uR6XB53WApW1aMv1VAD0D
BstzMNq+BIb1Sh7BP+cRZLO9S9gy1+XwnyMa1xpgYTM8IOG5IQeOpNdlkVYlL9f7
26XR9fqsGRBdDN26jlPobOihDqSyi5+fmTKQcktdDWfWm23R3Mn339XorvM0AjOo
tHQ9roQV6HoQuFu/162iB6cXVDSfZOtaU4FCADBVvt+KT+TpkavPXTMz/eLVAFKh
ZtVW8Pvbn87AYJPC5YOTqK0KqdGuSt2TVpOxLzwK6Hkbqzd/6n/iFa1k+sFpqhbM
7PmfuDcQUbMmrc3YzXyDpMWcMnjUZmM3vftFHrVIB5lx9rYSjuUpz5MJNTe3Tgtj
oonSCKoVKlcLYC31Rgil7wuInFMRHmxlbMud8Ixgpa7DmBCKTjqzHGnkidgKN/OR
9o+1bgbjkijJaZp3mIQbYXAIxDNvQg9vKx3MtwJoH6QMGfxVKjKVCKCHmQNqSeWW
Qw4McN2MVlweb8/em1NWF4TR+rpmRp/lsARy7v1h3JR7kOCYfYnnHwkk07/mDfct
6MeqwF9wKntYTXK0F1vYiRPa4IZs8kX7GxUReTRjvdNy88J9nQbc4Eoy1sk2KPHi
RuUeoWMwYjialMy0GLKQ/qaMgZeSauylrIMYYjwk+xTSNTo8D+yAwMQISiGPhZz8
IPUKsGiuCi0MZTNGpRhC3pOHHVoGivHKaYeg68TZkPLgs2xqHaHeOnAkW0qjfmFJ
SpSoKtHYVqfF+qSq5ROA4NII0Mngp48qmPOmF0HdZXqQKEpCH8r/P7+lpZC272JO
0SOnjt0X31t4reZP1XpMJpg4snG5gsdXXqZwidP4GR9U+PVtPjJTFlBzowfKHe58
kE8zHiW/k1lo1JgiTbCZNG5UGQLrWjRR3f2zPJFAvzj+laC3+nk4wzlbyIdUHJR7
KPyouJ5/Fzp2vDAoxVK+jR7fXYWfbrDZzy1eVF6Me1awHPiBM77e0yCOjGVO9DQN
kybT5bsig3wrLdPs3HsO8SpRVBeBYVz4Tqnh+O6GQbku+gqQtYmVRd6IPNB5jNjo
vW7PE5crZpbWHC+C8dHEUNEZqYslstvnmWBreVAPo3kBfQv5qaq0RemBAxqJ6CK1
moh4zWTWRsw7/NfrJii5XebQFIJgxC8BrtWY8Efh+qD/nKhAV0vj8Cny9l/HVEnB
LSrrIhn0btenm72xOKR7W0eyD51b4Ph9PUEN+o2lIyoxq0jVW/z6I8BjAj6W0zrC
jgQQ1jgF9mX0t6Kb1RpJwT1gfKvSHIR5rbCsINSCaWP1wX+Owq9Rs7I7GREWTvcA
X6GssPiHANHcjoMTQertNn7W/xYIt4C4uReH2hI0KF4qXDr5Iixqguqt6L2Z1kEy
QYCku/W77ahqWCH0T458ObUhHEDk67pNvs4OPpZlHIR51XhtXnRXiwucQDqusa7P
yGJhpKHw3svRH8G/zrOVHUw1r0ComW28o6x6aM74VLbHgBrWAiQChafGEnXL9kpi
OVTuRhuGBsu1iNXS56hTp1akjHZHFC+zjmM8TlWf/nM0nagt+R/ZNJjHcqKGzjWR
IXirxZcwbXjNkuoPVWclXxWSNQUDaxLggW3L1mhdSQc6T1amTJs0a/jVu7ErQrEF
4JwDLvewAtKdFVorPtmmWl5mAV+WEmxVAEBx9L8rUPnNrtp0po8UCybXdHHQEvHV
CFNFcmIdELBZlt3DAP+wM8gRiVpLGh4OpwA541LMWZNq0mPa0xQLOXcqqbmTl/hT
3GhOCeGkpzBjTzdFFs2ewwYEMkOs23E1YKrCS6fxPK6aI1C8WKbRaUG4safdo6Qx
gzToReqMS534EyXVCSU/dbz2oKF8X2WbbeYerbGCIKB87rFJtv4P+PrsjeMpIGXa
snvfCohy+k21dkEr/fOTh/txMke/lHPbTljeEl1Y4n26pifjuTvwfc0oKhqeVtuD
oFhlESnMyanHLUdZuKv2Yt7Z/w+PdzE41OPar6rUWg/E7VynSTNGirDEYRrIPMpq
9uqsATPfp8qsRg8rdJUVrbNYPAhRUqdHCKeLBPVf7cjz8lckstFCZBdzu4Fnni8c
Vea+iBqqylsW7NMTDQtGFSjPWphHsp/Fy5NLjEufOXFHm/klSFlz/bstiKZrJ2f4
WWEzPgzqYxVxjOVyWuxSLBxY6rOY4Ty6f+ph6sgy3GYj88BmqMHvhwBVkdNf2207
4L2AOPk4FAAgCuxUpZKnN7ihHmbytwJEd47nY2G9GFyqjj830vsqufilIT4eaZnl
qsmAqbwQ4gjUWBOxaxZeXoQhVdpQ3x89Gm9cGDtLZs7YNYm5DGM7fX8OI6hMwjv2
ugBgRdBCFwtTdu3AiEwSYbhVilWJJ2gn85AdIbUMhimLRqwQdvTJyqY0FQWAccX9
JOv+CKF9X/0e03R2sxxrhO9CX0eSKP2ovcbe52NB14zRdchtFDL6rrdTI2U/EmFm
S7MqYbvm4+SjXoPCkbDxwgBVPE2JCd0WE9CcJ3IE8yVDTt1SahbtkWWr3jbbVoIr
cfgjyYORG/9Gg3MENOWFfpHmYQt4ec0Wa8HOezjKYMhU9WfvKR318jaWA9IiLD1N
7WRHoJiNM42u4uH6TsVnaFsuJSLHzPMb6+pWlLlAPI1XE2WUFfuq916gr0mjADo2
OXcz8l07HigndIuG2OcV7LaDDAP+QtdhSFkXsT+v1MZPCFYsZyNZZVVXKgQeQzgK
c5dzQVZZUN4GqIubKUN3sVktxIW6bw8H6igxuXSE+Sal+5leeuzTmql9HHWkbLYE
EGY7u5tGwJhpecKg0FjAXZBs8m3v8kt4DOn4lnWHg+oPqvOR+n9j5s5pDVcWqMp1
nkJpfBjmP3nOqvSfElBc2hGYx3CsdDrtkOvhqSsR27Pb3AYjqj7V/C4BypVpbvYN
FZ9GAzrz7YZFZuhs5myIOod32CaQwCYnlQ7e77aUypKBgZcWUthPl88oNpoylou5
snVtFU8dMn66ZLi+JW360ipMv4loUxC1H3DarmAVuHlKpB++PBcyTOEqJX1fZfsG
qmjNQ4JcLWD/CBE46c3ZqWxr4K9/0e+fn0/GKMrb2y2qEgP59GBKEKax3gJoaciV
mZqShx+GUF0sjzi5uVaNjmr8/VNHWW86iHPlcKTAKL43DDhkFPCpQvMAmI+jmlSO
Ov2tiOrln7VDv57j96FLyi5IXQK54zXX+b3n1SPHbfSpAnojdQ9EuE0cM/oUc61u
ptAcF3he6vWxlhNFxG0Y7/MjoqRzXTH3zPLIw629vAYtda56zzJfIieC2I+0ZBu4
99b99tSHBQlQoK63rrBxe0qQhOqpwUmOGJOvge6LM2xZVIh/qL2gMiBzrWrAT5cE
8T3Ak2MMkhyqJuNqUY+l9sOoxWmB2KLGy5GuqTBciSGbw++86igbMUWguvW/El8c
HEgiakt9EdLMfgMA9eVogCLapcHtRlOhtuCitQkJzdQ4V4ei/aYqljl9/1HtwcPC
wzRLDZdIVfERk1LmjNtW6tQHcKfAmLdfdrO0DHn0N8oyv1l/VICkUH6XgyIL3gGM
jTsSbbMtT+L/fnRgj+xFUp4gUkF/Wj/3wRqBzQhjKO+yc2VqK+nG2ngtIMjI/Reg
iQIkGRQCnvj5NJXa4cfko4lMWjgUA9MdXNqsqPhtr60oMG5y6Rv40r0+gNRX3owu
+M8MoFM6UkTkljtrWf7plit1xi6idO59ds8J71kk8GumwOrJ4FRZPjF9WOQQnEeQ
yLnATL7b4KZyx2VCAayicnlN2Zy2pHXqdPTAR9svRm+tcDCSi9exa6awuR4AxqvQ
nfFrE2bymP72+fri9B5sY4+2cJfF21SuP62piNSNr6mC6ow6/ROFKmqRn88XwN6c
zKfCZ/Qwnyd7lpGm6l5Cjin/DGKP7PQ+zC4Juq6wH+lATCLusaGcB4NltNHmHzdK
Ma7Hwt0mJfGpPfiIp4AiMu6QnxzIRf7okhAtqXFcXIO7X0z2QgbrplIvEIuzFmr+
m5ULo9c1otQQ8enXKi7Ds/vzei2ZIjrYp0mSu3ZOwFmukWA/gWYo9s+awiOF+MS7
on2fWEkAOgLrl3A7j4mTa0ItfGzho3mQgshCQcDtKXH6MLQX3v1MhqyfilFYMXxg
0fPdpuMbJa/M7Nf9QuB5XjPe/KHGZ0CvCW0Xg/ZXANOzF94+rX4QYCgQ/5lS2Y4z
nMj8P9AUulbY+qofbxR18JSy7kNaqTU4VRqAc8Mq3/mnzZa/2tZLSAt8rZ3X5Lx8
46iHgAXhsQ2nJc0wdx1rWK1dknrmcYsXgA48mzOe6xEIiBDGOXgI9t4WxBTqP/ZY
CcUFN890xNjSVhyyooCwWbtPW0udaUxFLZ8oQ2finNP6YPihqiMJdLs7Bwts/6Xe
gj+Tl7Kq4ChF8IwUgjI7Logi5EHL1FZoMrU4rMIyhHsBP4zkO73CQSGln/rgRj/N
Ld51TLSBdfhsfjtLvMBO3mAldhfyWzPYgtFVN/IwR1O3EN1uCm1LdnaZH2JUQyaG
FyKu3Zo5IavCKM+O13lFUrGCXQHZb0JDtTVtYUqeCl7nVMC4/ALEC0PrEcBWoTp2
4Mf/AAdBwnX26pZh+qLJzpYdka9Kh+39o6EgmAB/6WbtrH+J4GPdlH6GEuFpwIMu
1xszEafUl6nACjqE/po6eKHKH63i9UqRIbSGmD9jybiRidQL9QC4D+UmXd/nWR0c
BE3B2QaJgbL+EO84b/VvvAw6CichdxCrVuW/b6ajJLm3Gi8riTpNkv4JXneqTWeh
n0Y+CZ3PhBlEE1LdvkvL1zRrHd6ytWrubB4N7XU2xsUYxfkRQf8bRcf/p+8CnfVQ
cJA/MWILU09A0n7xlIa7ixbPy35oXeCwpfWr+ffVezPlRFtCtxIP6BntVqMkqPAH
vi0G0TO/P9cOKZVUUT+UucIzjvh5RMT4Cinn+qm7doOhmn+o40CDuOf3YZGe8C/r
9fk7GSKByxMeoYknccaWN9oBpU34XmZd/4Klx/evVDfudoAENkW0erO0dmT9lwE+
UUHTcVZwtCW1JK3SYSRTDs+ca9NhGvozQsW1kOPw5FHVRMerzKOxVbdzytvSC1rJ
6+mWVmB7d4J0wrcwoJfGWDXMdLabH3gLjly/ace7xjVAkvu2cNwRmeALy7+U7ZUd
ZZgZL6J7Ph5ex7qCAOL3HfkMbhxjq9rASuxgH/eujP+LDyQuMYO0gHGTEPgH6zz6
zLiKvm5rBmYDbtUmEq7f4x+6eC0KUBci4AjJunn5s31Vp1Cwvr0mHKn6O0rarfdm
5YB+f/wuYNcjr/DiW5tZYEJgnWspveYMJn8jTsCxDfBAK40ayWzJjsM1VwwgZTIP
xgt53Iy+AOnPObixLOAnT/zVlCXL0GJVpO/or3+JKn3fYnM3/SH4GVXnhHbCfDMM
6CI4qbwszbnlii7P26vV28ZrlR7wL+ZbdTjZFqBBHjz+Zpy5DbHG4fqTspc00Qgv
76ZbZn4pKXkRTw+kV13Nb5pbqph5UL1Hqg6/JHDPDjEH4OMFgMAGOxM66joieAKN
gfNMkkFBeTe6m9bWq8+eryeZB9q6QTy5SM9UV44xf3cs4GbROLyHsjaU6uLYjMC4
5ovHSHbeFk2jA37V2kzocD2/afs89y9DCZu74gmLWwIfnVtAkSEv1v63WuH7H4kR
TyTIJe2rG1nFIlK0omN2NWNVac5/KV2CdVi6afu5Q6mODtzfWV9XqvA2hhCNrLi3
nRIKajE3Yk7ItVKzy/tiS+61ox0HeHPDg+QI9Eyi3paWI6PChcCMdyIqHeVZ5RjK
vA0id1q+tDUmzrkt8UdoomsDv4SnJbbvJB1F/ZE//oEVyr5iDP22B5hRBUz/KGPx
5SrFx7wc5LcZhFX92K+hmcIPPodQpUBaPkQfx6dIFX1IOGchZbObZQtnnIA6fU7L
dXVlZqaJMxs853OnfTuqVf4vBZB7uHaF2r/6QMg5DA7UIwnfM7SqP4GawTE+xyib
ED6Y7+ImqtP85PKJ9ZRwrw7bHhHEUHpV2FvhMu8WUv2tB8Jf8ampZD2TIa6dpQEt
Prbdhu8AUJqTtv24+0RH7xMo11sY32nMkqHqxEprt0I8Cwxe6xwSWX45yHjXpDmt
lxAkbugp0MYOLNxLUmQgMi7DCefDWTGdS+hDR/ixNzjvLeftO7TxWQ5uHYkFFd/B
kX3oD3cd5P3aLqdnx6YWjPQsrb/3mz0kKZuDBOlKIt6ACGLhsN/pUDMXkYV0h1By
9uWudXoEiFRbaElcsxLLt3k5tN5aW+XcdaO5mBV+NT6eNau8n6CP3UjHHKjmKtOk
wTQLLGO6nAgT7mxtX0HZmQNsmquBJCcn6MQaa/QoatFq2ZxRjJNwBEYxZichLOAv
DMl72RKyCbgYxMTHkl/8i4LjL00wy32DeSuvTvRfxwiwNNxab8Ci6YT6+R7HJjCZ
4U87M6W5IaIWZLYL323TnFHHxuRW51KRORO9ZcEag4hL44FvK+/8fUmmULlu9Qbq
ib1Uq5F+em0DhPkrlCeAmJ3ftBWk2nHfdfJ5w7Pb2fR2WyBFKcpV53xro0DMTn+q
b3ruBkLsvW301kJvkk8cyzFkdEKc4RajJFF8C9DJQMEsgEMZLQ2C+DVTvMBoqQrm
XVeReNt9PE7DUY3BRLJsrTOCXzgUAkaM9ZFAFmMdqoNu95SiBh0J0NgkoxDAmIiI
kbSpu5pqcbaniBwpfdnk3cUY2zZDT8CEuigRyIxNQtPDbtoBAmM7uFpuOBn/x+w9
jBHJDV8c0WpUW0/5U/3TirqREsgtqHrG/ycdq64gOP+jXy3/oRblT3cmMYzBADa2
corwThK3Q8WqdUxRD4oBfhrtIvLc32v1D1cAZ/7oJgbA8vF0K0j1+JILEhlwF292
3p76FYWe91aW3znaXKaE/7PgK16es1DoGYQ/UDWiSYoBFtlTAUQD/2QIz1ENEk2B
TOuGey8wHPRstbtVfELt7LJ69wf2EIVeAazn0sMEGsdzCj6sgQycsfDg47b1cbp0
2D1Hp0H+80uPqXjQ5jXWnBelpoyzZrpBk2iPrSNHIBZ0ESS0CuyazykcoCXzqNXZ
gW1OzBfIRvm0jQ5TvXVvSN7gYWAhP6M3mXAuiuUyNT8JKdlFh3V2z5a4TL1vapmW
l+rwE6FYaUNICDjGyx1Z+0wbdKI7P1HY8nr6AskLF3ja7DKCdY1R54MezB0I3rFb
MYZsjbotdpSHFYhceXUIc57rqjVE+bID2tnHjFpDPrx1OyCFsv2ZhWGclU34su9d
VIi75SPh/w1o1hoJY5hdFxp+OUW6rIhMG3NU2z00F2OatyEGQlq1TqK47Lm1fOZq
1mvBXSdvW/zPSCU1X0nRUDWxjCPB6bLrDJIlyl7HAQnzgrNQukWWMNpR7CHuqQie
5dDGYMkrzO8+ZRxEt9F2W0wwLZU+LZT5yFL3E7EkjZk64RvtSjKFbIvuhuLlmiVC
y8qWmtaH3NQU087UkGO37rDKmCq9BdB4hrccETwRPeHZUAggedRhv58rRtdu3t28
oA7wNrIhLvpSBw2A6o0YDC/PiEes97xBB8/7F8lnlW8Pcpw+MXqxQHmYaGdFgAJy
8lSArfBRaVh67kZhnASbQGeem08XSBKFz9K3rZIW7X9YS1tYn5KDp0hmFxom41Ie
6e6960vckhaXdKwkVoJSFN6ZmqggNTqlHg9yPHVgi4f11CG3ObBN/awRahumFc7q
PIoPJgKaxzWvI33jXze9uIjLzZGtvT+Uz1HU0b+Wy+jBuEaYc8PXtMkGqaafVGZ8
jVe0u8mUvvCfG0ku4u0p/x15E9ZHr+xzB8gCfnnkVJLj4z3hq+djObWzToU5voeW
9FxFhyWMqlnsCcEItzwbfqQYtlGwz44z4Nj/KqlreqZpYrvd877m6blg8jHT5h58
obbRprpoh3FQq7AE7Uj19HbdMvS2KiDfWGN2VQIVHsSJeHmFww6qNHfRprpCJogD
r0w/EtCRDLEhyQ0wZyCDLjfZhNDywCrpWESLQtCt/1hwltuuwJ/HUeHQ9LRntIMW
zPzDRTZ/KBl5IwmtdacHhleerYykZlYngC9fhy4ltDB6s5N+86IGya8JbyFLXpUL
XTT4pV0yjvy0e7nmDjPYYl2yRp+SJa1qsoGvunT+T8C9qVWVa4k99DREmtKu+5bC
LzTAPGaEZ3hJWUF285BFaJVadEGWIUlwV24PzjfqcI0aIUDf2YHvZ49yMCnHaB/c
mARUs2+DBnMvTvZWbDa6rfbxbFyD0BtgF+gnckm9JWXNNPvpX6cL7atWQmU6ORhR
HQBmXRkG3iKo6ZJNqYPfgY5BTXQDPsducx164McfJF/GtTDAnYjVvFaELC21TduQ
pNzXzdGj2++G3t9LeWLnjS2eJ/wF5z4rMFkgtPo9MpanDE9ONXmLPFg8fYlLBAIL
aLoCmdSj1ZRWgtaXMx9RXQNfK53x5yoxrK7ByqCP/7a2w6iL/quhns4NEkUeZn9o
SnHgXMNYvIG+DLKgiFNM8JpFV6O3THf4JFPzd0OSfwsLFTToJeRAkHu9yOYD7kR8
jA9Bb3OX+sImSHN80qO1f/NoLXaaMNtoLbZX2VSfZWK6+7L3jt99w2R6OD+XUlZq
FCrTucfKDmrKomnKmP9shmGF4BBSzjF4iOp/GW8CkXBwrXXncnx7I67hVe1o2oKG
+2LU/a/BBfzBValGxBqCgQ5zL/TPye/eIn6UTSFPL9LUZUEYoNUISI3YZZFMdPH8
rC9MrH6k6JNrN+hMVqSA05UpzEfUSPcfsg5l5JI2MPyvwSxRyueUxluL0ZLzdMf6
HEwKiTenhLl7hKD9O+eEwE/zkz6kXDrQNsYY/5KCrx6mV1QKnApcpvayKwRqGM2D
k23xIfk8Eb7Aor1sOwj9pq6LP2WiV0xG2kJtqADCJgSHsmLx/yYsedFdHJUXLFaO
Wx0xaydyN2cYBbD+nNTZhfVUCmjqCMz0ovBZ38OUUNBFAg0SD+6yLSVbXj4CwSVP
umS4WmKvfkaF5+YksxaX+yNuoqdo2e7pdL+yWGM9Tojg3tjo6tu7M+qIYWnyERfO
T7/hc6cANFbCr/ZviL7aLIV1lPslO069BC//0W2eo67rXpgLxi1gZOlN4HUVFTLg
ci0KsWlGeGifPTIYdSp3MOy+TEeXCoEMntqldKkDJstCztQxEN1wfrZzbSY17l5i
/dSRYnWaVfBclrUyfUcwzNhEE6rnWoC1iGnFGOBoO2WnEo1K/AGjZvZ/f6KTYTpm
rsGfsRHtEB/H5iLmz+2jHgyP4iDqXTUTjejkCYf+TWf3r+/s/OCC7H1m8XBLX+W8
saPARx/LaPYf3yP/binwD4wAsSlYSP2d0/QnNGtDwjg+tZevoDlalHYsPcMeszXn
LyPQHdgT6hka0zI7PQws59zhEYqIW5DZJebb6NKnzewZpgKMOufTi51smusTW+TE
JpmaTS3zsACaIMdzT4yXv1WIiwapsz9ccftaqZ7n1aSjvQaNJxA/SOyecLlXv2zs
BtaDY4mz2ckRfkGO0MZrrz0ZExmU2+QdBJUb6IQbcS93Tbu+jBCLMyXgMkiBf3oe
jrLWsoIGUAf4mIynke/7OF+ID1BUi+OqW+qh1yonT3y/lwWqOJIdhPpHKnlB6Um6
ySSbwXmBeYT8QMISBdtmDmzErVthyzQsJuPxplRyVw5o9YSEANdfgeBApMZDu6Lv
I9nU4t30QH7inuzrh0Z4Akbn+424UX5tQvN9s4f+XGUrLHWTMQskYlgGHzGXSVNw
QV2/d7WVxKiHuE/7ij8xVgSw3EY/pSZxBtaqyZZ1CWhjaEC0/JATCQbPyrLT+3IW
84oioZeXSdFZlQareBEZXEiQ6ghx4nm7iPNHJAx1kd3wCVoKgDlPalSAkENZbEEU
ToJfM1DRC63B4VASvSuIfnkdiDZzEpsuNasrs8GTachqviu03J+pknmDD5XzHAqg
BfJKAVbV/ojUYtcnp+Zl0KiMtoZVh3zSENbKHZ1WcMNobWo0zxHGfpl9riMFCsig
v1/MuX7+8t931cIJAKDVWM5qtmWthh9GxclQMCplgPamItgI3fWwMNWofYPa+zH5
rI9Qbqv5YCHAi9jNQ0DxqynSLkjUV2b/mC2gi+AwY34dL623kfi2m9eI25jylLpj
2Bx9BNDp9ItJviqhrUZ9isrUoBNIRfYoxNOTbsjUJNieT8dBlD1yWyHmcuzEVlkS
VAbt6BPk63gZmvZLxfZjycPrGMgTMfsYhDjpTSDWqZ7/J5pX5D727GGoFo75xEzk
KG7RQTt6WdmPsJxX4lWNgByyWDFHrRTPTO2smvfOQfHLOGAYAlmJ6q4M9ux0327t
D1GHGDHNh69EtM+OOQmrFnvEOC1drjAMH1CsoOD1urs2oKVnWviyaRHpRHeN0Zgz
N0J2PjFpcYpitLulfnbIPaA2Oew4XdriO4GvtJ5bGbAVKXk2HQCvf6lkzfNd1pG4
H/SXWPb5hXhEtq5DxjdciDV0d4J60K0gKtv35wMn3nJUIztG5OwfDH2QippVpFVc
zP4BWe1rAgTh9x85itPbD+o+F1Vo69y92nsSJm7neb85wgfJPklUpJO2awLo0qOf
MGmgiyelpkAQ+wN+lSS+Jz1ujcmgd0p1Hfur1HV28NRK0YRxTl+LPwFgJdAPR4fC
3jhg+aqdfTyWGajxLxtLaw5egRRQBP/14nmOSetmLXhWX0V64M7e+kKM+v0ootii
eNHoq/86ezqnTEeigzx5tuFMqLxBjjy9Kg9JT22B/KS5zKL+/P1QooPnHDVnvTft
TfmaWCxLR7PgIdaqkQFA+Sqr2uBJVO6Zss6wHUJ5AFcTQTD066Hfekg53Mkb89Ig
3HQ8T81ygXvis1b5S4jtkP5jeiYGPozJIBIMQni3wVNszz5lf7p1aaveKBJS3FSY
I7cMUalo3TnuG3x4t0XeoclLshjt4zhwOPu3gBa+Iw3lVA37NXeI+eW+52560MA2
jPUqNY617Gf/kRz3dmrG+JS/5miz1/mP3O7PmxpOwAqeGhJ5b5jogfJceVrEb2In
9cdReA5Ls481cuVdPO02mi66oMw6GDN4Ji/6gWNIBCcfDA6NHETyIoJ9lItB86rW
y3GGuFst95YJnDl4C7qk5pbgYX37oQjmET7NdLQcAb2ScmCRULVS5lDNKhYvCNZX
xXYGgMt5dCIBHv5pY4q7iV+En/AcjPQzvT1upTbIdMt+l4A5p6rs1tW970j9eER1
KMEwVpjaqcl0ISLU3T0bbE6iVfg/8B2/CXbeH00l6wbWl1i3x2VPkrnroAb9PUaS
9pvDFPrKwhDNcXCZ2Gkq5Mv1h1oP2SYUvQDxKmikbH46/en5SKbGmfcNJSS2adMS
K1Pkexl5kqB3G6WA7bxXVzlxPyXmnSBQo6yaArPPhHOjxFCPnHs2wB/EunrfnRVt
gM45EVt89CB781NvZfoCLM7O1U8n+D9x9vLENxH8tyzur5NAzDDupp8v4TY+TlCs
aq/V42kYqW7oMY9mGa5YU5Ykj2frefrJg8p0FFhceQalhj2Xmf3cWtlXla6QwN1o
m6jGyPL73P7Vi91888F6RGA6Jz52UVxmc8Mdwq5U9siVmDJVUS4lsoCNNtb8NJOi
QKYc39bdVs8saf0DhklRcIgj1NrhQLnF6QLUfqXUNeNub+y7ttZQXJRCdIQaqJBU
NlVRfmlwg8648m+OTTXeb7+B4MDAgKDYC2uBaeUAdZ3fwrgfaPaOUzdJfh2igagg
jMdC33QWVRuoeSo6WIg2GZljzVyIl9oUIWZihxbryE20yWkkxlkV3lDFWTRLqnhn
GIs/T3ev8ClTKmo84D2u2lVA2M77PLS5mqSTecovLcfl1uuShM8vvAwim7p+qLqQ
HrwGE+rWLm4p96vdz67BtkoDDWMyNOtVy2Hrpjv/XKb5ENz7Pk4rzvIULvaaqKfK
1Vb1d80MFb2aKQ7XtZaAgOV49dpCtZdxTN0IdZZkfSQlqKPzOCQ06T1EXPYXIaEY
u01UIhXPnG7AhQOstbSu9bEyIA4LqFlHWBvOO5JT/lniDZrbm8r2ikRuCkS2slId
Ayj8FLRU6ty5+JsgEGVwSyb+kJOADkoO0oMRt2O8I4p5qpnxBz2a4FCPCDbfidtG
hCl8ar14Dj5Ct0rutRnKf+VUcKRwXu6zivZweTISny5aG34n83tJsLxjP7kxTe5C
lX1//VrU0Dix84RAeu51mFjuY/xuzHsX0k1H73VzwTzgf9Lu+QhVm5PHXLF/+0Zl
k0NzaqmUtfCjEAPGDVoRu4YJKhbn+/Wx4CENRxJnJP+IF+nCXHtYw8iYOAIRb73l
38h7rEezTA6waujUHjlvoc1RC+95EVBywCpUbuPzRj52XMuyZwDqVcsUZ21Z2Mex
DMH1KgpYarLO5t5YKgg8CXzjqjElbxFyni/rfzSYXsiLKzVNufkCyIoBkdz+Ibl2
64tAmh788NQdZk0WF0aV52a+F40pRTKJ4l/86HtYcZG9Jvh3Xvvl7COdd/TCMYuX
inmZXdHVcEcLsYTvuhaGy9YsUvyoz37hH0UJIgLzW8rTUYUNpizDiewIG6+FLUWl
as0dJjIzUHkfFUhw2dpJnx9anBawuM9TgIHMNM7iTfxb+NWs20WSlMNnDnDffTpe
P9S1ipQxSc4lwImbpIGFQYojKfDuLz+no8Z9ZyGs+BUWb0Ectofm5mLwkJ60eG/n
qsLtP0JUVx1SYxxms1kz9OjG467yfzHxHjPMwVxpYPoK9LqMmVb51vgsBIERMIkH
rKEzFztqHlYLgph3Ddfj5aJ2rANjtz2ssNSVZAYNr8jmdNU2aL9yRB9+A6Hy1FK/
Ghtr63f5HD0txCDU3H2g2v3RCduHCswyWcssiwZV6Ju+LrKUNP16VNShHC0IBr/L
lAZZGWaa34WUH5Iy3npH/FDkBeG8YgOa4BcmzmNz0nlVRWnik3vOHFNh6CCE59Nn
g5VKHWPMmHE2GrJDYgIm6jpnYmlkUScpU6epPSVk6V1a6FgLQkZGj+krvfmB5gY7
GjUuKf02h8Hk12MMo8R3uICNSOQSyB43d0PveKzcS8BxpvCmtswMyYB/xc8dXdol
y9WES8FcaxCe5Yru2YvYlarAp4wicT9FtQNJ4/+CWBrnsoHt/suvIUPFWoViE5+u
pNGyLCaNc0UrEj507sODpjjBd4XMnKLQYgwkYwY+S4PRg/bq/diHR6lahw0O5EiM
S6Wh3V5+mTRlt5/xc1B3POcDtywnCJgsGr8Yn+iIJVyvU4wpRZbhRXC3X7d9sUK2
PxJs45VS58R1egSqD3asrgmQUFtCUpPKQTxsE/hNQ9tNoUfTXReRz3xa4xx4EObf
KJZL4S6FuqPOsIZVR97dmPSBze7P6rMUyv7Ynk+bL4ryazS5KXM/awI8U37sZ4Va
YMpxMXG0NBp4I4P/kmDb9JeWYNhE03bVGpGOaiAXVEaXQavG5oL7v9JXLNt4GGc6
bObiXYQ7Wty3ykOiuSKDaBQJ+A2I0K3XVWtvZmMc/TL1FIfbqSF9Bjx+gPKqLeT8
oJbQoqFx2TMGYBrjCWG5mYxf46NET8lXkJ0pCD5gujm9I2dOPCbzuqa4MuIRL4zj
It25g0ys/sT9ndKXvXmZ1vkm+QXbjPxruKXDBzZjT2SgpN/nRfJyhU5mjKKOsV0w
mR85UjHFwyZZS0L1fQbFqDRWE/V88RUSDzWANaPNIRHXw+1FfiTfzueH8XKq2VQa
izM5iI/OeCB4D4fk854z60/AWvEEkyJH7eGZs0GGJuvxuW2aurDNAixZFCBRCNmJ
LAxUyPLVCDeQrm6rXcjI5GzcAkBVbBrnPVqV4EvEyo2VWq3lfSqC37RZ8R4cWQw7
TiTEO91PCi9T0ahPFImWwS2u/JkkVN4ve597CvjnJ7Cg1mN4v+cdLszUbedErDbo
UvCTdMozmCI0+O+JN8PWC1eWj8H/V2ioNhjWlVoK/X4KeRYhG3d5Mf+BLp7T6thQ
/8gfA04h+62NucczqM0WQIsUW/dFXLP60NYoZdin+stxIwcBtVXfBRdcf0ZnsNoy
8zEvDjRKKsaMf5H54pU8iRlwc2WWf5sxTRaVzxbOA90L2fgU8YXFfHDR5lFWk63I
OxO4WIV89UC3udNYHhLU7Cy7yZT1CgUm4Nd0BEQrzrF8ws46VxY2VrMNIEsqcNfV
ATmBg5DFf8wGIJkXY1+OwEsCDvwtv5wC5dXFeFaNSsTjxrp7q8opXzc+isb9wel1
42NFELDJxvmby/t4y5RWFLs2vmJo8GZbkcDgipJSNbFe8SGyqbGM90SJf5BFTi/1
K6ZnjYD9gS6/DDM+v36EkVnX2xtXZocr+/7RLEqRXsXvs8bPfU5gl/XZiSupqb+2
uhiPiKmv0+/ieLnpWMAH5jJnv2Fvmv1a+YH3amEBttdI+AjEX2gt7bBE3DXC6LhX
BMUGDwOBch/dfJvbwyyni4aQ04r2obtprV/jty+9auNmM01hj5dTJ5ZofinXU3H8
LjwDQTDx3VbU+jPxkvBjgu5adwByTM0/GkgU0D9kIjc9xB9BFrKIkMbMq4sU6za7
UWudTtx9H+pM1mWkZ566c3DplpHNp5oIRowIbZ8pXJ02TQ6XvnZzLPzrw5RaAbNw
cOpI0hgdWcTpVe4df5Z/hJkoTCNEfrWf/mvLskqko92pYF68lF4KgzlXBhLYjL0k
Ycq3V3WmzbSwcu5bHw1874hcJtyrCM8EpqZQxCkI288mkisKIeNNtuaviThwpqjK
FCTetKOzUEDpXJ9aD1bAo+ZgraDef6apqvkga7ONDUOFAN0wpA+7CEc4Sccv6xgA
nqMB8CRBGKv91omHd1tVAxQZAuOCxqe24MPMorUZD2Akj2Eq6EoObK2PoUphI4WR
QwQDvFqVM1FtfVoFsS9rNRNot+ZqQee6DKU1/klR3M6eboTk6uFP11Qp41EOmhtA
pDLAhvvCLD4N+nEi7puBQ31wZJ6eAZynczLSXLvhxTRtJ5ZAt+AEUm1/7KtJlaf3
WvqGplo0LE4TmD9DXnUXHf49UZJQ44mGOJDcGxmuYkAONJDJsVIt5TFgwER+QEtR
EPEZlehnmTS/m8cjlsqQkt2j69hgt7bNr/Yz54+ASR51Hh7e54pfTKASkEiChJWk
c1EXqJiZ/TOOHkiKQ26e+QH2W+mfSmg63a1NmzwMKh5bv+Mw3vrU+OFP1fJSSiXo
JrK0+y+r1LYx/7lvn4HX7U3MYlpUp6sLJCgDFPmhCpFg79PUuoPhBldi3NVJjDzl
Vu5FuxLglL/30mPi4MO4IWXSUe5sarXg5PlBUq34ej7r+g2fNwbJstUbKmkH+Q6c
haC778SmeATgVxvmrfOlGjgUOyS3XI+Fb88l1ZaebxujnQjeWFMH58r6L92elYU3
6k8FzqJdlhEE9PQsoFO+MHGfvXOeD682qMNWB9wpDEfyQowUYNzHiBtGeUOl1l3S
2IzhUd9FdbJDCrQI21AD9NlIqfuQs8fMQ775suJf1UBjVGGgMcqbf3S0zHqmBNXF
wu5rfYTXU1o3hsIiHwZR3RMtyaeGxYCYN956rP0N66tjUjdTIhoeExoHZYiEw3w2
+mvNxALchqRv+Z06XRZZuHs4Jl+TNBUfun+TOfMvHp1RQTNcoYtJS68rXg++6QxM
EFtrR9wmO/jtPkCPo64EdJkvucX2yoxKMI/5WpUNbxIeRWmyxb/+DAgTxP0IWGLp
6zYkZ+/9Am/Ol46uTFfo/3MF1VHmDcaGu4CEcLx5Qs2+Sq1xhXvL0UH15syVco4u
GM8cr0pyXVc4lh33ihj7nfzT07qNU8vrqLRMtpTEKl3TulzDWxQftcu9xU5+xTAX
JUE+HjXQCmHyzkMn1OBJOtrmGqNfCXC3cgYQFRoyK6R2PxQF3YsJ4UheGFTYyqV4
Aha4MIbKw1ApZtw3j6R1t0wCHMgN3iBRj8J9J6CO1Cnn73cnNLXlif6KRIyArEwn
vIQhTWQqzJqnYLGvsAJDlboLQ3E/ZEm3oh8YUTs9nliOucR90NPNIS0+fgyYyMdf
z73PjvYsfGgmPf8itg2GrnwxMo3H3K8qEkMR2niLKjHPIL8Fa2SrV+TrTpFjMnwg
MDorUeuvo8jW6cqlzr7/L7S0WtOhEh5m2auWUJKkNSeOZknvplfbRCBeOzPdh1mr
ai3V5qWYbOURebDh8QElGuDMG+wnBntu3Fug0h+nXv7IJV58lcJPIeCSb+jLf9U+
OEGSyixb1olmcrXklT0Ho8zygj8RlL/kZn+ak4NEyVvjKMqb6W2iugOTJsFKIt1p
W9h2X9gDe45ti7yyW8vfBYR5D8fiam022olG3dG1xPsU4hRvMEO0uc5Pj+JAQaxY
yuJOBgwgEZag7Nl96SUYdYLZNyqzwDdxf6gu6T+DEw2QVh0/qHCRtM0Vt5BBqzPN
EP2sBuYWdkXjYlktPgijYDM5PpT4/7MDGpjLu1hjPaFdMtsIXUnQ3n43FjZRSSt2
PkYkDPE0/Piz1jehnNG3wT4FW/uA+xRl8JzXNn1iligMgmK+FX2OSTlEJPPMSHC7
SFRvi4sMAhZGEnO87M/FyMk4ssSP4Yzx6N7QRH6HeRCYBRQCbkzoKztbVTK87sha
V4o5loEOgNN3X+6CV1Dfd7UB9ymmsFoqeXkHUYL3hdTYShIkWx3qKRsVdI+9Irv0
3PHv7KeX4/8Dm1Z2AspPJmxnNEEXxQLNrTYIb5z0RPRIe1xgrezCPypY6uhzDA4X
zh/gwrk8t6rEGjjxA6jHOCeQ2W0mVRyrJcuPjiJjKlQbr3EDP2y+g39XKfXrKEMC
Z3FEQC9V+0FclN2FrhLZRKxvRA1akviB59CFSRn/FbEs32oYOpGrH+NP+HdkFhTq
pnTeEIHlhnerqWi0DsTNVncH8PvI+VjwFB4OhLeWPQJajeHVpbG3Jv+yl9hOpBsB
2lMb6elrANd22znQA8ZatngMj+om3499C3Zk+mlbNLKUv2EWPEl6OLFboMASnPva
K+oEBgX1vmvs9j8emLWrSwxxn1LTU8q4n8lvocXzxhH/so3VcM2HgJHBPq3vWvqD
oVlMLL2iXq+3gGdbbKWVpf+6c2W0rv+LBEzeTLbHN3MH+tU+TivPcR6dYlUDxZcg
QaGmu9lgjmkOtoQqm9YtKMDgVWMrLuCHg0O4BjmXX70m3mxLj4HFnv4a68ClrFhB
+R8KsOGr+fkJkD7nH7SFJDm2i/JS0u4WCjpjHWRR2kjO7iaKm67UYeTWemkE0dUP
jHq2z5DE4+e6/dLOaUnzVYNj8Da0+nUKkWiyVdZU5D9CXFJKHFhoFLhtT28RgvgY
4wacwbhesy24/HS93vNalJAyLs0NenPPNszWoQwB4WUlJa4zbRxzwqg04AxWvmmB
cN5mtdwddPK3GoJpCOoB4yJuVwj91Gv9Yj2tcU2x6j+8YKKyK+ZpZn9i2mR0Ql5d
wrbK6b+SGjOFoFgxPLbwOt2EDGkO23phMn22/DMiKRp7FzC+qruRLCroo/yIZBPS
3S+E4pZoe597hRM+n4MHqqppdE0lLybPK9GAVRJzG+uS+UKqUC9leSH/1rYVNrJF
a/unRMmnc1/yYOkIoZJ/f9HtDqaUMk1S19C3Oq5OfcWiN03ksQ5gioKLecor7AEF
I1qs2z8ZYidr7A9rfVlQIC5GcKACzClthr/Rp8g1bVGAAxmI7QitsnnJsoEFDcbj
HXPHhdQ4wCzuO4fjnD44ZdNdyW+EsaVmXEVI4Oie+xU+Cb21LIZiCWk7e5uPUw2P
aIFE4CqGUJHcnAyYC6T8RhfFtkGptozniDfpZzBDwAeT2OdoVhc7FgNCj6M+vuZc
EptWQuEe1SbXSIixWNpPjL+flbbOxVLKcjNqopcIZRXJKpd+tHyflPTDKZ0y92t8
HgPM/aPHwIjWG1WdB2qadw6DKltEsXuZQeJHxmiL16kTJXmOiSgM1DXFJjNBErRV
Pf4mxU0f/0UQnfW/OOGcBKWBeDITZOXFbYU54aZBWoUQ0tBh7hvManV9Pr8angJz
GWeQPXsX8cVVQwApnqZzySKqiOA1hL16WfR1syoXpMqzpIqono3n6m4zpZrBzqQY
Ul24T33eAMlXW/RSQqO/FCkyF8t0KJfyW9fuObPPAYFODqjR+bOUeuV28Tkz/g/P
MgA4UL7TWLdwXnjsw/tEVBcAijQbpYhVYbDgFnwHCI2540XyK/PxMig0gKEU/CW6
eOZn5tn4rikEgFc17lZBU6qKPgu4vCmi0syKhPsI6DtMy/q2r6elcnxTlhTvZh6k
gWXQSZsDmttGDLfgzaCPCYU+DcdB3D+yC6RLvBEKMxrktK+OYEs7LPcDm61rE+Fo
TekNmQX+Rm7WeinH+1CYGUltrDC6XC2hfkXaCq/bobadRjsgaS6LN82tiXrO3b4P
a3xl9ymF5Qotirwi72R0OXl04h4o5w3MdymtQhW1fCRDS+jKMpUX5SMkdbw18lHP
EWgAsnqWXmU6TCgk1o4HcQHQ01gX5h434adyE1TlBOw8QgH6R2lN162POFEuu0QO
CuuLnrJaaWOffMDIFGtUSLiNwO640RZ1WL3qTsyI+M++QC5/9unHSst6EzAy990l
j30NLUdrGtSTtFkYF6tB1Oi8FlS0ueLhdFkyCxIQgFJfuYF60FuXa3dGmUmRMJ8P
MuYVqrdeUMN0/PGILfmlCJDwqZwAokSiZeWwDP2DxPbBsF32FWUhmijCBNhZDJqv
nfhGjBTgTxwLAg/Sr4jMIxPcXHfSBd680F4yh51auM6pD6n1ddMk7LVH5MWWP+V7
5nADA3UtRrPDjZCmXIFMHMSyBLOBDfsErHDf/DX28T2TwMeyXjkpg+b8eC81CJYw
Bv8+PceCKZZNJBksiDSAgOWXLwhOv8TCbTk0TIkrQoBB4GclWTVyFrV4WZW2zVON
ZA4I5MIIRE2E9Ql+ekXaesx4sQ46JloxIcQ2dYYhOQCugdAxHGJo7mKCjKS95fjN
TRJyGqRbdx12uEkUVGVadOKmtWVESs8kBklPFCr2Wd5OOnhkFnRg8UNMFuA0k9kv
LueS6bI8SVXdyZjtKtVpPFW7CE/z23plvarmqd7PNYPYB+3d1s4ss8q7UiiKpHs4
q2O4ADBNzxhizzGrUJOLO7kauoV+fUbXdvpWh6qY+mdcuBY6J4bCAvbJ2scy5eeY
0B5cBj9LOFTHLgUd7m/0tUcf9nizd39ILwJNQlNzuhJ3ff13zt7V1A/Uvt9H2c70
c2dbjMRyEtRR+pwCv1qwfWTWO7KlsLMyMzpgjMTFvoNwlhKjX7Po33dF5clxsZx6
ZoZ8Dusvpysp7jXkmtHrwIa0Xp60TKNGGe3DWhykNFZK9K+vqHUUJ5uQp9DvdWpx
87x7HGZyHZIc6ntEO++dJfamFGYhJl+bxvRKDGeM++/2nsfg1uq1Duw6uG6j6p6t
5tM/3mB1EtJZt7jQYy8k9kyYUDL2SNZ/FI2/oBkQXfnw74Psntd/AfOO/0RlIpWO
1W/it44YmYRSQ0GXmtBSinf81UNXMUpS9FFd20GlxaRcbjxHMkf36ufBndExlZZf
Ll8dc4tiqcxgT4nc2cp8vCE8AO0jjLJUMZd8vZSnyIwSMA1bcgOJp6GMleYITQKu
F4zuE5AnO5x3s8zTGmRK7xgvXIfyL9MKBbZsi8vfOtw5yaYKY+0G48/iFYf/XrmG
lkVueGslxlYCsFKVokge63wqzQQJD0vVjolaFbg/GxOBCBjKUPEUVckBoQrdDDi/
Q8tF9RnqISkzdvDvqg4WhcwyayT85LRbMTtz2UtcKcICY7IAyR/jQGUNBAeApuyL
t/1to9vYgsRvmBOJdJjDEs4QZ8t9IPJS+ouhlIEE9Ol5zgqQN5yy3x2O2omXE1aK
fLRFHY3NABp3JZpdQ1irq/cwyYafAx7XfCp7NBQwVP4h/zAe1bG5jvwzJtJlDtFb
Htp0ouKQiUm7XWlMRF54vIyFQIfvSuFJP/DqvZWJEmbEXT+uxpXuWZn3AywS+SC1
2SKplZdZ5Whvn9dXpMMmXWo6QfR3yRtfHpBEbSDD4cCtsb6FQWHj3pMMFS9fiz3l
E62gdlw0mGlTfLWAcbTKRdVwINOehthHX6D+c4UvoTOdmoRD74I8RQw1UyBWkX4u
zEB0P0fJjn2kmk0yCpC+qfTQxRMmHCWM/KnAi8Z0Jr++CFM71C4cf2OcEHF1J64s
/d2OVUruqOk7A7kj2IiWWEvNPx4EX3/+A09I9UpCiDJzTyY+XjFTt6NQt1NxwAc/
LfPh7lIq89z9o0jD9MtyjcT+L++fcouK+U0d+G+kA6m+H3Qfh3trvBDD0w/OUmsI
DHOqZKFoWiiH10CEAGxWRfq8e9K1f3u0/KcG/okhwik6CijsjRp4j1jHiJD2ehwq
9dCT3Eza2unGnnCxBqbq7BMd7JI9fQJ7tUFBBgTjncgdHdHVZ3nw4tpleot20Wvt
vI46L12q1k+nOYziTGRwy7uX0wnL4yiTYV9wrJUlMGIO2CrjUmCEwi+SXVGqMJBB
OEjTcvx0oNNaH/mOFV54I7WlASvyz2ICcnBWRRRQtrpfGqUA8DpJEtYbthEdALDz
uN200Lq9DYV4LadPUcWBV9yE6n5q1wi8y8wmRnwyf+h9bjIVAJ+0X7Ipq41y7qEd
yJC2J1a48r8i9BVKgFCc6fdJWelLgEjVN5wBswHAgNTrWOaj9/q0Q9Aer8KMS73M
yySAJZbfSTRf4za7efsZeKtTRb9JNLfNi9arwGYY4NognlIzqd6AFnlHLG7dv0oN
BHcn+W5dUlYn3PoCu87CwKzB/M/wIfWUiBK0MksdoTNKmYUBs8yN14P1oeqSfzwV
okbytoIxTXHI2QcNrDP5KT5ue2vdWLZvk6rKX3yLnnW8Cu+iobF0nRfY/MlDPHzr
fwShK/j5dYFjzqliNjXzs6KkqyJm3Yv+S6twsl0tQwcvguN3d1UEVUIsoNbFITSd
syOokfqL9+UoNs9k1T/eyX7B2hl5aoaDfVZuyPgWp1zUcrNGEAXW4SIaFu3rqUSt
eGfhMVFp1rfR+antBMQp7WEooFPBuKGOXiXi3clvlJ6tA9+M5fBcbwVOwRYqg9Vf
CNBt/SdKTftH3QCr4pQcj/lrfclC5lVjX53Wc+lvSZ7t+e8JttBtx/e3ArESbiVB
dA5z2OPZ6wcyhju07ofDVSWCdOd5o51NHHtErMuobMNt3fj7pdY/0ieAtcEso1Gz
jeMXhqWiFvyBX316c+zGbN9YXhzaobs7InsU1vjBogqdiidASTLTGLr9NN8kRcoy
UygHWIBB1nL3hHlOBafENh2Dp9Qw/0197tfreR0WR/FAWwVqf+FPX+tq2yUZgo9u
OmstNGpiuvuA6Y6guirPyryaC7Ck5V8/Py8G091IyKhGPAU36JkgizhRwE+EKt8k
yairm2b/WpkozANkHYilCpXSM2ceLpSoFsTp8dx2ReOaFVyAZcaC+i4iRpP+Uzir
NbsV/hEQLTg90U1TQXwzQtbdrYjlW1pNpGKlHLTN32+cgjXHuVitfIyGRLz7mn+R
BYqC8Mtf1A2Mm6cgOTX8pvfyxJyBk7FCQLK8L/licwhTQa/rAyW02M0RRxTsDWOv
L4ygxHKlDnjh/PKxKOf+/GN4rVS4oUMCL/g8pzipTkI5ziuyupBg8PhD69lt6cRW
WNqYLe0candiTTKkJik5tLfSJMlLYIUodeZCUKnvD2ZXzWCFWSduRFOeArdOE5dx
fJVVhKQOAiBJQSjhNQY8ndhGqJar11VCZZDIoAjYJZFdYSlrA3UtCJZ06G2zm0uY
Upe2yScTeVo2hObhQTnu8sEghddD/JIK5JXlQVfVGgN8HNWdxe7kyLAWUYdcr3P4
UL2gL3+d2EAXD+Ps6phSGAgV6DuRHOKuwBux1b4AM0iqEaAEhBll85Ok+q20WKXs
zhzvjmXDwavKpA/R7qWPwbkk+GOEtEOCYIjLwJhbbiXPUSaTPNjNGAoaY+ZJPJLP
FV7N9kvH9eIlz8uD21aTqOMvO8nZv3+roy30tp1ihEeVEbBaFRIOEh3mXxl/aZIs
70gsYinJGfkmqQQ77+48jq1DBGcwB+v7ctQ71Imz/HZ7U/CPkp0wJ141PDp+Jde2
sq8zHKPtYks1RR+Xc1vQg/9UYaX0VKSLLT72OqTLsfVGx4241XC1hMq2HMNKbyzo
HjofVmZm/qHiIFoh14IjG1/aNRDSICGWJKJkye2BKKcsKovr5hoT+3NRZQB/mb90
ZPSZWwaXBkwkI0Tk9wDZqDd2n41px2krGpzmi/OKOhO/Fz08cCy3S2HfnJeXFifk
Ar4tDBhktARPMtmrqyzrZrv0+WldIt5pzy7vdpqlLvd7SZMTv6SA5YsrBgSNgscP
rLxBd+3g/giaJj4dVC0j9/3aEHzbYsSr6Wp2zjMZEtazxbF1+/qajHaHbSf26Y+A
sT8KubrfqKvg4IdB7K8mu8W+N0BFr1lU5Ruw4uZeQ0DCb4ktvAKkd/ggwSrBlLsc
1EO44pNkhYS2quEbJKmePQfvNAxV3M4mtMIfRlNCEvP2FQ+yC3vEfmI8NKSOPTTH
BWjgg9yeppcqJn4JpBtkNWI3ucY7a3iLcSOTJBtoHi9EYXIb/nm1yaGxUXH0iseO
yNTrTg7HHIyN8jokgkmbnkAj2RSoEK70bYu5I18uZ5BFSKeFSvLx7Dm9A9CSHBQK
pcSuJ3j8lAq+h0QgrKbOwUrRN7I3ehpLFx5dhqHqGT17vZY5dz6xemUGxs1Rk0aM
UKBQgYvlWJm78w2xTdxMIxhtHURqGmX5LMxX1ucEW/JyIJYT3ZOlf/WYVhcX+Zq2
tG9U3fsXfI69z4ZRUKkFo01xHqdduUaFigMu/Rj7XTl/z4PSOgsUrTMMkz99czWY
zp4ScnXltaZKT+vMfoJy46GJBxdxcdyxZEKWe9vcZ56eVWCvns5eadXFQ6ZmduOZ
p2N3aMABQqEzaKQZH8VW4fRzHH8U1ILVM1wdEye7OuS9GLOm6PcfxQ8dPZwEOt/w
SDh7qBlLbgenb+aaLF01E68A92y9xp/ZTaGB+5K5L4ej4/8SeCYDY4bd9n8Fr7LE
dm7qDibEk9YWeoI76Pn9ODDupEJg+pp2pUJbV6h1l2Ml8cR9QFTfv2mba6Js3Kl4
vp/8OG6RpPa3D5CQgoojNJ6ShqzD2GVN9E6U96PXRrOyJUyGGvp2vW5WyYzXq7t+
5rd/rKRRnEUtX0+NvkB3LGngIgWyri62vlLQRY4kMLJDiOYIEVrWPlI6kyu2mDVC
OWsjxf+VkfOnEGGx4Tu4gn5gxSP4y5WNSo77xOzEcY2evP8UC9AeRqJBzlR8BudH
P+HBYTBI/vl3hTKL+tnMDqaGcWvWwM1kdSEebwPbKHtjvV/vGEBAfv1DTbx9BsRX
d4hGRl/HFvkDqNlGPDUvzo6lWIXBrlMKpr/t+MW9uMl1+bCThFdGY4zgxxa8yxVS
baf6fyYG+hi5beMzjtLIuP2CLyj3AbS9jIKJDxrz8ooEERHA4wLKx7iS2nci7NKf
9rh1RgV6XUps8vU4odRiN637h0tqNbMU4NHrpaBC5R6+8Bp0KfwdEsvNDlR8qvsP
SIm2oVNczQ/VtHCDWrEPCYkP0uwW+PWcJcuPBoBWAVUZ4ow5pSFyrYPvwRpf2KG2
dBm80JK2abEaoh/j/wbjRCMJeS4tkh9Eny+odFMqNLAOpuToovE6rB9D8ppOqihj
tbXQ0viyY1+7vB+T2ubGCLazaMNMq6LtHAG+lXB3SP5tVGz8NWkol0Qau4pUg23L
QYwEqnN5Cd2HkvN1omHYzUIRUb42edaZwbNMlLvgGciD8z8gq0+P5kfEgAF8Usby
M4Xxm4pWIkUN+TtTheQ9ITNF56YFWiELtJ+XBVcsJB7aTBoVtHJc3P7FFInNo1Xi
nZ9acfNTguE8SvQ3lAw5BbXDTHUxMIww/5fjOLtMlCxxcmpHe6VTDePS/o46NYwJ
vx5uKm5RRoEkbp/TlPPd5hBceUJstFv69kvamkGuHHMBpdGAnJOlTZcbvbX/Vq56
QnapuqbGK5L6puBfSG5XhcNigvNRR0vTyacZ8FAx2hJZFHQyL0Nsin5ADatN2GYI
hy8eHwGnLNIadK2APgms+WOCuY6Edc3dtihup/TjmyypF+GREtCO+Nogcr+10dCk
47Fey/nY6N+UaPi4Tuk9zo+vrS/nYVjs230Ziu++Cd2IxoTD2MA0s1AZZusL9PBx
5ktyMWaY5ZYMvSz0goTMCp/MOYH1wh+jraEMIQMdyu7xGCH1k30o4wHW8xMbj6wU
orEwFZEHc0ZAJ/amfpoxef/y/7bUsg+hzyckycP0K6fqwi3RKVex5WCGlYMjWhi/
Ofv5ak8M0ZUHS0hTE4qO1wEHEqlIgDF2/2PeRvbrv9YYImkKSqZauAB00MIPeTpX
ac0txrSjMXUF9yPrGkC0rM9PPsOX1LoLNtxYBqCcdcjpSNZoHETMuPK8Lg/09psH
M6+R3THoveZZqGB3Qoa4tGYwFJNE6TG8uexE3WoNSELaPDmJOtoMRR9CoXah2uwf
NN45Of52GWopq4CJXMWInsL1n7Jo962OBCao7rFPNtD3+ttI4K6Lpt9y1JoICWd8
yilax+UTjJhBdb7ja0qW+zseC1GibfORkqqMT2LE/qaSCxm2F5qCruipJWxPigAT
pxSZngaJGWHz4c2qdKETtdz/IeoUGu0athnj4gtRctyLfRMKLl/ey9Rr//cttmm/
pMt5+jqaPf+4D+4HSD36ZyJXSqpX0WUDrs35apjXc4dm0rqQr61wqiaDw790OnyV
ezh4CpB4so3qRXaE+C3i3UJXK+aabeADEoCMOX8xJqPd6IdpDf0KKagAG4hWsog5
UNJwXaBbaUJIOpjCIHVRK3AcpLf/KPuY1a2EvFf9q+1OliCt0ZtQkf++6I7gA9Ns
Dyuum7bu7pR1M/v8yu61oshZVdBcAJgaAzI4erfgZivNUQpNDihj13AcXUUfBJyI
/YmsvbZM0P+FMC6d+8bm7Ev0redxyMLhMafQm5zU5Unk53DMnNIVlc2uzJKEEKTK
g/ahhqmuoOB4vQf9uCR8X6ILghUO+Q+V+KKq7+NuqR/d+q3njTNdkJftfK5KdZFT
xnfap1m/gBK9hnk8RPAH07QvBc+vXxsy2T8NMSi6CcCQTJ4UOShbzaX1HMwX63bt
WY0+UJKuiqSEW/k2utnFA6+ZZfpWDRmYLLj5RNFJV0PL5JAbrpp/rY0EPsNQVs3P
EI7Uxn0E6xo5PXOdOF8A6BUp5T/VfaaT6y2WixyS3lm4yLysuWZsi2PDsW4+Ibq8
bmJHXvLc4bAStKg7D1Wlz6gXLp8UZNWFnpZYGX0RnSSEMjGtoFOlTAWLDUr33Jd+
hkSZFTfF8bYuYhm0/iLXVilNAIvAJBiIhsn9WL02HgQZt6KDIjfm/o7O5ClMUP+f
8+OAB93X2oG2RujuXMy9AYgRmgvrGSu9arp7MoV2fVbcqUJrvV9Z3uu9z3IKgKJ5
e5Rjjd/vymid6H7xR3FYtIPnpxkUKBGMm7EgOVQ7SspM5bQo4mKVFktYKaIjLh3I
eqe1KNkRd6mcmWpNwdZhBJzDsNhah0FPWIK0ClhlGR2sfzhkvYztEL2W6CRzBIKQ
q4kj9U0tVyD3ATCqHO9kwp7n0Vmyo6sXeKrSCTcM2F7CqKTq+gmQL6LjO+UySj1k
vd4t4FzStsAD6d4+MsYs/XXZo1wJx3mjxDsgOeQXsIuJsbc5OTWdF0J23KvLqP98
9NrKZryvtoWzZ9nDbjIDuA/c6aYpqLjqSb4aZEg0qzlMJxxUfSn3tFhprhFmK4Lo
bPBoGvL7wlWTR41w0hGyV055verZAIURKYea0gJLCE9gYk6Dhm+b9Be6aAbwpWGF
WEzfb7snHrUiSocXbDQfvkmU+z87oBnJRy5P3oaAxWKDkEaZM1HH+Zwttr1nLY5u
vXQYyHdQiEKrUHc9ni6lLmiJ6aImIeWMvWxlvCE00nBGMg1cNA/sUPkNmN9R1rWS
uYd2eZ9Z8ftskglXkOGR4Vn5A+0yupcPprEE4IwnfapFBmPDdSj6/XqngEdjT80D
8QfV9qeBcshdYplmB5+oyuq/jBajAIrweY5mCzIsGxEkF1lAGj8z/qerz2swoHi0
6+8pDnD8IlgNhhMtgN5QqIBNZbbMgFc3FzXOls2/RZ2tFgeh5awQmQI6R+jKjmx4
50mfKkzjQSYBXg43132AinWxqxh2ccqtD5B8Qam9qTJ7vS5kylTCnBC83mdUzoKd
yWk6OHIR4csREZO7Kd/ATUKYcXgQx6Fuq+ZGWQfQXQ85wcZFO0nr6PNZzqHFAV37
MO36cqt+NzoR81U6NfuqmY2xLCU1tEJi3XXVkVZJKkSu4meF4tLmtCnk1d1Dbh55
5ybU92RqabAksMfIoQnTnGP2FTZamY7J2BB3GI82aH79AdLBczQVuC6gYyJzVlDZ
tKpijmACwr3r2lZgFnEAEfhRcOp0w0o++fGn0NzPO+y37in2xHb+lruhrXKDYfLy
rBAPXveGB2LT1uC6XxhjhM/m2jfO/XQoEQq/DgLnd9fqCLSa+7NFx7W7qRslpVXx
bI1hC47oVgecf9IQroYkqgmiAzmiMlyxG2KmHEs4r5DgiyT2rtUR4K87pyeMUV0A
P3T7sbTAJetBAztV/0PllSXtQfb9S6oLtEHAOK4XMRShVe9GZKEyXL2rZbFzIPKs
KjwuJKWmX+gq7XLdkc0M4AwlmYjI/6HMSQv9GdeMW+OeMB/5jYI9jcRqG8o537gJ
k5wNS10g+dZbCx+qmqOKdRwWfB3Sn6cLFVHxsVFNv4lLVA4FWZXo/wkD6ritjeYx
N9TsDcW5DFxUWg46nqHxjL/GlPWPTkPl8GryQGhyjNKdmSrRGFc0CTQ+u9IP6Q6p
YciFWvqOsonJiysI2wh7/Orl6ktwz9Q1nKh+TBLFn0Mcl/Ream2K2qz2rW3SoUoG
6Q/a5fPtJMhMut9h/7nNxmWtDIH1/gA0kgjalM6dgepihOmRBn5wUoz9KC1rAj9N
q5a+pS4KjpGVHvQQCdC1r25D0U7z4ARLwIxFza9eYFtp0+Ap27pIYSuIcCFaahs+
30PFHjepAqkAyzngJtynEyRKo2b24SHyaZOsOf2tnSuww+/q/KLWBaPXonnCGDnW
QWiUGUKhL67/c8kp9E01u/IhrKyhwXHvYLO2Iv5Zq2N1YXBV+CUMOnkYZ2s6GoRh
lrROx/llvO1gODl5Y+MdllS8y9lNa61C2C2vfLlW9LkhyY259eVPeOjb6OvEUrsO
cV/R5ehel8+yKHrSCqO20P4gxrrwBFmAa3OkXDfpTPvRQiRVGVCVAdzJCxnLHqsu
4I+hujXH3qXdlcdI4/9yp/BqvZW90CXSyRKorRD5xC50P7cFGwSrhZixcMf8kxH8
a+7BP8q1uOn64pE2OSwbs6ZcupmPxM5D3hdi6bQLz7v0h2qkItgoBk3rD8Un5acf
U1O770TKAGU26Q/iEyQ2zbPUuPmrUSEJrYkrwOZ5f+AcRqf3tvPXqK9Uja3xsU86
4u+hzCqjFkmXuXYKut/M2f0GH0KKgWJoVCPwmRAiDnm5/LR9N2Ionf9LDfBK1Im0
xVTvi/KRDfnDzsyLJrQb2Usz1SDojRMQz6PB7sx9xrejDm68a3Otz44obUAA0a7p
MUAIBPgPp8SmwtNSj7K+/vUXdyVT4mK5HGM4nbov0U0e1kgHlqI9Rr8qhVuOMwAN
gWD6ErnDYePxL5q2+hBBokIaKHl4L7gFMaCSCbN/hgAR5kT1ki9h71mE3zWsMeXU
kvePwYgXpmOUmJnG0WOWUOAxFr6auZTBlNjmVgYrXsctZgHzQLwsyVm5gtlWfvL+
WpL+NZWBgBKMOihXkbeekSmsUpzYm38ghfSLBo5wjeySgor+xmalOZqrOQ+edUiN
VdEPCoyyQPH1Ztn4MPsxTgeUKxm0JaAAF+VQSXFjRsL17mwUeZeKYTbvPlQnitJh
ljNjCNEX00l/vaMr4/bM1rrEoCSmfm/R6OvAoMTk93NoeocAqgh3ovLEdL89nqs/
oSRkSChZ/WsMlt6ih3N1HG7wpiXu1vMIyaZfwzAM2QXuRNoGI021SPRMtUgHuos4
qm6WiCzJGvU7eSsn1EE6ySqyDV1I6NyzWnIiaoN57ae2FfPuC2vqJQjZiEcwzP6E
u1TPoj+qWWFfAJht7W70Cn7nxa/TosrNPbYPmgWgRwm08+9Kx++kdbEMxZILEfXY
9PE62MtPfzBuakJSHbbiWDcErYAl/YenspTpsoOfP9GtE7ijPE1v5qEiNmpJScQL
aq5NH14hSsHd5Jptk/00iDJvNwSoP1VWFRpc7Zjpys57p3ZLykymhBUJyGAtO3jM
x1x4WWwKJRoDqMGHKzepnja8FQJzJeKRkC/cCaOtbq2WyqP4pnP/WWQN1GuUWBEc
YAijK91jlR9nIEZXrACOoiED/1uq5qU5BeohzUnSNy5Kf+yCrTT7nXO+kWtLWPfS
gG1Bcff0dlgn5pyM0HInvG++DLBdV/zm2gquEWmiSgFKS7d9bi+tHNgr2Mp/7Suh
AhWBn7dGjCDtFY/u00abz/xVashyP94Oi4hssCASkwNIaYdxTqeBlNSOkANhvfOP
N1Dp1zoSaSAlM8WW9pd5qL5vMoZ4wR57XVqYvA2UEsHTIdOiQgGLP+1skM5FeU/u
UB4kfilGPveFURxGELZeJLSvhZbIvKJ4aexoPE+uIHAZNCyyQ9RX+PUTZe/tUp9y
ioNntiBmP53qciY30Paec344vKIVqOp89YW0xAn293guNxaUcDUfdcU+adf/VWhw
jLO3Dpwn61IQG/DTFMHN1IltzD4qkz30p7QGUJNwu7uXwgmNmX72iAricJWl8upM
/6FnXUq8Z5ByuZXh4RdGzRjNDGYnA5uZzCBNXkSa/XpPmSgsxpY/nRQdBZBqporn
HFlj9N4fQqVKbOz0vD/N9ksEnpzOoXkWwhzFukIcoO4IxojxzLIvDYAxCagPv5cU
bcDQHr3qdX2kJ5nF3M6GJZRKrH9YJrV+WNuKrn3q3ZTR11g2B0tJ4tGRFclOKCzz
QT7983jnoOXyUuyuL1M+IEs8kAvhyQVCySB7BqTHhR1XVIpZlGXnY8YBv9Vvm31o
wL+eEce0YqkAHt0lQfB5+gZrTP834r5UavKFbbnb89l3781ngFCg4AcQ87QTg0kU
Rj0NUldkUigneZfSgDiV7U5B/9g2VdTdF3tFG4yOn3k2T/pTD3NSf0t6uzBaWtws
/ib/8ZRU2LmFuR8uPB1i7RVONo1a3k458PZMUk58qvcNeMu7LEKEiUwexD0EK2rP
aywVVPcDAJws+eZvHYGM1CgmgfILl22ebff++Nhhst/5o23xXfGiR4Ao+ZPkGNws
PZGQLbo4iRSzoAp+iVR0h0BOsf5YwaablcSnhYY+vfwRmaTwxZa9IU+9sb4NxpHc
ZIqXYbEp7zIY9PI902I5zi9FPjhVfJF/DL2W4Ll+b/MuuygE+29rEs6AizNiLUGh
7FWjI07ZfF5nlGiCrqExwwrRd2EwoDzvnR/AyfmXvv5HDr/6hgrED2c99x2tqJsK
k5yHfHVC95cOaPQGE8/R3VSA6KM8jQ+70vuji2LpSXDuDvmkmPNAi2Eh9ZgBKs1J
VK7vBjKDMJXmRZl+YiM6ZnDbw7BXgShzAyac/NvPytU5m0AJ0Kj1BIa8XLReECmm
rSTLyCqEW5h1qbOFDeBkTLh0dpHiyQwX6tBLMPx2qViQ5VjnzfvHOzzw4SqYvLpI
0uHLvPP8Q2NqBeAEM4CtPJV2icDsxB5sZ/rzPerLXqt0JcklKIAZExshoBP8OQwT
3QMTdRgtvI3SAkE/9E2Yg4DKm398WbIrzemtrMJl8OyPr9U9bZ1ytmrw4lJKrZSf
mzSbmwt8qFi4LWFiZ1CVxXlnsSWtDRDQHQxm4wIJEGY6WuUkE4ZsrvXt09VKwq8M
/DdCtwgF6O2LMQKxGZmGDsiZ54/9Mc/WJTwYx4zSw3kxM/jAok7GyCuKb4ewd+Hc
GNNieKz58iQ9n120Sm/PgY7o7doFzsPOoPS0TEnCjcKp8ctgc926WIMEMA42lYCM
xOGmFuryFSWYkMAgHafE9Zo98k1whLE9vaSB1vrFEtD94wrnZp1e0gAGiKOA9UAO
YZUD6+trRxtgJYnZ5l6xwgGzEJ2bX3zgbQeaaMfGUQ9xPcas7OMegltFWOw6ahBi
1DbgHzke3Zrn8miQuAwMBVm4v1GafljKMq8clPFHoCJI2XYJM/4I9Z55DjVt7j7A
S4D/6/tsFRq/q4gp/HhdsPIyGWxkOHI+j6sJ6LeKDEPMX7spdr6lrMze9+P7/kOC
BD417uNJ6SrudG8dRHJTUM3zmgKeB1KyWb6hxuIeW/U3+5YdZcr5u2A14CpokQiv
mYVz2CwE+pvA5GTWqaqpACLEoty+nwxMdGLW7oykXDXUZXNCAlbr8okKyIfBRNcv
xNn2EPzStxfKhsNQFI7FSGi/RaXPwuCMymL4DkSJaRWjyHhT0vjAWCpuGPaZUUT2
NjGAoBgOsYBcpTPhD7dVcjKCumovMi5XQOwp6l4CL7XIu5bu+Ho3YTpFBDl+PrpI
uxgIfUntsErebVHJGWcRnLGEv/chaSB0E8eNNkrWrhOhV4HtKoMU/nwmwbzPodY0
xE6Jn2ZicdnCuBxF3C67T4B5dYNJNb5r55AjTEY38N6ldFiqd8BlGAjaj6ET/+Xa
LocrYAUL/LnRjQOmHf+bVerUynVgLvaqfOVcy7EjKCPRdh+e+VzVKauynBXo5h70
IqOKLH4eHZ33O2Os2tb5OOGOLE8t315geONAI01CtVJyU00XBk1AUcbzYR7wIcoo
bmuZQMUsBJw8M0zOl82Rx61qdE9JwUDXjTxIIBFECGT83FrDQrIQmcqnDOOycawq
i+VCECcq3fw+OuSeGwI5kNDI/QYkMr9Sdk04qW6eFCQSY5hY03u/7OLoAeJVixTi
KCoIYr16VuxG7GaNkJ2wbjzlLWqExZN+KuDiEqPAFBQF0yrHP3+dAtiQd59WcUSu
uFQHfJXHqfwYangYiwyXP04qS7F+XftVzFSlB3tMObbFQI4xWPwxxfRtzaEz4b2h
aUDgk4680VBS8CQjqdnuVx9d5xHoRT6kAbpPJhnz7LGWkuNgtTqm5/4ZdZTVlsWx
jzy0u7NzYW/nRCRm1m0LOVaHga8qudN3p+u50i9XJxgb72LJV3EeHgRdpckyQcAL
a6xJpj9md33nc+Ju3U/boXYnTi6JLHbvTsTDrx8szn0Ojz5LQPqmJkRZtsfaSZj7
eXk95Niar8Rn4R+wcUncSyU3EUfqWG43SLWcWCUlCBr2KUTgvd+uCqAs5Okrv9X0
kgRPi1H/p7Pl+yfq+hB5wSjuPzUGuaLrWE0BEsyCNZBHhEdhRrYVj62cCTS5yF7e
LOcFMmYttIY7jsTFu1zryxUjjy4VNkZ2wpwIXsGofIqJbPlgP63MQWjfxiiWNjfs
Fn2/khTWTCiD4Nx0sDk7vacccyXq3Mi3GGT9/KWSiR6YE19YI7AogN1kAQi8uOoV
jMthgvRGT9AigjvX24waRni4lczuQ+DgQHxWg3jF7keD7S0nXADw7k8n9NFbDQ5A
gBudm8l8wNKMRhVDL/snt9URex/Wxo+FxcQ/JgG7Xtj7LyY7+Ya5hkqpzXdeyPyg
hWl1gbVWnHWjWpz5vC43ZEzEsuOxl/BggfYXDfvE+6rgoE0rJPI1nNgivJIIMVvF
DCtP8SLRepyBske9PuPJFH0NYC8OJPTzCeRFeGu295I40oeN0ZxT0FIvNEI11b3k
Gfu6yVZyYW9/C/LCuXAoDeMvc7/saukFoX1WrbZfwqFrtAQhus3oaEo6RQrNuhMA
NKxm/GTdOKFdk/8cvIzmf/LDagp63LrcgSG+csJjKGmJqUecGEbuMWOWC4QanjqD
kLwGXy2I9Htgbb2cGhPbmTsf7jNlPNnVUa61q+n5/SHoXOccHih17RMYw9e706AO
lrVDN5rL/jBtKj8Ej7Nbkg2Dr4bmRiz9yavcP1yiZndexp22uGpYATFrrBCysVhA
YERKjVFBAnXjvVYCFEpAWxuQaYlE2JDxuYg9IuRjOL6cVuCCvryN7XAWU/ATCG14
21DfcQ/WkS6vDmtl8XeqbkAvv8Bn2VNxRS8rSaAySdlQTFSfc/z93spqzncM6iPa
Ss/NO22N1mDwBucMr/K67D+gVVv3kJB8U4LF/22TBv0X16cVoIYOKXYlr+O8QiyC
wI2bylmhG/SftrP9ytXbH25J9BbcF52bzsPvKeB/HhRhnXKbhwrnexq+tH51nAhc
Xxl5C3NHxtlvvkUw9WXz5iWPGqY1R6Qz5nZNRuU6nE8X3Z1kGAHPXFGxzLRvRNH9
BWuI/pGGcvOJCp3rLc2k3+e9y0aStZBt0nL6rBoAqe5fGWrRLkhtXQx1dVKoqHo2
dLYWrwTfbwCgmU3Aimz4k660TM7Hf3eKZEREyBpC81GOBys9QLSnKnLKsihJYxWH
IjF9Vn32/MAmzgHKsatL69YserrIYtZAgn2/Wy0wVhIuFHWtl1wB4uXS0t1mR0Iq
/hu6K/Etm2gN8epGHoJlkdVuvwnLakMn+XWX2yiVjADMGcfXlB92oBP4rawPnRYM
cVzvmy+rj3HjeSekKinilFRshpOSEXI/Q+/h9HsPpCzLGzeZ2d7xKCEm3GvJjZ0H
GErwUqGHI06yAuZ6bar65H1tKj3cbSYlJTurrxwWX28AWVdy318OHUiRJcViDUxl
69IYLOOwelorB5TWvmuTjd/m7HP/nabn4cAsfnz7+TrXrDZhsJNOHWC4zn9kZUpa
9n9S/16h57Syh2WgxS7fusH0Yf0wVgjQ/sbDoL0MG/t9NfN+MEwcHZAI680ewVJ6
LTdQCIwRC4WMpb8BQ15YFNXompUo3p2bF95L4X/comEhqEctdX6A15x7T0bQbGLF
XopjAKSslR/lcIcIiSKGDGaMA7SPn0uyxLJ+eNRGNqA4v1EShqKMasGVm+D4HAMl
26RPV5lU+xWfGQG7hYDxVNFAbxaJyQhqN/e1DIWGhjGok9pA/oqJEHZnDuKNff/O
mf3lgjtkZJU2qwoOJvMkCib51pg3D+Uh6kbp6oEVLrnJhUNOlmrZzPGc/nGCa+zh
GgVNnzs7MxBSMGtftzv0DnoaaleKFO41JfU1zVCsjGKqTh7XAUL9Eve+MKlZXU9s
vzY2tgA3fAiLHVCNTmbBdzqNIcvfWQGpJHvWCGJG92ViScGymNOdb9AhMS69424N
vdpGgOB8sWxWX1Q+S4mYrh1cGBfWpbjTysycUpMH1FFIZDESMSQTdhK1DyHl8P6j
Ql+rGgH50ysg8v04Vz0D+IDGwjkAIhzSY9PySxeDxzxcv6HaLdEuFxpkMm35+3KQ
j5TCTFWYfrnUjmyq6b0IKNesQn7Sl47rijEf90gxSHnmNJj+O7zbOSwDUYZo85Ta
yA38SkLORSd92T+XKgo0T3fof7W1t2PkzEJ6N4oKuXdZw5CSOMQsGjtJF63hA8O+
R7xHB0hrJIT1U0e+0YaZRejyKbpxPBaYv8kEQm7E0yyUCU0SOn9wZEpNWpIGvT+c
Gc3TrDkmXQYO5/6/9LZL0JLh643eKkuTYdsrpqUhBqOXWTysBRMYj/NrguUy4ABe
c+L/T1u6NAMYywrQwVtpurzLXw9ko3I4ITl2UzbvXDC5oRjwTO3DzHmwANSPhBAy
E90+oKjFKDDMsdW9zzuu/Fg1FVpArReWcI6UieVm0U9sc9yfRMivm0RBJnupRU2U
bXMlftDRfaVOGTQWVBGP2UjByz7DoBKNYa/QOiiI4tnR5KQG+FH8kdGwHAFAZ1DJ
sfEFdOb08HFGT1dgINh6owv7ZjZhJt9YPTtEqYshODCBDJcs9OpFwcCRouWToVZe
v8ph3xN6FR1FBXa8Hefa5z3w+AC8PjD+4cwd9tCOLM67+H9yGgwNVxZrMevBRhJ6
JNNIMIgLRaQa0Q010+e2CAMwExx2OtPyAw+N3SPOVwNr+VTP88ZjMe7DlzKOEtqg
Zx19oxN3MQuLNxPszWbzFIKBbfbSYm3CL7Kldq87IYmXapG4ETLhg/VefLk9dGR0
zjEUwXgOKOzLrBdutyxaP/tAJ4P6d9QfMHoHv9PRadu+HUuOYMrBpK0PlcA+XOL1
xlF99gmsM/oEwitC/34IGdFJZbtTCD2mUEckmPjaXTsKAClA3a/xYHLlTzWItGEi
gqATzLFTJ9bqrwPPLGhGjXiRv86NYCNx2Owbjh8ayAW6FZvOJ6Qxlz5u1rVVKb+H
/hVsBwSKwkJ4PI0SEdRIMLn8JxQtjD8HMW1ty5+z/Q96sXvyrJ02BGsBux0U+8LI
pqTscxu1YH9EnXPRA1Zi0N+YtqKtrSRGxCt4wGzveEpvVXjU4gef59IeDx+FRxZn
/xaJkPj50ki0lUqhWP3Akty23fjfk1vNGGlrX8VJj4wKBEOFTY7mEkz3wLbjIohj
8T+yZYNH7bBbQ6jCKaM8FPm4moKgmMv9KysSgvPi2mdcDTldzbISZXGDcL62BR/v
53pRZcAcoOFhm37JMFD3JJLZSh91cayhkZnX5j7c6Bg0GHBnji7bOQQsYbTDsDMP
M3suMfag/iaDGDj/rVgSegmVHrVll/dxTFerKBoZQOk1EeINUzKhCj1YinY/5SgU
yLGeUuIuVPABKkKQvzSjntylFhRlZHWgSIYo57wQzqP03g/YIFE+/TdwvyOyNWLi
4BeHrloSDRtHPnMndk3WquHrT/dtrymVfN4fsWfbZUPiKTKrOLQ2WG/44wTAcvfH
Y3qxRbSX0630ywCLD4FU3u4rT5RvUdkYclfACDiR53xR9on7zAGZhfQQVyWw8Nmt
AQybrw8n46B6kWDPkeLdGjwrnDe9ALsVCgNSC9yxvDoTJlSqKxoBNKJjfzFGDLnS
lawcIhY0VSafe/pbzm7oFXjfGJ3fFmgfpm67NojN7+1EXGvZ/uVw5C3lGDRSpp2G
KMOF7ZHuRvxaW6+qWQw54j6Zx1EllCMIJQPzcD0FjZN3fkm/1otwTO1h1SJIis8h
hEaVfcEvlD1E3T6rFCw/iL1BIl5Mo9WJmaax9CAJ4ImbUdqzpIXkiQnNaCPejb59
iGM276Wo4RhKb+guRuUVnptITVgZJA15U6ZDw+2Guei2VFLeAt6ovCJ6KyICGr2J
LGWJ9lORYFTkJJ+oOlOrMsa+ZdJ+vjbfonI+rKmfv4fzfeNH7jjUTWhGqq51XHY0
NmHzJ5qwCPOd/eoL29VqhKu7zpE0sK9V+nvfKfjg4O1iZ+RF4fjkmEwc5GdxK3Vz
5bbRugjRG3qg7ZmFX/8exW9MxXLMFkLT5GB3WeFjEBAWynITNep03pkvWYM9r7GU
uyM1/EqOO3YRfXH4oFrX/j2wem2+WmhjS1a/1ifaQe3dmRFzj1kcjonJdRhvXhLK
sDQeHuvNa9JV5iOZGOfwKOs8WKR+P4d0FI/r+72SnLVI4WJQLBFMNbc2G+z82Mdf
qrhz0mve7do5anbfvuzsLlsQnaE7BuFrrwDOa6XS7IuH0t0Sr8HiaefVxG7TyKd6
yClLeL+4nL6JYQ3vX9w3G6uxc7pXpMoFjlwgAjUYFXZNtdwUYGCTeDWVOMaeHJRj
n2Ji8G5Ix99Eg472xQ7VghlFF5rrryCYhanW2oqw5Zy7ixjWX7i/xWtTmEuHdjyf
T/HmSbSmfc7lRZPz8nBtO0V2HFOl4j61t5EpEAyNhZ1nCQBYbZi3pP1FfxKBJ/F7
sDZEZYIN37v91bcLPmVnI2zaAKrD6oym0AdBCugVhY8Xcvul9gB6ZV+HloQbpMl8
s9eR6PRpM9T0viOAym8sHCuLJ1aU51cWK8SrVLZ7XZWp/YapN1130lVeexDhuv3v
dBKXNnx2/tXOovdCn/WMZPn+EPh2lWWJShjMtwreB56t/uN8OACM3gqo/GzyICEZ
plUOV9gEPsHRyH18FLBIeiQOabew571p+ev7k7dH9BG1Qlc/6G1TFazzCHq2L9sI
bMq8QqhRR3Y5t7PpvMdvLKKUAOIup6IklsDYEA7hltNKdDrVAQGmMH3FhuJ+1A/l
sphjO0VaxLU8INzS/w7SMynQLC5Ryr+dVFAvqWPi6vRYlTdyzkD7vYdw275AheMv
hPycMFrJkdjAnGTGTOSniJ3jO+Fp9wQhcOBs6sn++bp5PaNk7j/Mmiq7yo6PEcLX
JsSrPIEJc+5fL2VEGOnfP0xrCwLOJP1EVbprYp88EeCJ2EyUBqZCF68ue3mbCuzU
JwPI/Bd1yIn46Qx5mZJfnqe0vMbJ7R1D3UIb/8FhuvAE7f4KVsz8DABUtXjMHjjo
GfDo/s8ggSPKcm+PW3kZQMpIbfq+mhLPIWRNubzggkQVGAFHk+1xzY35np5Lh0Wh
Zmwz3dL62dvHuRd7kWUQl1YSFZ5rxaoP0VYt8fs2h3Ng60NBy6WgjXeFTYdk5sy+
ekh5gdyfU2aqwUi53xQlKLR3qr2sW+rx3XukkOMVgtbe/8cql0EuL1FR2tA8X9if
BSTg79SSCA197G8Yl7di+q8HRTNGmWX0nABnyoAtwqO4mLi7VR/u8kP9aDlrfjOL
ttQkvyRLFaqUmqcRc7NO0l76aP1QpOsQibQhU0pjR9WNUnjrr2NlsmiKOSHm6v1i
4DJchzCGw4CIbPG8Gvm6nQQEnD2KpLEI4OZ1ZoFoa8Lpgk/a5bXFefsbQ1R2wByh
BKmRKUW1NazVZQ6uFpFIy/84q2BtG4KLyt0vbG3JPtO0XL7V9rgmKiOzdfmjiUvy
gJ8WXo70VYGi+63KRlzw3k1S/G2gEKrDFPthlzMQJXR0rKIQBDi0S4VsNPW9+SFr
IO0AAJxzryby6or4OpoRsRr7VIEnD8+zsawKVncQ5ktiCRwUdyNzZoa6D4DhF8+R
5NOdSgv3ooPzDiAB/jyzBPfO0fWD9H1uhzWsYZybOX0YjtiVz8Qw2JqPLmbshpHc
Xg1iIVC8muPmc9YL9ZTq2mkZcSbziXLuDcKzpESpFh8HGHXWGby+qB3ZZeet/mwq
Ki0bv/LJpW36xVHYsMyRcfOabKdY55Vx8HHLf6l1V9L3k7lyP9Q0Aa4k9OgM+Rjz
ra1TERxX72BZiR1hfNNFfIROOKX1xhkfsngL4k76YcZthu1HH0MSC1T2aVRzBICn
UZfiybmHS//gEur6zOR5SvlMzIKrL74dZhos/NHJWFIYz1+msCbZcgtzWNaA0mWP
1bOcueBiwX4d3xPCG1ZdJRyosM0hV/P2bL683BRZ62GtIvoumQJlOtI0Ona5Rl5i
sVEsaIZNlQpMb7lXVNxYR591oel2i64fwXJ7VmM5O/EBLpZtkRzkYpWY2uZ+/olp
LRcSMDb6hxvvWvOUcw/mL+6+npBk7Qbji3vrxanVNFMzBA3ie0VL/FJ+ruN7C3Go
s0W3ppSf4uzrVRpZT/u3ZPatvHKu5EuEuGfgJSvfVpPhEHDUigD1JH3GiK12qmFf
3CungbBahUm5042iPQeSdjk5a+qMxwJcubTwIjsIN4+BIyPalGqkutrdMcVKMwRP
FwmGloeI2nAHqzGb3ElrCX0vsfMqxdY3IMJbR0sSBoZgRgo9er314mEPOH2BUREh
FhBF964cm/utQoD1yU9L/9uSTAwma432iVcCtxVcUZmv2jJb0kIPiokU/yaI1Q0h
YYfB/aLVO7nRm6Ycfd53YM4M8jcS9XWSgptCISZb+rvCjq9l1NyJykSVGnBQkYq0
MkMl90zXJRMiN5JG7OOck4yllqVQU5F6kkg9JFCVHva6Nh0RuR5OVMRZSXcLBLxF
g0oYsiythWLLbZ2ESOeLgnE9JHTouISQbxhNbNGBnY3WhjQtIpGRuQKMuKcPVixE
ru8ibXuFZTzHoprgwVLir5nybzNrO6f7OzCeBY+zD+6kNY2208HZsT4phY7SdMTX
HFlDCbjN4vT44xwB8PQa2WDK3MkT7696GB0aKVMYFzPe0z/4OTzY6zRTJifz7+oX
B7WD9B+8D3PCPAsOJsj3dah6rU4CMCge7yUDQ77C2v3s2yGEokivyBB2ZwqWWjvQ
E2dZAJYYYyoEeS4lh92IobCWa3c18lGsJ0T8PfNn5WtogGpvKPxAa8en4jlzY4w3
TrTDDp5pREI1y0PIEqy7Jv5sz6Rw00/0PB09aQR/s/tgLFnRXrO8Yj7avcH3grZX
oQPwCiYflI4moBq5jyWSO5Fdb5IYEbBvAVoRtMOo89IbYXKBtHgGRPP8tWsAdcD/
yCBUts0m0IwU7YjQWrmvI7CiTljMCCD92BCZ9rCfnpDktfShJgvV4PE97fJek91Z
bwmdNV28UHLziRHkl/nHA6sEFDR27Ugr9z+wLw0Gmcv15LXy9M5x2acIJcNCedVa
0+RdFmIN09BiM1yig25qDkKjLAQLnjBYnPCl8EiAa4MQQ7sFrmg0Qs9TMPnlG4Zz
pz8u7+gsISXIWJckUqBCAUQxKHHcXxdwVF2YQwArU4OcvGSFIOB8x/IVrB5t3piq
VRf0Wc6y8kkEzHv8SWIzLcl2+m+oPRwMZmxSMgd+4Pp65cOr98ksqd5Q5hUe021f
sMdUfF95S/ksS/cdFGtzSkGksIIma4kxyJrm9lccHKWhjl699m2riage0HOthSx8
buEV+HV8uQX4mC4RtQUN40Edgluqe1FgdT7LxhMndWhyS9dSK38PlIKSvtO4Pqql
tZA2Ri7AqiL+mWV+pwG+Zu6fp8D1M5uaBBLRnP9Q2uvMkI8qd3yYKNQlCnJzEaCI
XD61KBRPSVu7Y3dgJTfEZ8tB3IjiS/4QjaSzIsz6z4PTqml9TNHVDUXodRv7XmlO
qrserz6p2EhTtkrDVv/b0hw5YnBpO2N9C/WKi/90f1X8rERbKkvnRS/jkhBbZh7y
FuDAD40epEMArdcMGRuLtzCk6B/9zV4EugdpF70QzhEM28yxymFFuW4Sc2NgVrH8
kGn9qrp06Uz+RKqRB9SNmI7HDGs6IIM1E9k+aaC8f7MkBjaJ/5nv8N5Su1ivBswl
oI9hGhDaF0MYoZxIefcZC1Dw0QbWgbmXYUUeU9Uoicx5Lox+eioXJJx2ozMT4cd8
zRqnc8GAMtQbgzy+Ce6aTOzcC4vwiNy5oi2Z2Q5YG0oHKGhxCK90Gt6u4uCY/gMr
wpganforsdauKdbYcnT2ZXGiJN+dkAPhc2WTuD/7cjBKJBBSmxJbhYXVU+7V9/xT
agHe0jJpaYarEDCn7T/5Iz0k9iv8DbnCGicRGI1lzSNHZjBZ4YukKiCYjTs0N1OR
tZhX/IB5Pv1kXGGatKfGFWOFgMgO4s3D1j/CQEX10/FFh+K/hkx5yayVPN/nkRyU
vDn4V62z73NTAIqenlyi4SCzD0EjzZ+lDXZWvHZdGJ6ZQ8G9AaTXyYacQaRTiVV9
p5/bnA6V9iwHX8o1S8XQ7qWtGeaX+KgBucrKJU+e+HaLUPbHGECVURrGvazPoEwT
xrKk7LExC+9wbdECeg9svVwrhpRx12br9ndunFpiNB/+N2zbFfMwGC1AdZMWTT8r
UWzX1q2+yfK9GBV9AzbJeCVaiNtwgWkHgPr+rSyQ6i5SeO4Z2lYjQXwQpluvZPTs
pg62ZPJvT+L3Yjz0xs5q06kqeuaS3jfWhZZVyNMQQ4Xz0RU+Sbejcojd0Xej5nYQ
HwIbSqQfPrR3AdLd6pQEtffdw5RE/TqP6rH0OoIDF91XrN4m/WSizJtLBsIu42nK
7tFuMPUKDdhwFzm9TkKTP63L2/uI5Oqg9wLsZ7g6ZV17L66VsFDdOSNMEwT3JkGL
ujiEMej8GZNr7V+AyEdRbvLHMtT1MzZ+Noofzl676HGlVEDDsEaDMEy7khen8g/e
D5ubDNk2zKFLJTpfElz94ghUCBxNALa8hQrtVJMUGr6SjmveoUvsOvNa5fWQJ7Mv
fqoAkn6Pj5jXHQx/cEVaa3kamBKZWhMni6s7sFwKLyFSya8euOF2qTOuhJvD0SUU
9jdAyR5+IWMpPzDKHv9eAdzDG/EvkekqK+HNI3cPtBS4Z7KeAfyODGavdeVJsA7A
niG2DCaj4SDJTdZrEknUA70Dc+0keareGZCrvUgHtekD96XyrCgg+vUcqbYKPyb/
3233IBJr19QXJ6a4cDbGSqWRm2WQRtQuJOuEwCQXoXWmngGLODiLWnYSUHqEJJy9
kwsm/+JpTUYoiaxcJlq90jyOHejxP8uhzbVHxsaZjlM8sa5xLnK3o3J9Z+NhPogZ
8ITJdbCLRUodc4BviyIPlMb0XOIhH8o08wVYoAHs2lQ3kwg2KiP45XRN4G4vrobr
ptYwyMVxd/EwwXt7+2JLq7IpR8VMkNxr3oFLDg73Pmirs/c8iVXWOdi8LR8c7btU
gARCmbHy/xf4Jx5U3xttxT8jlzVcp3VTO5v24djWEkGtkdLalEBcdYaiRLqctNNF
PD+AsMcP+QS6nW0zy9ze8GonE8RxY/EVNnwVyABQFchLv+GIhG17cn7zrPQCamTl
jJOd4zmZLyINbTbPEH6jliQYWrNlYSRFEAiZuLT1B4X2u/K25Fy58GQvdpnrdU4a
ubiL1ZUBlKY8dZ83ZN7H59kRp2i82YY4/23i8MIDpUrn7wLKlByjvxAs7ov/7mLN
HsCgeAA11DI+vk9bb7+opRr1fgiUV3nrKXvzeCY9NW8fBLOO0y4XX+zX+s60py8M
VotGKeBsikqFJQTlQSaqQGXNwIongCal0zHoN+KA2mMViYIikptJ0tu2i1iYTkFm
Ygm1xaf/C8xfNbRZ/zMuw1KCEBvN1Kj0QiFQw1G2gxDlHxtYS4vwjx26fOXUabpr
MStFjNq+B4vRUR2Pt6O4LNUdgjagq7ECEC+hW6b+AUsC+V+XSW1PQN7W30eX4RiA
Bl0Rku4c8Q0dj+DNEaC+s3UsDPtLmGWx5PosNyOi2r9uB5nGoQRZdFPjeiDnY8g5
N5BBYTzkB9E10LhUjErI/WicyWshECajATsB8kky/Zsi53GWGFfdRnPVUx/dsEpb
iHcaOcWI5Va/cnI8hhJqhy+f+eLThjxstbZWLz07dEZjYPR8XeQtDiX0nMZLO7uC
p1GRp5u/NmjCg9OMJUpxiEtw3JWatQ6ZWG4ucQ8jozVpd6StvI9kdThibNN4CeRA
5CgtMvWQc8CwmY3kHPyDdGFO1wime8IqmFbELAYw+Ytdnu7mdoMj7nCoZxP7KpWJ
PMSQ+Z70jRSOkNQiPfC38mH2dFOD/E+k74qdDwipkC4Q/LifzD/qhcw5BB9rQmHl
oQqf8mXEFgWVQhEf55xf/wTeAtSaPbcXv1UojI+kkYrlk4JYkn0ZDd1tQ/N+xYIn
Ku/Ftj1J4roIuiK5vf6AcwrTzT4y+HyeUN7bHIWaWpvxvfPvbYLpd0rBby24gM8Z
8AhBzQHtxTbs622Q7ahIUcVu3t6LKA8AxtGs/YuiYQQ6PYnkhDI9RlvX2lhh6nyb
cvbEx7p7oVBno3NY8g9lPw/fF5negLOpvWf2y545tShOr1D33+70FwuycfnqcJkC
NTS8kaoWXDfGD/ic4dt5hHUnfj3s4/xE5HSyPOzcCiteWsaZC4YFlhMKnOtWMTGb
rEOEjtTFQ9upUF8BWVTWBS/qQqcSWYCnr2qyu4v5khdSiZuBVIJtpRT0n2T3bQ75
msHRkymhL3LT9ZpKaYcUeAOqSBCtWDL+rbZE+CXXodqAeDRiXeSkpYKJbkJTR0W7
20DbVbtqZoGkV3oHYnECRUeEuhtSJReuP9f4dGkyNT6cbikBKmYaeYeJ6mTmR/fL
OCkJ3VsCloynq76j1Eo+X987O9HN09bvSqsMJ3KoWT+e/zcXfr2Zwquy/I3zjWvP
48B8xBzciEXOvMALcEgxePd3QFr2WSd2bvkOmiYTorzSQB3acjQ0n7r4c/ok5YTJ
+hASZpt78Wk09wtD/5spPFdy3FF9jyzq/fLyaX5AEssakfX8UHu0z9jgg6gPG5V/
6UhU5PBno7GoCS8ZquRQF9LK3aO+OQ2TQ9eVllWIbvDpWgUY7kifqQz61tMNL5kX
H7qxqgAX6n9wH9oCNIv4JXqBa+JBXE83v+U3SyIzpAxqmrT0FVeHoUPAHE/JBGp4
mXSCXyyos8VYJsDy26OACal6BXA3YSPUvxRg9q2/zbfksNfu1/6QWO1N+BJ6dLhM
N5uWPdxADWc3EtlHfdRBK6ALenBzwcKaApalFEp9Fqnml/ltYm+aJkytja2tdLtV
RZUuZQ+YNVbugPAhacXs5dx377KiapGoNVBoGgj5eHYwslKuMjXVzUcrUemxEEAP
lEMIPeQxo6KW6MZgmlMV4l1zN+Ru92NL1i/quhTnZkGTUcACufqfUojtbHRasBiV
V4JbMDw+hqEMRAGi2/S7GhRgRWFrQ0nHvtWxPy1JpBajwHur8MZGXf8l0EpYUrkX
CAdKcS2lJ4gvF+B/f0eZjtZW4EYFMEGMiKI9wBJRDFBsLgNk213Xz/TftKzYu3WM
pH7RcHxns2lE7A2poyngZVZGsm/YJw9rAG+//4rcOBECvp8MJSMT8LypCkePd/BX
grJ5IE39aUev8Rn+TIdInG9Eol+i+sv98zJGF2aR25eMCuEESxcl6mSmFFUjpsnN
BEGWZY+/F5XCz4rMjDgy0Cd7rZ1BMfsKV3b0DU4o8Pb1sJBSZB8qxDPi5GcRvkH7
8s5uLR6x/0ZYhSHymSRE8MiC6Ii+vfx6YpDhw9EtK73t1Ic1ZNA+8aS6LbEQUZUp
sb9A5EJKzkvbq7Bd8xt9ZoGtMETKadNjf+VPCJ1//mOWQXozPAtvWwhcHKOz+O7f
p6dfR/nddcV7IUM/FzDLa1ElaUriUUyCWd/LV+GuosPOXZdRbgFlRRqmj0Xv24P2
2V/XDbwRnG5JKQZZ41edjUkx0Oo009CKeVn1OD+nDR7JEgp48FAdXCLre6O+nWKQ
V/y4KVs6sVY4b2MruMxsSdL9u8CUwcvxK23PJkn8G67/uYZ0+RrMupkwYEnQTs6b
HceVHvl7HtzL/GaNWzSkQoOMB4jKAGhZF5neMejaRUztfGmehtw8QpiVgTxpiVjN
9kjhcyd16dW9SLIix833GTMA8cCIBkHJ3QrmbCJUYBbXPGs8Uc1UKwSPB6Mb8if6
fI7IkLjuafTPWq9AzqeynPdlsi8/fOCfhN3+jt0uIaG1NlM46OyUE4bnk2JC6XPO
26Yc/7pZcFquoxHLX+M0eB/WP7S9UW4PSYni06zRa/H/+47R+1LLnRYJbagdijkB
MJZZzzppQpvvqqgyzS3JhxF0V6TYEM97aHEqZqJQ1sYgDNZquuwy9j1RnVckCsO2
h0d/vvXAh5FwZn1k0ILtfs8uAs+PfVnDdq4buucy6qlSonNXEXto6YiJvRQ7N/bp
U6yNAPpLsAnPVY4Zcn7beajrzGL9cnrP5c0X8xUsA/hLrhh6gPQkY7cHEdQz66IP
6hJwHu/RNMeePk38xJvsTPOuHQFdGMu9FMz9lVXSPyIgBu2vw9K+hAD9fwmECuFv
63yizMBaba8C6rSJrZb8maKbsX3aYHuUN0ec10rvNui8cz4gf0pBeT5i6CNbE0th
/0yWRINVi/5ewIzofcX6SlZcuKu19GrNBpKTUYgCsYA3PAeKY0WDu5++LTC3zUxF
PCzL1QPCkqWtf71touSoagzaEN6Hlyn1shEobKhaqS3UM3Jl4WWAMj1+TvLP+9Gl
q80lYhTIOtrEnEAFpI24AZT9GG1+67fmDegTqxIqxcpDyG3LZWhXQ1NjP6RGdesx
AOLWTFrrBaJCnW1uCwzxUmr1HwPjuV7ocucQqixciNhO0yY3h1LAa4PT4u7RnlUa
ZvmQBywaO0wH791OIPjEc0SrZQNncGEHU9y0h1VfCuVcC4z1OTaEHxLLENAkkcm0
MZnQ0hEr4fWzSSCkEpzN8tbdpwawy6MKf6NBa4Lu0b2d0faBGv4Goc93OsakUKWh
VQfmukFvdmtyj5jH0R8GZyddPqF4iPHOQtjLCuDMr0tpzjZHEYBQyTR+wuHwrWEQ
G0oGUj8ptSJPTkNxn1umqBtTJxlGCRnj8Lg8da1b5UbDHHaQ6y/dCzD8/c2JLopA
WXeXd2T9vRkwhClQjgv4aO/a/H1vlekw1XolE8VIjmDDl0FG7GVLiAHcBzK6qAfW
6bPAouz8pfobxDOcOZ/40Z2UJrdMFIsGsJHBlIa0kNTiFFk9KqfGhuhKcCceaZTN
Gdb14S/xuAzJOXQbdlK3LedwSb6CoAB3Imc0CoBVfch+Al8+2DeLR7H4xHvGj7tz
WCql+8/i9Pd9RYuumSUo329FVKd/vsMrHorCQJFvx1EOgKZqvhM7OquJ/MiD0MDX
S51jUH84X/E5rlCvR0WvXVNTJTBnOsW2niSUxEmIo3Bz7dz3K4Rn+e8hwNfPl2wG
3rNKmXktUKf8LGe5Qtj3/QmttCTGLp7dTI4UgUKBHs9Fva+Tfb14lr7Pl4EIoZCY
SpjD3kleL9sLAQ7ARjlQcIbYmnssykdGRO3+FdoM/MvEPKyh4E6i69+MpHHSsfEg
cpBsxduLo39ate5nhiXppYKBLVl0UDot+9+NQuoNvj7+vqxWMAN9lZrWo2HFPrJy
mPiL1C4lx3oltzzul7ciTYTbbLgjCtoUt5iJzz7NYFJLfbNKWaJmcGNCelIJaCsg
Y18mfJLtVeaqbqYNRovbcJTDMo8+okTwvev6hPm6aOPWnUf6lJHHvbHc2P/A7+/c
HDv1+u0KAcNVg6riK0H9KBTgk5Ui1V/9wqpMnlSYlbu9MNFJ0ywuvAMhBoOs3DKv
LjSJsN8jyow6dNtXC3Td/jQ1Lw5Ax5CJyc6NJaUqU9cucxSro7Etd89Tnb+n+d+9
6iyyhAa7/wYOaaABI7RN1aNwbpyWipZrnaqXwOdpRSavalFdxaxX4z4+UaCWuIic
/Z1XLw7xaqxhLVhaf62fjyz6/HZn9QQPODdFaNUDerPDfiMeIa2JtQtZWJ4cqgXi
m6HmMTIPyK3Qo/OQ2Mhjf3QkD4DFkrmdGkksFLPBWRhWtEbG+U7MX5yG04G0YrQ9
0bc4dYjEtW+NC2kXDOVkkmL2w71AzcU82B6/Ap41/FBo61NBnT8azwFCFy/AgzK9
mnlEYnnruwOKuMnU3bVx3Cz4pug851VLL2I3ITR9v67oa1xSHyL9HiQadcXi1UA2
IQaezwzxrV11PobUPzOZFiDsrjnipa8ezAwwj2V93cMFEsYJ5yO+3ThBs6KdnDdA
7E1vauA15YUy3xLFXSzG84HFFh6P3dGQR4lJEXdCPCVuxTvIIyD1ty3qYaq3qVQG
Re3hdGJflkYLvhZPC8OuL3LzOL1Swc8OfK+rCeqLuJ7r/563pWuA33zXfnZvRbQE
dzKXEku0K8AxvFdn0mIhvhFLDnRgCcrdKDi0ZjVxBWNCPkJtU9qlnhzRiejzeieE
dGzpLoR9BMQo+krmoNgCzcx6nGF7GLU2cccUMbQwgmM62Jhotgl4Mjm5mwbgvTKy
v24BLgee1I7rPJPGIqRhsuP2CzIDM2bXJHVlwHJEHw1lYZ/RswudTZD9O3E8Vls+
R0OHR4vof+DW0LS2tr6LYjf6ozND6BhV8O4FxDfjWbpOoNgRSYMQPzt5C7BAlr4n
cHGcAj6G30z6LNzr1dGh/gU9C3Nu0Rh7ZCplG/iyde71M8o5lhRjxEUMR7Uvl8DQ
AstP3FJ4UFdIKpgrRRRlEZUoWLy+YabpvLPQ4hqgYYeMhSld18VVrSA0iL5Ut4Kv
XVkTzcPoNesnK/Vid6QD5dSF8qeoK/teUsPLnQ0BNrTIpACyne5w6c6WAmhx7NfN
aE+wVAn9rPPrh9a6cQZWocM4M+4lnroEKWftz6YOZ7E8vf6zTVx6JByToc5vGfk1
Mgi+PfpFJ1f7fUeOET4R6XbrPADKbC2aTqA+yS1J54fLnl/N/ynEoFnJOfzdiuMm
IBRRFoIpNm+fwAe3g7dGjclgwkxRX8y4myBhsfqCxFu+KF48FC9CDAxLgjT/Jlpp
Mtv58w1J/cW7SNHR4hHtwIJMJ5y1qxe76aWVBIvWMWOzhqjczmO1upMSVEQ/2iSX
54rlrHdM/502/BIkzYXgyLfINVq1Cp7Fxq8SjthjeaQY3roOzxhdT7s8fiXZvFDI
wrpSxOes98uiXA8ZL/eEB7Su2vAFwZLb9LFKmpjve18rFiMG5+J5u+mppqNuX3Vo
sSorZlCB9zR7fS83xZhIerYhuo/0z+FoQAaY8N9vLKlaiMHiXUOgCZ9tbdJo1KLF
qQs8wLPR1ZOENHW1vJ9By/iI0jHshaCZ5acEbn9/Bp3hFYfZgfygnCRbEkIJmNS5
r4yfmvZz+AaV5e9T4nCaGN0yGTZo3dAzf1ayH2DUReWasDMImg5TsS5jvi0oTqNJ
m5QkmD+BzH8nnW1du7/yeq6WKHdtG6rT1aiUmczP4zghEpW9des6Fh6/AqWTJ0KP
s9wIpIY2hKeA2kvPdkoEIQJnJIO2pSYmiKdkANvR7rN8ao9CCac1SZstNRL/qtx4
id6/Wc9ngXS5SvW3xuDBKACk05cokPik05aWH1nG6qdnmR7GE6kfIBBAy2IfDTQo
xsn8wFv/nOZrDPwtxXGFBIY/YVUMb7TSc+rcjb9/kS98RKFSEXhFVB2iFNqEuZn2
aJah8PgnHqmpEDRiR4G1EZgkuxrcrF5c2322Q8qNsdOD07WNeL9tuJwNZlnuSoio
fMkGCvweaW+JipovMyb6omLeVU5KaVYNd6pHHsz1z7ZKf03+Pw4mGbUn1Ww5yLMK
hBuOb7/NNmACpLtTXchA7RunQiCSeO7ttNNXf6f0Qhb5xA19bD1DsmfmipToLKIv
lKdZhhh0HJWqdZtpLOj+vWNtvzYAzMLfNXQBaG2kOsHURY3rJ/+n/yLU3tjBKf/q
CewU35BMfbxLJnUSd0KJqXxctTR5EU/VQd44GX2C6FxL0QDMUTA58+UbBGMIqobt
V3scbHHUfpuhMMZ5ufU6j3EWfR44zRpyAcVmli7omQDI4TqGxfpzRIOV1EE1BVbS
eGtYlvm2GcNL0N0Ir7xW7IyqzNHomrmyAjr2rIaKVN1197gc+B08jNuAr0mojnsv
i2fCxSith0c/4W/ok4YWXxxn9RkNQIArnd5cP5l0nJGSxCKxr8lUoXY0tAgL8+ga
G7fOIQLIy+TJGG2xAh99817EHvLp1wA59vY2w2fb/7SXN+X9WUPzvHeFgsbiXg8d
T6Jqb0baGIErQNWazyH7Bgw3SwN3XfjoTrKbikNFYzN+1LhlTKq4I7dP6BdaaqpG
kmY8Kg4dFeE7KL73zKY9LQ5VBsNFQOCGcHA2c3rzzQYer6hpb2LKvenA4d7vdhb6
GXiGMM+qFYN3WxDlgFILEHhZYSQ5Nj7ga9yT7YJCQ5GfHKzSVxcfER7fL5q7arAk
DjmmjLwnMA/SanhHJ+Qf/DwMoLCbZv+7KI22NrTnFSE+vNhIN55EC0vb2KGLaDZe
lhpelG/ju7LvZLGhWlL8+Inv8Gtm3NH5ZFESqf5xcMbofHZFpAJPk1som8CxOxzF
gXrdECAwV1WtJf+dPEqr80ATJ4X9+/g/Rhyhfo5WlA7ajgPaDl90QgngEZarl3I/
pZBNAn3IBN6ga1G4V4eLwwHA0MGeodhOp8eigGtSjf36gsJqmcOv92qF4rh6q7Vl
RlzgIhhmcfzL5pqFrMmRI1BthecpRZhPdEcGTZPkmHcKNDlUsGxce/L/wiGQbrR4
Et134eqBFGeHUWG2Um22CbwL2zRlzMvRKt4Mg8gkmxAZRxngCKhVvZ+5R6wTiES3
ZrhNUk1klcmeFmRq8+Ecgb7hzMUljIjq88eIQ283XA8usYnnLK763KdlaCYlS6tp
wZR+X07UGirBH2T9Io84VzC1UmmVd9L/jYDEK82/diWTustYvhfZUFOZ8XpmPpBK
mOONSwdrwR8AXRh6sl9W8cnHY+1I0p8FbFbeudigCSGa6mAsc5VX1Jar5kCAvKwS
uLXxelpeFmqb9SzzC2Pgx1X+1e7rKhc1KYMY8kDmAT4tBD5NTfVr02vu2X3WJWNc
QVpag2m8g1b6n3wE6mXcc0joUQC0Q4TeTnd4S3ISV4aLDsSoB7+4pJl4DWHEyeqe
757XtWm60zn4PISPO6H3xYNIEEjhCPn5EbImnulx76G8BMUoyYVunESR8NhYRouc
XYB6ZE8YpTjUd2pMg8eSmEk/zxhBmv1q+BU7JJNBmK229UBZJqfJs3YkA6zKlZvu
wm5kILIvrJ4xo5vZ96XH4zqHOXBu3SDHXij7mJCJ7DhAZHJ3dRgZ5VyoIZp49x2n
ClBWVo5XyvfirYBTbIXz07H8gC3aOZwpIhpu37a1LMGcyWYB0oyZUi57dQiOKKjA
ILB8ijruTRP7INUW/oZzWdLOv7x3vDJ3bRPEEZswe0rYtAtg4UE8X8nL8wZnFiUQ
nodZG4AgEGfQ8NB7dy0n5hsW80KIdedkqQxlNJgjCIV/Av0x6U7WE6ZsGttA4FSr
+KRKbSUKQZw+phmw4YeEiBHRxwTAxV1CRsPc5Afi+7sdUtzNvXGEaDVvYGgMV9of
AvgsQG0etMxzJokUypwzQG06LA9niJ5JAZJy2kFObVOeWWsvgFGsTx9nAV26Irox
oDF465Zd55bXuMwP5PrJl/Y+JvcJ1fi6MApbQ53n0jzaMJUB12Pboc8OCLkJsUa6
UoXVW8IrTryHF+SISR/QjggF0I5KtNy1yKde4Q/7fcaJamKL0WwVyrkNcWLVKU+J
iTTmnS5uM2/7sgZWlHphPvX+crWD+E40ZFxAfCXnU/fBioSIhs9E0pwJjjxWDNV8
LrqYPVdY7Z44UviZ4G2BdGpiInwcy15S86fvugDcga9k16TeYdnOG9hTFUm15E8V
SN5YwS5yoNzvrpLWyr2f065KXOg8ubETUnU29+MoEfcU3b3y3mDyXF8Id1oAaoOo
AaO0zPmcepnwxPIetXS4aS8VuSi6XZxioLBXhDm8VVUBmuWIEkYzFai+9/udp1QO
cbSuGntFQTJG89MqNRre2roKT8LAk53pOa5H/b+gfefdjQrcOu0K9Hw3UzYxFmZI
VQdCfmO91h9So3HwP7wkLtHSetDyMTOT3AGUJ4+DsKfub7lNjYwtSgRBPSgQd/t3
Njo4akxHFCEywxum15jB9Exrnph1dk/qcOdGUTOn37C1B6Jzxz3eUrol3aBb0aaY
dYZPnnea+36hsvKt6T+eip7skA3ahBPXYsuqlEJQ3TTEgBP+AINOfznDvEoopGNK
vwuQJyCD4ORrkrrucHn8LUb4qE1GHhLYskCugaSQIoLOashWrUUGZRMJwQJZMvrs
QHKkuJF/JxGTxBJKTNwairxMSt+hCqwtaL+2bu3V5FQH7u01tzcIUABjb+rn3f9k
MKuwW2xNrR9Qo/XtGRMFZ07ikFewhdrtIzd/freGbCmAnT07IRCc08GF9yqqaWY2
xUsfW5taHYBM5hZSOZuTqIwlV5pnitZ8vTMmkGhKx4ISpGzHotDvnYQxCSoqFNs5
FeUyjOlIO/+3n9JtBoE0YDCHI5aKccfwZ0s8TGVd5K3s0Ca8xfALQnYu5PF8C+nb
wCiTSCt9z017/1FuQo/C24dALGyvT3o4JRm1LdHwaMaoSBa17AB6VCFv2mL5d9ge
nQr4FoVafa0TaQAXtU5XrlM26dKwSjrhWGLfY1NS6yTWBcuJLk2jYVbpAK/Jif3A
7sy/3mnmAkjPo1RuE0daSlQUgqjbq8PHvA524WvygibGXXV+64LX1VHnljLeyi9X
Wr+ljAY7FIVzXZCHTyg4e96GCyvjyFR/2EAss5T1Qk1hgI07/jdVdiNPrOTiYIbn
7TrsYiKNacIBX1YuuiRnocHWpOWXHlEsFnWjwojAqJaISLrVPmX58Z89tjY57ks1
wyDecKSXrnJVmyIbxg4hqAWbiHVvI6roGSCEZmEVNjtVJsK9aYuf8BorDqZ3a0iJ
9uNzuwdNcnrYZgeOW1SzftyKEre5H6ssOtDPGI/dAZX8gMJ5Lhkl/A5+NVvj5wZr
TQSh/GzDlIWEC7/xv62jRplz/D2CkXJn3rnbAH+5He91FqinGrqf/pWO7zXA3cxG
Ld4Tcj8/Gj7/grk/HXrIKAptfK1h2ASXQxFounq6FKGB7D9Wxuy1Ivk2ablfHfsH
f+dV9gxsaDPS7W1yE8oQB2nqL+CS/JvaLWEuxkORDWjJre7KZfuCjvvk3jctOsuj
6zmXcgsX1VCPXCemYAlAujHQ0yODW2vc0V9Sgsi934Ye0SZEV6+a4AmHnyBYZamM
b/351WuLVUPFsLFEtLS2QUfSU7od4va6n7Dtq27k7YrqW5GM2QLwOuPpkdwq/5+a
3wACwmPcQd7FHHmiU7t0+IPOT/JdFO5ArN7GGyxuVnntLymC9lZS0ftgp2tisMSk
K/jiBQxmQCrj8IHvwk43cv9RH1B4+z3XcW1PgsEvjRQXB1SvsttOuXsqXAiaRQ9T
OqcE/MVhdsRQzV6fujwCqG8qM2eJ39mIREOXtVs8R1JEDjPdBiRyAmDpVx5peylj
faEJrLvPp2HP+B4gV6ghUQTeUFwG3SbdPtfOOWrZu2Wm0FtDrYLCeu8GbUXu9gfy
jL2VxnnAnCoNSXYDHOZ/UtydnU7pHaiWafCDDc0Q40d32zMz1hX0CPEXQckKf+Ut
6AlA3kFNFlGrzX5KBH1hiVlCsxzKPL80JIriyEwYycxUFgf7It2Hzi3/5m801XM1
1GO3QW7rGXdIR71O3/UFz7oHz4VIVjLYSiHF8BiUq6PSoA5Ujlt8m0+h/Fl7eIPS
gvt2qEVbYHXFYnq+RoUdCiZOXRE/8ptqVni6OOilvEhMdiAPY5+eOl5gM2qg7Wec
hNESW9CDXFXyydBZ+e1tWdNp2quD/HFxTGOKfTtVuKgUXgkGLo3lHojvNqmsGJsm
IONC4lGLIJz67iXdrXnctRFRYnzuRmXJvmJlti0fs/M5I3gsWaFkQGHgUrp1vSeg
X+7GgB0aUAoBXN1ARE/dHrKMtyMOYp0IuzZ6Pm93tNcDE9fQJll1wjP49JeRafJy
wCLTt0tcH20WhUSl1/AljW3YuMzMYaebo3y0ca2vuVTw1tj5aWP60xQZ4XLrXFAK
GFVSqVDvdiYEwkrRARPua+C1E87spKn+3nncIojKFvaHqaZ4k1B4H4eZGAu1Y0m6
QJhPJPKAToNJ10s9G+SNMLNOjGFXth959sBTxgAULakFI/xHwi9fFTckBLvTyytu
25fWKtTF639yYLtRVgQPB4aRk0n6LyNbRci9T3F3PVAyjn9GB58x7QGo/Q0UBHEz
T2iFeMC0DZO6EwoKf4VqGEW2rWMKqE2GONR/Bv8RF57r5EMhm+J4Osc3SEBuV0e4
PnTHZRGCR3fRpl8PtL5E6czZDNfnu828q/JgbiEBhsm3y/q1g3RnewpNwE16FbbM
YPS4Um5wIZhM4gXDCf2RX4V8KgPJBm5krxb/QMKHvGEyOsRWhFeV0xHteSDXz3fG
8dpGYqqdAIwsY0uYhWmXmyMwI+BBclgobcR+7B5RwkWLZ7vNOwfICL0VaY8A2O8S
6e7D+aLep9Y4IIvPOc2TL1wu8ZlBDL3fF/zQID4kTkwRU+07MIcImYECs54YCwGA
+k/raLKszv78ZvJpB+lZsKvt4ueJSmHSbQxf3I2f1ifJNsKNPkCVBtJIbVfjm78o
D4VxGbxT1bsT2+b7RGIy44OeucHam1em6thHJ9HFlx59+25kLQBbAcuvVqGSCbnt
AGCB6b49Nb1E+bDL/aozloz6WiXxi24pORqPnXyxA3CCO8E/IkP+ssfwYI5wEt0/
Kpq0aVVGyfWGh8wE6DAfczikw0MvexsN+UrOHeXXklRgKzzvGVdbr7ydzwdw2wGH
BWnlXlqUy4IHOJTHeQ1Pkhuzti8D6cGSRnWLUU4ed4jtsTy2zKiiyv9SgFo3Xk0h
XkLgIasvoH0ksXw80WhS1x9Zciwdq0xiYuWMdCPnnS4MJPyHOgVjfKZM8Nvkvb2c
2QwNey1Y5vlFm9O7UIjgyp+cKdiv9tpdQLgJmfoQY7J2jL9UTs8rJnABlOFydTtb
cjcCThWFvkxyvIZ/Wu0vt9k3oQogxY4Ca1df1Tid2gyhUTajx6SNy+CQ/KC38ao8
EPKACuLuM8S/L6Vwm5LWogo0S3wtAZ9o7RsubKOoc6gX/VPUvBItVrQv43IJrooh
aiWne5BDUB3v2JoTuufeeDhPtVkeyV0cjkgpU4I7XWt0FB20VY6Rrg11+u5ZSWwQ
7uiwX/IzcrdSkgqzlI2jI91UqkmL2nGCDUjPJCrB8grhWfHK7kEh/qbXLADQITL3
fc+OSGfa+5V44ZWGw0vCcV96+DFe4Qr5wX17NjPDGEbo07zlFSjVZyycRg35QNmn
rg86KFtn5urtfo7/54RmdwKOxSkMl4Pt1lJGbuP+21GhkLiJRaeJt2v3hEh/34Qz
MfYDVbFpAl2HfeLppliC+iCpCBZtUACJumm3nkBy2yBBTcI6ojBiByCj30Pdc1kQ
iAhYeL3r2MTizXU9fYGaETwQdOtfDKzJfrwK2lo6SL5csuq4pjVtQ45Uehoa8Kwr
EekSsdxKYqq+LZDD8N6uAGkohUFH6O6PZw2Eb5nVl4m4I0S5sN0tWmgNuSP7KRrm
zflmFV8uoffeWaINz39lr8SYZHserftMMHQGEOlY6p/0j4Ef/zQBmQoWyjpnmslt
QEnQ600Sy5V37D1rv7vzHPXypSFArULQrmMNAiOJHklsQhYtaTDzY6HcedeM3Dck
UNk+pfeLNnUDRXs6QPC+kdYRnFvx2gvfZFePkfkbxYMx895MQC1OIkQJJ3lG9rX/
ahHtClOX2Awu8+Oya8oWT0jQgDX3b/4yyziQC0wyaLWqQAK6/qYEfR6cNMyisimb
16VMek/K+unN3jsE49+zx/L5YV8dFiyzEYmkCWYFCa1FCky841c/Q1V6vtBeUX8t
R27NDvOviDnVxEJgZu3/D6YWowp68b8Ee/bY1PYpbrF7XJ/3RHkQ9lFM05BwP2Dg
ORHKmCB0BuvN8hM7QyEPVqFULw4tkcIzNtHWOsZ4+QoX1z6U7J98Odiky2F3TOjf
eYWveZTnx2cA+39ZdKKJBHE22Em4BOiTZHWoi3+HxQQnsbbDqvkT0hp1xlghLSNi
EuTZnh9ditF1lGivQ/Z/FGkKSJ31jbkBASD1xYNKIRm6EpFZDRVxiI6qFDaluLEs
mgUWxlDxERp7pCdl5ZHwwb6ChqirRQX4Sl9q9hiojcYte7bV19IOkW4pM78yabCA
JsBZgPBgphUoG2lTUBdS49qYiobRsCWry+DYTZbPGtR+fVxJG7sEFtfoKnnRzgFZ
Pc0xvmqr6OfDxcObvgN/CWetMp1EghyybFFtroEPX9ebe9GU9Eikp1YXklcOeKUh
jCEvt/X0q2lfLYSw59ZC17LJYVNMfrMt6TiwpkO7rdSZDvKiVbgJwUz5I2VlfBuz
6OkbpsvK6quAxraJEPtWEc71NEmgIt3hhNODRy0Jt+EzZL/S5UQGNAwaFAxg27Wy
lVt4OxDNuv+KwWTZAuAR8RWBC1c7ij5CCkYoq27nDm7bWlQM+HnT/SlyCnT1lUv9
/XjNVdF5KeSrYKGczKk4aNWECn0YkFtiv7Is1TU4B8g/T3GkUr3qSz+K7BuHL1JB
ZNjHgs+adURn2BmwbS16FTqSli+oGRZVrGGqdoet3H0xktieQwUlGfoxueO/sQYu
GWamxhkgbAcn0SkHlUr0raQ2P3QLUZGGYfYrEn14x61DMXK8oPoXt9vDwJFHO8fe
8X9POZmfOZg8ueE0U9jXgYtH4FhEMUgzt1XCta6cTasO45R5VUgDUGPZTj/wOJS6
vsxwGoRR1gnFvhrOpiveLmQ6b8tPeYxaBeGcrYnzF3W6xYx/PSO2iBj6emRqR8cK
wsc+iAKNzn1z5yFFJoiZpRjKyBwuKQVvqVe53eP7dB+N9rj8W8UbvqVtYM5k9+RV
pV0r+au5W04vWtfSozIrN655bNK5YE4PuwwRY2WZy9023Lcjlbw1aQvenXkcIEeI
VS5YoMTSlHXfrY/5Aa0sv9wOP0YveOfy+MKdcaoYanfGIlcrg2VyGwbIHYW6hCvp
ittiaIg27XKBrMyRK636Y9lGBDZOqr4RGQvb3XKMDhCkgC6JoVTPgUezglXmPf9H
s4dTzCiexsFunRs9ynYsbV1UmZO6scPbH750AgZfAc/a1MIthMHQ2NpEO+VcHMo/
kg5azUSeB1I9jGmQeFlzV2JOSIusvQ4XcLme7S6qbs5KwngEnffjE5WZXex0hRax
3zVQ/rDRXTfUPdABi/34+SBMM4vtagutNpHZnHstH680x81RomxbKxZ5+imlegEu
GbGQqUdhSmIJ3LTwrLk7MA9iEJ3XK7WGng8nj61fkQsqOwkC0Tgi9tpNTQDbQ9dr
0B+uSNyd/pq6l2D6ItQJxytwhSKOXga9QkLIsbw38ubJWiONk+RTF3gyw5X90qAm
Up7V4ZFWNH0mSGevGIubQ5mXw2xE8vqx2sCDxfIO4TROjY2bMgM9ogTANhcGuvp9
q0PgwEWItvx7ybUIN5CJUIXx/QCVwzdMYpcghDkYuVhNOl/XV9mdI06tt3ue5p0d
EAsUt2M9qrd/Vxi9+ub5gKPIAHFTTtv/yJFjYGzJs3LdC2MxtP7EP009YDbHaroF
BIyKnwMQ3HDvE0a1J0XnxapxfOc24GFJEtGvo7syjs6pFlnr2/pHVj4wPrtu02iG
Nn8NP+U/3nI3SxEHGk+AhHqa4PBLq/i91UbUhw9nrK7o/U+O3zDLyTs3b8ruuhwY
96ebYpUcCgJm0WTGx8hcT2b0M0CXfc4N20ZwaP4IsUwQB8Tdn/aR7UVWymos3o90
Epo02LCQOCnUtoJXQ9nUW7tQY3utJipvdtYXSVBJXBZ7FRV6deQtkMRLxVUXQ8H0
UCIxlMIbyQF/12BtrJebaPoP6ZX5uCBkLpNxC4e98mc3YILJUFHhhBsJ9CZ51xDZ
3pQIKQt8sF3011SoPIPpKFJ5CDfUMF/VygW9ZPovZ8tfVHVnhYzR5ZDSfz4XXbud
2waujabo3GJvAOXoKJ7jaPILaKTeXMvGxOMP7VKB6KfZHTjvOTI37TrJGYRBiapf
LHwti0+fvdgKj5dX4RT2oxCCKLe0CX3O1rJvU4iPVwMC+tI59IQbz2LicCvY9BQ0
rhncaEX4zHPgQkC1yVQwzlsynvu9DxbRrJcxPyowDqUud0X93Z9frbtcKqgGG+ii
DUJCusPsU6W04JBuynYRzr856HTsOgo+e179BIrMJtFvtuLIp40stcGpZBuFu7rk
NHP+EiUbHE17LD3LuGbua71rPHBQgt9hxEQtfMtnpnelTJsQbWR1hZJeJ1Yi8u9P
ToCEu87J3ZGj/6lKA1xZrT63GcvSRW+decnejC1Q4P+tuuAj3tppsgj9k/TMd+Cw
3IoFfn1eEPw12r2B0h2GCjr+LVr21778oTxa8+Xc3xgRI27ysfktVFpQ5276fL0b
Wu9Ah04lSSXKt9yjEVDGHIkys11wDzFIlZ7CIC8zY/kXS1/a82sHXV5L5GzUwC/3
0ANkig9ujrb5Wz5CIb/xWkyF2kALy3IuU4GE8x54ImDyZU716Dd6VyP/yCS28IPZ
g1EnEiP4ABK/lW5v2rz4VGJvIo2jwwr9y/6rXbrTCwdMxZGBLPwDAKPyxLY1DeCO
uDPvD1v0fWUGIVPsOdzEXd9ZbJNgb5d6MkjZ3iO4lumvVo4YqFRoB4/hmXgH108U
bHiycCopIyvnOKHLRH2zwJkcKBmAhWnYD312Idt9HKzk1RA8T4+lQS+XQ2L567jg
0mQCPAMF39l4ElxgpRMidSMv9WNzYk+UYuQNZIsMCuCmjICG65nJ3S2VozfBSA21
7P8tQQrqboyShtlvtfepGguoOmu/GmtOIBFjNovuRQoPdV/MpvGgpFCAH3clwQSq
CtflVzb2F1u6HT1dQJPMq1bpZ5A5rmrqowFdw0jzRuN4NoxMfm8Tu1kqUzcEePha
9LKJcico3YKKX4VkbQXalbm5vVKkAnFNAvLYzyAJqC2f7WDPqj9ERMRs+mEpZbWH
5JYO0apcsoiqpp6Tdb2Mwk5d2f7wNuJFiIzjqhxxSvOpN5J1AbhtqSgcPsJe0NlE
YGZwFV6VjDj6W6Fp8wFVt3HaTVLQFStc/yIpS4YxSbS0wzDKpT8QWC0yZHInbixQ
x8gYokBJBBDL05MyPMbexdZQQ9q/YoiY5jdG1nA7mQ+XEMKB4bYRc4Hv4kBtdu3h
sigTBcxXDAOtMPS0YgtwbLBGRCVrXnIcFopGPvUiwJg7xKJk0P1kemZZ3xyIZWQJ
LPZnApEyEDhhYKWoIPPd6ggSglnIvq8K43Zoo9g7R4DmW5KfKEgcSGrx408M2hRN
NE32HhDi/taapO3D0hLSrEmTmgyhz1pFBaGJ6E61aursDyids7OAy8Wkfning55D
mxJs8VZzCKsQ0qs+B/Pn1a0cDupEvOhnUOjvpq3yLH+Rpg4lzq4+T865pup1uLlM
Jta1sYQGscUD75LON6jKui9D8RztX+277WHcdF+Gvc4M/ssxrlb7+nVlEVhtoVMy
mw1Y1YBdG9YqSc5uPUEWNgnbR9d31+nUUVF5ZV9aTuXe9WeCAK5DGodb+Mfi5L27
eeuqPdOwHAbmleK9+okJM0y2eXMF5ROm0Do64WK1v6LLnX4Zvs/Zrr5a0vWPDtuD
cJZSL5I5yotS/R6njSICXCT4clwChnqOjtBeKhMBCSH7W+8/riEtZJhed3pWx3Ni
D0T9BZXfOdwksBs3bYveMt0kyCOSI8C9GRfjqdiWZiIQPlLWnIp9p4+HK50EyCAb
phY696IN0WTAvbE1kOd2t+ngvJKL27DvPmg0HJhlA6JgujG2KcCa4Pw9tFZJTWgI
gc00xQNJE/kR3d1FIavpgjMWqspnm/kY5jGhBjsYrge0LfKzH40L1LchtjhhjwKc
5GWxTPXlCnq7XLUZi8wGAr5Qv8IdjwT+Jxr1vUmR9yb5BWRsld8O4vtj4yzqKd8B
IR+M1cLYIyfji6Wds/49mChrefsKcXPlcRpOGxKbJxCHsPn8CLmIoDZnQHpXpkQZ
t0XQFqhJ9/07bUxn/+gQN0icovTaTi+SEnLe3E4MFrRM07ZtR7KaM8lHXP6uFMBl
00+UXDNr/dFhlym7IujPXPgHci6Lg35/224OMi3cIwX6lua5aOdF6rOer7kT6G6I
zOZXUAw3oSToNlXeFKBIlT8uytfWCnVauPvqjN2AUwH1vbcGhPlJSnyDQaJXzah3
+FtWGJgluwhZKoHFqoH8KVvZumxYvPmSY4RlkIc+tpjNECdZj/9E3LFxCQ4TfrdM
+5pnxthznC2j863ChyIiUI04/QVjAF9lJvYSsoZFhj6J6qj2V15LOu9Y8Qb0BeNU
ALuBkMrSMl6u8vXjYAStbd/fQchvPhBB20g+ifdTYh7tOoYwWxPKRIonYz50A1fP
MXN1ThB2obs8TImrYHLG6y79WFUxP1GdM1pWujfEeNirv3NtnvcPzN9Mbs4HICRL
OmnRJXMLdcXCqw1QU3HQ+AacnqVerWZ96VOmYmMS1F86uTDiJ+y2Wrx6OGZ28aQ+
jFyIF4i0XPHsaKl8XKk35t9tTXzprkpFCdnKXUdkrHFCOj6ZgdCOIb6bwBb2Efx+
xOYMUaO3bP8yokiOQ6qdAKHFGicxmB/kjrRvYhAd/RJPVT4WZOmOePuOO+EDyqr+
C2BhOlGLdylRCmc19tIQvQE8+RfDvjoKP/1eCLbYeJ0jdBNGfuHrlAHsdH0waqSS
ET2nwepLGlD0w+KsTBoHt0RBppp7tZZPF/02X8Mb70LVJ39kdEn2Pu8SfcQZpUmL
lEeVk8A7RO0V1XBdUTeMHw/1ORepj6bN6hEGXURtq1ojq33Fshwlvh18zFMT6woH
idbuu1I38iP4A8E0co3aVKipY1aEXJ/Ew7IXSA3yBHEAi5bs6r3xtO5xjKw9pTrm
ZtIAdLiKEQ2V6ZgfWldTI9f6NF3yPgfP6m/Ah1ATj+7x9jiFF4IPtTK9JOnWgT4J
YQ8psliy0HW5cdzjL6/0gUwEM44pEU8B7dmzd1xgFsxm6VgmjXpAbdv0BO1hiJ4t
wf2XXUU2/78G6UIZXqKcGkRFrZhlZI+e67zVYa0h5W00UNHESpTaV8U33SQ7Pbh9
Ap0VcUNXMcEdR8oeoAN7F+gnc/e5pnFc/wDbQhRS3BKbpEdRQp99JOefBOExT9t6
/5p3I5Z5ayW6M1EN01qdM5w9Rpb4G+CquRbjGOa+81Y/I9eQQuUiVWb4U4xBvK6A
RGI1idDvFolh8cj4nyjvEjjXuDU1UChrYSKdtlIMbJN3o0S+uKvoAjzwLVgjeZY/
cqt1z7y+kOIWyxBQPWvfIFIGTkamjdt0mL3n/HJcdG/0MlB7FzImcrW46lhJpCum
rl0aZNeHjU2OXELRxBtaqCmBRb6Iox5lPrRCj5dGRwvhV0oG4qQxo6NrBciZwDOn
0+OLuSugUrgZdENhy9uhHR4vXH3F/6LYW/TGzymnnPTQ/13v6M4xWApUpGK6gmx5
jFBrXh48vphzZSZu5dl6I2DxOl9H6lSSUQpODpt02SwZNbaSapNtIGILKyzfz90p
/b+EGkiuGymNB7OYfIDweAJAZHBLSKUbFG70m8dQ68R5Dwu8e6X2Mt3NCUc6kPxU
FqYA/8kop16r6pBzaJln2ejBRdzEbuGVnNo9h/gTdNvnleK4KnHyLnWUr+8vS46Z
kk31kP8GevFDxnTW3t/M+FpysKtuWpuHBY/vE86hsFnl93xoyp6N7e2OVg/MyScZ
bXAP9NlSpAPBZcRWIoNL5LY6qbdAwBc4dLBVuig3V+2hJe1MnOlBAoih8J8iUYw6
OK2K4t4QKxdnB3HZ9gxaabYzF7qhlYJ7mYw/PWXoFlEckX7C4XQiTIvzH2r4TY4Q
TuZj0ptWfWphy18+7spTvff+fNnDxj8+n5wo1sU/HVWamPh/YXLrZBSGrtoSyzho
6hYkTyotZqGXiY9olheD5yYldIh0cFNtyfZgl1HpuqYLtGeRYHoQdr0ZFCt96Cic
XmWVZMhTBcb52zntf8IfGG7NKiADfgyK455JJNN9Mt0aCIVhzTHrZXEvqN5GKWdh
CcYoljRlAgjDRN9MD/7K4rNhp55L6g253izR12NxN5paIlRoqnRgHpWQ5HcVxos1
Mle9rSLL/hOF8tW75HyUGs1UabvvMKGMKCk2YSZNMpopJNsx34TImpOALjpsSgaV
3SOO+K/FyKY94pGyJeW0SHTqj7LXeEtaiKfRf/Y8SGCSfLoP/F34uM/Cy4hXIDDI
WlCq3cgAVwigdRuESGol3X5itvkbe9gK465AAig9fX/fn2P1XT7H06BwPtwdzC3/
JmJ02ibxSDJfa/FAAAMzqZhFI4Kreg/+4rft4gWpxbN6uSR0BrbPR1yjWzOQcWne
2EQbjIUDUL5Q6q9cIaa40DEdjlySC03/09680LdXhDaVT7ecaphR737JlMtSyLEs
m/zKDlwpXigzwAbbYud+RL/E+q6/IITqFiYtTZlT+p3p3gzMMuLKxJqTS/EuFUt3
yLha+1QfX/SDomRtoM+W5CtmUfmJE9FokiPOjrT//MjlULpo8L+QUdPXcQALTpAa
MWh0aVcc0UyhsHnLraycF1FHguYIrj6aSXdyd6syrmVKNwBX3zBSO5He08iusk+I
QMdwEnn57/4pcIz0T4AI6RwyCKPhEACHhMsNfWZ4OgM4J3A3+0hfTtt406VrWp3g
B9WHvOFQY/5MFesb7/sGkm7QLLX9qvsSY3ZebTAvCtyJtxEdnKbO7HECxAp0nSwR
5yTKK+rbjVfaZzhcoF/Qa83VbsqlUjr/aj7J0i7XRNPlZ9y8lcUjXDpxo0m8Accz
KHlQugVN6pHqBx3RSOcSFKLPie3EgoGKjM2czGVxwiUGMCnjWXVdg5e0W4THrcjO
/imdg6aIesynMaAWGSjgZAYNAfkikelayZjJaC5wvw6wIlJbPZeesDHn32ZfYPE8
OzL264SPBR/fugGEAPiNMj4ljW8G7jyJNBjiAeYtTQYu6VmmR2/AL2wtUhfekfuT
EatKufQBZFtLHQngCKV2DHRUtCgV1oTL7NlckPakUrTJNqiusCJja0ewt3HOVNms
iiPTl0oN1+fL+ljwrk6gN7/liqAhliCXLMW56g54V0palPtL9Z/K92/5zzFZ3yun
H/6mLARDeaDxuJ3U0ai1xJIfV5WtOStadDipUW7WkdSCwkK9KdZFxkY0RhxMxo/9
b5w/Rj1/Gcnh+eHJSRWazR4FoT7hEm5XEYXM/O89xiv5Ur+dvtDVJo1eEzD3ehk3
0VxXfYzJDKeralSnWj1Ybf09fDPhWuFOsyay73IS4E6ZTA/i42toD0nHp1iFhSk8
tPBG08Buz0Z0Jxd/BzBYWjaAg//PSqRkcSQp30syF4MRRYHGxEUskSpWESm/jw5l
pOnJHXKWemRo8UUStkzt3/bh1Mk2xSygWPEQpe5F6Pfq1bEwwb3g2hyafZ97829w
mvWY2BVJ+hWbM6pEVfSBkuS6SRgwpW+6dCyVbFbIjgbjCqzSnXGkgedO4Sn4H+4d
z7ugVVUnYG0UwkDFTbD0iu1hDA4VNLgSpH4tY+cpsrFi2H7EvnkEGHSZUmhcMlHj
YPlgnjT6Xt32oxE2VPwt269pjGK2/aQMrMfBor7OXNqFUIyLg3DTzWIpRGbsRxaF
q6kfvuPET84TAJj1PuEaIHQpMDlDzXJmWM2o/ssWyEtIEpYThejO6yK/jjfjVxq4
u3lgl5EXeWGiQDh2DXkaAq6ar84wcRHIdoNxPPdX/MbM21f4Im3y1aOXFkDXy8iB
hUK1tIippOwSqKpOSSlvLAbfYD+sakA2EyAuLZ3LPc0bO8orCRqNBqTQG/KAGuqv
BUSwr4JT6yZxemuiqL++wcs0AmNI0rxfcQUbIh0OmBKtvWoI4HiPUdp9t8hR45R1
t0B/u4e5ANuOYjNLutXrOGakMHa4Fln9kJC/VI2CJlG29dK+c2vvpvO1pabezz+L
n0YwW163nBTivjtJI4UpR7Fg3cK5LgFhWEcKRWMiicpbV6v30ecdoLb66WxosWqT
AKc5gUrNEU0xQtr6S2RxBJXQnlTTyjI2p8hSexlnp2P9PqxL2YTpbB+6rrN8+bsR
5LvzJyHtZC/46EEXJ3f/gOTgRAZvAL/OTu0hX+FvcZIt0tshGjN+eVpf52EtJSGg
AAp3qLhjo1bvbugh8Irq5o8R1kqo7EOx0JRH/UR8zKhc/CkRrCzEH9iX9GSN9npr
xFfYSzAuKkMzxtHwfnxKLYF+Ex9HgjQ7d9q9HK29pV/1gYPARpgK59tHrwLpUxLO
z0q5WbAEBHyUlpt2YCjbHvc9abWNfjUQeCBuWJgv8NDZHKaJkTFXj+/p0Y667QBi
FDxDZZdOuDzXu3snM28PEhJBZ8DQxa/NuPsLrXCu7hMFNnJnQL41e0+zzDmtob20
ZUHcXWcLdmcPutQwgBWasded0So+CJ9RawBps0pavSY6NJuOsRPhfKSF/ShF9hzd
Oi39isY5jZ2V7lNpjWOdmi7SzRHa0sKcBGB/AI6PUdmjaTbHtKzjdkEIlWmj//BO
uA6/B6BcwZiidOWSnnL1G517DZlpczv++dB7n2DIDnoy5Or8Vv8vmxxwgEQ0m59g
PNo8WJQ6Mi2i6xoCfwP52meD5AlxnwM3hAXRcVCMpVRwW28gd9WlHm22oSOlHHwY
EeecGfxq+k4Oednvwee6lhJQeEeWKfJ3Xu64l18+FT7Fl8bs8myG+/ZtQ1/B1qfM
AknmBhSjeiuBNCvK88pZbqZl2Axfv9lu/7m9rYOzBc3lRsNV3JZibuwZp7uigxni
VKQhaOXzAUJ6d9skgQH4GpnROvR19Uvz86Y592JbEZKDwMlnvQosCFzqargia4BA
+czt+y04Y0Ru1ObiNhwFEF1HiJZN5GKsrYQ5GmGsnvU7e63Fb+FjevteC0sdog/u
98t3FzcNlaFL5dyQotsaAAdHxsivky/s/ApHzozeVCThgO1eqzD8EL9x8phUT1PC
8ZRZAmQ4qd32b7M+TqmZlsQx+QyEd14PKGeXhC0u3tH4Zb5TCFFuh7w82WUQ87Gs
Pqs/B7zkQWvP3icC+x5F+GaBqI9oBzUYy1XPRCGT2RUB4L1FbMb3b5KSTqMzlhdy
zuDO7Thh2ZRWnQQGDfFfaxIDzvYXWSIoRWW4uYZI+3jDb887UUZj6eexRmSfLvTQ
f6fxS0Lw1PY47W/X7K1zz0oyE1A/wsCT/6WeB02CKb0tpkN1O8tH6aHNSZsFahm8
gXKlcat9E/N4n8GA4PPi7aAFHZxTvKgl9VBxXpwXhj8M21TxjOOVlSek62SgUy3H
XzKNmDnJvsgvhwPLV76WXAdbTnmKZH8n8L0jo2mhPNFIWUC46DECNpPuDWQUFyKj
Xf8thIACtblIOJ9LwXFv0MDE1gphW1P93Er1lvXcxpNrBiRB5cvUkHWvTjkyPnTE
FuIuyA6ewjaEvEevdvsP5FQ+bncUMVE3pAzlAk8nYmnVo2cssI1cxkGKdUo8XjPM
1slcdEqADmDyLqLeDK6PlbPjf+XB0Yun/lTCKEDXYvKrVmHSgZwdvm+LpUYlXbjO
VDz9IbRUITiy2Gk0Sq9k8Vtrp9JTimBkiPx7UsJ7S2d/kM5BK5KOKlohboNJP80D
Pj4rcsMDJmgHJ/q42ElxK/cpHRJYeslx1E4fOgLU0nFCVyAtHVyuGC8meaht4B4T
9CKaCJYhz5k6uiBEDVl6Yo8PO4dCdEMfwFjS8RKTOK9c7HsEq/htIwYxpvjP2Qhq
v7fOeMK+v2MDa6kwXmSLHQVj/Lu6OqyW6OFNuTHCVA1iZlYO9HKxJZ3aAjrdrJF6
pfqBzEpOLAKZfBPSQBI72741t4pi80SSogjmmDqDerEKv0ui9tPbkIbLmgSvb8GB
tzqqP9bdmO7wiAHjnaM20Fsp/ayn9IaDJ5r9E4jMdGJ56p8g6ybeKX9e5o/Ejk3+
lGPxWwUxx3kp8vs3zW9AyAqujWHfFPDRbatYVSihB6EW0IqJxJnZ+bmud0JY0YjJ
HSd2onH0Y4thaPslSI4SCPWEYkikl8ERCIGcHMN2jvgrd7m/MLU+5gKXDLf5QfjF
VJPudQDHJdcCRKqkZvbhR6h1jLM4z7/jSvUuDTOWCNVSIhMh4A1c83Lxo1OdY3c4
8MCN9qsD/HyI340MdZ9kg2PxGWZlBgIogeoFGimp/P0RXTyq+7g3bz53WvPm4g6l
r12X+Koaa20NmTJJcCHrri7U75jOmTqBA67mNWtczX7Xn/oJk5jx2IKbor3Ks6kR
zLJdHUYXG8mQUhqMo1APqsLULWFB2atrlKMLay41I5V7PZ/Lumqs8jpcCcHO+AE4
BirGXP586feW/jDD3KRDO/17GxNAjCaYQmYy9g6rsryVLiP7TTDUXZfadg+myOV1
jRoDx5qwvx/D76f13EDP6HjP82wjgy59UBO9hAwWSAWaAzxyV6rNXJ93iHjD/AXp
GJW81U2sEZ73oys6eNLvTralPOg14iBW4Ld8gZUUMtPTNFRDzLCPFFDzLrdH50bG
uD1SRL1pIXa6IE2UssrueKJ+Hy6j2TcmSZHAxUCkirRj+e5ZZMmZD0d2A+5mXhoO
vLyUnqvEOajEW65YUmZYbLJKGZ7Nuq9n8Aa0OWflT08DorLyjWm1479iDNxFyiFf
FcuXE8hKCTfqObAG+f1jSGExdBFr1IMSCAaVqUzDSYv4mzpL6eiXpbS8BISZWalP
YeebSsSI+VGtalRr0bHzLxSwKK6JJuNyVldVu4R1xt2ibGZHtd6hrFZIC9Dd5MgH
NH3ISx+o/LtcNr3A6X1RCtDTuCnPJx6FV9TJQ8oAgQo1zWGV+oMHaN1E9M1lnv9h
4biRvoYXLl6mcEuVig1NI/pVROST9nuwJhsdTnYUl1F0s0Tbxs95dIxsl2MNIf1P
YGp0K3R5Gnd99z0Iqc4xLHQIO66C3VauTrXCUaXS5kqIivp5DzCxflEBUDeeB1S+
B5MVQmF/zW+w7GTrEddCJgwXdB3ubSwLGMxUQTZtwV5Dm3DSBDkD2fO0wg0KVkWR
NAXr82QapfNo+RzTEZEFlhhUhoV/kIh0xmIJnKyGzFVGtYIfMRgT2oqlP1f33rMx
9GnXrbCp1n33ykEBXcAVn3c6hMTPkGsw8wGoTe0Ht00/usa2sqyhAF6d9Bn2tDhZ
0C2m9UcbVSNBU5tGusrqw2pAFlLViwPMk2g6lS9So6M9fHZX8qzCoD+TAy7yxuGd
uutj6jHyeV1KJAgjiGd5V2uabYU5X2SZpLfl65Bq1CKsmnthjre1ov3Prez3Jy+2
0KYZ0SLZ7KDKXVil5bMv0V4B3j6ww8l2tboIVaXTMaXcaBVEK8Ofp5NqBQ3uupEv
ZTciQD9ZEmFGJvNVghc0VblarNaXW010VPOGLriLjguhlDScSGURgcQ2wdO5BW49
SnDR4DSmJ8Yjs3uqTsv/RmriWNI/4VpYyn41ijQZQf2Lzcjl4wv00r63/nbZ3U63
w+l28LD2FDkt8anNx0mzfdb50yTRbKla5TvRUryzXMKnx87BbyoT2N06KVg9aIbM
j8ayPcxgs7CccigFOnS2AB/Z4q0WBDoe3PkT7VyNu7aBVqd56PiKLmq8BUrfX0df
QFIqYcLeFWuCYzDX0htDaLFc9uUMEGCeae3fJmZxwJuJK3My47mY2Q5aVcBZIl++
n4acxCmHyvZ08OfJlpmyt5i2vD1m+0lVmr4iC59RqfcGLSw95t/HAafFdEt8lGu6
YnRAnUTysDXgfI1In6g/vr0u6rgHCkQDDu8lxXNLUsd8EcfstI9QmI1jdC/V1Vj6
/b4nbhJqlLxkJwntNSDrbrOdpsht1FYF1UxVhtx/oil+gsnutix3vYCQFOrg5eQ4
KtPg8nE1xH5XGUjjH1a/5cRbBfrmm5q6zhDOq3Gjdin0RRFkSYo+gRlh7aaagBEh
gJLJqK1d+Qo4jQn/x60Boo3cZx3zzGPcywJLRiRjU4epY4hC7/NACDaa2EJc6uZx
rkbeT3X8iOpNsOf1H7rxX1bhGaOHWujr86AwIInuwlp6f6NiU2tW6PSVHXyrR637
LnPA+ohSacYz7+3NqnbycvjEvK33AHqPiQH1NJQPNdDq1TI26Kpr4R/AUQabG2CC
iu2i4FKQ/yKkYEMoWFN5laF0G2TspPHNBdgXq4jKnoSzyluZR4puCJ2/2Poea1LE
ZqAapxgMAocmcMGQWIQRFVRH9yaKHCfj6G6SlfIrARzibgcjuTrQZ9xpQi+fhTSv
aIQFbugmtLqROO+SIGuNjt0eS9w9rv+3xYlVu/G3VucMBUNaoU8HXoSQck/yLUZw
Eg2dQJLxDTCUGZDGmC2pg5516PISz3uhZavP+w0pDZ2ZbkS0jNM8sxBIECUtag+4
MiaRlUJvkYxoCYWA0KWF8mEpe8pwKoZ1cDmaNZO02qgceeD4OEtNpGSebyPRXClx
Dsw3/JTZ5jnxTL3RNHT7MxwDc0bQtM9P7BKn/MuATBqZoY/M+3/wTIC+rjWzCqTk
WdwLLrQDNrMFvmIGoiGh3aBNAUGyZz/8Zp8EmSaHFVIlMcXL53W2ho7ggqFw1ic5
NErxGACuuJ77LEoRK9KXz1ablTl2xA7fBBF6r7ikbEZFtPDm7XLtJarTyTn8dQVc
/xFnQHYhMxpxpZBL9IcbN5dDkP98xtTP+Y600o3k3bqiX4wZ3bGNRpeAFkPwIMP8
lqTE+ad5NDrjSbOu6XjM+Lpa/k3Jbmh0lpUCj65rKqIngRGb7xKbhP1fq385sIIy
y2IeoJlBeuFgL0pMRR8zKLSb+HkVq8kzXWI5DqfFH+9DZBxMC5lwptUQMoYo5TDZ
znOqwTsy5F+wLyg6U9hSz1cORIq0i6iuLt2QXWOnFSXvDR5M7yeMfxIaJJk5YO4z
QQZC0tVVMaH18qDAT21oFUVOPpx6EiQ9bVXKtY5Wulvig+NVywQ8+VmxGd8VI7gA
w9SP8UynC657quzjY4uIwML7qMyWbnQEAMulS1ILZYQWzQvmtYywy+ZeIV2vfa66
RzUgsrnly+lmUYf2SA7NVinGrlw60jwpjE9FboM9mUMQK98nMtofN8Ja+fscUHFB
vxwyS7q/cSkR27fiT/tSYqF03Zry3HcnDZ28d1PpZORmKy/3uMTVtaJUvoFWELQn
cRJffhQlTk1TI71vnDvqd58vmBhVRkyJVpGFGsuWCgKc1AqEElZqGP4XZllWnZVl
SwC03OoaoMjyEN0ZmA4eVMz4Fubfk+V1RfF/RZJhgGI/k5P6jANNKdeSJZA1vaRd
TTJNi4kgv4Ong9KlzGN6ZtPyOkLuBkr54e4H39XWGlFiWfIYegQwPZ4MkxUbUTkw
Q4o9vSZVKejfxg1SSYO2Lz7gncIKP8WIXwW3uG+FsQB0eHC5Kn5MTAyaWEN49Owr
4INmD81nVHSb4iYnvviDEUclV7TvDr6SVd80ObhdJFLdTtx7OHOvy/5J4FnkSSQh
EqYiF0SQdSoCsvYolpxIS76kH9IO8lGgp8ZC2puPwzSkZ1iwzmlXOp0amCks/xrq
oiew7U2/dF0+Gp/stDq42C3dYI9y5avOXSMiRodTNRONZ3IO1HK8wNSd+EJhxEDa
dupgAuivNZNS/dgXKOkiDTlK/oESKnv+lr4zz+LUv8YuMILcqZi2uRKMXGQvS59r
+RjgBUMdhq8uzMViwul7jfu3Sd6EKdI52VQiUO/EkKaR++PLG7OolTkEBitVgRHZ
a5cLwSGcGt02ZUj08HZFEsG4WgjleqUEUsoYK/mt+flJxksxBm9fLHCBv9aE+bgR
SA2Umvgm3MK5gQ5gpmBH0r6YugmC1Z6pEhv66dq8/Yc9EUucfJoWYfn2Sm7ua5NE
jOoDz5ne2bJU+Q1VihX5i/I04mPjZ+SI27zMNI4xERR3baBe8AJFCUDEQ2AEed3n
8EqbyZ+zCOGIMtn6bwNtaUlqOpzlK5KuaLVCC0oQ/LznpB/8m0JyxmAOYa8Z1iT5
5DMZkhMZDKzDmUCPXvPy4PpGrBapOGO8G1Wh4LD1p18rslaH0Q76ugwrUajSJwKH
fTZMn9kifBqFpEiedmIcLCOLHCRn4Cu46qu9a3Mxhq2j8gv0SWjmHXVCEwmHZAuq
OQ+eOHS+vYL4jNM3lba7CsNwx7IVD5lbxWNhcPVV6Lmo7kM099NV7zg3KiC5AqZx
e7wDOANQq/XMM5gGZW9pql3/s23799N/mDIBltG8kTezmpdVsWDdinFLGuIVvKdx
8rfZb5YE/AaNoqwjlhXqa7yhf7/AHjwXSW8FQWbeLRpX1xhYuXKZll3x07JNR6gP
CR5pkrVO803bG8TSbJaSPQ6u4Ne+KqFW3QdcHy5lpUXN56TgVKDK+N+RE881c0bO
GGUg0FM0mysWZ6Tp/oW4EvLXXFE7XsuYYBrXGfn62ciT39WnMJuQKl6fQkfatNJK
AZD+CYR/sBHn4eYnj+GIRJlx7ItNcJ5aOQCSenF/TGE/My43pi9ihw85asIPxZda
6LnvsTMoEmtnhB7r+1N45sG3XerrJA9fxwQk7YJAZfebm5Dol/ari/cAlXHp+7j7
sOsFwwOmnL3Qs6uRe9hWZHQUzBvPh+f7bS2fSZ1ZZ18A/4qpoYtEA6h7vX0Pbb8M
TyOP0toxL7/8oGN2yICTaVlNClaM20zPDGpKnmsgtZdUpmQsQif+E2wwxOABTp6O
uyk2sXZm5VuZZ5hbTTeI4xTQ8nqePOoYbWSRh4qETUgBoEaJNDLjBV5gpImsAblU
5hUoWxx5JvmVMQ6NT+Vp/oo0llYuCjkKhBNZx6NKgFyRRy42lh0yv02FxfTCt2Y0
xjo220EudTxvqLlvh6MeZ1OIUJ1EoVqhDknOGqEoXjcSCJl9U9LHH/WZ4C/5tRbR
O3vhKspFyfSkPu9AdPXvDXfkLzLJxZVn8Oo5s0iQs1sBSOf9hje//uALK7Rqi3MK
FmC8Q9o1dyq31hIdydRdOLRqbIcpwzaQVR9Pz9WGs5ZZb2pkfePlWucQbTXFKZ9l
10SbjV2mwEWQqWMgBDOCZPiB0QYzXXX/U3wrl4Fq2WNjOIBUCIfVTgSXN9L3ev7L
9WvEoT7apYktMzvQ42YU0mgIjjq2GDp+cwWytLnCxB4WgevLL1WdoUyOUSGtyQeW
xxoxitEaAtx5wMmzKy5TPzhhVQwvzVhZEkhifgS54FvG+o5FzULDEoBY6EonUpud
bpaTzEEFaTG4YWLdy1e06H8xRslBFigotAvzyHXLqk5nezaWK/8CcVtGvkV7tYgW
74J55TasiP6TMsOXWga2c4IZvcn5rF1WNmsTqftADZ1a4q9LEL4bgxbRl45GMG4u
Xqt3n3LGNil2G/MRxwbx27KolVKSzScZ7deQ/AKVKN41ZX8BjhRsBjLnYNZMglSL
4xAE63Kk+eJJ4K8VFInWOAx9Ki7b7H91H1CkuM59UlFr6ysntaCKKwzcgWH8tNy0
0JrRI3oUfHdguViVIgsBavKSbp6BVC4oNp+j7Kt6LRfIRH7PMX/wCRJfUgzGnAnx
qAAsCfN1mRqfiNSNDqaELP8uc/SgqrzZZDDUgEGlJEQj+oeD+iLBqyFwPSeeex+A
Hveu5JjLh2nAfvlCHhlwRfqfjuImXNUwkkFVKspyk4tUluPpiT+uuNenm/ufLZ/Z
RuZJdWxzeu9Q0cigpxIJRGXylo/ULba9jpFPoAkrjjZEbno1TZxC8eOyy1+AR6+D
CN1jlY0RyGMsuTvd2X53gALwXjEg/A57NMKERWqMO0vKCfXmIjw8jghyPJc+7gt0
iq5KTam20JP5Va1sFQbmCTi9UeOeOHvQs7xsKO7/qlGXyi4BirUX8m/H7qeMkyFr
3CMwNb3rM5VBbbeuGc1LKTzqbfjFiBtkhczvNhcduEKkgVWKJq2EYHF55XwcAyzs
bk9R4OFuKx4VwJ8qLXGLoNhrX59aY0ejU+M60wxxup6x3DrEPviu/4TlQy+4ue1W
evjZ3DKq9lZJqRjM/N3q09c5bZw0slIemwsRTY1fScicai8aZ7osWWgNeT0XhYO9
Zsg8haPjXh6qW3Gy4SHaN6xoJo2VujCRDFIuSZz4Z6YbPUw2bilPf4znb4kW4Uic
Z7Y8q5cm+9+D8h4ITeNGy94xAl4Vx6VLJEEOhzTHSajfIIN06PMKgzUgTp+46Pdt
YRuUjKsYgoQT1AGV9hGSB9qgEHT2xcoVbrh3u6DWxf/p2xpkO8rP5N8Torlu48ZP
xcdsmOVZia3UW0ttNpZecl9fsxthb8at0j65Um5i6UdE9D1DPR9UfHKlqJ62AFIx
MWJ6AMzC8rwblwQ7xzovxw7b+CoID2Si2xpyNcoT1hj/1pAqOhztA2puesUhNITx
4Anf6NrwhrkKVTJgfnWr8wj+3tQbJk7MZ9/5A/Dmqzrtdzp34f/W+H0Z/ogstd7y
vxtccRFYu8eBS2TVYaRBx4+IRQjt08+kRBOx1t2D1jS9JMlDSrcqclwXcAyOLijY
WtQ6VCDtNQTItpTwECPrbUMPlkm/mEy2JRHr0mY0Km6/cgHi1ztHzlB8lJ0eQ8eA
E/qY7iwB40wgqHCN3oSVZ6WA+yci2DLGyzcPkYWBiIU+RzIruH9mcnH0tUjUTcdB
FdnsjezOmWxWGTAsgKC7G7qwBd3Y6b6LixBbOS0bb2ohAKTqvE8G4sBV/H9ZS2Dg
Pr528U6I/vj/Me12uc2VocECLnHH7thNSgbsvWePyVULWtfbRB+zQZlUFXnhKOIf
NqHMKPKieis9wBfFX3lG1moQ8tRQbnQFGeaWuV4e+CBy3eq8QHTD+eQbThprtDxw
qfIIeJmUZxjzedLJlLQU7aTFN2VUfDnUNh+K1+lftP5SXfLknPKA+NdXcaNdYcbG
QYFTyj7BMj1uFTayWAH2rq5uJhEnNq8O3gCPJJz6jXT//42jRnx6MZ6H7muxZObz
Zo8fYyj9+LJgs8m/pqnaMCxQzrwIIaT8TYA94tim1OS/Xylozib9dJPgVkGvbJDv
48y+yOGxmywfwMP11yEOs+6qWrywybQC2KcSfw9xTYb1ss8ELcb6KURNPkDC761N
brTmxYPi7zyDmU1xHSvwA2WMhW2h8cz9eKwPnu7875UNW2x6LCRlAJovcv980whc
Dv0YYp2C13Yr0VgiDnjbYKYHlz5MT/V6F1QgGzpJIDFfWSUczSKYXbjivyGhNGhD
nLA8Y99KRnm5far2RlyJtMmWLJqWu8000W9K32a8jCsTKHmsQtbTg8JOybTn9Roc
j5EBVCHdbpgELO9B5vIs8Mv7lEB79sX5pFTE5+WeNO+DSycCfYiuCoopgA3EcQhM
yGOrSliKm4d2sZOXnY4ulErn0oQ2CIQyHJNhRMx0j+IFThpzPJaGvigHNAp4tjoU
HT8JKP2ZJY69RPOqT6/mA/7WUwVxAtEBkqtx43XO4dT3bnrJ//9wuSp8eGszbZlB
vNa1Pbwj2VhIJMh/C2s+pc3RXas/I5/OmXJ4gF9/nTM9aDpAhjWeV10gse415Q6k
LGHsdhCZgVfZGOBKgls3V34QmJbfoAKqB7tjAjteYa/ljduy9YkQh3n6/FjCRuOf
Rh+/3UZgJJJVHTPYlfhQw2q5MuY1RLxH5b8fktLRHQKfJFtQi8UXgXH0jkY8CLL/
pqKyt2lOkvDqmy78jbh9nG706bxwE7VC04F+vsZqAazSQzltxs2RvETb5Oveb/GL
BPLEjCtFh5PI56QHtrZkFzAU+gLANtLVRB01FcILUfM6wo96cBYxhAuFzl5TJSK3
uGFCaVzGuQvlUH0raUFKRyVZxhc6YZvnoJ53xorYZWHex+yHTZxsEazG0yM0+YRS
P0tUloWe1zGKwxzHq0F9Z6nYQ4UWwx8rgg3udPhbTyKKxcYM6O6FNLOngINWNhVl
busSX/YWZBJWmFZBRMxnVSedjn7obGr796/FQtPmBnH/S+W/WnBWCy5hDu9Dic43
ujpI3nJCiHaQIkSaB/sMKYezYnJQijttWvX+YA+Vjcnc7u0Do2AgPctmlbbLjSd+
Q9vDXE/k5w6XbG6FCtjNz/F2R7exp9dEFwFQdYXOQKfnaXT31z06b9oszaCTzuXI
xQ2MYzDKTBYWIuSiaiF19vY+N/P5PeXSV8sf8aRU53zpGY8YmEmA0kYoG7eDFO7s
tp3pMVIulXOYeWzZqK36b5ElP3ksYLSWUXxWU5M3TweUw4HwYIEREKNG1Nq2Lc7J
7M+zEWYBjT/iwh1PDT9bZA/U3lNIwuMf5Mrp5jejpgJKs5hWJI1v6SS8x+BY2+fk
s0YraDSJkKFg5sf8TOBPaDKI3cpim7xT9Y0R4iRrZjH0PCDE+s4EsjLmlpKsFw3N
RynId2OTaapoaioYHVP3zdYxTc99xrGUA1pl82noZHFO8ITJ4WkR59yj6JMMUisl
2YkanQ0WgHI5hrznshLLm+Hc04lRWTBV6tqgq8zmG0kSm/FYm7Hhah+ShYuV0YJn
7PlqzZloo3yEiMjuV5L8SYxFrhXuDDNDCYnlqP+ma9LfLgEZCLKIstaRXkk6HlNV
mAQtvWveFmqmTOrL9YEAlICXqfZcbN4NyXXmvOWdQ6T1TXr4b9SWEIX630EpZnog
YJ8dxxh41Eiq6BsEWqrnzSU8F3d0XCCqIN6x2wQsDkmJbSrIZow3FPh3i728EO5E
/GS+gNr6KTZC0nUjWkbc5ZXSBbMQCgjKxa/ICZ/a6ikZTE5K3j1OfpJI33aEJDTT
tuMkvq1FKR6WJ9D5qXc//mChWp75nX7r0Ppy4LgJiHsajPpikQy7GXSC20DuyVYn
TzK/bnf9xRrQny/myp7bbZTS8JXI+0i92AY4EblzKnuST1TjiyoCrtytiBA90t5m
XYGYuSGz1liH9pq0NQeDQZ978sTs9VxsP3Ml8GuniVBZjye5X6RXt9+D6Fdedawu
yXfT1bu4H8MZoSZBNawzkhhbKB9Fr2YFqIQup57PP8StYLXm1tSMWBVV2kakMkts
ellhoOBBTvlfA/NW1EajDFcurMpwV0Qo+88GC2bqCHZghTP+uch6hX3D2rtMFm0Q
ZOjxn/mPNJBHZ098niXRwsoSb4b1cSAq8Oy+x9oWHIwunmlcU+E1gvwl99Q9u/C8
92/6s1mzJnpeVHJTCksXMA76I2mI7hO04SLkQSR+ToBliFzMGrgPeyzHyerM/Co+
spbttUNgcIWUZqdSSElyFlhWO9r1V3uWtnnAegUwHtEQj1iJgucY5nmUos1mZmZ4
GgmtNwvwoOUgMgTkXW/yHjI2alrlWeQ0jVQYZf97yAq+G24WG7q4kGZTcD3nV0NF
v08mHubKHZ5qDMEXh8u4aRMgfKIJmb5IedIIATaZvTlFTBfMiFxHQYBi19Pb1H73
XfuUamsYG4P5UCS0N4S0hmqbBK7du/L7NqTDThSj3XzZV0yH5x/1sZmlvQpsRzDX
VaKtm/sWtA4tWpmrZst1Dl3ElaajeHwLfQiBjPtF1ppW9HAqByi7oHQDheQuD3ob
T/uPlC4sRsE4SVV3wzm3HUL/9QHoaVIFV1SsL6pNE9xW9FhgFeBeJ+RH359MP8Qv
A95ccHQZFJjnzfuOn+T8L9t71u/3w6l3uC2fP/5alfqLaJTNSgH2f/B5t5h6WBhK
uSq2C+5a6HzJMmG7qE6YZ69h72xlHljzqps7SCW+75YzfGjDp4ifl1BpDItPnyTQ
O2Lx8iN1r9AlPww88awHMpllbtwGtRV4lm9Bo9OcDn9tdU2nbFgqE1W/cXwSS9iG
HuDclYdLEjY/znLyLdDohDWW2ZP9/qJkgIHHLwA0NH1GegdOZgvwLXpCqzcWGtrD
Qo1Am02PSX92rCrUqiCHcjQh33EfGvJkS9j+yGXCzYXafLC024npOTuxACUveLRK
Yup/oSkynIewp/NDKkI4mvBSLpegsJR98KQVSnJZJqgTzCN3ICptu3rDuky8dZEh
oZJ33Q4bcz7SZxlIJZiw5z8youYd/K2l1pZ7WWm9AvSNTbaIMLBWrnHsYipHgUl9
W8y4s47gigSCN2swXmWDPXUmSY25XioQnkjID0FhJ8lP6hhLGnvr0ZjLIHoPRqvW
1cBalTWuXZvrpxGzhfvyX9WlU2xMsQ6VPO7i3ei99qEe9hjklVAcc75fknhRa31T
jyd4mYye5VCluT7JeCfwSMpTElSjLt1Go+7nAO5+kg1yricObkYeGAwBe064yXvQ
oeQFoc9R9+qbVL3jJzyB3kcwW1FkmohGpEc/ehNxAjd2+rm4CWLun6hYU1XPfCYB
y00OoLUPnryeale/LeAW32C/8QyW3oUH0IxSJKnajNc3zkHDbHZLohN2ejuUAXol
OWGFnNAIvgrD7Ygo5MMOsbJWfXVCPpkBRSsWT/4M7NBYZHySQH90mNMzFO2gzgd1
Nd2f8dQOxm9yHd9goQ2gRaQ0TrY4lFPGeOsdyCMaVyZ7DqU4/PB2dmIgjNQQHTiH
pLH/AyRv3GDawZvOlI1ZdY35TkzHz4NBRl6WVXmOEdMl7LNxppas8TTxjEHP4gZS
2gWBjAPeHt95As87JPPwXnShpEOysa3W1hrae/lRH6yG9+toMGO9gWAbaaj+0Yiv
Y/3WZ8/Plu506kHttuVAR0kCXhDk9xX/oE47oyzmFv1h8KKpc9KS58LMataBbXcx
QbI8hsLFbmihQf2r8n84HpIqeUw4OuFEh4U7iP0mqoYML4uDIbHQmK8++yYdN1ZQ
JV6gnl9cJvt7Hdi+UbATNCdzp37W4boRrs/WujCxFmbB/BFJjWSSbT6P5AqvXhYi
YT8aAyWGLGLMAdf7Nhu4eelt03jskKFk2oIxaa8m3ETmQl61vYVCHQ0PQrvK350C
5q7NR/Ms02uzj1JvzBzdstsJM5Zz+RBKGHgyiy0TlLmAOatRIXOLJDH5OWvdQkCv
Zs0amhfEugeY8qRr8+FgD+WiKAAvZV9Lw64r3ilozJupsjIJJQCEYDCMngVDgPz2
LoZFU3+X2m4lb+a8ju1jHXZ2C+5rhPePKeX6ob1sT87RnYNt/t861UCOH9oGAbrv
z+Z/+TJWUNtkUT5fX2Bvt2HxfGn7LGvsown+GJ2eVBUd7S8v/ELaIFXUYXA09vxc
SjQVNGJIkzVV5C8uO66E6rRV/P/I60zqBurzhgUqeP0LQoJdQnt5t9sQ1MLBFYUm
g0EJ3E35InmMAHwaa0uLEFw134nmtPhsgEqnwYKOUyBdvsF4cM5JR4AswrqDur/0
aCXsMtW/HqLnqeqrcU5SFQ6r6WGoD5wNPo+T182TnGcEOz4txOboWoKHJ2D6LDz7
6HIN+eNh9eTKHxaLIkessM/giPDiUvAnwaBN7WhY8Afd/QwysCF/OXdWS0eY9DYq
ArrbXzMyaPnGNeCpL97wyyc5wpV+SeiZAgL+U8lac6cBsCI88y/P7dtuvsFqvH/m
1lColKROHdKuQZ12gw7FlEpCASg+yh4S6Ex5VFVB9x5sbK3wJ/L/APUlvcERnVYJ
9NeR3kYxdRIoshv+E7ShvXDXgQCvS+gtIoLcyWfKXGO0DfQXUiw4XYm2FWkyOJRO
EnKFi1QRs/zYflX8zFFk24cJIxES+RZcyqpC6Ny5DoOLYWo+I1ttO2Mke0DzDaCq
iHtoHrlP8QnHv/vyLIj12SV+VMCCjotfBf8gmYZTi8jKQg3Hc+mDCi6F8iL6ESDW
SYBiQsqsHp0Tu9EpXgR5ICglrq6GKq6qjt/xif5S07Nd/E55BSQZh5wQExGOmXj+
Rfvy62uYw4Cre5TYgyjuWFs5OVBeG+xYJ2JQngExGAYr73QVFOlkLxknUtnUht+c
HHuNX1Lqy7ZxlMkfLZ9gTIhWBjXE7zrG19tPbQstQ5vKzJ5lUQTSvGICHwbGpCil
H+6rsT6QeHHYkCH8TZkzriDRt3q09zEWWzJdYqa0JU78NbwifX6I+7pnPdpC8n4U
vIjZRG2ZO3jeCQFSJRzp32aj456Rilh8fXt0kWig1/zNQAeuqMDKwL3Tql4g0PuA
2fgWKUS9WPN1iqNtWh58uaD2LNGSWYYVWMqwjIvx5cV9qJ7XdLFWmB78fGGCd9Xr
zTOtVipaTyryN/iq7AM1TEsmFbNi2NiaCRMMHpZjbacFbfsMgX25Lge+R61NcapQ
jQckvNG3XCOS6iTY2/rXQP7tSGyEoyLX25RNxOBgWs6USuwG1I22Q30sW8UdX4Aj
ekiYhjD9hWEJmbrKbZxTMgIWv+oNtVmKfI4GZtrTF5JNieDMd0EP1Dxs9CuIBM9D
EmUnUA1E1zk2rbpAnUfPTEEoGFcbufGFLO+jOtOcjsQsbuOQaVKONA75uEC9qZW6
veRtt7vZbEOldYY02e+ufVUifrLXZcZNreRAqdIX4YEvzREb54UZSKPVLrwpJ/Vc
/4Byx60JCiAR8J0Dbh5XgnvDOVWDZVP5hF/gXFtt8otKJSp8633njJOKsInQ7s/a
+TlQOy6Gw4yvIMdQxmxeDoPtupgUfs8pslLlIVIV+/YS8dnxiKrAbcVR12kYqILB
JCXHp+a70AOGl+PErkBWOBdbZyItKAH1CT0kRJKmXNWM4tqvSLZ4RIjBFkQZJt2H
1X3BByaH2+E0O3/EhKqjpvY8a6PwXQAbl33qiTQy1wViKgYwiOYaxER0UbCD63x0
zGP2SMcFnGrDcnbyF46v6FEWLAScr9/uGR+62bYW2igNfKfZrEd05zzEU6F2+1QB
Kw5CE4tWfreJ/Uxrznm7fLaZp2pbK2+b4BLZK0TE5C6aQED47NSLMZylp2eelcKw
0aexeLK4EOu5otKOcWkaEQ5+vEYvwzbzUMer+EVkD/ma0SPy0nMJagsHeEM9dlT+
sT2Xdb+YfmUADmKeRP4iqiP7Ob4UWjf4EiQFMD6kRt7oUL9SCIJXos5QGrzSUML+
iHplbq/cStp3ZL8Kdj2BefmernYZWXC4IZgm3sEK5mpYcvF7eM+l+PdBNyVqT8ns
5BaHYQdFGZSQC6D7dovp6xdr8Fx2cRImlMMGZM+A7GGRQ5N+MvahnZ2k6raoYSnr
PHz1bhU0CUsUaOXAk58qvRnvmiwkxtmDN+3ONusQrvVFui53QXrtub8tQSP1YP11
cJhN+dNXD7CKwsF9vyTjtM7GtZbvhJEarMbHuFfwkuGN0AwsCtmD3bs60CKiJ+Lx
DuSZB5NHcwwL/31dc8YSj4K2Y0IXblttiXvTTgTsfgbrrNJY8V79SuV66BL4fYmM
EP6Cn733mmz+rG8D90f/pCsBnzIugpg92AnWj3BdAGzGiQSavBwO37dSEegc1I0r
ukGCXeim3NoJQDdFV17HX8jjQKauFEEt7LuJZuf4AiWdfa3OU7UYrmPIegAkA+4A
OnOlaw73WcQgdE7nuZzH1GUlDdm9FcR97/M/SMitf0ptg4u7VlLK1TAGjzFVPKdz
BpZJXgMFmYSG/7ldbI7TnTcRK+SvVoXByBn305e+mcJUOuumdqKAbXP9iI5J64n2
l/7Jj55UFKBIqqKLDtrvpSkGyCmK0LOtlhNzbe0zVLrVvjoQYl3eN5qRYNFHntAz
2KRrf6YYQ/mn9sHaSvlVHRAt2Aw6+czE2ollKsUqIhFecfV4XuBYZcprNQAEy4ve
G7WCVcSyAdik7+J+H6C1UauBnMyufFe6hj7X2YYNwF+2y8DcQuw/+SBiASPlHSvt
nN/K9F9c1j2oTWOgTXOHn0OOnBLIXEhIHnpSGNcInM0nJlcce3Cy1GeSXNlv6pMe
Cv67HcuEaYTSJuxx8UeYnKSTZODrSpEK1ITLWb+uHEMJt0+jKsxOQ6uOMyd1r76v
EHbRQq7faPgcrC0dDQrN5lUsWN2b0wAlRnj94ZYDtjOAlQE2M4PMvyulggIGECSq
Tto5udM9NM+kHlBWqGyJ88cCBD7lEtmqnM6RKDSZo+8zVvu6Gp59xfqrRhewPuBv
0jZdDK7gLGE6OSwf03aIXjb75duTKkpaLSRX+Zp19dqdmt33UfioYV3OewBBMOfE
GVwLbcinCXtoevHUkPK74nrFk3GRx/RYprkZA5c81qlJd2k1TnCgKmzgJ78rv54b
IdoDOE/xvtQqtEn67yACgD8uYr2Dgc4jqqHXB97wYOe+iFDp6VcXyRdky6EdMEbp
MUSMMEgFEX+eifsVLyk42BVdhzcxosi47zzJvUgL3JWwj6zNaMS6s6vwLtedhDS/
8enrRvskJ/JgXox1k7hrCKBbQHg3qIKZXsEj0/fVh4KzzB1balngvxMS+Khpqn9Q
Y2TqwAJ0WrcmQMZ5uAzKj/YwdUqCg7icpSEwCfsHLX/Pmfm1zFCvfeUvpzjGOlk9
aUwSGIhjjQOPIiYuUP4F542klhdPZ5tsFYf/8Tw6M5oZH3CVP5xndu8D0l7w2Oht
aBV5h6RbC7yOoL70tGGPj8wgMHEo35wYMQD5vAGCMDaRLIk6A/izXvuOegF+PYDr
I4Wn8qosSI9v9Ajc7872I9Ifg4TzadNKACcgUshUqBzYvHlzxq1x/KfvgCrRq3nB
8OkWVl5n0alr+qeFoejHfkw5A5VvTgwwB/SjEGq1/+UYHTC4QH9TFNwkmO6ymPRZ
j+imSKO2R7Jxj7E32x+eygAK7Wxk4HuuMe2wzhS8uhMqgylxXPgT8jqQ2fmopzmd
zB+5xLDHVpdqiwPPSIeIYKWs5fsE8cZH9s/w5tID+dZlYvhtOjS1QAot8iI3uhHn
zpPDGVh+CvwhrNDxTDS0MbfWYOw82/C+1RuUiF/AczrrktghDohCiZs5IuuqHrSg
+mhcebUjytvWeqzrQK8jUl9rTRBC2BH4rLjF3TFI+3rtL8e1iHD2r6Ed8LqaoMZK
iAHGSXJHGHD6l7/RXWsjK8KuLMChcplFoTUAaIwg2IxiN1tVGhYZd7D0TJ056nwd
Ddc5AH7BdWy8xjIZcAoHlQOuk7TixgphGY1PwcFke9hNQVRlxr0st+18ZncJyrkE
Bdmlu49j3tCq0rAYqY0fW66101mcUZklRM1ggqz4/8wbIsesOxf6QRiXDlicAOLK
5xYr9v0FuA1MNtqQGGqtT8udXmZxh6u45Y3UHORiKTRAII4PYZS9YEidOo5XxUTS
bZ+tueRNms4KSZAxcm97X7t4ZsjLfHJBoniHg3T/H2SRm4xOJTyLP+li41I2W4Hm
1KqQ9gw47NbgqNmpbG0O4kkpiBZgq3GbxLS1OmuzYnBArJk4bC20LwaN04V2Ispl
dVgIqaGuYz1oc3F9j7vjI1F94gB+DT/IuLLyS+uCkhgHA/8r0pQhNj+zmjy/mmxR
3TAhkZ2BzILWuNDKGbO2qOEe4XzcizwlruPtzeAEhvptxpwUE6KFxrll3Yji8jeB
Gfmo2o2fuOkvL3leyTLjGEUBQOftZy3r2sTk2BUouv6MKVIu0aAbJwvfnEbm3Yii
/eHdQHDPUOPA/3hxIQMc5Vh5mhzDcsdNMv5vDFHAVkhOsNPgYhYayubYl5JzycG2
DQO4gG3WpZxEdyZLEY+FKZP1Zvmk/jaGRq5izjJl5rv8IA2PWbZQgar6aBG6N7k1
7pbZxoQg1Dx7mjxm8eAhtA0ZFP0tbJNOGu1CVoX6CROXqpylsrihifTymSrypnC6
gGzEGi4l71ran2gpGL0xGk9hWM9Wg3rJllzhP5/Agodrfiu87RyF4U6sIJ2d0cKd
OQFcOsy9Oq8Ed0y3BGjyZ20rmCg/+5aS2vJ4Jlecd1zuf3VY38dP+cilrLOozREX
0XUr3XxQqHb2yYmPIyyheUAFcB8gRtBYWXWFsSS5u2CxbwBhCHe3cLZuX5BOhVHp
UkgvDsj7qNEtS1Vj3SK4Tlvt9RP/BO017xyQWZxOzX/o0edRRZ3LJlRP2ojCepJE
cLF/8UT024iLEEX9wvDPXaGOpPBBF3U2w8g+heASl2qK+5oQV3DQS51+p1Ri5GPZ
WE77k1ze9/rLm/U7VG9Q6JSgO7yDomiNPaGbRVyvnxoYByf6BvyYJQ9yoKkBsIQy
8xZv5fKqguQ++l1Tkl1UxfDAJxlM4QQ3sutmP5jXsXTYP3AWnshVF4xyfe0NjNJG
iUZRlPNd1eiFY9PvgyhzwgobZhYk2WVlHWC4g2ulmdRQtzibN5yxq4cMp0/RCXpM
WposVcuGRl8oeht3sV9aqHJtpFRME/1/pzqunNJTy04e6lpygPT968Ku+q7Ly/SA
NAVLL6B5V+2JxBHbzlOvzjigSxWbLqHHJf9cr0bi2HbGitcM6MZasoe+4hZ8hEVf
Qdjx104CO8wLEYxSn6GmA0JVCYMEsKIujDWVFBLR3daHC9xczLZJ9xCJih4ujOMo
x4fxaccnU6s10RtJQNS67n+JhdPHGK0g1ZFvn6m1E39xU9bRJ/T7+G/ZXks4J0ur
3Vw3zeckqz2lttxOJCnst6pCET64LK4Ob9w0sGlgBCT+5VY5vwj0EZ5dvfltLec7
XgGtinnDL2fEqCZbC7Q7D06q2HXaaZM5SJaQZ++sGrAedqGRtgxoRnA4r1Hi5ylx
RYNVXcOP7p2ONvfK9JqfRZm5XMnlYo/vcyjmEZQ1qFyfyxHZZMJZ7XfIFGNQUzkd
3uXPGZ22Yu6F6PxI3L2LsxyCiFKaTpYOi10sWH1cWAXEKHPZHiYzGe0+yZ5U0FNP
ObXPKuJtyz08FIuDzhgxBaMZ71IR7+J4nmV563lIDgARmYVG0CWrhJDHVmLRrNje
o0OLD3C639W3pjF1VH8e0o5mTCJHxyXQmay9JgLk3jssPGgk+Y1lnMPYyuro1h2L
m2XudocBAq34FPP2k4IferAbUWA7lyAFPv96BtFjrIDn8rGEjfjZw5vqTwJcYmrM
QWhdwp8AOshlVwwkCxbgaiUbcH8olOMnxWM73EJhy1SrZsLBS97nfouJWnMYBmwe
iUK6TCwCMHntIde9N+MpJfDKk335+TYyTwuC688xMBsQ5Trrd4S/9UoYapTn2iYy
YUmnsD4QUw7bo9MRd4czOoedRItb6VW/ILdbCXklYTkJY4B06Gg8Tru1CnjiZ18Z
eyxv2YJz3OUKl+4HeEYjiDT0t/AdEvJcf8fsI30s6EOt9VZRjwEQ6F1qNDyhN93B
1xMrMqMFPEkDPGSH1pkt9sBbTAWNNVnF9iSnY/t4EG14o7sO10XhiKtZ0YZou61O
ipF+L4V8lHvRszLTTt/bACGPmSghkkeEA+F6GkaUoU2jDcmm0FBciouAfC+yTcRH
TKp1sVCJpTdWNx9uBn0PmMwoTpcQzVI2oYfuLTxlWcmStWnzmIreZGE8k10+OV2F
m1AoSZ5+6SG3a9XynMEQz0ed7ouFK6kATPSiia3PB+1tCCksi521qJwyn7nfV3tr
vdEH4rq1yfTz5hbQUFlJZmtxsrwirp8VLXKMrFAreI+rIsFZ90rL6sBUCJC4nxBz
XxGrMl2I3QW7wOHqQnEbX63M2OkU7WnPTC/GqUkWmwSR3o2FQdo9XrcFD6uRJ67M
5Y3Gm/ithHIk9k9p4F8IcaJdGB54ZuHjiEQsnwfxuvVhAlxtMJXa24pfcTmGoPPV
Zg4fLUQqi56a8onnALnAomeLX1bE0F/PQsck/5vZMvOET18/thMPyA+rTbiEJdbj
E+4N+8YiV4ELK+CS9BFfmB5yNYaAADzZB5ZQdciS/qou2sD9/R7iKfgetY7qEohZ
5JIxrhKBC6lv7gBL6lnq2KGmaufdcUs1fWNdH641g8uw0rZ2q2VKNDNBV7Yc8hr0
yKhJGSZSBgvRDTMPTx3w0ZcmkLMGmcWcA5OWXGEJVIVpeAtGiUrjEk8ZU1ksIYaS
hy43X7qZul7ECv1xFUWP8f/ao7BagHPzQ1veTOg5yGdP6QRF679fnisaB84VhO7T
Ywxwpj6a13oncS+8K/XyNqVYc03arY8WpxwsuFmK1ZR+3mCDD/BcSxiR80y1ZQrX
1896Qv1JXyPNAoZAckfAF3N2QqwQhVM1tJi4uvhBRvPs/qnVmgI82x/5I8M0Q8EQ
e2FHD9+SkDehd96o0grRoRp9v3OyUkz4Bw2v4uNt0e2oLQLmWu5DGGOd80a0c0Rj
AYpdYIVQxgVPI/hAEBl5gc7dXdr2Lj9v7vyqNZWklmeax5VxGFSipd7EgqhsBfgV
FeVOSgX4YayKXuoPwJjbiEGjVCY6cZypy9+WTjk0io2l9lP8ICWAUI/H3UtsydEf
J8TYoUX0x+8lJ7+GwK6+QRTuGexBjbr2OxVlYnSxdE6DAxps5Q5bzhIOJo1uH0ey
59Mu1Nno60TNnM+GvqS8iTSdHGsqkvCXNsvztqZpFafErnxzB1mQX2bF1PhZrhWs
NVZHgKNiwQNwP8ODSON+gcjwuYtqZIyNWlT+S2TRc65wdN4E12Wl0hOlNO//QSPO
vL7TjMngfF76NJiFpOKaxK2QwrjmTrMrjYX9sCww5nQRs8oc1nG/4FFymNJQY6yi
f2/R61rjPMXetxp4tSswbRzSm64oMft57T50aGCES73568ZkrL6USOReDiOemn27
k6uQdgIyjgAbdSCFUsgseCRVcKvI+kdjIxmHewojulOs+TjkZJ5OkRZ6H1981W6T
CJvy4MmGNgXLsU3elou9cyaiXV3C4aprvRWzkEtgls0YBrG80/VoI3s/oyCf3AAx
ek89LsPL7IQ2SsnbwIG9mbg3AFMl5qh9kosOAZUFfEwJWqvJ2y1LshdEta4DzShu
Kmkpve66EP2PXv76KFYDHIEn3F6f2b8QJols/myMkxpScF9+f+3TGviRj6KMG79H
5e5W9EsNdhgXv7dScJAeDILHpW0nl1tC82g7MMP23ZpvDO/7sPNm8rxjOCw4nu+A
aWwJ8WdGAVgv3OC9PkjTI5bSay675eoF/eOdGJJn6IrpHkcf0eKF6FMx93V9mKpa
pU5uRjcGbjz7YsvLZefSqDetvJCcFzVLzOXw8Rs8fzNUF4atwzj2kGy0jXzs7BF5
JLJXzpILkWK1mIyG2caVoHQNvWotrUiERYRPwePsWB/tKphq0UwVxfqhsZVdl+gT
U+vA7oNLvLOo8b6gxPeor0rYTZ+g7Ho8QwEWSHSjCm8UBIJjtJYIGR2xtowL2LId
YMCgg+a/vZ+r52gCOotgzTqlzYTQ7SuQfQA580kP6BTzM2ZJ4DDP+qUH2tPL9VOn
Nt9DVTmZPVVKWwv4msxCnm3hni7i/v9FEpirEBTaJBQUnvWQb/fz7Ds25bDiJ2wg
rDvevizoMIIhMJrq+3wVITRp2IiSPqEC8LAhD+BIgAR7/3ao6tBHymdvBEoNdLz9
B8EsyzGi4FeftdbvDb7BJUDBLgc+/rNs+9SJVluL2Fmncmx/vEnYZnL9hIIbOYZA
IlH8KLvbXhvfmLydWDVFur3CBg9kAtJHp8Ul7OOlYml/WDeVz0wGVU5yJFwQnDdj
R1R1r1C+5ha+1H0RrRdv8IyuaAcIFVwOJ+u6I3rC5ofTrM+0YnMeK+KhQZ3NzRn+
iCx7iBgJ1MCh5uOUGv4lHRGiWjrtqWRDkp6xMxWWGEnhrZNqloexvIgVUxHjUc7f
ZucX/9lBZ+e5LpK1enssqdjKNIQH04KZnUq6e+/0Usgo5FYe79lH/foBpeVXV9Q5
GHMky+rEb+FW4hnCO3avlLW2Rf10sj+0JJZ6wknOVB++Z3kNLhzls5f+d3eBcwLl
V0l7utX0OnttjHKPk568xcmxz1LbsT6pCPwQ6EHE62VpPIXd4jkljQ8bIID5X7qO
PE1rhMidOzkQU4WJIuIlS0zQ9sZSzx4n/NQJZH4mEPjgwJqk0H4FNcz0XW5Q7Cqr
PxJw1dYpxCyzDL50QrO57jHQKfp8vS0mkLy4MeOZ0HbJ/BQq8N+vI75j8uz8l3n6
5xGUk71mJViyGJOI12T1KWT5UkQZa+s7jNzH7D7OevYA5CJZP2LmTa4bGhCoYd4g
/YcT9RkJ0rNjXOxBf6iYJZnqjeRFR8qCngLXD/1WBETo/hH24OZ8bRXTGlCQAeB/
LTuel9NUlUZzPr/g+NcdAQyMQav4A1QxpE32BX0cNpMl6m3dMcn+ttW2wp/oxhqF
5YSjCMaAdpBs7kVzJVVRQsU/+ol5j2mZCjEod6aPDcQlX9cSt4P1LbaVrPsuPhIH
3DOOM9QLnU/epOVaD1oelA7GHZgOW2GDFhBlfjvYK0uPEkxmNc5hZqMFLPDJyWHo
Cx9qeGtYDHe1gcAnW1Rv9ws7aIt9rNuTD+1DfyIXnmtj7xrGUtW0jCS2RRt0IFbK
ewf6dCcicoLEqH/2WMcGI2af4vDRsU/2wFLKBujeel2EINKjVG7Tov8YS6VS1jNA
QWt254/gGnEC5ff7Yupr/fWNfzxFqeuxm1uUkF0TdEvPFKXkyb5wt1alyMlBqq0P
PiNY5biipFIsuPDsGazxrzaCN72rWKHtI77BktJOEMab6IrGMDr/Fhqn2TYbAyGQ
WaPp7e048I6KJblyUe3hyT4gH9HTQqw6WW6Fj9XNhvlGvmm600jWi8MHLwKgNDuE
EKYiBTHQHkYse6JdYn3DetuDfU3QGpQSWTUMpu4JxF9fr1Rmgq4sj0KX2RTGQeCM
nJe71PyloA7J2enCxYNqGKfK3sV9NMGQ+GuzXOafHMfvhL6Kt2wjWaMmLAv+hRmv
xCgMcyfYIWdG547FNNkXlaLDY7saOB88KUsJKWKWRZgvQQL2SYljad7SwTu+pkya
8o9V+FyqSSb00+in+8lsSCtIdlJQvjq+QRJzR6Zq1lecoaVt9FqgjOclBRaS4G8/
DtvNLQirKBQVLXnldy087EAANDkR+LgXwapT65OZY8qmHbloQ//X6Rgb8k+kqg/H
3rbwsx6V5dWdf3wQz9f4XklCuPDEI+d2LsZ0O6ycAC7unupT6cLTyUs2JsNmsR8e
hC6hoy+VfokNifLXQg/vV89waxACGZ/ErhFYVji7WfxiL8nCXdxT8tE/zQLwYt/j
uvwIgiMX8S4onzvDSLFwdtYy6hevQrfSMEvhtqhaxh4ZrWvuGqIg3hfUA4mldh0a
ObVdjQisZRCfRBudpaJEuT7yiKQ5rhVN3UNfkvRcoVvzBNVDgkA0ybgn/9o+i95o
M46cdUPdWgcxfzy6nGnl8kREwCOcb/y/nytbez4eCaENUmZmaLt0D8YflbegrL2b
hNLNbPQS6HtlPt273cx2sEChds1pWEUIWtmrkTkCwEe7DMs6kduNAjqbPSk70ENC
xxFhSBKtV0awOb+FVIyN6eGd00SGP0th6W4EWieHdR9svgSxSC03lzeyf0MDYEia
/X83LP+ewak+pU067L2zKuReyN95JCk8bL8p4g2S7I1+IURx1rruEZJYr3HH5twf
wSeEzC6G9oiJDNdhy617jtJWhXptUEk/WEZvyWbFznsumvnEBUyrAK2TvYUQoz3u
QJeVeHy5MObJ/fz7kOPoqVUkP28/TUi2uSZ9If74FmlfmaTUpbdptyWEsGsAoGFL
a5OdxdMnV4i19z6pOSUpCscVwBDYQ2es41Xu+gqYlYtl/XOLXKiJymoP+d/wMSDt
MMS+iSh5LDYw/7QQ2+qszTMJ7mNykezH2l643NSTqHL38WMuafBM5Z3qWDMFzbUG
bMax9DwqbH8U9BltvEPAG//Hto7/VFA1jyCTANUX9AlxhkxUIdruL6WP+wR6E2RC
TgJmnhj4qhmdYCb5Swfw8AERf2tmLKP9xfU5g/P+Wq5lHKlXFuYuSv2ibf+X1tgK
Nr0JcA0FUQRfXOxUvdcY9uoD+V8T4iVkOmSoVojjz9AItQnWKbutK8bGTfwVHch+
aRIkUG25YMA6BVsrLgkgHZS01rEeNDDsG3lYQjNM5acFK+I+1MD2hs7zTuxW7NIM
N7NyCAm0jQfER8QZakgi+HJiTajvbeeeHFCXSUZxbo6wX+jvclid+NIM+avE8Eg6
Quo3hFcqoMrK+ysblbiNP/Elg4xSBPkNL4MxEvyEaFVwGjcDoq5+BlnGoJY4yrlu
RADjtzPxGztrayVYOJGl+GZF4qJAnhOpT5Tw+QRnMS+KZSJ8TcCr1DmDod2Xiven
1kvB8aCT5GPOTYdZWr3//hkQwFPfA9BvFm+8xP//ImGJswCD8MSwv22btfGUcaev
Z62L3gtxoB0ZHQbtpCEIg8deA7Up063EJc/9uvyoAXA4bW+dzoztEhto0L9NSWjM
KVAi/tczB66vMA8w1ErqUFYgDgLO7mSb9n4btl2/rJBVK5lpPxEhsbQW8fxqFoQS
ut4MdQbjgg/o1Rqi3g/rMahYJjyEjkpojYd7sMW2ad/Z5k/oyKTjjU08c7PDfZRQ
0XLCZFpDKbNfN1qxL3q+4vNebYiUmkelX++p8a3aXt1ZROe1VCzNEDhzro4ahIRL
s6bIc4L+nsLhNF0QmiMjJBYspXw0HIy/FcrlzpIKLU6kONOKW+Fus6GPZukKswuh
+xYApZku4jOL6Cvl8thaBNUTw/UgkcKEBRMHmY61EQ5gOa3x9o9yP4SYyzLpVyri
3a13rLOb2dmW0bbNJ58lLEjc4IRX7x6n4OITXKBuvQJKKTIW7wYFDFe4sMy35Spp
XP6SbP0Bc+Md5zKtqqoVpBeANlD3XqFaoVT3CaHr16nVkFjeFAQlqim+aRsS/Tjo
QfPT8HMYIFa1CDqrNHU3MH/Y4KBTAW/+92N14+AsijAIU7Al7udp7NinZ4P5ioem
0MSqezgKnFK0PC9G16YfasjuDX8gh8TlXnVuJ4lgUoXRPNdl7K0YskYDYYRoUCM/
a0/gQ7hQNHOZAvOmoWfolIfpmH4K2TX3La1fzWcAzLIWKYDjdDcXAdk9U+AUVEWo
pD2ilAFl0XwbIsaUZiSXVvyqUqpEsMbO7/kIWoHqvpnNlqT7D8lWnFTDLHqr4H10
y3Lic3Dh9ZSocZN/YDMd42V7LNX+y4yix8wz6BVwxqo+caKuoFHwgEFtAq+ScP2G
E2m+09KMgb4b8D5TykVIWwWoZSEq1jqU78aQ3bPXZiLXMaOW+NE51Z0RPHil/ojz
fXM7nO6zGDjziTH+IYrVkz2SGLrVaDYiBVt208d5nmi3gDU3C5z9eP5Gk2QIEWle
o2ajc6B5NKZXcG7FzM/Sh21RY+IZs271oALKsYv4u/auG3eV3IH180YKPrWwHHBf
GsvWwyBNH2ZX/3Ua69wPO1Oarq3HylXPqYlS6LnyGxkcjsGZu3fBvTM5B1b2dF45
n8ChZrlhg5UHJJAqkCITzJvi3zZqs2nT5Zaqe4vlqY2dQv5cIjrXhx0hUUIiwkT0
gtUW1uuCGVir9O3F5M/x+sHL77lx84r0sRw/26q1aVC7dxCIVS2R0s94cdqK7eL1
3GYJGae3p9r8WnPTbhLe19WPUNuxzPK4d0AK2TTIksBtUL39GyzNrdgk1K0egUsR
Nl2bIpdeIf+DDGMC1KQtto8MGfYNiwur3w8r762itXP8Qq2XtXMMLO0+R5Kfku58
KueqED14LKYy7xLjNzV9NQ1Bb36uOUhBu0IpjESNeuOxccA4+loVLyjexwsVXgLg
w3HJjZUk7LhqPPWf7cUSbE4Jk9Qlf2T6BD0flakJ81AQ+uWxcyNKg8RiYQoAbIgy
tsAhsrh/rDUXLahyi+DIDp7hYiqjAKByl524q6m/Saup/Ih3rBihGeZy43I6322D
uJaLb5RIU3KP+c2DmcCvM5cR15qU5e3JI2CoTVirsrgYN+LlgAkG8HXD1DMgxFaa
c/65xpXCdoZxqXpG46IXEHJg0D0L/twmi0uXO0LBjZ/i9HMCplNQluwuEOs5QjmC
PaXe4GmsBLMOtWZXVH8IvQadnt4A3F5bH2B8lb2qu0wCw0oeo2bXF2ex9MahReKX
nLOcIogxoSVkSxfv+uzAmagVjimYHOuKvTsUdAn3Ac4D4c787DkBk+TKZrhTA5mX
NS9UmuzgbHcXz9yIfiNPLTsKEOMCYGWvVRq6dDVcMkw5GeI88YJ3gDNTle6ugNKA
eoRLmjIiCCPn6mPtbhS2U+joqbXxSuclHjdHgP0/2J/JYImhjL3/XdS1O81J95Xm
jMMKOuak20S65DsuCoQLUadZbg6BQMg5gUhkLiA1FN8AGFTkM3VzgyZWAWnKpMss
8I2NqK5XByHabvZtOjYM1YNukl/CcVfdDp1vxHZj86IJQBR5G2B7qhcOtBqh/TlD
KFq6Vw/hBlxhiJnmSwU/X640vDjcr1gA5IdQge7CpOZdWMZsZSo76jHB24DJpvrm
GMrcLYuA5cIkE3iT8RP8+MHfrFDCfqKxTQo51Fda8nzzJcFnFGJQ33ffYaLZfLZ7
g8Q+Sd2j+hjmIHNxFu3LpO3w34AJq0m7Wkkq7V3l3fR27ASxK3njoox1jYhSXfck
NepPnTAxUOVz7e73wfKnnwoFWVcKupW84oJMzMBBYxf+xY/DPgnuf7OqBzSRHZPc
9m1sL0YGjCcVUgLfcbzHIE4ar3oiiI2Tg8gm/u1c3g2FTY92nD7L3Sbgnch9l+Tj
4m+zscoMaef47Lyf7gnoD2e6z3AtOoEEDRcdAiph9YXb60TLgDoKtXh2CdXBGEd0
8NB3XJsaG/k6k98ZVG95EtwDr1Z8+u+PNPBq8wOFZ/K5Wbmf2l4Lh8KJj1FZ0se3
CnFvfT8cARUGbTDieHZSvgDRzvEI8y4LEpkKgHAYhnMp93drI8V0L56r9MXR5xTJ
huuWvcqicThcNz7D3dzwfQJHul5KNuRrGTAiife+uOS23QSCUMA6BTdSBSgxPZLE
ste7Knn74GzqQ9AoYQ8v0Oprb7P58WmgVhD4nHWEadFHPXSU3LEB91Mgq6s1oahO
0FtLtMYwAHZupKpVL+3lsypxqNa0+YHAQ019ITaPDizJgGrB7s0e9FXHcwo3ODuL
Fs98rcFfemD/rB5jYVppfuS7oHmJ9UF1lcdlTPfDFWApWJh19/8MRUmvF5Zhn2li
c2bplz23kCT4jaLeaXQmitZAhtLVBx6AQHac5ithSkAMIJXtU1a20SH3uBorJK3R
zTHSk+rh3wDltsy1S6BtwFIWZgtQqq0vUYCTzkIkxFjgqivu6zBorqD0a3zOs0ZK
ar3tEWEwK2J6K0wvBkwNqVUSZVPlHpbL2Ci++ST05Q0NDV6iswVCSLzrPY3gIi63
Df/XR+PeBU1ROTBCi1V4it+b7IyS1NTnTCJ5fA+wOmnCF4E0vBB+tecUjdsFGqr+
cLZH6KekEqMbMnhjQgq6RjjwTwdUxXxnEfhA6OIgk3XqrCFUm5tjOcIwl5mxkcVF
cvVBQTXk4VJn9D3mz04stsG8wUpE1TCDnDpnNMv5t/q6YCkaD5R7jUWGr9BOorFn
O+taaCdiIPXJe/Qd3okaRf9e020ihxNZY7ubZ228F81lOuYetcBmFR0iV3Xi4ZQ4
/OsNjvPpzNtpBMQrqP++gRCSmS+Hgvi3edulH+w9KXLigiSAXpOIFKXLfWd6wavn
F3Xkcc5jLb5ydGNIKG6GabdCVkx0rzdg//TKBl8MW4q1n+TQphCGOlagQah2qHS5
8ceyfWr95rlHdjEVyvif+2CET/rbcBeIxG7VCtOY1MkFU5AYS1OovpRQrpGPV6RU
+dTBz7Dt4BTzAkzTSKmcspw4u2f7OVjtne+hH0OOrrNuChoh0yC/KuKbM3ksGsDL
WGpzGQ0nCu5grHH7RovD1wg0mRk+R3ZmTk1VHLmweMOMyXK7C9yf0RhPB85o4P3/
ALfbHLVriI+VHbPW2IaND27W4pHKRxoOdvCIK7qB33IRNQafudw5vzNOCr3lsAfR
wmVWebj6NWjPI8lpZjVAosOJSpHHTSLzs2HHb7ALQvyFjtqL7zf5UdZZQW37OtBP
SROswsLUAcasd/ybf0bF06rg++yS7DL9IYv5NOB2qUPrWiVapIE1Awp0VO9CL+je
mYRLVx+t+KTyUB6NeYIE6jwoAzTyAMIfc/Yj8BoKP42tYl7RqWduwW+dNObpmAOW
VnjtvwEWu3QZziekEkviSa9iT6FXMKyKBePFX73GaGZ1MbMRgYQgyrETLELOtvEL
cJ4a48uCxdRtfYLwKrCMp4WSeXFZfqDM8r0BS6qRwQcE/L6pk5Uaf7C8CdCaQA11
jyYiCLkhrimL922OocmN6R8AkAdXhDv8z80gR/WN/KffWlBdVl1mhP7Vh0HGAEaD
HVmQQM7yTPdVTlhgvDjhbds7sJFxaF93K+2mUYidc95ucnyIG/SVhZO5zT792E6/
jnITR0tyorgGqOkAg2Lf5RzrD/w05IO7ODfoWQ7iY6dgCbs53p2kTsaMmgezWn1B
TBrXJ7P/nQB9Gqws76wdSdgEAyeWoc8IBJepXPPAyY2Ef0czKA9Kza13coeoYpGd
w+oCPAdta1FDeCBOXMfz9/wptpTqsDJTxlq7cuf7uWaYenbWBleXUs0AaE+QtE1W
QVzfHHf8eEDzVojsVk23mRZfM0/DqROM2+3mL+8SMrWgI9ki8lltDknkrr3adT0U
Zy1C0KKX0EAti/z9xnmEs6m+060KMR8hZha2Y2IwaXifQAFCbt3PfL1n1Z0vfZSB
KgQydOWp/jQW5gScV1l2J1J3kG86HfdnSMoYtTy5LxgIDi7Ck/PRM1PRZ7v/JIM/
L+sO13OSHlTB+R0gYRw9RBenW6NgrhlQUpr/zd9NrdW6M2hfBnLlw54dygy3UlIo
eA66yPqhn6wvrdxYSzBCfG9KVexCWcH1QFNHcP14vJGZNkgOQm6sDSAZLENC/0b2
o8uvRpYVgIRNImVxC/s3gNaCbyff+HnCj98O6ESDE1tRGfU5JBXbNwKifDB7DqKb
jwlxt76lAKuO51de/5mKB/2vXDGuvdXtrA2zEGVUfMFTq1kfVvkWMqBuBcUCk7HW
PvNorkkQZXD4m3CeyCUZWKZ8jrzKwqUZc4I0Pt2+o4aPHxsaiy2FCgSe+6anBeE9
VHHYg5hAKM5G5ou5bQtco2YO5Tt/vDG5TfFF985AD2Z6qWGQHQ+kycA2G/IiwSXY
HfPHMX6N7SADjflNNWmvM5p4hth5uwTH66Jwmv1UCh046eSm2Ju6kIKWosle7PRG
hSbcdpQD4pqmCpSQEupyzM/qCxtAvTq6hKt8c1PbebVznfi85vsIerPFQDb1QGDn
1otFpw8UJ4XVd80E2dI6fAHOLznhE5FywE98EHZM0hnMzbS7EviulUP3NNQnuhd2
31kDAiALQxrF2Vh/dahnN7GtnMk30jtRlBui9zyplNPwGUsFzvogpUSlngwJbD7C
zKmJMSL+Ynu49UDb/lUEADXt54mEbYNlycV0/VZQ+wA+HYxcjLHeK6I9e74fTape
jd8HvZ9MJ+9mbvvaN4Z9EsWjSdl7SMAkJCfe6r8GKq0dTef0VJ6UBqM2gaJh7MBU
Q19Eywqp1uqT2S0vloA0BkCKM/kpTqRvGPcGZaWoYBvegq/jRYEAtp0xFjSIkG+Y
yFDWll5oQ4ERB0YZXjHOaxPN7yiZBsa6PgXTfz6gUy8ZFMjiAaptadhF9Ksm840K
IWfHOVGW/Fq1UAScLGjFOzvFBOoP8wvltsJIeP/tJNqLYowIqLlUyyDW+m+v2jpV
swevSYGwQj5CXjtYUcKofJQwIl1cmWrkpKQbAnHvEa+AHeNjXAt+PdzKauJdy2G9
B6N9TvXR0uqWAefzSph60U0a6YF6tu1Y24nBjC+FUKQELm2DUzSIgmAN3fPLN3gh
JHdJzKMuviOiRMXMDrH9iksTzBVRJmuXiZ2uOsEoOtGKW79lr9j9y/8HaCEfLHCo
Ij9JnuwTWoRlDCMR4hM2wDfLMu3OdSRo+BMp02AVw+3K4ThKCFVf0Fk+6tOf15Dt
3HEuaT3FOA0J2bJ57pNeW/bgqGkfrkDkM3v+NfUSFP4uDBz94gUoF8N1wCa+Hamc
e968lQGq/2js53q9Oh3eRUjtBTU5yj5xfuNHcXcabF7atjHw4CCfs3wmuk4cUKjL
uXjviltqJ3o/wQzGiDM6zCtn5NJ/xyq9d9IzJP6M7lfM1FA/nhiBccg4OOmImgtv
eDfsjRBx0RMIQ5ciN8HJd/6WvgR5cqa2nWCgRj3AAedHI0hPPNdRKrwtIZFyVqnK
7Bxxpm6E2kF8ZRTGVO+3If3XckZQ7yvKqtJ/pAA53j3vhWLpCaLCzQYTt9rC0U2x
8OIvdz5LG9fMsGc8OIJgKJaFq8lYhZcJhXWN7wwikrUO7nwhZKJ3TbLumqlzglmL
z15vOS68WtvfoPEZqOm5TOxxeRGdM+nYg7EGkecxuXckcFfNYSA6GbwJ4Wlzz/Ut
iyEkLaWzhElw3HiOE7w/kl0NPZM+tqMjiw092LrYKAF+0+oeYdjQlVtFyFovmJCK
y4Pu53yM6jw9ltFBd58BzRLuIIi/ZN9PUCWPdCMVQSHKuaw01oKkCQdfLTVJzozt
VgcTuwiUpHieFh0CoTh3eiU63nn/2jFeLElPJ2eB5QGcbxUQfZ3GOwukn+BvpWdq
KKojCt7kjnd+CkkMB9caQadpNQawi24C45YiPZF2ab9ySJ5ff7TRJO1QKLmwpFgv
Jl+NZ1S0A5O6/hrbB7ihpjckrhhpEwlquAg92Rt3iVk+sJzM8HjUuFMvM2f3luFJ
knGpBS+b/XIWHOd3D7pytdWBWUThZiv98vtI2+89Xxf04GhXX93ElERZLmgfTs16
mqZN0xzOj8kwU1ZIc6mRyoUqB/+lJiqcsJfu5tSefGkc8bipF7IrsNI0Tgx/jrkO
SdwaYHKPaS7u2tXfeAtcDpAfyNIBj8csqx03lUHaJdwu+vEmS0iVEF3y+eh+KjeO
0edpBw5zUWMGLomJakxfyKv55HB2EeGrCmdFdNOc/wIiuIiDfxDg+VSAc8vdhmcq
0RF32b76RPu2j4e9OYJfeu6XYSWq6fbh3gI4xtBZK0vfxhj2Q0lnX3Rvr/k/bd5U
Ly369dhJoS0/r1RgXmdfeQjFhpm4yKR1mraKkn626OkN18+Ij++wE2QXolKRowa1
L6f9QYYJVVK1UvXU3sCfJo6dVJPWLNdVjo/aakePb1FC2AwmGUd9WBkqrU25o26a
fTp57bjZVO9CZaA8ucUhLeUhYSloS3TS0sUPMO3HdYA/o4nNrwmXi2NsLle+ngkt
oXN9ljtaKSacGeeaxf4h8cjKQH4GpQvTa0+0cPQTwI2tI68GHk9lV5R/VZGpGA1E
j2n3Rb9u3APPVd5+ll8wvcS50fVB+72g9pRBz5KTHVohQX7lWuyK5/fLxgsESYBO
yh0KzQdGWzfyY/tPTwWkanWBM+TiBrs2KDnMOLyorixXulQIJHFyuFK+tcMIsP88
kW3D7/Q3SqmFhol4EMPe0YI58yPh7ergWBNdez+QEyH4Nw9ZIRDgrCILxlmhiOvi
dzeCzwxh58xeNvgZrmsK7KauUFfzBekJvNroQ02BF6EI3RgcvRNT3Mrt60qnZhg0
1bp4SVfuaLOfxsgtjSUwPTrNGKBsPqNRvdSrgXUGGUH46ixRrome97AU/ucL3OLm
9PygZ1gRW2guLLTSTgltgXXoQ2NjVMKDmd7s28zO04P7F/agkotoiJRkl6Ont2J3
xonpvO5By/nTmHDJStUrJawmr/Aplt+8M+tLtXpAQLYaHuTuqqiP5SG7occaEHrF
M/OaNdGsf5lJ2u0rkDlv5Ttr2VECoFKqvsGzaLHvdyKwendGv49TDnKnDLcyQo8m
/aspunUbqzz7vDX7BU7ZIQfRZiqnuQRO7Q6sPPbyiwS6DZOOCSdCluWnUdNTD9WG
xtUzjwfaYo1gI9fO7TjVPrc7xr8sVu16L10uiy9x3y3tO1CrZOh0R0OW3yPyzv/w
pgVMS6BUYH0Uk+QCuPoJgFRTDU9cyBCBGqgJkem4PfIpDYMd9LQ0SJdjTy0wZ1rS
mAdTWFbRjHPYEEgDo4RLYmTxJ4g9MQoXOZ2s0qQzmwCUnNlWCQxRD3XfmYs/VPGK
DN8w+hITowBaLRgcxANhYAkB7gnu3+rPSUEOK+rzWMd/BDGQa/AxADZCZgwoyUIJ
sSiWGmnnHWkwV+g0G0fIeeq64QnSdUBG3kO9k6g+5qhKLc5EC3Tc/McMgz6E7gbH
rWyIcAlkr2FHhSUdDDcoz9bFZUgs2szmx8dn3+6tO64MAWF1A5EsD1ttXOb+YyWP
nXQQ4w8dKlzMbWTkrY6RI6+Quqmedy+ulT6FCPinK2CWN4aJLJGd1EYm9RiKc5Yg
zWANzRdnDJhG+/8B70X8I0O03Y8v+hcWS7ZMaxlciekMSB/832ugBV9HxYBgXZa6
zJAp1rdH4+fZt2rZ7RW27AiPMPZu1F5XrOp9e9em5DSIX0uR8Z+8kpnh4coXzeTK
C5M9KsOJPDhzBCQSNs+4WoINYwq2q203vsyDNuzW+MNWcxQoTD5sDyl0qSaBuiOb
6A16F1//Lu1nUG8WPp71TjxQ0kRAdJHgbfcF8ZCAfeTnxY94SEUWf7i7eXg6YXvu
QNv3OEoO0Ma9wQeM0t6yXOCrZHk0mnC3G8vGnRgtqmB7bdiXtRAHCmqx/EZgL4wr
xkrQu8gEQo/e+38xQWxlM9ynZTztpPY+pKrtWRTwzy8+S3pxQUZR2mfyT7dNiRGU
bF5Dog51FMNjS49JAVnq6sGpM1iRD4mSrp8TFU1uYPfXqvnzUAz+UuEawsBoGZai
2b/LZQm/3VGuREH9Ldml1G8Gi3V9jo/rAfXxI0SbnukxfGsOfqjVdtwXm1SsVydH
NtnZxlHqx0kRaZFMO+xR2a9LHsOybY4ht/lT8wqxwC1tMf9dAJD54ASu//F84OLb
Eh2o7s2a7JH+eUH9Ffn3ikHCnNAcXQFG1e4L/2PHs4nSX3aLE2pegsRaTUMslou/
+tjK4g6CqXz/NY8C4zLSflu3Ppq9fAlatis5Lon3/b+gl4qzbSMyVKs36vjnkgNB
11GGgJjFzrEWgl4xJvSkMXLP+DBQjKBmPoOPseX1CvEc6y6ZBNdh3l6WA2WyC7QY
+0u4LwTEVweRudn78mYm2pfFTbtw+flE+8ul4ijbhZ+1sq1D3D2q9BLZqGctfI+z
k2e4SWiH3xNc0AyCEFMEAT4ipAFktpXJGJa9Allppv59phO7wBOdBx8vXfJXg3i3
D24jkkoUO4nl9crP9hk3T/BF/HxpfaaCK/+7DHms4axh8z2wfGqJ+rpdS53S72om
3Qmms7UIAZxEcf5Vr+b2Je8FPqqrfdjNEdA2/PZHRh9R9CRfyLCSUpFD0rpIP2C1
lrDHajQ1dxDbbLvJ70UuDrMmB3rjVWeR65pzhKkSk2/xU9+hAS9lk4n4ziV5ijdc
ZaepDe0UqUsqZnXTOsRzA42THxPV8GpLZnYv33y0p8Y2DriBAsLF8TTcddGbBsQK
RXJXUBCg7ftYgnQ+Z54PzzN34+hVqT4JpxpZwDJtFuWC2zN3Pf+8MKhW04/Ykg2d
pjywsNFNlPEB1wphPvp/hw5TGLp56+kAhkaWeOQE2eWKuQ4ynrjw9IlHpHyC/b/2
IXcXNN5kMBuxNISaTc3WsDFmdxPD/rhpW7/1kt9fN14jcC/jrs0HwlJ2bo9icAL+
ln6PdsTcVc2dxHRQvtsA4GFnSupLgLaw35ZUU99DMvSM6ojTXPJLyyr8qq4WDAdb
8XlCkV72/MgWWg+zKyQYPhriUb2Wv/bocYIgIc+sRGECLLU2gtEOX7amQy83FRDO
tVn8OBC7wKEHqYfTbOrHB86zojtEaya+qv1sZEdYvewylZUPSQBjV7VLV6f3K2vV
rjpshrBE0N6n8raPXKDaPVtBszpODWtJ6wR6Ua/G1PGMdMLkIiTL/e32x3QQrxBD
B+tinjrxfMeQY3vnLb9CLDF7fYQHijL3r6AU8lr/dJ7WRx0Pd7N0uVvRT3EiLKrh
rywiWsl4NGjC1T0/niax2wPsdZp3uZwJ9hNZve9NDxoXWPutIbYRQaXdORiA+phm
SYivPRWAnno/ONPoWc+6W1u5EWSx0qvd86ek+NcRKHusULCCf9a/AHLZXE9EEfmu
vNqDLFG2v0pemkOkQO9xP4sACfIfTgdg/HZ0DW8mI7wgQRsAZPXXgkqvWyj4fS4e
xxawEOCNTLCkBiv+ZoTmZRsRvnvNqnpGKeBFhRPl8vWEWW/2swjzVAIYA6l742mN
IDBWmpymzPzW+pZJzl+0O6o09h1/Jqn6I64fsVW2t23yPMWt8xg6VTYuwGQB3tIC
ovd9FLdvIunAsScJfk15w16QxUI2H7lxZF9pC2jPFtydrXs6SMOVwhkUOLVtE0Xr
BwtMIMQckIdalmFNrn+UKLuOx5wbUP29kKpfDmwa7p+t7mZ2qBLG2+cnGj02IxVa
Md05nJpkfTZpUDjiulnUTkuEiYDPH1hAnnjvpnWq3gbUfNh+jyf4Tn3RPd0+q4Q3
0Kui6uxRQNygcRaEC98KfVlkcT1Fc1H3bCU+ZL7IMjC+ISVehAYj2p8xiGbXAl7a
hInVdyapaaD7FHcVavPz61tSJk9Y8oUDi1995CfYQL55S/HGTm2KGFuEcHrcSj56
gVFjqHVFt482liMW1Gj0stoO50ewEEEwOIUfe4XO+nFPr4HkYLrtqE6kfGq0tzJ7
1XbSh5DZ7aCyFq6Qxzd2o2WMMKBHsepPLMxJ9AP9Vc8eNNSiEuwMkt22RFQSC3bH
DNDXdavfwr53Jip3jfslQzTwR5RrHKKJbwLeTuUfl+eY9reYjJNrhYjb6kzLKw30
bI6UaK1Dd4KGaLB54MHcftV7RzVbHCphuqLNfKc4pmU6J/E29nO/ywHgT6XyZev5
RxPQDgJFvzwSI6/eZ/7riynAavqtGD6PFTqcfWcirP/XqGJYE+C2XHugUlRgsXki
7J/9s46BPFp/H+hv4vSHqk4L0VJYexr+Bm2g7PLszPncunhAAbZ6ZkzGAcII6aBx
Pm5gCc+I+cRj15FYkDUYqvBSzNmubTXblBTjNuTy8wMs7UhCLNQRn8HETl2McqiJ
FNT+M2TjFR4Ktd8NqJF/GuTWvZZCbrhfnPY8Ow3RpWXfnpZTB60XzLd0nq9Fb5Hz
o21xicVyVYxfjEYNQxNF/F7G2L7wQA/bvYQ4NgbEJH15AnFZc3x66cKH0I0C5a+z
EDb7TwxfLwpX2304L28RN8yTL3f4gpKkfuL+GAu7tY1vSG90mls8HfJMPI4TzLPv
FQ0OmtAnG0K/bECiHLBM08SC+srTPY+NjMt6fKcKmzx0fCQqIleNWmgpPjhHhXnE
h/K+gXqRfIo+qSQiA3ZUtwp7QjFdpf6EuMwv5DKWZJsMeqgQt447EbZwjoa01dXJ
fWIjGYqrKAatYFFnUo8rWUGjqTrrk9cCRz0DxFz1fjeJnKBRIZFLG/Hj0l+/iy/9
jlEidMA8ETT7wlS7Mt3m92bGWMicc2TWpS2uhc6//oBOadCEh4pwNWuTbcedJNov
vgP507xel3/DmjQW0YvBbUQ6pCI+vgAoGSjtjP4gW0U2lniL72vzv4jQUzbiqHmG
FIeA/m+jwkuPJzQL+oQeOSVE4pnmGVlSjP3eY2KLT//zjfurIk0xv4ReCSbARnGL
Zbbb5nAg6Ss3nwfofQxxonmRJ6V9Y+ddNC1DVCqshvNhp4QPZyUwVUdV9HFMydp+
M/NFo0eOWqwXCcFBUDYIiOwzIPvPCdBVW9bhOlxZ9lW3P6PmbYsCARx2kAkRcTeJ
SXRaifurMFXf1k0Osotg3+7yMHJVBkYt0eeLD8og1flRz0dA8VfcUbsv8Iy1PVai
gjg0HnIAd+XCgJrTuB+4NFi1Q3cwbtshqp07F9Y5qEf3Fu/PrvrF2EXND302bLoV
yf3F9EDAjwp7/O5s19iRsDS2MbEdIpyi+E80wkatj5vdr657xgS6aP4/FT558oxj
gQRsFttFQ2H+rn9J/saP8cllVq2lvx+ewRyI2tLaI4pP8JMLFVdMdZSV9vhVeUCc
VStxNCowzReKKxPnilSiJdA9/hpUINVysedEnGr+oK17gnj2iFVgjgrcw4j0Asz2
wpwRj1u7+ZTZwSRq3hrBLWeAoE6swBgHZSxC2Uyk8BUJaQXD/3tUomzYfBwqkgKF
JyaM24xDmb72PZolfoPHnIf/clIimKZeghndWFu8/rygDMGBIl+Vcmjz4wvBFuKa
7bDu+7cLfDvJjE4yrE3yz1RgqXGatNyeKsX7qn6s3JX8UhQy2Id5joHOu83VrxFC
O2URYDqg19KICg/LQh4MjYQcUyGQs1wlPS3Xg67ZK282FH2F3k/WTVvJccYFBvue
DLtAm76YK0mk6hvsl7jk/ckhzLD3HGqZqEL7nfZu+e9Q524eSGkEEooDNReYfM8Y
GJdeLkq49xYAP/Oo8f2j8ba7FRubnOg3z9vRiIleBx+kAhB6FBkNAqht1E+eAmTw
wMW2fGnKUzprT2iFF8hQabRjkKbeC8NgMq0eCZr++Fb8taV7FW5ldIVcIi4Yo5ug
H0mUx+RMPaZ7KEW++B94DmdinYYSzdanJvjj4IXtuQV3I0jHOWmPYN+fyi8VJH+h
Mx3uBtCycpGn56K13/oSvBzsQAeE6fLF8H1JRS2bAf/1MSCKGH4i7pUiNxQxVb5h
v4urPXko2v0q2FH60MKbPc6Yg3HNE7Txq1BWYy+hx044Ph+6JLiAUY1/e7gKraLb
gZgXiEXNbexap5FwGvAg54y5NjG7eMgjTo9Uc0N8lZreKBHYg30bvhiKy0WLFpdW
OVj09THXlFV64yZH9AChUr3bxUZzgklypGF3Dc3/U8lSQV6zq9LfgiB7jiUi0Dlx
AyasTDVtdftmMh4TeY+YZbY8OwwDE2FJ+kfS1VwFfNc+F+0Sr4D6eu/6BBd82obD
oawuwXreOdVPzvWQuMfGTbvc3OLJTLkuf7PwOgAWgQ0GR7pD8ylN8JNF24fzBRK8
Kvg81pNhC9tItEB3+cki5PUm6a0V4hIUGVZXzI3+gzLl3zmk3N3jFWuIAF1insTT
O0Hu9+/RPnxlXGIZGBzN+kgfhYbT7QoqmiHiZObfchj04fZfzUmFlHEzvMizeily
Hw5PAX9i9FKvbx9TDQ0R9bnm5dWduAB+l7lZpNEYNjhOHFyTdpFLXjx/F+AJb8VP
CWwyw+TxGvi9oynPGkGWp+oG/hjKqj4YK+b+QDV0qIBPNRwq2TiuHo1xER8LBQRU
tj3DJAaf09hhnH2AxpZJWMxxt7t2rD24TvN2C6CTej2YWjj/E4rDOMRvFmWR/ScV
uI1DxzDWJOqxQcDLg9s3KPDDZKGO+HX/xSSLqQFtExJlHQciyvRE/DsoIqAt6ato
6yaP3XHbKaSiKBAbmkZwf3eeCw06beQ5Cflm1XLquk/98hBiujp2lS2PoWYVWU2s
CWk955K/Tn5s6jp62emEeM3CsX+gkXUyqcoK4ciao9Psa8PQY1++gwqvJi4Awaka
PN6Of3twy9Ci40iUwGmPsw3qjH+4fjKzLbteoroFuzyd4lVts/ZBJgnDiTINt9BU
BHd+CgoaW9dPPfv55IXVAoE/b7/yLdpIx8ssyY4gjCbWwUk/08kzzrTq+5QD8bWj
mN/b+TWGE4s9kFwSFdfIn0D1V2fssY+I114uS3h/zZDOeteUxe5iBw2699opHQKH
/8/s3dwCfEfRHpO372KPDGrNseBiwLikTJVqwuxrjaU6hQBaASFxdN5hcf2V1RfK
5YVEWQMojhLkKQcExbLz2rvpxscTJQ2pWl4OLAtsiTBZHCPEj8uRSCRMghIJcMeb
dUoJB5T/3owXNwVeIPgfukRauu9pEO1ZA/R2leATC/zcCnNZF57OSkMhQxUHye5A
fwn11O7WKJlc9BmD4ptVJR+A2+5t/TljEZRu8vQ+814IB5G3tOuTf2BclYiG/CYY
`pragma protect end_protected
