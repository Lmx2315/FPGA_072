// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.0std
// ALTERA_TIMESTAMP:Wed Apr 26 13:33:39 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
RF9rCUKXzM8NBrx2kRMnzfms0Va58Oh87gvI/NK9LPGdq/tZRbWKPGsKFA7JeXNm
3U90Qy5fif76nDjMy7qFnWG+TE9HLimMGWXQMm4M+FpalYPZODSvTiwuMNNm69Dg
tdG20uF4F+rbpwvFiPBG3OQxUBYKBfuykR9SC5eqZnM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11632)
7BhrgAwpyP58Ca7Fq1BY282O5O+/D8kROZvrqidu/kZjguM8gdOFEzXGOsv/54JP
tZLl11/Q8MVrd+joYI70s32QQwJ+J8g+oEzA0lpuB0N7XJIAmrvUQXjxVvEHG13e
p+Sidn9PKbDpdAMoHHclxrH4XAhURS0OXlffV4DtMfW32LQl4jrL38LHnif13CHD
msNRGYuZ3qC+fxF0Urqoy+OVBjekXPCmrylegwIuKKuv06/PbBPg7HJxxUYtEC3e
LQlcN5fJEmZHfR3w+xel/GUSsS+QPCAtGXJHtrnbft6S5rIbnkrEP3b6zRkVF2YV
d09Zfg3T9KvUSyr0u1cd9oxW7Ci379Q3/6Kt86Vb4/puph08LQvs7dOhH6OgSBi8
ROhqZUiCNIopvB6QiJ2c6kKJNYnz+DOxQA5wGusCcjK5uvGsko0bgFIT1XbG/kLG
EtMgKtoEF2YQ+91JGMyfjER2bIXLLSzAxV4MRLnYYrSH7wDW0Zc5CcXwEPx9WmyG
29MPi+kvfTatuMNqVWntP8cf91Ccb6qdusvmDvfC7H6fLuRSXyTVQQpYiEC1uLJl
W3qHHvJw39ZBrXnWK0mGPaBTYnVgWJt6Q+fWZBLUcpEzJ70iwdFBxur944EbSA5w
xGlhVjuksUiyR9i0mWiE+AkvQ47SJfDBNla+iM/3OoNxlBUaFcd+ZSYAYFS3j3z1
nQqMsW3CIyRzJfiFQSn4DJg/KqNvli51tMeb0mrRPoHKFzLH5r+iRnSo2UJevYlP
BRU5lO4Fhk7wL2BF9XnT2Ql5CvC3YLndVw8ChN9tbgFb1EJBRQXHCi92InK4aCp6
WznWgntDf/F4EsLTa+a0ViUpGOrYEeFIxg78+VDNgTnNRjsq1I1yUf9OxKMYUay2
qgEZVT7EqSSxkNWoqDTcomEeZM+lurjqS6HQBqqOqN0Y/IGEemGIWZ8d1VH1nm37
Vf/kIahStkyU/jl1cK6mWCj7oWtWUsQDYgdzSvO8dtYcV46EtlgE5ldbBSInXsQQ
dA2B2RoZc2OLLAYID4MYQQIDzxDf1YMPnIUD82wyyKmCIWTKav79uqJFCceDoBMN
1s1gS9QFgTr9pZEsQW+pb1vwjsDawkC4PhxFro4oCub2gR7k/x3CsjZ9KRsTvc/j
eMsYyRrYrRJ0ZrzlTAwQJOLQTtatYoxuqb5/psk3UL1FgK1hNJC/wBnE+kniAHAd
ociX6cJzt/2raKUG+HbZTXiTnvOky081kiT6qcOJ1e0HbCtoQIOMTf0NiwUJhuOe
1a9ZePRJuRSEvHG1qQUoEHJeAfPFL9bbl4PQpTvsEC0tUXEGei8NViSxaZsQ1jB6
0e046vHe6O80LLo1DmEhgAgJwCK6cweSAw6jDcbHed2qIlTa9Q067qtBuPtNLMAz
kA4OX+D2qs/nDp9OQYPyXMVmQimYYGBCE5IjNugbDy0byul9ikIW5AuRd4gna2Xi
dFnCDNH6CkfeEATOmAPt4+Qh0lbyXvd/MGTqdCZ7vP1tEneZ99RMQSCLuPusaxZA
87jyrxQ1A0i3MZN62xMdt2TGVLr4ghO9k9c33mPuKkSwqz/kTlgLHhTm8jcpro/6
LiyPkiFuUzYct6zDNcNx4D7rFf9TSNwX7I4eNCSh0aznY5CCxmFNbfU8MKWGw9a7
lcCya3p/Q4jEw69aMvjUlGy7Tx/Sa40YkZ6pnTM/c/pa2NHUaSwIzD9A4jtZICDv
GB0mvvvQ5xCvPHPE2USfVkg9uGjRv4fvlUxbabnQcT9jOa4yklqpzsAJhf4/u3Eb
fROOm2Xs8daJA+lTno0Un8NzNehR6dF5I//UknLYdV3s78MUlZ5+9AhNCJg2n11U
bnDb0l08cVkEoZjEb1HfvhvnqU92RDXwWijfR2dOtFlsCRyFC9SnX8utjM3StWOh
PitPY9LQyTUVfwDksQz09DAje+pCbOnpAttxgBpvmG9kpAWQppqNVYsLo4aZMPJ3
8ox/zIgSo9pmDOeSqX/rxgLCJRkZFklLCajRBnxNV1Rx0cwcgPo37sjCaF+lI/Pq
ZmSr4NNHFIYtg820A6Ll8efrQ4eg7J34FJmS4yp6YQqjD0MFHR//bXS2Qd9N33Tx
hrG7YMuggl/pjkwQJy9eY+VUTMowjD+aDMpQOh/Rw1rnJfyuIrZirLeeJd7grobN
i/M5eKoyOJkznlE50+lHfgsZeD6fbPPGnEQbvr997a/0MDpqagq9SWk7QYVu625f
+rzPPWLF+uOHgBMOs7QbJdDUkmodZXJ27UNnMpOUpTCwwa2bjNk1RsxmsxUkkWB3
by0VjhIaU9bmhz7hoESzXROV9feIdmfY+ELiqPjlTOuWy8suNhciejcEufPS1rS2
qHiNtGaWYAjEeVRiWAmJtWFBPizUOp9u1x30eBXbxLAc++jeNpz3XhR1Kp9LA1ty
CcZD3X6uXaTjno84xTRaVyQuyQMmDJzTUZfPaQVSBFLItYe4j/d76Cz0gpNhpPTE
7TUbMdyBbUf914bIuMIlkjPXvi11aFa67JAa5xheR4WlKTLjP8aVZqRrkMY7GUtv
/9TqLg6gTPku5BoX91KTT1NbSqfZPBM7TnbuXM87TOD6M0Koz22/SoUWp3kDv14C
R/3e8IjrvJ0E698bjyGTvY89cKaCOsvetyEYxon5bfGyiKZmeJjtPq0dBNW9M41c
3lJh/1+MFag1xMPwAZupTugCseIORY+uGDTLF7N3L8e48QuU7DU4j3GICCGsssBy
Lm8p2gwDOBgrjgsQ/v5zT4s/UOtlIAriRUXIpTEEGyTLFjMsCGnOeHg42cvIAOQA
hX3F4Ll7b+yAqUPXpYwu/w9dmH8TBSeINDVXE27AFZuGlJkAX/khv8mvxro+NUXx
iKNI+TVaOlnLm10J4p0IurRo//cT+Fi286P8Ad1YKAkOUz8IG6kXvCwBjgYK1rmr
rhaZPbQbRXMxT5+T+6k4Q3+Y9LeeKf7E2KlIk7hSa5IT8Ez3/rGS9RFhw68l6+Tg
s/no/YCYCg4K3Ep1g6p6P/Onm4Vt42Eg93ZCdoMogd/NMukZoG6UkCbNK4/yNxR+
mBYOXY3ex348ptQtQoFUJuuRJ6FPp/ZwFps57F1Ba+G4Ew+sjgujTmMzaGKewZJH
C0lLtIe6MmmQgi29qvvOiQhRkSLAxkTJhMRA6ZPROoq90U+TiNigZHDFhPkX+TZ3
vp9X87de5HzNiWoeeL9zG8+ltjWzoWhXp/bgJnD2PLEw7NiBOORhNyTK1jhIchVv
cwtR3btefkHKn3htVD7MYNxauocZFqPFSY23h7h2vRn6Qh7qkV+MARcuoFpwUVxs
GDJFaOUBOxMgNQmgnsw/lsp/Q+Y7bL6h2FzaDFSoQd8+4rWjL5OJA+sS5umlntoC
h01+RLYB9OEBI0swZwkar3/Ssjti0q+MzzsJ11t8l5fG3I+K4563n6YEZ5Elwuz1
tiHDozcmasouByEOrRo13gR7IC6/JkewKJZPY200iuw3wWpoPI2RWr64tTTtZJ1v
C75tRvVTTgoWNFZtYkWUizVKttm/LCabN7iYNtpNKViiGxNRVgqyAcZm8u6QVIf9
pKENWwLGqRlL+4USKxFMjBc9ErpaaThP7nCa5SbYycABwXAsIWvkg7sWa1GZk/Pn
Lh7ndk6azqbvWpetjrBMEXA6EXh/s/W11WtYtX8GQz1U+tY/OGrXkL0JXcRdS6se
bkG5jnHYZezUeQ9ulbEglw7RiWZ0Be/3XVa93yPRvpdc00w7nHHZ/dwv/nSYvWih
M8lMuCa5I04azk1ryRlQEn2oFLgvB3c09QCuOZqhlZhYAYtIUd57+aDZXOa1NcmY
vKP/iKI9MO1UvWpvE6kADFoxm7Vk1juK26nq4SieoDWeZjTUhM+H/J+ujealv/oi
S84uOmF3wdaZwlQ5oY6IAjNsaEaEtCFJYboOkzqMqUzUSkKdCp/o+4gFesPrC+MI
o/QPw85TquzUBtcuhHoc2QN83NnAi7o0+UDMO8lSA3D8N2b5pWZ3nOMEJtuvIUzA
9PTndGX7/Q5zg6HaOfIywg8rZto8mWVBHeYQfNlK/HJD07lEFVKXw84wKXtQYefX
Uemig9jfBS2JKM0+B3YDCtH0Q5w9KyX5LdFEFPBjw/4f6mi653n1cpYunCj5NN/6
oeMVJVyK6TOs1HCB666CMiRAcaDnVQjv71P769tMVD6Z0eemQwSCMac9sUWzB4ir
Ua5sK3hdX2wF36cGFRLXKAaavpNWeg/scV5FjYWzhWoGIp/WVuUd4mbGOrHt6Pv4
mtHzDpRsQBP1HhURBbMSjNETelW3emIdvX4qgEolJ/o6Bczn8k+AzDW7YfKTqnOg
PrJ6LYrFbSv9bPtMuQyb+hAntQ0qy9b338pSFIfzCriwiS75AwvenRweGZs8mS6E
C2BTh0qCNCZlxg/uzE6TZ9nJ2IG/By0K7sFH0dSnn8xP5cMtuMt8CdvVLU1ul0DB
HWlaPrqonm34t4Y/eSpG+TGHfVGk9nbL48Bw74WyX9NSiO3DiCnNMTpu731VjKit
3QgULz1cfzAJVfbP5a9XPImI8gy+95AoNAV1IlrKfVhb2dcPDj5xuKy42P/eECv+
4Pd1J3xcYx6vE2RFnzwSQ80lCDBx3dRHAw5GDgiBHpWSO92BAOqxECYEeC/O9LV5
utmVRNBIGctxpnF/6nstdjhMeNeX34vI68BIcxDYQInWiwSoFMHE835YVOroS20K
Kasr6iUMXYG9K5FV9+ikDNzTlWR7aT2rS7OYWgd7aNWf2C+NMaJRSj6zGDb1UZTX
VOFybHosOxHcTdHQ+0Us6bSKZGPnL/T/qhuli+XEm5Zjuw2WpEfermfQetUfv9H5
8hRygVjscbFCLJNpZmHgTJ/6ZP+E3xBa08D1SPfC0C/jm/xAvn7vvSv3lyfv5BZq
Jr9JcF+04fT9qrIIn8zAi+n7YB38TYtOomey9KeusflPwyG7EdKkzm3V5+5pIFkY
TZZiC4GwA0ZwVbHkkjZlgqu9yeBWRDOQIMTIscs1cl5OCprEY+mxrk1HagtucUmH
/P7oMK8YpAlww4HDlx/yRJK5H3yCUO24I57vrFWNbvB6YhfRe0JBzP9/mlsp1jRS
8PzEbCzVO35UxvyWg3M13tN63q+AeRazFGFIDhiH3oGzkjLGg6RSRQESzD3XKVgr
IEATdjCWQW5B6oVusy9J/ykEjdeNuhxO/AdILflGQ/0hOMsCZrXgEbRPF/1udiDO
jW8Dd6ZGvb1cCCX61Dk3O2m7L6CHCT2oOIQllBxnTvjYfD3UEslhbKeXw55u4HYD
YYjXRH4XIiSVis0dgW1Zgmk2tG0HX3HMoKy94buKMZD80kywDLgzBBrrAemakdTN
Qei/ArqTQDSFbadFcZ2eVvk5rqYPsIAEIATM+FZtCmjdUrsb7C5egKvCC4xMe2ZK
qwdjzpv/4ZrZS41UMv0TtJNdch4Qp5ZRbs9d/1cPnGKPk6R0U7paFbTzP9GxMhzt
On17wIzh/Ah/aM9y3uY6MZx7wiOxBIhmBapsRpZacTznr/udKQ/zGfbfZf0I3DAT
f9x33vg2paOgTjXu3JfufbgCZjZNMMtNFcjkg2Lua0VGaKBL2umgGY+clT2nC1ZT
asaVGHDKB5PCRjJhIOfsiKyTC5OufuP1sLT7ZjQmpUYX9A3+8ChIULux59NaZwcS
5fUnsxsR/f2HFUmzgOOQgq2TLqDaSaVdl7tpzuik9z4sf+RIX4kri1ipupdtsVke
C2k3bkxBqt4TuuFwufWsdAVARtoyPW3Qgos02ZWjKT0bh04EseEclvva3Od2lS0P
R1voDf2zcBknfp8VY7Qh8OzgLoZBgXPPMW9d7Y419+qDF2SLR3cdONmd2MZr1mVP
3rIWkOmTiNyknmKBcWn9GT3FwF0EyZaoIV8ZLAnx489FUvO8ql21DLAk/PPn1pkg
eAc0F3uzksSkgEzGgQuZLBamnPCiVkTNZFdMbtk1ByTJiMj5xF+V2Yf1WpaJ43vt
P2GxKDnm7ohRxwfL47/mM00KiuXMtnet7HLSBTkyUIp1cY6/1jTX4H7QuaikAoqz
bqFsxpwDhZY3+hfNkgvovVufUvR29+utfN3SU3e8pNw8lynTa6Nd0aV+/jMEa6lU
r6ISh2ftuTz2JHkx4m5ypSQEuY1YOmb0EfmrLYqbL5+rxhMT91MGygnuOolMyLnb
0aCaz19m9nB+HH68dcSAcXY0dv2MnSFSEVAvt299SGaT8uzNAl1xVHhjXTGjL1yZ
UP0ynzS9rQAr9UIj/Bk5yn8KR8qZ/AuPk0/r6qzVYnWXuB9BH7jBU0jEyme5iy4N
LDtyTGLRpQT7HwO0TuptM/0s2fNBNiV3pccH8YB7I14I5W2zFRoEkEqgwkgSA63A
M56TSyd/bV1L94uolrYsf4c2deZtH+OhNsqkGTe8IKL4WPN8oKewe9qJOfgneau/
WtnrT7o6uE2IDiUodVI4WOGAYORcPqb4R3CRF6BFjZZvoJNvHMtSII34D+Tjo+wq
rrFDXpCH1HcVAwLuF27TrZDgjd2IZ4QzEOdPdzVsVH2jJCEs/DBfa0oxLZqdmzVv
0lI6LISHi4wBlkdCXEyXv4izOPZmt3Kd37jE14r4af6JnjL3JwDXRsIaVpg3SaZZ
wrsZWqtjoszSxCtRf35b8hhDaVV+mvROFvIrhRvAiOApcBmn4OlNeXlbgXAZSLpn
eVDsfHt4b4q63iuhdvDVsPMqvZ9n/8mKMl8CrIalObbJiPXj/YvONd06VIqAweJF
GY3ngiuwCSRNwQCbK53mapA8Lszlvrp5cDXEN4NWW3+2pUPhi4bwfNTgsm3hfisF
zJEymhgFP2TMys3dHjlRpWTdEukcIdTloGd8aD1epHlN5VKGoQ9cZYHg1rT4eN6Y
5BaaOEcUEfnl3v7rlICRZ2liax/iB3UCYnYPB2ql6MEqE73IgZzdlk+z0LgGYEuF
12msJfIe27/TfVqNj+L4hTvtgMezAuTROZquigkA7nPWeHUsuJ5FcsQHx1zIKmQy
panSGHqPVNvohSdR7dNDCHgwkl08Xt7m0xYd9uBXwAkSJ8ITnGVrUCT2rgPBkLvF
kvGAuKxyRyrQWfBv3pAtY2JR7nF9PGHkvVAKPAr0GrRr/73LfBRn65jY4X25y54U
ksaJpho3DDAV3vGLJw6yoB1Y+pVBmU6EHySGf6yQv/amDqZvI5oI3l7v+edQfIHq
SCXWplJPaficCspDiSByllfpjMRaKFCu71tuiJeQ40D6A/V+4PrWrMpJ4gYEM0aq
0HXYEqSsGzcXcyqIvJjdbWTNByuBErLwlHwrYBQPfyajvxhMJX8R9mBe4mQziirx
mAtj1b+yomq7d5oHLT7A1RRClt3nOqS8dR/sj/bfldPTZf1rsEif0i5qUhZnUEfg
CP/1/AbE4xEtQ1qRkZ7ucMCpz9zi02Mql1ubZX4nkPR2UZ3VtqonxvNkhIsEd2qx
s2m/jDgQB+8pMCiUJATMIcuudvaBTAW3LnPxyHORYLG7SAWTaTCvKyCPp88kIMIw
oZnZnwYfXXi0VJTw9kW/5SxnrFmSJwFUavIzgVHwEwE17G1He1qQPAwsbw9hI2WR
AVx16BO8ZN3n0JAgJWuM5YuUOoAqxU4qy78hsSsLQ6ptDslDMK9IfWtK2j3gM95x
yQKyi+TvLyyMgdrYV2yD+eCx6HBqrzE7X2wzm1F8ex8oAhq6uKsF3vxMZz31cUpZ
nyMVV9hBrVWlwFejTJOxaPRmJLuH9aM/qJsd5ntJXcYkjocURdQWUHem1mFdC3B9
d4PGG1wt2HBpG9cG161m1TC0D31yTZfkKoc/cNsEYXJYCy/HchAQOtpy+D1iYGaI
3Q7IEAzYmaseWkk+9NRyULBGGGqhHmYEJxdtI3ROsDBTcYsYEYo6SLXJzsbCsqgT
tKiavkJMAfkF7stpOS9u0iUIwD4el9QQzadlm1mrz96R1O99dS9DxC5W5jYYTInV
VkXqBx4vE7/RUBYefAxMS8Se89IjgDEnrT39Tvpf1wnjgv4tE9Xd6bKbusCI0xx6
7rdIokBoPcy7+o+c1oplDWqQloPknNJOtSrODRJ/1SZhUQitxHVSbHPJHrYrsnB6
1MWRTdahZtq0POmuA0VxshvLHYgd3XzGyP7zTseBznFLuZQUW7k3clXFlJKs4cef
Xur9PnfxDbSS6Mo7rdKKcfwlnlXL0ahlpJfE0IaWVwsi/wxtGYfJP3Y55BF66I0h
tGISUQuY/s6mX0wATFujW0Yqom1dZmX6lONE8nR9Ef3Tzs482pfcS+542ieZZ8HF
4Kl9ms1GRYfaHjL+zu8PN3W+6TqjxV4xXlGNND9gIHyQqDWSD4P/vqL1+KUp4LLP
0IeY3KA8X3UmGaMnnNE9/8JLkvn7wLSS6S2HqfunIEkfuHSPOIqJijhiy7ZvRcFN
kyvQyk0X6yOxuzVMD9b8vHRzDzRJI7RPswBMbygIrZ06B39yvssKb9hpGI9bD4eQ
GCDF/RGZPMVZoLShoqUWfoKHxYchA6KmZomGxmqNRsZe6D/H0264/2++7CepBpXm
KDtdiAh6s0Dlv5X7aLxJZE7iOGYGO8FaApvs2bYIaPCKTXAmNH/u9/ErSMujmAwI
u9fIfCW02vJ45OwrcFCP2jxgHNMyY4kygh0YTA4kNRzDNA0muB1V6L8NXCSYQ2+d
194f1KtxB4rI0rJgXRrDlq2ZT65ZShmp7lRx/MxzlFc7+a1TNDq4ngEiwioRQ81C
6pmyGZwhRmoCfOHCrJ/ezJqtAf/c09Ii/E3/0nT0ijIJxSp4jxnetSeCxShA5ePH
eWkizPuZoWEOrgty1ZsGddb+ROloRysdDOE8uE8ps5r61MrutUMoJUr59wC4ol1B
xlpHa/gLbpFx/IXzHIPrzfPXL1pgj3myVPxNMZzMOLrV9y3F3iMo1KptV/1Z9mra
UcGqryxzzW1RHOT8mIsr3ObSl38sTLOqpMaIqCunbsZSsviAPbJ/VWmaPDeimlZH
6SHkNU3a6CKZJdjapKCHyABrAbSv9kCO98GIonNvRXkvqz7OPZfZVJv4blScr9m0
EEctdRfhMS5HNU8EIRDfves/WN+LLfCkF42t0L7hKmHSzF3+xwAV55FIfOPhOE6G
o1jPMvXHFjRb335dOHI94n+OKfPpz0OkFyKRFwZimvorM/FyW0MQdVgip4BSHGr+
O2yW6llbcJ1ojsy7gKq+oNGw5A1ttxXP2JpMwqiPuNtwBIk+PN/reA/suCZUUimZ
R+uFoje8yJSzz6PVS9v0rEer1cprX7PWP1xFvMmSzsNxaplKdJnHPp8KIs2uQZq1
m5Cmk2IBElXfIDYWEfgk0Qbr7MexVa5nbJDemBg7LidKZGZUr/y2/MgUnI3gBKzh
U9TQxRzAvDExjqhjP6GwQbpY3KglD3kguejg0kAEtwNthmjdpLLzWrDWlADKIjPF
J6SQYSefxQH3Nmj3WZGFkdPbxeLvvnAmdqOTRv2/68IRdXjDfIAfJPPnEUsEwEFi
Y2gY3LvY+HgZ3GUp5gP1bwlmzwYLT/7Xd4X74hGlIV5+P40m1nOPHfy1Vx5C552g
s9FSXzTjXiavYNoYNib3L1eUT3mea+IqBDZL1km7eHkb/9LZgRWngLVLeKV7in58
EZzUYxK0uD0kNz72IMt9W2NBHQx/gx7isIfS81PanKP0HlNvf2FlQJ/usfhT+8Db
b2ni8Wd3evP3n9wBhL4V81+2YNQ1gwq46X8A6wsQ/Jw4Lk7fu3Fhi7YuXzqFpMjk
ObuCrK2FGpPihjhyzrEu54bM5k2fb+m5H2zoVWH01mDlSleNHK191U2EHnWOSx2k
E/FrcEBed17e4mUvD0lmLHeNlzOW5NNBJ4ti70eogAE2X9rH8Oo+Pf6cT44rk98Y
3zSnQiMSomE9xrT8WKkBRKpHDu+mtc0npYmNqqkM4O/k55P7yzwg76dGIg3FkDUx
tUNf3lyLtjj5Rsey6y6pAzjf60BurRPet8lEr6fxAC9Fr+HfXT1RLrs/SBx87mmg
AScBf4C7s6lPNvDjv8yWu2Ta5Y/6+6C72/zUlkGb3RAsg96zbA/Z8110YC6MLhXp
hU2BwYl1dBoREOCK5tY9853XkvjHgTN243lPmTDsGr+pXNwUJf/zymz/QGZLN4hR
8Owkxxo5zEpOV25aKKcTiK6hYpOx09Eys0PHPQ3Q8fy/QPYc7WMTGOXuwdz0i5zW
P6BlAKUrl9zm/CHqO7GmSWzQGysWCi279eML3HgHViImKkvN766ayTTMMAZzrlKC
we0JtGdDTxBcT+Pqswtcui4etneeBBGzRsiAuVNb+dvGsNSpQ0YtO/RtijnmIFQv
S3nRFQPGfwIwlL31XBAAxqm08vMgfErtoiuJJgdsW8oXv4CMoL5STLGXlT7Phv34
3eN5Y5ThWEaI9VesHJVngdb74TUGarglbSd2ybfsTSBwCncI2WzQdpd3fy5Tr+ol
EIZtPZzQUhidptmf6FGX+Aw4hW+X3yVCZcFQ3SGC9Rsx4jvbqK+UiM03LulfXqEi
8TB5gBuSgfHleEBvh8FeA8da9obOxmWWuem2rCMaJ4wUbJI8vot7gCtUkSEJ6mY0
VDQTsMIML3/ZK9DJtjNPZ+HsRDT4RZde00e63PZtjgzznLbYUiJ2h/dK2yeK+H2h
QNcAdT4m1uoNzI+IsEDXoTYu8972cgLiqLh7MXxDA0YtmS38t4AK+opcm7DQBtSi
+8q7ycVUdwHp7OEf/AC/yqgRPS8UYksq560kS4CeojtFwwXYOz72Wx08uL/rjTtv
Qrv2Eu661EWzG9RmSjzwHJgYkFteKmH1fOZjgoMesT0YgwCN+sEFHFe3bjTd0UCe
tFyGV8LDgdQaUWTN94OEey0j1wn6HNxbEA04Pok9VPGeW6XYiYBe6EnxszspKGtP
L3t7Rl34n4YhTq4QUJ+drP7zQjj/wGRjjW+7H4g86BAk0oFWVcNAo9jcXjDydFOG
RDqALnLknKhP8emxcx5ZfLkJgnIEcpn9lPxHhxZt1ftzEolfbkSY9H+RnPru/M2W
vD/gkYMmjPrnvgJ1elyIiGP1Libk3r7uNHuqYRriPYRuAWr2m9109uIHgWaLddOi
uFAl9lqpEZnVm8fHzLd+arE/iaxiig2BeYxUPz6lh6YDIvqm27EqHiMz8ia0GliE
CMloE8cbg/Q6rMJs6QUClYs0TSkT+QRV0+JTpzHnYO5gVSTgZkmVwpr4ixLCciHa
bDMEdbSmUnzGfN1HlSe2x/pUw+RRdBT63zR2DB19SiE/kYCEFOE7UIjZ0eGMOpUS
5xdCmymtELvc2enJPkLAtfLZOl9f+USPsmH9lj/1uaAws41M460gCc2k1AKW9O34
8dVohTIqBNlbafpYDnycvbODcZjPh3I6u9Wb1Z2PIHmz55S4BIJ80fG6Io5wOOVJ
ixP9zYqSmosCkwARllah7X8OOhc0/9ZQRAyT4J4VfYVD64W4M6BmjNfwH6BGw++2
OejubOUaEpe8wCAGPSoaK85HA4bBPxe+7cERnGw0Uw6dCsJPkSb2XdrctE0GtZKi
nmKF3cJkScCCrf6aLCo5NIkAd6riq9NcVMtv9ahazKL1X3EHqai/W0ey9IpoKdIq
9xpeapVywdMwiG4wdxkGGNNE6rSz0rurbjAVWJNFp63YSlq9FJhv02wc5vQtyLN7
+v6h91E3DiM4KCUGrtUIb6P3u+uG7F7v4IFjLnjyG+eC6kMHqvBMu9mNUEr0GiMC
FPR814uH/OreHk1aA54EVUZjajZ6hsFI6P9n5PkTWDXSfQXFIMH6Bs9d1uvaNXbS
yPjRpxNs0t0WxuagsMpIgvQda6+e66U0OITafp7XR6WIngMn5ySt1nr0UCETe5uF
JtZxrLOU4YjkFhQQAzJb5khBqRrqv2dUODdIbLv1Lzu0yALqs/dvCl4uMhPwmxrh
4UL7CXCpMVRdMo3J7ZlZCldFWDQneZLf5anQv3uNpIpC/CEZD7jhO5HtBSp4Bwws
O2tSM7ZlkasTZ8rljBbjopdftUyXVA0Q7sUHks2g8ZuxFekEcXFtMYZ5gRtDu6GV
6t1THYBjMaD/wTdzbSgwwI5IXdwtvKMqCBEU5iytMm22ykSceXvcRd7SPzrwnGcE
QFA7k/TYlcpSvG6UCkg9rbKuZlwnDkjq8DwxX6UN9JqvKHvFeLvPh3CSUBeNGfdx
zuJFokAluFCvJgphhOtjjiKPp6OVq+C+KZnsDm9ohR2rr3v/W5JzB6utpAfrRFh8
BcVUXx6vP7AHkhvZ9ekoZZq0fnfp1wXMfUjvdC6s47c4fvoYs3E/S5tsHrNxOU9Z
3jmlo3wxsCHeSH9py4woudq4EXwtbvvL6a0Jk2TooLmyIkJTHMLkOLyXsmakPIBV
1g+Ne4rLHPRgVRE9Lepp8iBQUg5b6XfN4VqIqjkXUyM1p/SFEMkK9bq15SIDgs7c
uQKgqOydqfIlXG5OdaOR+yBMKXDWbpnbaom1PtVEQbJ2U0h3eDwXaG/9VS1QaPvY
A4Q2unYq+x9IWsLOdOHvr7F8ROjY6zkLb7dvzDw1lIQWBXQWBoxyq4ZRQKM78F8K
Lc7PClut+3giTh/DGDXTcgWOw7nfgJ6haM9qkSwitYT1DqWPqw1Nn56rWNi8lDMu
rduDpqw8ltXw3gTByqqii577pJZlWpqpZUMbUBFt2cY8aU4jNRRR8dj76f3NVGb9
6K3QUw/S169sgQni0ZFue64/8isVbx86M7/112w/U7B4SwqD3FkQtb3yFXhZbfeF
ORgFcCTBa1c2+bmLJHkGgk2sKWVuizK0U0Sbr7/Q4GrZBt4R3lInH7vLJXyeojAX
MBlN3ZSLIba1i/oG3Ev9EjL7ba18oqlRN8lnY28qe9XERK2z9KJa6ri9zJMObs7S
YQ/A5mzrT6BuXOd9bSypm5FMz/P48wEM/RzsVVYgAYvrPAvl7tBDgxPQElI3SR3I
iEgXjqXOFfVl9ef0RwbjzMbPuXIPmELDl0Lq8+zQybJx2rcCzHI7uKWOp39iG8PZ
Pxfp8oc7AWTYxtVb0617vI9szwmqU2mUyuwvUm3Ka/Uq/e44gRa2lEQ/4Ylk2uSI
WLWHZfFKliAY4/p7O43WdIaeyOCJ61nakjfoYdLXdftAkjmOP+vRsij+srGjQeYp
HtzDoQx2UvsfiQjXjuXVT4/v+HPwPPAe+CzpB88V/IvKQieU5c5NnFI66yxLiaiY
3PcFYvaZyLBILMG7n+ykQUZ1SJDfk/Aqkra7Justre2jtWVqzu1pR5SlExn1gsJl
47ZnhO0XfQ66p2CJhwnXLUzdXhilU974eS9Lq2jWV1R5jyb4wWh6t5T0BhNcxigB
L0gU0Wty4e32a+Dqu0Cybd6FBBW2A52ZDHAqAJchbfSdnVMm+JbVRDngok1PqrSI
YYcRQr1UWVNeP1PaQbxw3genWMa64N7t4AD6Y1fwowB3fCjXGFeHpL08tI/5lAtF
l5ptuE/TQWducPCg5dFErfY8QHMOTHiESjj+T8Tqunc5jFMcU7MR3j2w50XliHMc
oGWhMLttCB9lBOfBj5tSoRYYK6AjAz4RwCQAXxqIgUL1YNxP+HBbBVTNNOH+Amoe
/78V/qzQnPoCQ9C8Hvwy3VWfUpbHgD8f0dMslBdcmgFc3I0jCrjVYRXOfsKemxn5
nKngbjKXPATwFlGmJJpmRpbcB2ckm2o3HDNfMERvoJg7Ucp0yKiWfkcEJkiHO8uH
hg7Jv/5ckffiiKem9aKcyQELoE6+Np1ANvnt61/lAbuEMPBFaE0V9DP1YH0eXtif
JTedZ9e7dwC6EzjKxnDK7RCjLKGMeZkQzUfiDXaBKYhr69z898z9RXuBnAXJhroM
RxnOR7mH5jUhIz1geFxr6KyJsIG/z4mZYiXUKl45SrXS4KI2DUu+PVUycseTTAEe
RT4bsg7XI7PN5G6TkNJxmKfLSQQHFM6IKAGIi6LsXnauuGvl04ZR28o113BNJRWt
BHoL4VmnwwyCtaKcwVyEE6scDEYrhBQz5ATYw58pjrajTDDiEwrpTwIO6W6gbdAf
/uY25ovIksBQ5W3DkHafohnjKZMDdy0jKUcZOZ4K3sPXD2Jbp4yzzAWJvSV7We3M
NgXMdjhvBkIQK6xabOa2bQNWx/+JORq0y01IuWYzuKur3pWG0ufKRWI6k81hahO9
KOHfE00TENwWKZQu5eaoaRhkT934vABYtSaChTTEkBSwMdJDitSOaf/IGIyhBSTJ
BX95hgWFLB2Ii7wDwFg4Zc2UkrpzIRR9yE766xeKE5BhgLT84sq1wThitFVbzJv9
J/UctQnlSDOT94EVYQyO3NS82jpOQaimLu0R2cLRpzy1TvY1/oyWVcITDGViOFu+
hWEjsjpcyzjDMXKC6OphU6OJzmACYB6tk3rD5yvB3c2GZuJxjR+KVtUWwuyJSuGL
MHv5Xm0wblJA4ssT0VZJ+jCvgdBWuOALqFnmyXbA9HZlhkWNguwglaxiOhn84LE9
jmuY+hzdLdCfGlCUZpoX99RoYNqvTzryVPhCeqWJGxhlL7aa6x50zp8sUehMUB96
EoRNcY84W9ggXnscKTO/yg+bRz+URZdeKNyjLXIf2/xuTaL9mPAjbYUyi2/CWiPu
bIrvRQaFSnM+KnFRcoyrMMOLdQbgutVg9LwyumdJbhaaxrsyRoS1Xc6J9tD6f0Nv
7fmjgpenMkycXPx4guM1Fb/+A24ZnhRrupLWpj17uslEhuuWy/d8zqaklHWLvhXA
dQ9+Bc+z3Pss7n5B60LIClNiZnsc5sfVK9aukd+dTVOv4EwV2fLjZiFCLWSamCH+
xi7iAPHxm51FqlaMmYy3V+q1YAkOk04Wx3X+hrxC/d4JWdvT0PFPCOEI1KvZH403
xER8qemetiRc4vFP+Wx8v7d68a/+H1c6jtGemhQjtRWgzQYKYASeRtOJLKAcax6J
0exzzInxX2424z43KbLeDkCWKgewFLMbXO6KmHBP7ENDOJBjWF564hwTzb/CTF6g
y8tlbEDdduNrryDgCv8yx/XkNytGW5Q5nEB+1seRCf2yPPmOcGpq02yT/aP7PE9I
KZflBuJiVcoM5+ArVyKgOdZmTTmvCLhbJydr71iINRTHuqSCZpvHuXqjpPEdnMRy
Ms3KmmLYnoQgkzd1wOTrHOGp3O0nBnxmiAAB7Jbhyer59Jotd5Q9j9ELoR96m44c
rXpOCSdZEUia7kyiIdkTsmlVBOrqgTfCJ8zEeH8N6Fm3ILJ13fBU/VBrvwDIit8J
H13S5BEBz59KFw4c3Mw64tXRmPKX3KILiBSJ5YhpdXDyEKl0Y4C0wx26NzzwwBfs
zvheX+IREnFMk2wBL+nD0qQD5t+Rm3tYIcgyKKRc/giS8/xAiMFwFKOWFiIf1DyT
tvVI6QSw6/2X0WcSrPFNziYz0E6giKOWyLn/SvLAaxYykuSGixemkmQ1jUgIZ49N
7pFgSlBGYV7hADGk3sxtKg==
`pragma protect end_protected
