// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:36:48 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
UOWuW10WxgpNpg/1DhYWaZDouFCZIF0ihEyeZdDGPWYpyI0vLpjz/FW1bFMryLcm
XREaxTsvddiWJID5/revf4btWaSMXp70DH00RnsG8sAA6ujnqXrFiIfg3dNxO+mD
8ohMuLxnIFyFE7OdvwILNIrOeHYZfGQdF1aAz3RY0Ss=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9184)
E+p5Xs15gBzT97KJVE3gNg2rtAoNEWKQwsyoloH4F2crCoaPIlNxHlX8moshQFAL
q9+Gzg8c10I2f4chG9+e3mK/xww/CSDj68eZqxwkyeiDCPNsGJgND5vJhfiXq1ar
kIJeVJNKwEoGmrFtzQ2IeKPgJPdUzZhEYykxuhtDS2VVu1wiqZqFLCk7IkvcaMw6
ttq91/P4lohe19R1lU52URwCigbs5CqhY6FYLq8UI8OJ0XCZlYTWrZSyd503FXt/
46qsumEyt+rZmsPGpFCt5hLLAGKqYgV8Se6JBIlTzjOxsTOQnosXNnfChuGS96IO
I7sSOts5gksfPOwp2tQhdK8BNnDKHf9ustYfBEeeHBPWgNa/lpEM/kgo2buSeEK6
Vq3ww2tPy/DHNQ7YbKawDnMY/XvHHwpT5zFGWD9BYitUdy8tIVno6JMwhtlUM3N6
McLnL1gaALm9v8BHuYKxm2kmlXpNwBsVMnMrcgtz+3aLYEjAeuVSVcBLVahuCTp7
g3bJOWWgEQe8ii+AMjsK+jWjCxe15ky/SGiaYtda8pTK9FHTyd0Y4e8sqdR5b/37
hW2AOMfP7TE8xZQwifXC17Ua5utD4T+D5UlOjcT8PVLv49AKluu0oVJZOecNMx9O
cTvEDLs+k7XvVDASh1zAm7T8GlZcQqSvt175cVQJIMJHpFQnRs6UalRd5tqZP0hu
myfEJOcXGhO12UIhoiNzilvr/XyutI2tVJ09Tj8rELP2hk9Wl2dp+MLpdRNvUMfi
/k98EFNy3aGR5aKXgv1mW261bWsixQGA8p5GQKpgW34K9XNrCUtZK/x17ad7pP+5
SKFk7vVkNMjgnUm675PLT1A4BCzLb7TNJW8a15jmH6q/K8nM0QVugbIQEVvrl9zF
rKHNLmPMjtXMsT7Ak4wBmepkWh4RLmESfFDOujdM1pYGTLqJ9FkXTl1r4X348gvK
IZNKVUlHgKz3rycBtLaWPIWjPnvQ9optj5mceuJ8rK9Mtug1jcF5ZwuAxivUle4S
RVCrhKy1xF3NctaAl4YQoZcpmnCQc028xi5tRjZKQMckmeYyisQEcRigd8Ci+nuX
2DF7TdJvxca+hoy2mIvgQvF8pR+0+xawE4HiX1zje1Ud7ejTCfDEEppO+ti7pl8e
ngOnp/DJrHxrnEt9T0Y3ox44Wkkx23cbmhTbI4iqAogvdNbHCmGLuH3AcH6tJdVn
9DMZJDP0DAse4FtLyK9joxmrwRBfnWAKwS+hq22ZWmH9uo9Klq7Ld/0mBNRVzKrW
OGWkpZC3JrxAO6pMbeYTpNtwvRi3BGS1GWp3cx8EHsbP9CbGL0Ztk7gL2tEpqrE0
YzvYJLEvoL1U8/J75Gox3KV/x1Fkm3JP15BDFz/bw8/AFziuUvYllwQ+cCvyqM4d
HVN1qX8B9Qx4kkOjLdBzrFz/yaFIgBf1YHbrj0sEkrRDeR4hNm3VABTbehQMKtuP
BkGKGVCkXxZYMvUsdZuzb49NVtyvA9n7ATkt1TvnUL9ML8/SdnkIa+WqPZ23SysD
CJ3LoqVGL0WNQ8ZGYJyxxGuqAEIn4vapO7wEBUGw8vvbKrDehElLpqhsfxpC45Q6
j9WlITWxi344LrTTpjMYItax2HkVAtVNI0+U7f4Ddpq12sfozW7rg8WVunx+JhBz
1gsIJ0eKgPmvHc8uBh1UrQMGPSq8EacKxXJmgMX5/WsvRr09qKYEnatSkPX862yM
KCuaxkQsE/M3AZv4VThkiyLMW20PcETfy4Ssuyf76sS6V5rlZeS/aIGep+C4adPK
66goXL937RZ0pLukq36MA5hQDKOz7AadWn8ZmfWpW8+pjEb/Or3cTmXQOiFhjp0h
kIJP7p2I5RqFjNqTBL3RZoPZV+GBLIZG8BuWkDUNmG43czccNQTWL3+3oCN3Wla8
jGijOaOAi+HtAgBh2NMRh4J7CFVfU9McG/Y7JqH89h++Dtu9WfR98NVRWrXFb/P7
fBrOXv9fhJO5eCksLH738E9lED7TeokTk4At/xGUb69xvP5KwnPMbi91z+AU+CKu
A5MR83dm89YYRbmTBikZ+OPVox1jo6yP66+HUYvnhGKuLJ/QNpaB2vXEuvvZJy++
duC5GyHOB9s/xhwbmR/B7AgOPIDsrCZzDOlirtvOBVWdRkRQ/vzTIZ5kuhQpyObS
/5Wn6tT6Cv4N8J3QSe99rkmyO16ZaqkWZ455jgeEPhwQHX0xhs19w38QK2ut5CgV
C/fJQVJ8H0/V8VNxfWi/Zuse+xVUWmVxo2dd4weta6zZkBS4mAW9NAW5Px4IL9L4
HGJdlBOcjxMB+62TKOtEsXnMfkz6lb16aKCYqiFt5QW6qKojn2YcP5URpn1uBTrg
g4yQsHhjPiuvfTaPa8GxGz/toh2u8S1gtt8Hvorb/vdR2Q2bCzjNOfEPEmWdZ7rR
aW76kHdaykMoO7y4ZxFO0GqgE6sKlJX0L1XbbmeMJJal/tOLooqYVpjAAjULXNVg
3GiwvZ9VcPdKtsQrZNR/bGSS1sAXluDybYXDFt0wf5df9gIx7B+7BNyfVuo1/8vz
LBJSh6GNF4C/49oRV/jyDHXMeq6VERBJknHZ31rhEobVy1jiVMafHKs3oM1Sn05X
cyTbHBQoH1Hee3d5SDl7FrLBTRLTvPdLxj1IQE+6Uy9tMfMR9b1YKwMBYlzWW/Af
jiKE9u4S1oVhBa0UjxXHuM6onLJRLQAvIAPFBx3/KeC5OaKRx+fUl113T8MoM4qe
6xipZlUFGjTXNxUrwC9Iys9ZUBKKx5uqeut4jDhGwJb3ZbR0iDlQPrIMZv1g/pIu
nXNpoLD3iTvhEXvCo/mK8KweVPqIQfDlw4bqcGXbdtW4JLV2N1TSERD3ZLU5TKrk
oASFLwxErXr7N0vcbVqjNnpfgK1wnyC3d98X5wf0u9D1EhsykFfDMyBjyUB1kHrg
gJO1fDtMCXmsr/qReSbAqn17G2UWFFAVBs2Brvmj3YQXTNfiY0ONP2Qq4+JazlEu
tQTHREh9m9dtZp/yjrF+dCBmjG4X4BalT+kr2wHVnR6LfksxXlSo4elke5gU7D3+
CFHqbBDIf7ZSuAGX65HQerXI9is6sAtBb0Wn77TNIemvTWVj2K8PSfQUiT/9SniB
gv6qy+o+00f6qV1gFPu7Ols+tEHw+0GDGt7+92NXJk8FYJtLwgg+ssKr86kEwCaJ
qvuQLJXc8NIXgia8gbigLcaztXQPvmDOh+qhpOad0ZCBDj5jhiLPu/sUzq2OOur9
NYNmYKxRYNV3UkOvCtDnsE7mBE5XN4FHk8FpNuEcxUg760e+MRplhR8O0SjdUJv7
Y+iwHDO7+/3RyghFaKJME98qajHhUjb9kkvIC7ZRBk0pCd7Fs+CObTpx9xtqGDTR
SYWdFsxfIFzO0Lq/4iiBSyVsSi6pXxgHC+5il2ofsQmzYU+AC9vyvloeM41aHoBB
b/c/zXvC8qu4+odVTTxFa3CNv1d8S1XN1ItUQTOxYTc7KdZWeI2CVzhVbkrAPt4C
LygflpLUUBeeNHY8Txja5PAIJw1wXFbs4c+ll3Ar0sQ8oHTSbV/qv/CFyyOdDIC2
3kujQxP1qSmtWB0U82dVs7dbBkfM4abH78zVCDDA5skxpDKFqScfFxU+KTJDsDC4
yzVVDTotj/mIDxII0Jl9HoBHgEnhYOG0qcFQxgZpDbQ5FJA2j7Xl0A5WYcLjeuRf
CfMh+DY6seBmkJi8+UmIzqJzuRz7w7ccGtKuuIJJ3VOMcXdpVRtH0d1FMbP0BEJK
ZCSmddSwr1QwJBHucu0+If/h3HSZ2OESf+4zV25yRHvC/4vha5ppkMHpANx2l3xU
+U6D3qe6N/Ate7hWsV0a1cIihnsWTZ4d2Dhv/ynrvPbmdLFwacQgr1fXgDEGjjZB
zu65fX0wIx/T8+ivd/C/aXwaBfsD/WfOQZsOVpZIBQCz9J/kIeSYmsZ6nxKhlKTv
khpgWeJ00ICXnjyFxg7CSgQuVnKVrwW/6L9ygwWY11M4jvD2EDlu8KQeR/CwRG/W
rE1+ndh/LAYM+l8xP+RjKnjFh6pa5vxFUlRBgcEqLqF3Bjb6sMxtpnf8PHKxQNIM
GxkHFJuuSR3HMrmdc0jYJcHt8X88oMrgP5LWueTYMq43LGQZRYw5WT4WK+fk9jEg
jq4nwJZYdLics/5Rf0m9Nw8KWXQaylQY7L/4XSKHBMZ3xvWgGePl7jBcuX1Jygeq
itmlQafg1MHAFyh2jZVzHIxZ41JYZ+U5cgilGCLbRPzB/pQNs0A1/THlkyKF2E+j
YM5lWR5Ic21zSdsbYe6ul7+iNuVp40DkVGCSYNeDKBQVbmn6s8BYFGbu3yIPyU6V
VA0oanMcNjxNLA7iCuvbE5BNbLsQSJPQr46XTF1RFPfrf01JDteEREj1xDhYAUin
UMuBPN8IxUcK2SjARuDv3PBzxmhZTF7BGTIiGw/xOmI96lAjAMRddI9naZJI/hMq
1lIR4+nXzL7iwzR5rqWNpD/CoFJkbAf7yD/tUDD0LvNP/I4uWLCZDHzGqwnAXNwn
6PytZExG6jEGg6BH5Ezx2d6Px5OOl/qu8bkG0RzCY7h/vNzULLHYnUYDw7ZN4C6k
XbJZUTb09fhkCLASDQ7WxH2zJ26iKVHk3P/H5S96wydCUzqlgB7Bs0BhHMiXtu5E
QNWqGEPTkp5GQuHeYjCWiwFWpK+TJ6TBszw2lxyWA2lAdPAubaSgpxvZ9PG2+weq
uI9RgrIevUNQEC/3nL4oaxVAit/y6NpTP/1akwCN5WCnR34ZdTURf94KsZ7eUR1E
SQ+yURuoVuLqkNgTsnf+hE+4aYWYm9FV451DDbaMoQyyLrT/+ieiBZ3u3cQMeMI/
6OG0L6erzNz1Qz/WyXnwWXcfWldDkmIs3BV+gPTstEoge+JPmXg8vKEs1YSpfuvf
ep6CbfIf7fS9BAzce21TGMRSZDEjdb90WOBQ9yc5MZ1aWF7R7WGq+n2DQkRDQCzf
Q7um1cpT44/hDDI5H6lm5hRIK1vYpz42H+VvYJlNH8MRJ34KVXH14jnO0YEzRY4I
69SOKdj/e2y/JSZMtnkUuLSaD6VgDlf+R6LzHDS1tmVgMr3zoFyBtTtLzrosVF9X
iRuCTm1/UqBEePm57S650fSOC8rgffhU32eUBJAwufS/QlyilSAZyFqdaiKHq5cp
cvzuD6bZL5jPb9G1UNEJvtXwxs77dioem3s+sJagSxAxFy6WAv+MedI3Lspoez/M
1ywAEpk12w18U+ldwqd2QEsG5vFHy1yTrfbd9ZobgWvMzFBvqbxVMb/t+fWCAp/3
JYs+Z4tF7TjKTgnWGftlAWBEPRZPWbT2Ca43asDBybGQTullc+H8ukt5zvxJi+1U
ysjPOy8Mh79aAabDXkXb8qaGlPsrHY/zpbjUitZ0uCouvpQMuJmwd/eI62Giy8kT
dCEkwyUhZfhmTvZMKTg1PgapaPv1lepKJOv5xDSgZzg9sVXyZdXbRtDdrWR9vYj1
ZL6tkWgja2k/8GGC5z04q2wv6bvnGYgfhS2JLLiLhoihu9FemFFvdhTLngXWuaRG
dELaBuxlkcCvpM+zeclqm5sCl4pNl5NDitGjDSOgpzdeBxv1x/PXf/a1zPs/09eZ
MJRrVJQW+W28Q007pYMCDD6FwVF2UHOIF1WjpJtMsl8XwNMT2XmyCKtDG/M3d8MA
FUKy9bYViY0rX+Ahh1+BkAygLDAdSV/wtsoLOg2+nC2EjqV9tog6g3EFp82qrz84
+jX2xtWsD2GMDvGuUvOoGZRUgArduDBqlBjg5Z1NPXgTyU372jmGZ0S7/xS15xBV
DfJYMBbcMxSru+mKW57h3Bt6jU+yo4Kbip0sIczbaksbR6nrFltiiE9JNcwq1tp0
tMqZt6BF/SZZaXn3D8k1qBkC7njmF6Dsn6YrcOKT3JcdalvxP7cRcvMaK9lfx6RU
uQTeZMVxBGf9Q1Kjgn3jj2/3mbaBLDEHqh+JLQNPvMpfsv//SXSNhwle2rJYXSww
BD2R/YCw1v/0NEjLmut01LvyG6oISMHctOxSgYU8yTmb84qkkYy/inQ5IUACOWNL
dkQyBfrROZaoWmSaNbQYHkAiFn2qxuWSpwqX0Qo17kBk/2bl4OwlZpc6A01P75fd
B7RmW0ShOBchLTAz5gbfy6QbINWJMeIEcRne+VJ0BEULnQ/KhfIrQBEmNyqgFJ3V
bC5jc7Ov5wg4Bl2j9ZtLl4PsPHwoamVEZTeAEL5yaqTkkY+ZP8ndhMVVHwPL09kl
si3A6RgfWeEMPgRqoHBT+n2cbKFeU4pGCGF6ZaYMgsRwCKiiC3je8VURkPfBWYOE
0HMNQhz1ZZNdQpYdlTEC+3+eHjLil7f4d2L4X7mY0nmlXohoUoH6hgMUzYi5iMD8
w5GGWDaSf3Zqn5Czhjm+RF9PfbCQSsw5VeaOufaaIJKTrYMaNis85bOlb6b6z+fo
YN5BNc50s13vZOpClb39wW+e4D+HePyoXIP3D+nT6cVBRW/Th2bu1i0BquKlnR0N
/YrrFgdSwqFQOm4oEAkTCn6sbIHxWqq7hHVkTpRdPFD4QUDxCEgRra0Zg2Aau0vd
EnepN1cfw/4Kjg/IhMU8o6287f0jKqXsKc1Y07cxK2TTFXtRVYnVHZY8aaGaaMwg
YWoXb9sjgEkTTMuRmESHPIq6+OqfodE9PGYPm1dVjVds7knkV+5OmvWllt+nyzAe
oMq7ou1nweAI4cNZeb4WEAh4wFQqS/wEAVZ3oVBJm8vSqSQD46LYsN8+Y9L7VwDM
TaM/XfA0lvIN3xL8sVIfECcvuJktxwgsf8q924VTFlDPWwYfGBsO/PCEJDvtravW
aOiitr90zLbUbF7IF8K/bnLzccWBHIESWaFupiCUN1eCWtgX55jDYLEmjXFvZ3JF
H18sJ+TkZrLsldDYoELyFYfAxTGsNKYjkKlEzNVZ1h0PhGxQQTwGsU9EXh4oZ9qf
W7bX4FG3/sO+EJ4/aambN5C8dStK41EGiXxs3BE6Wwip74hsM8xrCsHS9U6GUOHC
NIUicJtUmTPpeUYeDw7kNOXcyv45oycL9oxjz6nqoM1EsuGW7kCcXCP4RMueZIH6
9BAwxYHewJTKTir8oan2B0GAlRFdB9H8lcQXoDYW/OceggdsajViGkqpYc0NBO/X
Gdguz2spz4mQcrhPERs9+OyMlmKjNc/2RmoUi/QsRvfZ6xw9fqzs7ygrEm2N3tEG
KeDvmMTmr3AcITE71ks6pSVmbBjuIqeW5h8LFPTOMgXk673aYLd/R5L/ocZvDOvL
euB92LCiVRSzN/J7iwAOan5Z3AjhsMPj0TeD6Rc4ZiE5KYkHbhZA++AN5SyyYFVz
x8PDDUhZN+1W4R3N45KQwJtfZXJljDliuqVJNdzsONk2hAVVEEPri7RBZd/mzB6/
ZQyct7To8ml9ZmzB81yKZmFZB4Y9JOP2qnFUfMznNfH7MsCs0DDWJcdr8s1KRXp3
VyMtC0hhipqPR1l34thBdCZVVByzX6cL/0EklCay0IOkmhbFXbj4R1KYzN/dJF6d
3o7nggLQFQ73xoRP7GwbxOrpew1dTHc/i+w4oXTpawMgOn8A2aMsK1ZFKROz0sFw
IREDmzYGDdGoWB+KhIdOvNhuTYHp3JeRCawHr1lrBZq3NKaeYFSxRtvNyrtqlHxj
KVblwbbIDFO4R4Viy9r38ixvTEdAht1b8tuCb6kA9nLXm4fw+YMMmwl92dSGW3E6
FhXu8PsKuozcxkvBvLTjyBAHZ0TI0h5TmcfHfyZnbh5wERMdWGBV1WVez67+KmbF
kBK6WzCXt1nUY3hWjydWtkziUK6z/IVspI0ZHeSfYN8EJsa2MQT8E83M6E91KdNh
nfhaDHRWs5wVRsSbyeJXmjXrqNSG/IsgOSIvRoqYDrUWorAijHFfr4vD6bfp3aBf
aC8xUERaZjersXK9sBxBuD2v/oxUO6Drt4eXGw/a8tvK0dA3rtGFSiOeUt/ZE9Bz
SkNHcSLPqdhRkcX+sy81NOxEiqfDKv/2do+q9Ikt4SR1z/NnHAMRmQnBUwCEdsnU
VsIDygW2Jm8PvKfOzYYRTakr7DTwUc/axZBcY8PA1PNyMPlBg5HsT0Tw+mE2Verb
WSTnlxm8rBwh0zcJLYJSanFNbEjMfax4g2eZcfA96xeasG5kqUZwJ/56K1h2JyPC
ndI5BZeejr2GQcAKqnTlfCPB3GeDM+QrmJSLpQepMAt2UfDj8liKU2cryDTPJTjO
F41MTvOpwHMd8pgf6BnBa4fJizTPerr3kMwgJDPV6dI9oEIUjd8SH/loQR9dTLAx
4zs3LDb+luxIQcyHMlaxbUX9ah1YAkGfhpZEpv43EuWoANhwDfUJULcrA0QTanAF
+AwvM5EZ9ern5abDY99KKr6Z5pOgsyLh5oB/X/nuI4jPpfCrnNs+QQ/EHlhJd4kb
qVk0qyvY6i7DMOHXPOI1J1PIX8dPD448CMk4aA+pu/O4btRG4wrNFFoojC9lh8GN
+b+Mv7QmrvhFmnzVkMwp0Oo7V0agAYHIRchvfOZ7sNnUyT6kByxwGHErvvG53mfm
NJu61aEqRsqInyvGS26ashKORNqM9IHxetYlxMUY9laY8mgrDRJGWh4FH/6kpx6R
BUXtVeaN93YahmfLBrWxASYTueGlN1PxyXMvS0/ixwrTmZwdL/K2VPVrib6/Qlvu
heb0PRVq7VVsiJ/xYoinWh7SqudXZbjYbCgPxsm7sQjbeLtihlk+WRciOxiLzRyu
wRU2TApEkKogqo3vwLQMuT8evUdEYN8p+JIbFxRM7Y3x493GkP/oomr5Rbt/G4z/
YGNP7wx7RKXxvnPETeJqet+Ry351CILBpIMCa9A+6ezYY/VySSsCgFe2bTs9BrZE
owJ3DR7Ys1WeX2QQJbEhCjdR3mOwjj6VA8TAuCERpQ/N+HeV3ec1aEr7w24kV2Qv
vijVLHsD8w+nuuwcP1QnZgj1yAjIjAv33vUpi0fcfrPNisC1XT2HkvDFyayDgBD9
eCFe4zSEmZ8msJygFsHZ5q+a7NlM1JT5ESsoFc4P3fQO+UjzOg93Gacv544VdyzT
fiEhgok/K0Jt99IdJwRNQPLrKaO6ldlHZH9i8FM/mvt+icuFgSgX9FJlGnTFZDF9
SRkNwfENue0b2yd3vdJZNp9kfMEFpTbh8ojkBeJDnl549CSsjjN8fN3udZm8ycBG
vU6fOrKM2Hq7Q8X0D/b0+1EXqv+WiGsCpfUQJqi6RI1AvBqIt7SvgDlC56Aok6y1
JSVpVfHa+JmjESEayzq4j9em15QU+DWfbwXf+blPbYMaq3qtWplqpxPRGVgPNH9x
Viu0sNixsJktoQeNaVYy+StcmG9rjl2+4OJPov24hY+AS0e236/fepFaHbbV8VJM
BCAsRI622aKt5rbEpW7uYcuvhSpMKx0irXu6onIQga707OblGOkErkNRwQ+xxj5H
qfT2KGRNoJS+A0cAbuROShSAZ8jWqGbVI1qesBfkxcaXCTn9szpAgfUedDO6FqT3
MfLAlMJSumVDzMUAopV6GLQ7Et/XH8rtemGvry3V5MWtE6Ivw96BwYhvgTMAwSFu
ERyGEF32CB2msMjGunArcbdMlzdz5x5mZXueSE1TIO8BgWx25mNmOH29CaRw9fI7
uNsLT02cu8Dj3c+yDxluvyQJFfepxWIEbTDx70q1lmmEt0buox38TTlj9QJ0i8u8
3KsHUmaggFa7C+t/BhcDg5VxHBpSKH/3eyMyeOh7jqiOZYPZyOtus3coOFwhY1P0
S40k/tIkUhdnoun7FpKFdnxgseqiO2DoVHWowvfaGWyeeDGx55wkjkBRRqSTFIO1
uVfZeCsnRqlbc0iT2EfTqSrx9OO1oH+tX6TIX+52eETpTc5sLJrbVsvn19WwqxIG
sw4wZrn3hAt6v34cJuW1/e/m/fRusidQCKRSU4G9mWiBO1ie2FAKThDOBUAgKCst
4QF+tF5f/rbOLOX0i17Sp52SclCkROI5AwyXBew3maDsy15fiUrFiTZW92O0/Klb
43spVTHexHSlve/2xhieupNBG0cdeX7HEmjNf0PMtL4yL3sjsl8ipRorpvhcpWuV
mmDIkQuJzjmcbM61nF6t+8jtZJjHbxqGFS4CCo2H1GTtPRsoqvILreNc+xjjeAmz
i0EWeb+zlGjFQROuxcnrsi8ga+xBeQxrnCd+vmNmEB9T6z+1w5jnVfWpaYkPGzZI
CERKgjYVbn6hzIpR3g76trpWgez5Y0e9P2JPaMMQjrzIknUOiJsVjBmKbW0i9gUx
YLbO8cWDZrWoJCiQ2FS3b7tbp+bLzo3Ky4qQgNHl4iD0KiPTu4lVc8ZOcKwu5IbF
pKkdumDRZ2EIS9KQDU2s4X8XwKaUeIr1IJomp7YuQrvStYaiAOk7nn8HNUsURrE4
jZ85oxVmQFQiy1xfYKWu07PDUxqVgY8R1AziHYoqMotYBesZMJjdRQppQIL7elkG
pXJ9TVuF+kxb1+ElvrTHoJwS8gS2L041MCT8g7pR/xfFEHHSFkH/c3LUFOb2Yp95
MhGLLvDqVNmgGuI2aDgtKjM0jGoSNJhDfTkFPiiaC2s2BEYEkiUvcOZn6YRkCqxM
84AEqWepfhAOk0dyDzOIi12kQ8+4TD1m8a5IIuN0AWniNy+taniAT/+SrhWPIYNA
EX5c05iLyBV0QEjYnvoXPH9jQCNFeI9dKdX7x4uFJ31R7Drz3O8njYO0CCXZCoqe
tWB8XWXq2nGAL6+V5APOn3NGivaowcvW0aHilpBAbpQSl/5ZTMGCnbYkWfX/EC9Q
cR2GNB+azZ4YTYDohh0VfYty+4qZv9LEVptILMAsrx5KAFcgIwO0LakenZ+rcGIw
2yc4v9+exAV8Nu3bOm8nbdOaLkDx3OcsS3HPgzJHHch7Leux6F5wdEigTj7Vl7c5
D+9Q/JvrC1gnANn/gOBOP0dAst4t4xVZEjtaXvSFWuTI3JBoL5ifk1jYBAX2Chjc
e9MBlzBxWGTdVZRGxhaROitMs5mWtKmZQTuFmq8nfXtXCJqiGo2RxdPHLqISCPJe
ZbFJFpeOQ9j0/AXA5FZUM30CdqCnMTTjcdrxmav/5W5Dbx5QVKyBYiPYaJ5leC6D
0toR1N88Z/wG+1i8wQ8mEIMyM+QwvMwV0GngfZWxIneea7QZ3Xr7U0cCwtt21LGt
/uDi8Q9Jkfv6cisd/TvxKyzQvUU9r1CqZRcTu04oBuayyf/wjJp9FMz6eKVVLRWa
RMw01Df3Fgwsqf9girc1Z+b14/yYi6Sa/rfX4/nHRhJyV8zp+wKkLbKO8zCuinFh
dAnGhP5eUduYNahl403033aQFvtEfmF9DGjduRGYApkpMWRI2bht2X57x0Tm0hIA
GePyFiHArZVA5BDwJvl2gUb14QNo+i306257evb0xStvy20j8ru2psDKbZIAzWPp
b2Rm8BSl/ckye0Wp+5N+VvKESiwoGMWwYORHGAkx6Z6W55Ce84yIk0GvcF6yo9DV
Fle0DYWoHmTYpuMyStdWA5rqbnA/p/Z973wj3eFpBc9MOOdy8bvyuc1fwwa2LwSF
QZsG6i7G9lmg8FfxG5HaQcJXkkqSjf5i9kYeCt/BqdZsqaXRL9C0igQtxHZk3l3L
Tjzf1I2q59h6TxNaxqYjmevmmxHFZdrGSuaADhEoVD8aq2Q8qDUdzcH91KwdY3ql
GwHUIFJO7+Hjvi0vGoPGIbq/hLYAm0nwMphqm6lADkmWPjPEv1+l7moABDktr9/K
cROEPaiqWbnn+qXIr1v2SdL7NqzUQvFVj/88Jfs8BO81R85Odllv+tusQ8F8nE8M
tr/lGAM1BhO/uAAGEcxZzzGxNmYYlXoExGeUWGaXAYjcFYX7ClOPbDL5H2Gf5ufz
AyPsL7NQFpSRe3PnPewzY5pFOpMmrvVwaKVD3RKz9HaPv3umMuAsANEoaIJnCR6Q
y4jh2AvC4ne2ZiPQPKVvoajLGljCv0NjxLxfsdEFdXgEl6aucsXyBQGNA2PhJtAA
aWa/McgKUw7cXR/EOegUKgNCA3M1dnd5L1WTLhS5tfkF4URWgdGoqlcaSfOkKxdl
p16TT++1NV0wZYsWpbt4LSmCH0dQ459tbtWBGWfg2Q7NXHwXIZahdJ2ccPjLuPPX
7ZNBoggyeOZBQY0Jqtz0Y5d/GyFv076cOjcRznlAPU0v7P3dxt7Q1Pa48VgiCw3m
lfhLEGIAJJyj/fGM4ztpzg==
`pragma protect end_protected
