// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:32:37 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
AbAm24WQsie8bUWmxlZPSM+KGEY9YcEHREuXTrn2GGpDegCfQvItw3TzEX6dPFlA
GXSuRBb1BvrOpSKm4Q7SYw6lsuUY8MAQLRjdUiZfiklEFAn1pjHR3RWlNB9ecUj0
JSjZ+PUgmkeO+E5iucooRcPcpv6M5pckLVSNLHU+LHc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 22368)
frGd8rKqHJkNaKU4LQSB0RhXOt0EhaeetHf3nwyU9jRAlRZ0yItD+L+ZylbXdlll
ebPfBnYHYeEUI1bkUViKkQ3zRiPv+l9AE6341lyTQ4eTpHXOfEFwEJRdwxnFKPDL
XKfK6Yj3b985ZQY+MGn13qro5329l1N8LUXnAUcQ3k92MOSfi6vhJwXI5XVFwvnN
WsmKVFUbJiMY/vG7GGYoq5IHC9l9LIU5C4MlpUkP02kbeRbaJZ4aYR7a+WS2TMCj
Gltrzik7yfiojQ6lN8xs5X+cNQuxlMf/s0R2DDMG77mIt0quFu3vcO8fQbsDgXax
oI35dIQDvF9dgdYDJcQ1D0XtNm2HtL0X8aSY6D0hreeitI9PG5ef17HrBFfE+ZQS
vqg0JvfSuehqAiJ4e6q72kQSe0Ec7+T6pIREAy8wciAV/WsMKSiwC03AgwNkfXwR
lVtWZlUyHfk9eaIODVZ+n0I+dz7vhxkH9T8+28AW4FGm1iLpEwyl/qrVUxtw1kpV
h49oiiBypCDvPCUxSsMbD7gnWP/bFHPeKqOh8OC2JSJGY0144e3zLonY1oUdiwjb
4ZSgZvxmYUBSd9AmMnKodgBw5jM9MrF5rUHfv/qqLERrBjhRGwuDkfzE9cM3PyrJ
qD5bMnm70rugGmCTbgMXBNWm8pYSlGF5BiTxbiD8eGx3FLn/SCxeJekFmFAxW2Jg
8i+ZVbLLBcvorTVb7VLYjcCRkr0BfoQDjX+YReKK1dq7V9TVg+/RmWN5V5tp1erv
8CCvaFPsDUx0/uBGSL27bxvn/R1zB0eAtNQI3SjwmyFaZNN/3uIRtIpk4CtwLRej
7EAN4hjdX3iZSQnik739B7kqONe/eFzdog7cO7cFlIhbnPxmuus0ai5CaESL5s6j
Ju9NWigqKufN2R0GeDoUUM11ZbMPwMFn/yqhiB2SGSl02xcoCYDJb8o+todcNcpb
DjuFwa266U8zkCg23EjZgjVpirrQ6ebe67Fun02ek31xyJGNB0/FcFBfUjpTBy/r
ngelsBof50vkR2bkIr4dGuH0i6DiIxbE++3IjPtcU/s3PECwmqgKE4ZJ5SYdS6DS
9cNGHhjD1OwXDy8WR23lNembqi4bQRuZfMNhDHl3aqGoLAzjFouPmxHaClV3cnMZ
u08Yk5onkLiU3qHqdBsg5HAEyDm/BaCkVjti56VsuA8f3ST2kV+B+qzkUEDyZylm
eCffo0bbzhmf6pCFkjb8/M78oLNqfSPtGSuVO4l6K2NklnYA6H/emdiYznP8fkL9
hz4+GChMH9JQP1/TmxuV35ImtbykA7HPcu9Q+Oy19haCiJzLsCAg1Zp4mQgU9xaS
Zow2mA7ZqF48RWPl4liNfNmgg3dSHKjAaW7jxWgaFhd+sq6vbdtuxDHCOo86dvdA
wbFDlYr0HxHPX71V5fNhVHYUnnKY0wQWXmUu7FM9WLSkVU0nI53l6MnY2Ysdj/RF
YuNs05VPmUEpoh2Gg+9hpBIngLCrxmFZPTbvl04r9KPBrsZCTKrasVm5DpDBS0jB
LKBzWzCS3NOL629q9wPPNnUZwOhGVaC8SNtnTP3ziC95LWrifsgo/c0JaQZP51OG
LZpy9vNCe5zUv5qXZcECwY8YNrSTx41E8j77sPb8eZdSYP5p1iZFZIpSsLJUVARd
kDnWCSHrhBqyPe5s+2RJNllImTu70dHqaJ7TGtXHaCT+VnJtM8H1Afq5KBBVlIdV
qfGrIPpnRJFX+vx/fXRsaTYQxEZ94wjuKpD7BQ8AcWJz9Sr1KzIq7Jin7fXn41W4
tyJEVHFrGAEe2ORLuptRHKBSmpCCUH9iutJdLg7j9O5JcXFzePTXxJlIMmcoAxI/
496LUy+4H/92QVLKxk/CzW4A5KBhg6t/rGpKjZhdTyrvDxMvJG8NxCNHZiLfYY/m
etxGaHEg07APxipAWMHeau8XXFqrPX94/NwryHTFo7XfvfhJj2v1R9QLD9MVlgl0
HLR8Wu12aMKfeKTrDG1vu/S0MneQFbB63AT+6rtsIB9Gdn5azLykPkG66p71DaAz
5GFvO6wohFMI+rnYp82eSv5g1AVosbL4W5By6UgYnKCHQeU/brB/7JUUVFfoRul5
+1GYKKn5ICa2o6mBIQULhnGz+6VAZ/ETwGf6ETe/ZbUt3Rw5yXRYZS7n7GSTbWyk
U83A0j+44BB0TfDBW5kkeOVynzJjNJ1vJph9aJppiyMcIVGxEqG+wy1BwvwewZOP
y/ru2mvlC9702IBXezxv6M+WbrrlP5KC2lqpAj6GFKGqS2vmWGnBJrg5qJOoebyV
YxMLEqM/addyMwVXmerjKPLDFi1O8RK6Cw5sgUZCD5FCAvVwOdv9gUCyABS0eSIT
hs/XQqZyX8yiaBvY9Rc6PYDtxKT4QiJbu2Cbl5siMfT0X/NxD8g6YRZfR5LIvQQi
FC9AYu6bMWDEIVKkq444pnYQWLUiC6/9ujgXZs3ZYl/JC8ygFV1aHODEaqtW8tmX
7gNEZj6Fgq2HJNKuhueaJqqRXUuIpJBExeXW1VM0Y8vdFf0Zh2YRsyq995bX4sDX
/IpdoGaqQwXCue9qKSzwy9/BIOfXO3JTzXZSIN7gsZ2h7uOENoJ2z0o/Cqqz1V12
AFgP3+Yb3Df7gF3hRsj3ILXJrX8mx/ZfaQl92ZOiekznabbWlucVT+cq4PpUA8Ku
nsfpX746PlnSTpjVKEgUYQUK/pIAcv8TKZEEAjGiR2wypAB0pTbQ45Rm4B5V78+C
Oi5bJ6OdnPoM0HrBVu+fYpZnvaVPT1jwGJAc3Ljg8+8mWIs9E6X0OIM6U6eez3co
D3ZvuwH+rvQqscXJcghpZ0zPCv0REvYTIwqazUk8c1SHQjiQnPKIPLMAZk84Hkg+
LcNYWKcfbY+K/QHci4axykBNYgh/poLTlji8QeYUwFjfjVn27V/nh68E2/0nKxkg
ayM3rO24QTk+JsvEoef284J5HtDYFojp80H2iqxk0InTlxbPBq9UrjRieU3DZkVB
xyUKmg7cQUMvYA2WfGeRdVcWZ27w4lu+wStDTl0eiwCbyNFUZPhhTVQcbWPqRI4s
Cy/KnFXrKLE0t3mnjFHvJwPJGufrlaD1IKYYuk1pmxnF6STpXZMweP9bhiGdpWrW
XiTfDPrdCFR2k72FIMe/rRxk6N8TpiktiP5RVP0S9X79qk2Eezgr9X8r6lBPuBVG
PSAbaZOYu+vZgDAjD9m0hHuSv+eYRdUDu+ofBFS0PfOyfnx1bDBqpvNHUfePZCWz
h5Bb7R82t1FTkOwR6g6enzHIkgvqebTDfEnbIDDNjrnHEGWyFlTf8U6SK/op7+95
sqPm8UpZ002u2orAaoTUp9lIXl7u0xfx+ohBVR6Cvr/rfW72imFCGnIajVxsm6rK
uAZ77se9bJQ1Ni+kaZSuXTouifKd/w1M/rh0pEU+2fJfxE/JfPjm6u1+hu1RpmFv
3YiHE4lyA7DtvNarRmYdSv1XGHbw3YbpFX08g8SERzBuejdQBmQrX0tM2Bh99NRW
MkoMBG48m3EDQdn769HS8UgKSGH2QFHcopKwjRQYvY8UFAj9n2VF04GLFnmsZlJt
fMRFu4R57GMzTwI8SdLvypnQwVhmt4qWEuqtev4VOcyG0pdvzMI8pxagPFWYHS6m
NCIa/oivbL+tJmhXuRw0J4LrmJbv5gP/jFEtZQRstJ6QxdijOAdcvV7xBwgT7bcD
TRt6yagTpLdraCajNk1UWjVL/Hf6Dh7PEGvi7uNoNHG1TZjcpYlZ4C7GCnlbDUkt
Yifw7gqUbNG/FL1fwzz0cv4syoFm9K8PREHpNNTqR0ETFdSPHr3r/UlCHpCjksV7
q+ih1Pyu8bHwmrDEk447OzdS9H3ZtfGE/OX+kPS8bRwLOBzZW9O3HHvgsSi4x3ga
GgODZVA09v6UMF8QKQ9UmHOL8IWwaXjBKI2oH57fJeahNFFXrhxaVoVcLhRTM6+x
fJZaZZ7hD7vSA5s87tXbSTjf9xOSl1FJf4D6ZvGKtU8hklXNdbdZpdA4X6BhhvO6
Huql43RFeQK9BXgpp9hBDYx2mWPgwke3iRlgwxOmGH7XwaEPKUQl/sTCm/dPfaKA
0ddbM6OIoY75M7cHnRxD9MUkUZNB2WICvFuH2ImxWiVuKjOCv5/SnsxdqrY9bQa0
bUb99MDsMAuNAc3JkoLhW9cQr6Q+PxmDJ16ZHuDJ76Oqwd+NkEbleT9rOmgs3UJ5
yTGlahP9+l5Gslj41ijhGPC5+u35hbvqbq4oIbEvXFugmgdwhw7GVz1sSgxnRgeB
yaKaPKy6+Uf3TCEfn0ZXylCPQ1B6mOQPKCu4BvllTVrOYoAdZhi6ywBJWmuqrQyY
tPIPPa0kbXT27T6v8YZZd9wGIPdDA2X+TYJLLL3yqf3hkRiihqOkGhaN93XAQP4W
1IrmnZgcQht7+wWTnwHSvop8hI8XHCdpWaVZFQaBJX+Uc+8zyU6GkQKAHTU4L2dM
6HghB3J39HORviAQPQOxIeiUSLnrek8HIlNV7cExR0wEw25uV4t2D7L8eI39V3q4
X5a6bZzVW8WKKURYAF34poly08DE/V/J5MFXJVQ0z0QZ/ylYJoMiSXwK8rf+MMh0
uTUMhdGdDjBi8QPFKu4287CjgnN//qpjS8rQ/4x6JPiUA7CjGZaywkbEgDFUV1iB
qvEq+gNMIEjv5b293TnadYcPldLN7lHOuGNDiefnPI6XZGxQany2z1VM3mk7H2GR
Y6cIOOlFUcC2G1uhWdwulUKZ/NRfJid4mL4O70Od9npITyALgcnQV6MdmAz+jh6D
bCHGyRuAlj3L4k0HjHPS6Ci3GUVhq8NnxtgxT87jWTO/mzsWkXimI6n/E7IR32xC
4xvvPwWrLHTajl6CNXoDJXUXSzMNNTh04VzJlvsA2DfPCuTYv4GsjuCLLdHauLs+
T6chGiXvbcWk1LRQoH6mbiU0BTX9r7gciuuBqp156Ru4HDQrV6Kbw/J4Y9TjB2Md
+pcu/cAK1aALpEnRwBDrTgHRrMcBghw2+igurXk0AajeV6tL+jkkeh+w9dhDsSCa
1EW0XveHEdpYnFu2RW/qUKItvw6gB/cyA/wNC9Vja8wfCDQFvvuOdWmkiXmtqbzh
BtzlwMvY7uprJPvNh5u1LCz8ayYfofqYsrVKr1u+6vh2+ZcD28RG4WR+op+rDXn0
gnW6Wq6I53nd1WnVqT7cXO9PLNElME8Ivciy8TKoSunxQy4Zc8irpB2q1dzgyupx
RsrHKSfqr1DGnleRCjsr5d06EokpE86C7mXoF2MZQiE3INfcyLI3JfBvrNNMRgml
7BNLMfIV3tcAfRHx6QzH2FNlb74UUP5f4FUYl8u+tTP1tFilGdRtPW+5XMStOA3Y
7AVELDrdKZjQdj4ZVSLjllx7Vy5o2BeeWsYEEMf5DkQC8o+Jythl+Fo+3hxGf2Qo
Yi7tetiLixcd5mttC4neCJ4dBCmpG6rnu/eh1hXhromKlqYBBpof7jle/CmJg+9x
616Ux1y1KNKUYsrdr1RVvGVek/Z8PQG5nuENPMFVrPG1VTDcZffexycH4zdNHMbp
muKEtjjBAALRPOhXDRIsScH2yZZP6VsGxM17oYHujKKrYoqYygTevVa7HKPnfm5z
92fRL3qGZLfhzicrVUxwkzgTCVKZrwvSKyzA5yfR5LPeDmpjU4TudOkee96i/lGx
QKZO2vULx+kgZELhXrSjEiCiBfF3M4nWNGX+09HOQeuEPsYF9eX8eC6c9BTH4C5Z
Hqcfc5lHLsnLEP1xcZGOIWk24ChvZvruZt9h2zx+K1pYZLBoN4atjeV+CoGiQX+C
B/5EeCTdVc3kCYwxdtyeGU3xHXs9aou+ZL1MH8mGUfprliRObTkG877wBS1Xoaz9
iR7wmIMxDbliY+kgMjI5BRufUCpi6ZywTjpB0iwWR+wlEkMW56i/MRltp0UvmYSR
skwZIQF+7Y6AKl8N/nUTT88ZLlAn3hmELn10lVAP9J2K97DINZhbp9xJqeJRTbho
keMhyozRjVr4JX9HpigYW3rryQ3CyWL6byLmjubBSg3u7oL8EawtvG4Vk+bFJsS1
+V+vKSWFRm6VlisiBTw1OdCZCliqrbUylEeyHFiQd1zFiPHlWy+Fzn9Dj8BXOi/2
Koi1f5zRdeobr209t5Oqdr3mAtx4hgqGIVRTKsDk/mFJ40MzD0JEPNnmPuSdZse6
f3zpa4iAfl4wCm3stijdYYugymr+v5kCWZWYjIWi4G7/mBYbH0zyD9YFtQbIPDZG
cRnXtFYvayDP8JnPx13jUaugj5YWIBuhRHj0nDXdF9O7PYY/sQkoX5P3v1P6Ey4B
RZsydNfiZF8ZyiwEWTefSAcg7pesS2wrFe4AGcJtEa1NmAACIf2UjVCzYRV2uFPw
geMbDEFg+YhM1RD+NfUGg24GZoYcsDQM9KJZFPR2uzDeaYehhHxwaxM8Y82PDs64
ui0Ziv/UfH3rLmYTXdUDn/i+yXOoFN65adnAQyFVhdx6gPebfgFl5YD00+I7ChUz
0UtJ8aVGeeWdii8dQMtz6JiTutExTVaHy9NEp1JhescXc1vRNVjaWT24a8HUyV2d
JvGbyDy41AqeIFJxk3RSr9XyTv2EY3MXBIQUlOZGLFgGNkyq/Tja5kZ1tCa6U+DQ
mjm/i8mZ5i9J1m1u4tbYcQTKK4iVwiY0ySgDZiCGYqCpYwcl54cj6QiYcvu2PbW1
Of3cMMoc8nRQTGTuIhCfpscFlAHl+FGwng5s4oRQjL1Cd1Uu/okAvtRSY4POGWjm
aYQ/f8UNcCixsx5LRlt1UyYFj14LIHr75XPrhPtuMw6ktWIcBMNDAHcaCle+m0gB
TCHi5MvH5SP/4Z0l3hT2Y2HdvWjuiiUmyDmmQtjiwZWobrkfTqlZndN2HzZCHzqK
bXnI/Aej2TIlOlaambC8oxxxh3JAIItWLrB3SJ3smxHV01u0SPvWYrm1tqkTRlNy
HHTYZ/GNDsSiOtTSQW7WDslsxfdiL5HlDCT3IM7vy2xnkgubQlM3XoTTc1SjmH8K
fxk0dRTHR4degdppOAECzMU3RHcDU5N0myXUasBAAiO0WXXEXSL90s46dSjqVCca
8GLjF3ExD8PbYkS16RhoiPwVpIuf5fxjRqrEhBeZ0/WiNGRYcgf8AIkwNizjODjf
MiLTur1kvgQMn1o687t5M75JaavOQqd51wDIVLAoWi1jod4/DAL9kQJoO1ZvjexW
GWndCJrNc+PjlM6YAMS74oabCF+g51LC1uLti1EGQghHy/w8BS+jdZn0FJgBjuQB
LWoER8bbg6+g1ybxFDWYc7zsaL43TK0K+uUGhRWEHDZf/J86YinQ0n7H4wVzhL+N
G/ntxv1m5iVbIuKdfNHKIb/OAmO/0vVOYZZfu8N7rMdfPlHjRrtHnVLTZC3Zkb9C
jl/ae2VafOCvqzsOkCWs35PmHTQZmCNyomyLL4gK5Lo+7YT47q+OMrAY9Bgqena2
dhnPs8Fa7EwkBonJu7aXCr78G0rYYDFTkIQgRGl/lDt0ho0s4hr3EW9MkOqCg+wU
QOuKZe9lV5+nPRetCGgcfRZ7xH+V4zQaju4odav4FBLOW8vF8IWEp0Bus9NkxBBu
ksKP4FRJP7b6a3L79RT6vxsEjFDxcywJ3Orkb1oUjzeulAeLcgrDF02vPCjnmJs6
fGGCW6LjpKtXQRzRJLR323CBPPFGZ2bwOfcVnwypi12gx6vmjwh+tFOb02uO+KeR
DCCdaN2+Z78N379kx5pPDkJYPAskicikPqtijTfxVoJfKkV2Pa4DvuVidH4aksL5
1WknFEm0S7M0fHplRiS9aPEL2lEvkFh6p4Qdy5po+A6Y2NWauRc9nz5zACXtNpLu
pXX7uiEuUXs8ZRnJBwVECRYtGr8RUYLuVp+UUgHUcmMlfYPvFpqDKBcfeU53LD3h
S14HqIm/CTfFzbEwLuUWplkOFtQ+Mw8NIAjmxpdmjEUFAu5AJqAyFRd+EPs9wT1H
gBjBWCoi763JHDC0f4IDi5DkybCfcPfhSDIlivtyspHWduXbQ9gpkkA7T/58NF17
eEd/fDXO+zE5H42A+D5JuB1KUnKVIiTfmhyPKsyNgmNWXN85ilhSP26XVtjJhuTC
UV+XXKPw0+mwUNmegJnyUg+c8SA9MYdl9dkMwmrtrTkbCu+xiK9bTprbS+FSVfjm
M+dGOL4kKwT0Ct1Q+IwIKraanXikq6/E9QMdX/VYs3BkYs6PKB8P/wDhowUAe5Ev
EsFmRcIYIaC1OIRojAbU10ObHwpq8a10O6qUILi03GuyiKU4sVpUPtwuODwU5UZX
etV4vYXX49Ow+fmzn/jSYgNS48YaUk3y7Fgb8CEVmOUgVsvjEIJ9yotqaClj3rYg
iN1tUyF2SUziUfMQR3l1qP9pnqX/nQ5bxWUq9f+UR/aPPLQ6Aidk2mVZqRiQ6rAq
wly0XXU+qd3xTsUzNkSsRmB39lWnKPVABDxyqkTXshoD/CBah3lCVnWZ7qaipJCr
shLdd8/esd/F54VJyTMpNstpqeR919GiLyV0II8j4QxrOgvcOCpv/H3aVeLAO6yd
IWrxIaNBcdVcYVBeB8T3Y+5jZR16sdjI7pxIHUNwyL2Yxw49+yagDQB8x5uWbNdE
nWaIPyUYSKr4tqzZbwGpH0kzX2RSXkx4QqtqynSF1bQOoG8nSiLdoXzp8YwQ90Hc
1mWKbsRUpIvihtUY8tPLvajYFOjRV/Lh+SWN6cdYAGGvKJ02zbf/BdTqTD9WiKQt
+NPdsD/L8QPZDaKi4j7PjKM6f/7U/FMSnPH4WLs1TY7P06S27udCBDIm1EKdl2l6
VdNDJwyOtylDPsxEAChgxGQvvULLdI5tS0w6cs+iToCfFEfDQwcWTYVN4LZOGKr/
7Tpltc8zsTqBGPou/vmQENPP7pDSM0ftISK01FayK6Va0A5ApPEPGUomryikP61s
VDS9SYImIsP/MagKm6WOvBa0NEyEYPA/LKk07JrxQ9yGG9vNGZnblIEm1tLL/ibf
3HoIwu6VPHe2s9z0R8FOV1vAJtXdGkfA/0h3uIxrIzFqp8WS3TrHtS5dDDLXWS4j
ECICsZkjtAz0JGnpBCOj382xUZTaAldyeKNT+9gRXat66ZvIxZdehfoKYwbMydJ5
2Mbai8PIcBbAoHtvP/kDnVLJg9DO3YJGhH8zDoQ5/ZxudVa26pJhlUpNUtQyVBbT
Xf7Dhlgwmc5riAxeQ+dLuD+sSvpY+A9VwcpGGHNmapD/X0PxluD0DPMO1MwR+1Sq
ZM79765mkW1EX5gXv45H9j2dM1YWCu7On2cojf9ToxCX3Wny9y0PFL95kG9eYVCg
gF18Cwxc/kVfbBfGhOHjNCNyvnOX8+ZcDRdSrDXXSevqJG2EQhZRtGEh/gfWr98i
EYYaaXrP9z9Q4gH47SJrW3wl+GN/1IXkwsTVGdpK1RID5pYYHrM9M/n4+5ATi8GN
abzK8JsJ3yYc6aRUhoUcYRtkv6FWcnz5L9SY8C4IfINuMfaL75AH/gtSWiX0Bq6f
z9TjTxj/evzZSg9zhNFOGmrF5q1mX6YNHwfD7daT1E0eVB7bCc2GH6McZ7Y1GKIb
5bMqDXiJV7HOyk3pLiK7ngyLOo+Wib+3CsEkUGnqas8Ax+VvFcfJ5LIZLcMm35Ah
8WVaaR5iJZtwBPkVH/yYVIP+ovYU+U8Inq8gkx3SX9Kk94fPz6KJISKk32RyrhY1
t5hrkVEKFXAq4hy4pSh6MFVK9UdHTDLo8LQCCxTe3FDbC2owbKugoIZ3GrWxiADN
PniY9oYQhcIPLWh6SeUx1nivx7OJdk6NM192YdBurU+LytkiBi3aymrFedE4Hzl7
YL0RNcO3DZVLFP/wO6bPxtn1ak1deSSM241PelxVSf3smSkfv5/iRs4salTzq0yV
sTjqxB4LRQxWqYuzrhE0EAE8zbnjJxYsv+VSnqAkJrpuCn/XXxxyeXklhnYXwvje
IYClSEr97D028hfvNnEiDHU7lcKQWyfno4RUYBy/y3Fecotx1JwzZKZYip0jaGGQ
7NVGZNBkaMtSQNVN5xN/7z+EjNyFD1d0OZh5LCwfs4RSXrJUNVOA/jjP2rTU0DJO
zN46dCabpBenCh7lKhZxhqTYNWdbZ6q/ow4JQF9AI4kwb19bwKLnHlmXwp2bzV6z
6Xu8Nvdg97bV3Vcelq92t6HqQovdJmm0H3toCML0rkPHtti8ckS/34f81UiELP6I
sC587/Ot5yfnXfrG3NFF+O9R9iOQ/+1uEAQ7QasBSmCF0Ykp3G9bYwxuojf9Jgnp
CiIKv3xS6yagS38a0ROfruaYXqu/T+wV3ZHSlaUHZnOqGvQe4djxHyYdGShsqI5J
MGIJOmEfIGeJxDZOYVcMtD1xU8dPoJcIc7T/PgrW4m8bIHUKTB4ZrWn6wyv1dEib
mN2tEi1gqHE1x363sJY7DjGvxF7MN+S/Zf0y9AfgfpYJvp/AAEB0FckL2BCD0A6L
asPvtoiqAETJQu/qXZCv5AqiOfvrE1VasHQinm79ZFfL9DrBiLN8yYDpEA42/Djy
VMfJvN8W7yR54tVjgout1vkPfUPGqcCWnWUp6BWxCIFe12pOFm9g9Bkod6e8a6MU
SAsaNofFzFOht0N60dFtyFeX9urUxP74zkQEQ7MywwL95p/ic8oL3twrfnS3Vpd6
SN8SBaJ4x00b0aMASXg02ZQIwDFybR847nhvX9F6igk565DIjZpnhP3OWa9THupw
Ro7CdzO9ywbDJJiRLjH3UDkm0mVP7TUEpEaTWXlZ/wt3rEmc9p6pSVDPsVR/foaR
3a9rgsTAcPlZ+O//DK5ScyGCTPkTtRJDjywqcBDOwylWTPfXC8fFffroQ5VsWlh3
i4kWmSGI8kfuH7CntAWaFweRK+o5w7afvEYfrpd1prd21UiVFBMR8zhhp82mUL1M
ZYnQwFDmyxaJnLt1KDic5rVA5VXKQgu8GXyzA8VP//gk7Jtxfi2N36UVsO/b9xpq
0pv3fe7JsWPNPqQWtTeQv7OuTEMOeC7Wd6Dj5uKfWncTdT9npfowuOctg0p2g8y9
Dmqg7AWpEca9l1ye8AnY3dHaN5oLeFb2pWzaXkSlXAVl1/dp2ZTS2AkwY89c32um
QY1UfaWqqNC+GwQUVgFUXl7t3MGW4D/dNii7W/hPZhWtfTa+5KkKJJLUlYSq/4jc
h8crFRhkW7SK6ZiOVEnNpTVR/WM8RlPCZuMuKGgxwOzmGioaSEMcYNFuIIfa9fAt
9p1d/ifAXsPFffhw7+ovQ2yBKtgWsMGAn8I9VfapN8nYWw7dh6nNFg2ElacYsnZS
jo29BDI19rMFLCnHVOioehG85XT0dPfw0ei0rjX2OeD9xNpjeZppl8rIa/GbUGA5
x9n3rpA7bGHDAfCw+RJPmbJlt0TNACo7N+cYhTUH4hzstdYyLfGXOGYXfq6Oy6nK
rC5aMs09fzrpiIJwQRnDIM5HEeu6N86+4CM03oU5a7BcoWpTCrVU4QiDYQIEYwpK
hKbu9D1RLP8PVxjVvhhBpbYfDoCvSztTjOBE6mQgTt+g+k2ndpkWYhpRUaJK/ogJ
e96cxPxWcXOdY4usDRY+qyET40nXJiSInCjhKWL7AXz786/5NxOVLDTCV+HXp/p6
b4yzIRZEvKWCEXZDUt/IqBvFmD54K9gaZ0VPUURaQsor8KJXU7203TbDb9Wg455Q
tGC4g08RiivmxHnvIx/Zyyw0EfCOhfPYLjmB9G8rBhgW4WhNRe4E4bmAJ/qg4R4Q
r8PHcvHPlWnivN+X4mqTdkntjFXTV+6LyHA4wgRZMdsdCQ3XCF4i54A+rvW2acub
8qVbo0mIWpFJaLbmrlY58P1kcnzxji+zQWKTsgMhLD3dRRSUC8GJKv6Jrq2sR9hV
8FbJjkcglbA4zV2GEnZiHjQWCufyWfRNQTO7TEJZTE6wRKjdazr4mbipRtPBUsGz
usY6lLlHAxmZdlIHc5YmGVoxOdX2kLYrsZAy8FV60q+6wkcIvCUez9ctbez+Sqdr
Bw/e9ZYf+RUoNC8/Bkg6XfTxzOV97pmbKpfiKSIVi0in6slgKg7cNGRDASwEWb/A
hS3FPmrmBUl422tWG20hl3jOPZGnCKPohu+BtLOR6JsokmhcSKZOrpBo948hWYnP
xTTGhBNceX/iGsgvyyEhqNe5H1d0dUUAfh8LpmheATOQ+sxFsMawNWrT4fBZodmP
jK+E7QKjYTx3uHbsT9W9aW6tYMdoCU97PlKW5YMd1u6+IrxCsi4iwfLvt+ibo1ge
IewQJv3ijPC3dXGICzmKAkRHG7hE+ltLM15bPQJjBHZb9f9reuMGmx9egejG36yO
w179m126erIMK88iVV9TGe1Bm5YMk13Hb73YZc49PRfYtZYizjyXsIIAoh/b1yzy
UIuiaPg7echG22E83cbo7/jGILN9deYBtv80Xh3aRotZekbGcHTKcW/JlWBTOSnY
McMNC2ynwkSi+pNSmfKfO3oYAAj3EieKjACTnkGoTl4YnnRfKtNOP1IBcFoNGLAs
G2hQ6ebUn9F3v6FJ8SR+s+E/bTAk5XMIun3E6inEa/KEV88pqJMmvLkw5iYeFdmj
pyjxAp+wPu15tS5LWoOsluG9Rg14AUZ85wiexYJmITKQTz4/URC5W+Lhb1b+E2PK
Zi/dUjzxDxV3jtoR7oMtNZDHab/qnQEamu0nZmKEEGFuywMi7I+pw3A8lC1FjoGZ
4re88u1cABQDTMh2FsrT6wTus0E6d2Mr1IAGGMRaQ/ZVdRHE5a17HasmLA12Q7e9
vWWzXmyv/m5s2g2+GNT6nsmS4LOfs8VuMO0fJJyB/hmxCjwXzO5rPFmWAhz5JIbX
rluZoVVtXgbQOehtJRv+B+pKK48vPMyCvM610KaWnXqqKDq/CaXL0j6UwuS++ata
TuD6czBpAPMWDE0VyElRnVzatl6OI1IS5puur2fzGtIYtaWJ62hE/GUj/QQchl76
GuQZMKkRoirB0q5CqxU9rLx1OHJZkMLDhOYU21QIqzYVeu2LaWiYYofGJMeh7KcE
UrleeYilSWML1Fak84ep9TgQEmRNyQPtKLIlupg1Ge0F13i1bNo7lmsdF4zQeg96
bqctlvqXIwwCyQ06lIoyMWf3xLvDgEWEm5z6dzB7II75JofGmx5CC2sKjmrE2s0F
Ck4j2bMAv15vda8mLXpzhcp/aprrumJ8L9NpSxR3U9LGVtpktKGzamPz8tkUB5M9
2FC1cHYPzFcceNE1kpY8heyUCYBdzmJNZqBSfLXKPI+44d3cMt92rBIfqQHmHLac
dkJEcZlDg2XTDjx4IcYD/7jqu89ahkisSHCzoqiStUpsGcfiOi8coeA1DKLCaeyh
6bSO9hpUM0SGrpFnpuwwS0CsYdr8gvrKYF9QL2RgZIh9XaiYvmZCiGkWp2S6bNXp
2Jkc3dyPdeHtNhp4TRbj/qKeARll2NJwimi2CjpjA3Y2ySv1TSn0Dh20DC0a0zkL
eX/L1EubmAmnLSXI81x6h6QKkRt4f/3u5I317TEh4syKihIgpAlmb5Jpraq5rUzZ
kihVcGg+MP7GwZrnfuaSXZCgb8ve80HjB+IkS/PHpMIEtdray2A9/AZWMhet0LDQ
ect+6JOc/9ZJRvZC2Q8dl7XF6IjFSNSssiKzQ+j98WyXHW6xh7Rui9lYwiWgHqYZ
hp/Tv0qsXpwktxDyyPorTNZFbVvR3QiBkgopnLCIp1FG+TJiXivwYaJX5qSjcMQY
nkgvBm8GEAXXwy64xOQWA8XFlG7NZhLs0JZUknJkHXDFIkNMLI7sYi1pVunNe+Yp
jh0Nh4aAdC1e3JqOWxItLirrUxrUSByXQC4nJk6JdKAnUzQObce0XvUmjoAd/8JN
J/s8ofA4ACy6D3ZzhjwL2vy0wkUUA9nInwOOfKXRwydj5zPJCxRnvzJNHIO5Zloi
aFCroaM1Snf54gCNWkpIMvjL3GYFjzxWiOW61Ui14VrG8FCpjJRyEl2RZDID9vIh
a6ioCf8POJXKMPYYLFtsNcLuyoD1YlQ8d9piVSxJSIRVnCXSccdpNICm9V51p/S5
x9wWwXVeLP+lxVGY5HKtrhNpiXvCi8UqjhXPHkgdMJte0X+BJYfF/7d560dRBLc2
cKNhFHfX0tF0RI+7E7yPjfD/es1KUS0pKiDPHjpF4S6JUTfOzjnRHP4XzfEsA23r
q6fDutBp7NLZa/QzdkEwvfaOhwxBWQNtz3XaT8hPu2JY9ISAHkjjuyX9pPLYMlql
pEyeZk4wtsAlbcOpWRTL8a+mS6cuPmxpKNvO4vWG6QWK2+hy/gaEezvVs9R5OCRv
0Ic8Di3H+z/aAoUpYzDa4IdfhrtV/C+hKXxgLTVDe9VoUtqQyXj3RfL5g89GqdUN
ENrkMyXHbDT266McXgbFd6HnlUx2JjyiFndUqzIRikn0sm6U2c4OWb6RkURz3sdL
cs9hdNJU58q6rLegLSDsjSq7p7+rDPO3DK8UipQzM5s2RL5TBYahrlhUwhjSFTFd
dT0qDQGdTUc3dShPNzVK5Wpe5Jv4wwQ/GQVcZ0K0wkrn94RBTOirJQtHyvQyMez5
fRbxyqayvKIZFL1ZBfP9V8G1XkbkL7bOJRQOYJcJBqk0sa84hESa63DX+njjv/6I
1jDE4vJ9YCoN3mSNvReYTDWuCisqX/aUD6qltdv9cIFnBJ7sSQOg9YInVARKctAt
QJ6TC/6aFZ7ihXGHgMmPSKc4D0Q4ELi+36dPH89wxFUHGTqVGqCQM+R2QeDffUiq
RmH3dyIZi9BuXE47FaOjbN2+TpdP4geSgm3AgfjbOgWqLNGs3y+dSgMXDgLM5u9+
9eXv+IgKZL3gzcJm5Uf4i/o2R2dVS1JF0eB/m4qR9d+3e/T8Vq6dcNL3x9J7RsCK
hKW1a1y0QZXXyQ6jrmY+33sXN8a19An4NkGEXDhotTXjDUEUBSPdeicrZoSorYUN
STm99DfM84fZz7Rq7gz6pEYgWObt2tDSd7TtGa3Pgkhn4DLQBYpFX4RFvw9mPYid
jgyMEaaq9lA69cW+qL32L14eoLjxDeaJEmzYSModuNx+bUHDYbZT6v6pmQt3ij3Y
WskrC8vis5vbt7AAoTbaMavdPIPDz7QSZ33jIfsSizN+eaAYoSww7h+tUz0SVMCH
kp1fwjHF9YJc140wz6e5PPLXxYigOfOHXNKXD7x8v096pTdhADnXvczhG7uoRTyO
MVyJOagWItvkBmhUMjhhezOtwPmNqT1oXjGIqXJvKXGFzgQ1Vy/CKtVlYQpJb+e9
y6P02WlN7+VR7cHtwM0mAfpliwOI7lSlv69UPRCtfHWDwzDQbFLJaEcydxdz5m/c
NOJPP+LpnNaWbmopjSA9EU5hUd78SJJfopbivdgkucdSqN3yDvD+MMFbXHJijYit
laLKcbOy6xyk3TyUo1Y3EFetv/L+a//Z4Q9J8UFmE2t/3M0sPB7hZXvF7FuRme6Y
ETExgv5wnaRELNOqiHPCxUiqZN2IoNt5rkiGvKZ6DGWJly3ei4SA7/U5MaPZSvzT
qCL5KLM8K+32diy1x1pONO+51VvHGwmoxMaxKK014qdvdUsalDoZWYQoaOJN4Wf7
cmIIcWu1NVTtY0f4Bx6RE9TG9sRWLQ3UDIpRDWlIcsbBWt6uVhj04v+NumrPxnYM
S2ygQ322U7wVn1XwNWNo8Yn+FsK4RhZ040CZuEqbGUS0Hr/Qof7lR1moBg5FrnJf
eWWxZwa0Fx8oqaPD5Yw2kLKOLR9MeLKaJj9RvGq6lh11durd3TArxlbZIEcESXDA
IiT+0Pnf9jxMO/0Md6PHQFS8qoyqQLA/4/aMIEImrSpu9MWiqcwFjtFOxXqYAuT9
ZhgGw95P82zCtvg+RCvO2R+5OeG7yNSUbVPWgeJxra2aktikLRm+ZSVhMprWbNVF
q2kcx4xGiYfXPq9pQdYuFidjoL/jxfrY3c2tfdeqB7Y8WfHSnw1imqf9PmWl5nrZ
u4BU11DOfQS+M0LDCxjGkHtaApx8DqZcjNEnCyZSlPEi/nds/QAEhHdBklGPisQn
9CF4pqpSW6H1+SJ+fQ5Usc1havNgfgL+d51bsjVES2N5cjTnV8UWyqkLAjND0ocy
J+kLa0HHXefTtcohSTTSj7LXWOQ779uSeNU1il2fXwobUjEW3wh8uXEf7oxUOM5W
mUkPkQzeDzH5Qcd/SLF1U/mKOq8zYvstNqDoPl5MFtNx9MY7m7r2EvdnWZzGKGh9
dQ9UTl/Bh880mQjvzeUKetgB0Cg80nHm5+Drjaf8uflfzSLHYVNhb0LNCWguf1hq
2EM4ymckMwHxVIZzL1fpSY8SBa336V8QwjvmZ1XJLAf3EiW2V53jsWZzzaIy6S9+
/doMEB7ES+YwIJ99fvZsibP5c8gelDFFQF88phvImVrzesgvs33ASJVC9m2QOQAT
09HhM8rJbiyMN+Mbt6TFdrLv2iV+wAzDrt3L+YwHnMZlF9ORI0uGlfLDDmlSFF3n
po8VNgk+kUfzGLZr/s0p2Cj/SKHW/GpHdTRm3XN8eKeLLoMl08bdLE6rFE+uWTjX
Rcv5xGKWz/20ImXuXJmlryDb3iTXdE2kp5Et4t3nFWOLozc4XJFRpt2qByELM+Y2
m7bG0WEEyD4x2zl+0l3IqU94yn/h2/cKTYRaHoTC28FI5UlayAsX8FoSibJ5Rk3w
/mCj984tql3gMnGz9Ea6ZdZhXuIehPiXzf3AgcDGn/TnJqHQ+OLOk/GRaxH51BmF
PW4GrnW86ZwPjdMeHK8GBpTU/BAMxflHtEH84VPzVQPfX3jUD8ungTohq7ZS6FKH
WJe7IENzt9I45H8zLY8pMHGQspshXBYynXzEBPa7pbTK3ScLibdYVg2To6jGclvl
SejxADDbFydfLTYeBpHTaqq9Qlw7Ye7i7t8LdNAUC2bcxAXY/jE3RxIfJCrBS6a0
n1J/9Exizku/T740GI6MXIkNswIbfZxZGfSJuKCDqwH4jTTwBCf6rWlaUh3IvmlU
oUU6FsYY6DhLnsV0IAl6nbdSMXS7eJsO+BulybJqnB/623V0dwDyaSbnPa+0afCT
exMSSZEZEIS6/JmS8VY6nt92EM7GhgKGgEEjdhXtlc/si7MrETv+/G9CdTo5rmyG
/NeHZL1c9g9giGUBl/g0jsisLBSsuwQ0We9VolAfQ4uvCxWNkWtE7ddI8LPuCVih
/DfC0gF/L/b/ol0vJVmZk04kMwGNJWvc6xGTYzuPKW39PnPxvMSZSFX+9WRbChXm
rYd4S9QzGuvRErMZy7ti2VX1MKCtD1vZB/N8pdwcVne72Wkx0Pyg1c28mxZh8gt0
Ia2vyy/xYiariznDUV7/pBt4w5bTPSetCZmkyVgfoUsORTgUpZtB900RPqQ6e+J2
eMycu6ucclO50YLnG5rv7uOgo/MSRtoSpwtgvCHZg2PSHwv0sc+l23LfDvB2v5yj
p+2azTMRh6oz0DIWxS7Q7q6rPVyu6yokzh94whZAUrTESq5vWWiLJGWm/sXsScN1
dVC+Ff+Vbikw1MQFs7tb6wHpCwqsF2GBUP47RYhco87sraqz3bNnLe2KqC3JMZB1
QA0OK/HPfiVBVfFu+UvwH7f7ftWuqretbQB7ahs5jT4OHYP72JbGQPAa/trOJo3s
La3m3QDztMOlg6eln89jAnkemG8PC8IFFO71xjZSkjmQdr+35j+p6SK0A5hWCcVf
NKrqL2GXrS2RHKafhO1wE9vYMcocvuUAMwwjqSKfDglipvqDA8UeLH1YeV8EPN+g
aS2GMY80VWWIsUrWdM89+poM1+ghKA6WImb8QuAx7ivYZmoow/wjw3IxgXLE6G9e
3fdReU7V6X/EsJTib22lk84CpDV6meluBkpv077cgXCigq+5zYISia2ir8iR5Lcw
TY0FDp86a+gkOVex4gYDvq/wWr1GnAQ7X+2tq0Uv8zNpwNE45WvkBaiybQLcO+50
zEiZukNuBTuoafhqsuhHloIRJk9vrjFLB7AHHJdpgCx7ALv26n25tm5+Jm5zEQey
/nH6Gi3ScLQgzuKl29g7/5bXOEm5JsusRtEGGJooYwj222tWYA4AthKTo3yuP5+r
w53Yua1azlK2T110fgy31AwTzMVOAqKptznOyWNj1n8HyMgqb64on757xHJ1lIMF
VmLGzsFM0oHh9HU/E70bgpd8rdjIuMjwxgXjU9vkDlRXsBwbF+Gl3DhmehYChbDC
Q9u3haa/G0LNMBxsKmOE3cEAMf5LF08M/byNhi3Gt5dhFLCYv9pPOcWHIxSe1pdK
7161v0qC/VK8l0p8QczPTUa7G2AA8mG6R+17b8vqEy2TOKOda7CiSH3Md6nBCG5T
2fLbJbAsDvFtBftXKVR0GHB4Ws20Im3ytuSwmaOgqfWgPFhvDSwcK7J2IuUMjtis
9Fmjhaxzq5NfMAFPChh2+fqJJFtT479zWOItjuD49vZ8Loc5elaGwvDRx4uboDKH
juqUWQ3D8+Er/B/KsGkiGQ/TkKmPCSJbycbaGYM4xDyd7yH/mUG0zvvn1iBiufkG
KvSFCSqAZ6LJYIZ+k6uoc58ZOFVizapXQZQfCeVSFkn2WNujrgqtxGBJ52R9wGgg
DyQvAFyoEHBe+kxIQ+td03i4kUzSKUgMzmHX0x76kXRZDmjOu5n8mk0XuUWLWGjF
7/bfXwEqz68RxJZIwABN1i3mHUPBrA1BexhmQZn58JGlI6EMbu1+Se8nM6hbH04z
sOt8IzuyWP7xQ1VPviUFhboImsHvhFeLNLb99IJ+52KncMDX+N7O9gWF/K/lbR4K
+/pJRBCkI2NJDjY7ZhIllQDSnh7nawmhO4CTv5eCp3d/nYEU+CN4fL7f1SusMy+o
NgPgsgHiwwOSaV6LBEyFYdNI1HvuBYyf/cJM+nZlASGHpcjxIiWEeDpawSJbCTZD
0SAC6uC6TISUpW4Jr8yYKEd+mtmGmxpCdW3DnflvCSdSv0qb+Elr+xcVwIzzow2O
8zd5emJ3BmCyTIhwMUy1+fZ4U+iD/QUz9RDuaEd7ahWnQ9JpErd4rjm8VaawTaeb
p7yevoRPr4xe8j8s6SSvPKgenuGIcg3K5XuPukE4xkjayc3Ale1P+iQCxGTXpM/M
FNIZvTXHjbKi+5kskO0Orh4MI0CEc3LQNzN9O0hknaiiaHct1Baxaet33CqvSdOr
366hH8R6J82kabI35Wvew77JlHYKmmapSqxCmbYSnF+FpftXqO/B9NWrNxX2PYu/
cEQWFDdsliIqmAhwwqvtksKFl8qtxUO60ZmqMaIq2knvxELqzfY0TuZ8m+ht326U
Uuz1gfkxbRuYUbM+eWhZcT/rxI4POc0e77UCt/tLYdljXlGtakWM218dHQpD0r3w
XH/5yhiqO+jkAJLMELvQpeRxfCexk/ovuWn6QWIwwNj1+Kj5KKt7wMTKCVdYV4Lv
b50b9wFd7QPtXjPAD+/hPVxzqxJvlaRMC2VaAbXHhKAc+Lv3A595YnJwl7ilhSKX
y3hPjihLTmyAeVZbUGHRnN+Bh1DyyQ/9BSFwnfRpOdyscTXCZH3zhCnIagHdg0IX
wzRxYZSRHXrNJXiO8VDPbOoZdLtijb5aFIklJrpt7siYRyK/oUV2u3Ynx8zGiG3w
W34UYCZpMOZPK3H59BpiXi5NDR9W6p0T1UP+UHbIDYV0VFBPvIdniJeArA3TTw9m
+hUBbA5W/5HERBZ1wo9MIbDNI4LSv7kFU2PzfGYaImEyUW7KQ+LDXIq9usAxI5Lm
QznBePo7dCpHearFkqh5kkO5QIopwWRIvx7ESkRWI9fYy3ukKI8DmzlIdFbuGrrC
3UxnJ8y8XA+Beq+o8IamFwZSyfbLkPFi5iy8+kLmeDBp5q713tGplrxiIBE6RN44
di6H/uUBd1mUzucYJcic9f7mnTGrX6N12oQelS7kIBRacy1cegR1wO5fC7XJMnHN
9ii+1RwiOBlbuoIy6GmnFVrce95/OC6S2EFp2VrSybMVjCgdYpClatIITSZeZqa1
WamzrbIvou7+1LJbqP/As5vac7Op169+yDhSNhNlQOZhy/PkN1nVSlAPl1Sr5l5W
tg674/nnd1RKBRlsDMmtziPo/W1wTSfTxn3EmPK1WqNG8Iv7xUSyxvPXlxbcA4Yw
0Ot49NcjWqYrWeRXbOAkCq+BSqIc6qmA2yvjhwRou0fPGZ+waZcbQOgKJ0zvU1b7
VbFvlRoaEfoFWb34e7Xarq90Z4SSlb4vuFIYoJSZW2bNo742K35VflnWJPe2hhNb
KAEf7JaIEWIKu79KOswohSZLfk2XzxyK08E5oHQJGAwRb+2MvaFzckGYi7P7xCuz
qeozuM9sFsCos1VFS1VD5YUu9O5s55fSvLoO8ja3PybqtMcL+mX/YwXu1nok0CQ8
WA1TBSLdBlSQdP8Uad6sri0b+AM3IcrphU1OkOAA7M+CdptO1ovqjCPVsBNJ1ncx
Ivchx34w2v1PDGRL79LyEwMYjDM2DocqxerMRyJiafRwIfN0tPV559bqD63hpET9
tuNpGgnw5wGvDtTGNrRbcXam05FSAeqXw0Jz+UzWYyNB+NlP8mw+WJpFOU8T2MQz
j+GIjBwlOsOpgWkyu0y+7DBXHylKiWixRTlNNsHiAKq1MTBEdPoS+NOpZjFKvndU
s2j408AiwDqJ0S2VmWD1Pa4/QO7ncFbO8BZjSED30K5myt4CFku1GdO4ei8gyMtO
OafKoqVmqdFLLcecZGuXgIgN4P1efR2/iNP/2opR7IwHsle5yrJoLCLc3dAqmv63
hfgfRRihXnO5MKZyWVXyDr4DNhs29M7hkBbIzu2KdQVsbtm8v2pBBZf5brM1XPkA
jMgYeGAckH6P6foite0WpyNECoIxSB24FRiXCkzNirifHp3f2WrU7jYtFGaQ/3VW
WzocnPR6KAmB8NL5SJrRtyJu6he4x+fhT5PN3X63EEiKeYfMUuOj0bfLJmIUk6Zx
lAIG4QpdFeDOImllcePc7H8mSMfuWnNPRAf9zJoX2FMKTDjZO8GJUFkEqwm0m9iP
BbetPVNLyNyTfEzAI6LpP4sT3Vpzzud0JGE9f2SsRVJm6z2uztFYNgzWtcMfpuhk
bB7DUX90Ot2hJ5MTyLu+FQ6JSJXs1gcxOTvpF0divZUOJtiVkWor2Cw4ndhbHq0o
XCWzUz7cvBIcS2cXLFxsBjKp6n8vTVdzaPU4+Y56XqXe8PnDfzqwHDaAy7yPsfD3
GYIJR42414XLnOxahsEkpT2Qns5ea0azbKb+AVG4u7HeTYJbTPiQ8zD4bA3xAzI/
XH16HdnRonKkL6ABxOIZ6iNSYt9XBbXgHhnRQa0FRIGR8hjGoVcwvChJ7OWcWw6q
0oGEJVJLWv/ySh+6j5YPhmdotP9KP7otWeHqb476QpTAbgeEYL+ZN5K75fYHaACY
tlSnGUrMbNmvjS3AiTodYqMxYwM2MTkl4Qpn7kTq0sl271xgh2dV+mrRh0pXfjn/
ubevJ2KFF0GcHD3N1NJSKJyMyUg593fFC1cE2q7gTYOaBL0+yBMMdvJzkMuAsqHD
EBIrnI8yUYbiKEakmgelNWPjx+0dDUp0ecTdBaRo2pXOOIVd8wkYDemWRtNJJRbY
9VHHCHxzN1bHi7S20iGKr3hG+XmjMKITKcqU4YKysv5hgWJ5q2CrKOnWTZgCn3/8
wN2iTVGO73Ik6+q8pZVP8Y7JJ7CJqtiQ7EketFAZL90op0vqYfYpsRz3E/882Xh3
wgo52xI20DLnka5P+AWDD4oNmXEHkeMCNfuKiQ+jOVp4SKhLt/qoJLbsqeKzd6cv
IFkS+q4VelTfy1uxHPuwy8H3M4IEX0Ufd/lvjk5/vHukvs3hXS2+huDo0bKGQuTH
H8eGKL0+9ZrNmCpFVq0+ZCc45i8DSVbmireLNuaf6u9TR2Xpv31ENVoEqM97o7cZ
88RsDzP9F4GgKKrry7JssaHP393A7Fsl4IgeEd7wxYz4MuqfHA+VSaou/XtpYfp4
Kgc/EDLWOKy5dsBIEpIpcDM1G1XcFX8h9k8DW+mtVeq7GRnypDbwVTD4RW1SGUW/
4i3c4OutWRsojFltKNrupY4rnylSENlULVD9hNBVQctOEgR/ln0zoHMXazYTF17R
tRjNBwwk72VJ2epXgDejGUDk4oBaDOFZWPhP+Mh+oMQyP98ul+RPP+xj/oRS1fA3
qywsrnbEDD1+DevBXqU+i0PW1xoTF3sSnZsT1irgO7e8WMQCkQQHd8dKR4JwHljv
iZ0hdLBhZVyHxUfi68KaLLWWgMOMmROQ1P42+lEhU68cJRv4KU6FzSMP2C8DylPE
dnQo4pOQ4VH9+bsBfcSPq388ObQaPN6YXq4az+KjmXhpgOtcd2KP1I78ElmkAmcy
Tkaobyry7mrIn4Xtsrv4TxyZKW5AJJPMAZD/BANCXu8PzuzuUd/sF7X8mSr50qr9
QrrlO3I8Y2VS/BDz81JzZ24Re2SkxpAmEHTW6ai+LRa9NGblkyz+8vSEEA9ANEdb
ZeLNcjQuFRKzOB/54kPHb8xdhw7w3x2f/qC5XynM4tTz3oqhCb8b6O3M900VJtrj
MRnsav7V0wZtmownO3xEiYb6QNv7YZk38BsDv8eJmIerytmGiL5iMw9YGHqogiL3
8fnAkyxGjIDmY8ortkRHx2E9YkkXrCqVHM/3jo8OaPd73D50RSUyRcCld9Oy1WYt
CyWo6pdBCW1o5Zw/94dIYoOKGjkEsZ2jwBJoEKGM+f5pPrruT5m4IOs1flfsWKKJ
eVKuR0zkW+75kVECF7hrkfSF6azM4zU55ieeihIsF9nDO5Z6CjfIyGdR8dhz4bzG
wXwsf/Z25s8fF9Q/vUi5Z8X9a5GAICCeojapePJJTfHc+Gn9771cOkxpBa0gH0LK
sxbICcgpuWC+06EREvfVIMlcjzb+uwaNNdyYU7VnZvJ1RqgY74KUie1W44wTQNDL
mNt/UG2Y7y05PqUOWCtdHT0slqsEeowwW5J+wm3JlLfOfeR6fUruNaNnHp1XTPeg
Nzevg1Uz9tZnURjp7lMzim8Cfr5HnxYif7wEvBbit+IIBBYJIKA7Qzl+P5nTc/Dw
EZbcLMn2Wb/+sc8jlgB3sLwLq6EV5IAlFb2RwqZ3X5n15fWuCFZT+N5vwbHDTfWZ
+N+nRUQdwtIeBEJoN01g+jLTLB4OZjwwp+z9HeeyqI+Kjo1J/llYTiMiHt1LIJSm
wMru2m3KvZSr5P7MooFyEM1u3/j5SUcDT8SWv94T0dp3/LLTfyHplxNPc/cDZeDb
XJ6gF2s7NjjZllJm9amCamdxN09yQiwaWEU6WFE1AlPpmTJSUNaq9yeuYhtp9tgb
dGECSL2QM3AXpgEzIhfnZ6UlcQTHGL5WGx3af7BjB94B/60gLbTGjjpESRl6iI8X
MPsH5KXBJLvduNpUOMeMfqIyIBbd5jQtZ96N8JpLbrqU4+adzoaG55qNOcJwTOY/
vj74n1RJtU1V8/jfpJxDBJLKHyiufmUx4hTP9AejQXF9L5sGZImdf7v36CfjeUEG
w6ajfbG8fs5OdvmIgQu9SR+xaA3uZLjHWZWVu6nPR+noyV2xCUQQgbPDUAIDgXQF
2O/NjwAHYU67z5y5nnBv1PWS2T/hTRK49lZkl594I5mJhiL9zhudBRubtFuZhzms
oOaoYCAQ27nCCCOXjVOhxgxMOMMclJ4oFXCPPMYHYY8DDpfvHz2SAkby3sHBNHEq
AH8CvrKQvWuzx5nQrUhTg5Cn4DeNiZMIhCDzFeN7XRRqkh+TS4GgT/TPDMMcsinj
DetjAHWHv8/gRkw3FF2ihnVA9kz6fWXBpxQQs476+HaajP0ul5F8ZxFyzeze8xTZ
7iZt0rxwOVvkBj89DnAj2OSNaSfLCxeGY3ufVfWSsZc0F/B05YeScoKUHwTuYneI
DsasUTGBDyY+p9Iw9NNkbhNUNKBr3Vddh3+mCHBriN8Ia4Z6qv57sZwcx9FDlCDf
mykkeciHEEM4dVET51Dkc3uqNHcZbUh2fOyt//+czBvI2n4q3RhPE2ycztcppt13
KwoNjC5AY1aC/KgakEjt2gnl0Y1DtF3Vsgw9/G8i9NiUGTLPTvOF/t114fjo4bqc
a8S9pZecamlzWLBAgXRjeYo5gfk0y0A8h/SuGkEG3D6wArcG08mlyBWU4A2bW2ZP
Iq0noBtjEgB5rjyVaWigptpLUAEA2WFXLDlXqLyWIKAC3A51AQajsx89uotOqCfn
mZJFGOieyF7drlsHniXE2nTPlw+EVzYL20pBV+o7SiyYePPd8Pal5IxGNzY5Kobt
J6Kty1yewiDno/wOOQS0eoDbdK//NZ4alPOqLXVx+IfmQD/Ao4aT0DrJKd+WmOmq
kYCHW4h+FhepBmV5FC8vdi2BRPfgp2O5YLkLrmuewlpmOnDirFHSjPlrZmVCYtn2
wQxCc+9SYwWcjB7eMM1aLyVKHhJeUjOMwJ92SeUo0NMDcQiZak+4vTEDGR9RLIbx
NeOIqBk3KyF2AQJ17QCU8Mp6IB6JSdVq8BHq0J0yMuPMnkdFjbxOYE5l5TF90+9p
NEPLmXHcUUlYKb/C0On4CHEG5jaZhy9Rnj4cYhT5CXyUxpt5ha5OAW0kouN3jJb1
JnPSU8zG+U4mEwjGTTz6FEq3IFKxL26WQb5kK7fflKFhBwmYhsG2DN+5Va0VV2ZA
ytSk2ZhlZv9YOvpXpXYT+JhwXqj8TW8nzuK0aWCDvpwwOkAeUWql9V2PnDXJ7G8i
ZXCYca9shAxfxT7u/OrA3Yjv0hNT7xir01qyiyGoU5fpceP8KAVbAZvuVex2ehKp
r9qN0onfhzz028dyBIoYLWbPEePj1H7IxU2OyEPilyLthPmdQ/f523jFZcrj/JVk
ijFZTqVfSlLGkwTJ+c0ujeenITy0da1d+1OfpFiMDUJaINbxWUpKiAsd4bXVRmSV
8FJRXNHqUMOYxYOVna1ZLOsujk5vrxq/l257tvRfy6EBZAxHWJsiNauZ7QX1c2Vp
+1v9xu5RN8JnugsyIRg5gwLQIONvBk86/TzAHckeaqeAk2lSrpsO8zehtemCWk2x
wSmEobpqq2pgWlxBMYc7yaElEk3GRbIhEQ1zzz7fZmS74+20h1k3Nk279IiB8/+H
+FirsVfi3z6+PWPyiT3Q+BaO8Cw2Cb5Ck4lZxbPngFwBh2Q5SQhN8ddUdW+s2/AK
Hrc9Yqo2TMafS0gWpfndFLVPoorTlrj81UQN/+ptkpGE9RR3w9Fnvt/XIp4pboOV
ynDUtRmoPCinDG7m/wiKalHWVAcL5yJD+Npt8IDzFq72IipGwb005dQxLXfh6N8o
B/a2GDQgNbF2azMBG7Xhkc76IyB5/IZcCqVdDzweDod2mEYDYG342glLU4tATXVJ
NOEy/vctZnAag0SFJXkqGhC/ybnd/AhyiYoShpyr9870KUPqT6T0yI3PYj2gr9O+
tzH9gLLjGA1Y3vyiZYsH4GP8Xu27uBjpwRt5idKzhnU9nNOi6Ro9SjcWZUn3hpfI
fWDawVc6FFoC1OU+HYpjOjAzuPiVtMcR0VrpHhTcrEQRaM0LijzgOo+ZpvK1/N2j
N1nwYkaRBwx9oHoaLzyYgwo0ftIs5DI8Qx8lau8YQ0VmsmLLw40npIXfpqzKwdot
4yN5zGwg/3SjZw3LniPk4FOYJeFO7ZWHWqBdImumHyNhUSP33FawEVevhgCnyyVr
Bhc9ShsUNZsqQQIiAflvkLhvDvJ9gzxEG0dDfNRUEk5LhUzG49QExMOaJw/i0Ans
GX3raWw0qQuFJZNJzL1pXxHdhJO1+QV8LDBpMMhQ/NifztxK0wbmIFfuXBd0tr9n
0I9Ut2zPSnSwXVQ7GUWC7c1SID/VC0u6DJY7RI95zeyy3dwP6lqoH20HsgTKWSXo
LOrLJH/IGG9wZDPn2t2o5Zojgqa3mkB9ILQvNOOFl6/jneh8vesjIlklhBqll3fZ
YdGmWxHvG+1SFQvFsY9JOSBmCx/zBJ9x+RJ1ahoD2hZsYE0pC7oenGZ3bGACOmfr
QEOSMVBLXz2vI7sM8ajteuC+RrdwzHxIIZNQKdTqT6Iu33oITsUITDo4rtwoAtro
sGP1KWzepgRGYKPED58wjNwD2SFaf1qOGyrIyBL5hbqpse/1s7Hbk7ecpxrxjqQ5
p7rHOx2WHwSAE6xhNtbj8zaq0KUCHl/FBOcXVo8VdWXN9q5YH4PpcnudwWltFLmW
mamwwvE1RvNtQA92CYdEXUxzRlAaUtUFf+rUMW4qSI37JlcAoImukokj1cgjJhTu
ggogXnW3+MmzxGP08fLBUmZoOK0c2b03ExPWPaMfY5Dk4l4NFZwYj5GrINA3SLOe
jGpDoFepRjtb4hh2HmmkmpZlmhO3qldrCfGn2Qr2hozTRD4AqE5drqrbMg5kebSu
jrrsBbEz1Uer6tBiXVT5/Mkch1LkrHuCupOQXUhxJ8VeYRM4yyU9RaFJHvGFrNkC
5nIt67K2HxZqp9A6XPiVPMJdUnQgN6SaLvjr7Rfxrq1iljw3k8JGI9lfatMmFAqd
SHtzdTBjLc3RZKVr5yc28qHCRltbMQaM+vacwAAu+UU3qXuyBd1egBOb+CrIeI/f
DGhhmiTgjbkQVOTDDQQEuQy9lkBlLpOnI3OGi6opaIl41q7KTIJ9N1NxPh0GUVlL
vcfXq25l9jbnhqqXG5OjF7vNTOVux7Y5Zyu9jfR6+YIc0BWv1NXHnfCoWz97rD7n
pMysHEgEBZnHL5o7uMh7TNiiiwkWaSkJpxkcT67J5q/13rcMGT+sJxyeOHuKevYb
EZJH8/ae4LIUtgrQxlqHlykERttmzz/ELu08O1C8O6NirArckwryVKoNVnDeia3m
/8nwIQY02ZAkD7fNDT8OROBn/QAmgeUwRjLILMRVBR7oqKNN7/ULNV1VVadMVVsa
V/EL/4NmBKv0+FdNWui8tilROBYCr7YPO5jOX4gEmoYT57ujbS196648/TE3OQrU
dGoY/OxhW7oYWrO51fjrBdqDwF/XHLhLzgDnYQeYsXHlm32/utohQZjNsPjKPsTY
plSY08JjEbu+De2rp1439HdL1YON1uY4Y4tRMxoEZzs5Vr+sFZxnTn5jZ9gKR0Mu
2mTxuLKPR6cY1G+XeDJMa60iy/v8CNqt0s93U/TqI+n9tQQmpG7b8cpn5S+V5Cll
anp21TD/QCFf4r1hXE8hUf86xPZNcBp+sENv+XHWHwKhvkeeFOZHrrGyxG872PA7
wa25Mh1INRa1eeo1OsyTKVPd9y5pVflEaiuRcUD64bb6tfiC9rkRRJ5m+1/R13SQ
EPNzAFmf8vdmh/krNpaomtMv62Wij5oUED1Xw710Ox61TMXSlDWp8gstzka6bsZk
wiNoXH4mbkgtG8RWp5x8zbxqEXMSb6c7HP74Jk8hFM2JiJUl+0SqH3Ep0XfX+w89
LbcrSUREhEPpQwhiXOcNSxjaknr2NEDqxsUtoKZu+zQ9Ol2Hnece1iPJec/f5rC2
2I9xykODltAr9QXuI3mIiXaatxAUXYDE4FbnTy5MbptBgmpp0Pcm2xgmCdBZ6eAY
fjThkJcGJVg9z1j6Fp7K/wZU0/Y3s7xDx++p58BAUE6Oubprh1idG0VEHrq4E+JH
ILLTb1/6mNHlhOMJMcbSGc8+JIqPblBWQQ8yaW1d6eRIhZ1+QuFcXuSiDI66rbEz
Xgsrq5AHoLeI3Ti5N7CT463Qyv5fclf4ixTTMlbIUeQDu/L6VLe5ygpCUk1wLT4j
LSNCfFRp6XJAVIHFt0dubuhw+jNhapXMbhBQJIsOxWi2hFhsuy8TnuQE7npoXrbP
lMF6EAA/gbsaAacKPp51/orwWTFE1Uh5df/7bQ9HomIQkxlMEUrc7A2bDJ7G7hlM
yRO842uYjLprGYz7LdcaiXDQdmgQw9xrDXBDUHiON7kofa3r7y29pXS++r94358G
S2DRzbshhvS48XKASwqosRGdLurLn2ZiF9Zez/3yP23JLqrJeNtMhEuzrfeMpRIo
8skqwsBQ/PgdNYf+uh72hN9kz8W28Mctm2nuriP4w+f+mpR8t7AY+G7eafgBBjX5
iMi/YOiVcGjp8SimEAxSx6EHH1oxUmM7zQm6ERrOEqM+jnAoq1hnNxfpyp2Yb/BP
2rSPYjJ/RLycWuJwYOhcw6lgk04RDkKfJtfCsnp3cutu2IW8LvwAQsgNOdXn0hf+
SBu6eHUA1/5DWlvZjYsRPWjLLWo2I9CDKSKQq0V7YX69LahEfaPsijVD57I4cgUc
KT6T/ocqydp2qVEKjEZ1nNaZDiTW4d578EKmzkSVjIpY4nc8N99/254U2KG+BzZO
90KwyIhBNOfOGqdABrjKtTuMEwMvH8NQCvieq3z5DTkjhQUVlGAmibN+vk5YTs+D
7PiJal7/vVpYpL2wnJ0JGlpjPXa1606U+T5IkZy5XNRR18gQbYUqCYQswdANV1XN
CnAFftJIH0Wp+SKTGJ0fM7MOrufCgr7ZukYIGXe/W22CP0VSZh1qPch2jDtd2vFo
S5CoXntm+hSc5DyQLQ0sEQhYf4jj289FaA4STpWRbnhxNqrtGhK0vOZXmGPc1zXm
v/J6E28uCN18gYCo/2CPwmdWxcYuNgbIUsKJYcN+HOYJJE2Z7KCj+9NRqqhmVKyQ
y36HkDG92/Mxdjsert9vLfmoE4aQALxJDYIck39vxeIsSF15OEml+ozCyZQI4U/D
LDaDmcPcDilCP3X7vmNArJ9jpUxsPWK24oh5F7jWsH0ZzWlSwUvxoFkMVzy9mToq
SaIMzMlSYhyDlQL9nK6bzg9ruclr332uUy8/JCcdlT1m5OJkvhsNIlgig95o3szE
BATrKES9aHHS0Bgw5CzA+B2lFIZIXTB0UqJEI8fCYNPWtWA/TQpQfOaiWdp+V5iz
UGBKUZC1YyDKPwtZWX8Y4qz3tfHS7JcjlEwqWeyRAPI4adjqD5X1tX7rll6g3riD
G3cVg9J/NKRVpA//ZA2PUZe2bt6M+SzpGiDeMzVCvvWBg2uy6BbnMdqWR9JuW309
FAE8I7h4HibA65+6Y5dKhUPnVD9PxZ32DT43kZskUB1TPNBcZKfTrHqW6mYCyStd
80l4dboNaO6B8+DF50cg359hFByoaRJP3f6xmUbET/TSfUwk5vHghgqiXYcqNZiN
KASuYQoqUJ7aONCTTekAPuXTltss+Odw68NGo4RHP36lgTm8d4U7YWk+5jQoPP1R
sv0ndaxhQ78fKlUFrTDnUNokNiJtzMxPMMaNz8OWcBbCgWufTlxEZ5bgytjJ6+eI
TMccUxncxqNP+alFnMvx/naIQDUEJuMq78/F97WZVrvF/n+LlGcTaqHioAsOWF30
YlOsC/CXQTiY9wRzhidHuuxxzoQ5ckhmnR2vLXKHNehducY9jW+jUSU3/e/HsWhm
+CRjh1JKkkIKsdJCAIGOpnLkVJRbMNd4CHYM+AZLH7HRfOxTR59BKEx+X9KJZt8v
EvEa2MbY9FOXO1z4etIJMkN2xxSJpFPKdD0ufvKwQ/PoZqFKZmrBffZBtLHBdBM1
g8PDT5PNPruRlYJsTnJ/ViSP/hyCCMNICVJW/ZZM/2PTTNc2D9Q58PtBjKKI2wEP
e7f4u7dmyDO4g2xCvhMDkPZlvdOdeRa4ciKivBksnn8DatWYgD0I1dhWGUp09n58
s3v8cD/t6mn1ofloB7vOawFEMvbQjKFFYq0C0pm36XvfPMihMjYsQGoIcc3hpBmv
stmpu8T2Vm4vTmXWG2g5YAhsCtjtTua/4YX4a0XrpbNmCTqv5Nu7H3TerySjDxde
`pragma protect end_protected
