// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:32:31 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
cHnjtxnzSBilLZqXia6O+2wzeQcNqk1lettxNkqHLdsRaILwvfwa9Qu38cEnidgG
wxc0dxwbWhlSrNYi8QSJhEBiuX292oep6WpAevj7/QmFC8IJ2w6pJ2iFl2Bwp0bn
1MCODm/ZQd40HnYU++UqoestVrCOliTon0e6cKPZRfA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 48656)
cMOtXcKtPTmwziwin/KRq1ZwE9rsHKhTgDLGfmmOvSt6FsrZoZN2IQJX3TZful/5
JpPLduRp3lZ5gsOGPdVd1XWpmIqCIzM4/unvuSu470LccqhhDIG9KDtazBXx8uoc
8iTOCHP2lMQsKYW4RA0nci2wUX4GEC+Ac7ld2ekxvR3K0S/BmlgGJ/fYdI72U/tt
LsQyhg/5b0emM3DhE6oPF3OUcx603tnas+4EWc03QqM/uJ19qmgsaYZ3qQEVUz78
4HTFHEOgPcKWiHgU3yYoGiKb0sGTquY/KCHqtJbmFmDIc1oLM2w9af/L7q1p7Eh3
TaQrFjaxuRe2+m8JRFVMeYMSIEUvfd75KXr+SHFgjYFHKDb0G04OA3NnySbj3Xh2
UgTwCJLdNgvrQ74IWLDzku0N69w15A1XyodyytseSBcTOKbpCt5sEQPH0SDKfJX0
5wr2u3cJ5IxsuLzU0Awxk2ytTaqdFakFUaO2NR3D1yCJl6UdCl0UihaMdsH7TsvB
rVVOs5d/MgkVOoLeRr7V6Hce3GpnAsQQpdGjQ93+FxNNeqrF2cmKmWyosqqeKljp
fUcHPkGQaF4PUb3EApfimpx6jnoKSBLFtho3nzG7mLwyBuHML58BliFiABX3VJL7
rU73v6Qh4QRkPeLSajDouNeEuSpLZzoCSM4jb/axxhaNEhntKDM0H6FKh9XSGrw1
p97LA/wYGEOulbeZIijBitBQDRYQDRpcsuzSKhYLc0DlLUmIyzqW26zJazpLHIHC
P4jc2ag2/nxKG+H+vv1N2/JM+r24/O/SGMvZ2W9Bc2FjFevLEV7hjOT4n8hqPduY
7a8JfF5eVMzr/JTs84aRXDdVdNIHSzfUtJRK81lA9Wv0/OXz/t7iySBN8ss2sHXL
7ymSKR8T54otL97iJ+f0537s3bMaomyMgud+AMO3DIxU4AczFswn4XtNjKX6LDnU
IulHdUOo4iFDyrd3qN2D3KgWbQOnDmS5xOp1xzTy2+CidsRHYRPqjsnUp9DlO5am
ZN5NEEiQvamJdb1YfSbasCOwgW0GnaM07lUtYK5f4iCukzYN/vr7+S+EI65TxeiR
zvB3Cipvudq9N/Ft7LlALc0Jlhwe3+zSIIXCAK9Xo0YyFRvc9Z/OQxSdaNZBgW8y
i/Nl/dHmMD5JfEeizS0G95ND8Z0uYVDGY0l6hYtaMcDugOSNHJ44aLRQgFP3+JgI
ydysPyhkaenUU83c221I+23aBnRYkeO/dus+J/ZYZv1UYtDNTRPT27CjEpc887ZO
RaQqUdyGmLeI1iDwe05CgwhfRuZMNdIvVilIIGvWif8MkpxhWidTEW8eeVqBGaVS
YeJPrAlk44VkVEzx1y6He6uruckOF0DQIrkRSc6670ShAJQVZTwhOhWcsPTv51GH
i8dB4wAf8KUCMQ0pKXxtfuCYrAHdvgAYnD27nQkNPhOewqprU80vox7yCTJ2wH65
4XUrb6nux/6aQnTdj50DgZu0BeTdOq7vSKpQZhEtWnfLXdXhtIlhmrPm6ISB0EQy
nkZLli8ByHTXIfRpTL7bKi3HagEpbvMa9hhsZegJGp8NeAaGi+PlGZr9icC+GCWU
1SphJn3hgT9pDRJiMv9Tlo53oT9GTP14sO4lQxwc/f56tsv+dw8sN0/M4zkm0EqR
03146aTnnOizKpqZb4tViYt5xI5l8phPw4cc+nstngyOXXU2mBUm7GWXGJaYuB73
xq19KW+IJRsMjAKQAzR6ZrZrF/XEEc4abj5JUKA7dQCmFAPHamhDVyYn+uZQ/VJc
ak5+A/vtyCW5olS5tEeIfJXKtP+KoYEe9sJiAQKfdlKzhKoRM+v/olNzxH4xs8+J
zMWcSwMyoTbj9CP2et4bVzZ0+RkVtlqiiOeXmGMJsezB6Gh8JGlbNpZam+EiR9B4
h8H+sXBgHa+l5XfFI9wdT8wg3z0PwTrv8V8t0JK0HH+oeY2MimegaBbUmOqublme
hn0stQMK7QxeVrwN2Iwj0l3WpDk1xCJas+zqrTZBYq17k6WW4sktYZIKIUy8FaVc
ZALqxjYmFbN/8vOI4nf8yflPW9HCVNCTYFeD2UYP5WgM5simXxHQvchyngIOADqf
OpB+chxwVyDhy98bTjpI2PqWpEav+yrAI7EG3jW3ZXm0TqlxheCPiPf7KQ+BoFK3
RweMlk1g0UuK0nBZag8qVxsp9U1ylg/w38pet8vbrZvcbQbjEBWbLUFsWA2hZp4P
AZwSrXkvv0togOVrhEpL8r7GoTObkXjbXtHr/XWV4SuL55X5qfux3oAabfoYvwrJ
FQtx87jqHu2iNjH/cdOJ2ULZRS53j3bPTcl0RoOK1G0juj6lZbFLqBRMz0MHh8GY
IKzP23Bx+M3sF7Oigk9rqqPdqia4VLaf1yKlyFtkrv4GnevlykPOCTD9jTpUzTJ0
qV2uTWZ08j83dYN5HQZO/v/42CZzmQBB4z1gAWz2o53iV1NaAU+UAXL383hFES7e
DMEMM/LI5blxs8c8IhtsNRHXZlm2YWb63XU+vP5VyKR4bc+xE0nCvYo1j+iNkaCL
V7Jl1gWlHgZdn8zwMwuQbXtJYHzZ6oHL3Pdu99m+yr+tiBntCRNmwiTzAeQe2kQs
eS4Y0wcVgfh+bbrtuNBo79OxvOUbb2hvCv+x5ReVOMqN1HwCGZnds8M3uqYh4ywj
7Ui/tCOcaG2SJhYqGzazoJUKEggMr4n8Ksk9eCxzZCbRS1B0tikjS5U6gK4UiO97
uil1UApTUnaTiJ5zruKQpFirjRKv4VAPRM/c6vUrRJoseuR9Q9z5nQB/4wTCnEWw
IgpbEtz3Ye+r3+eCOqMPoNX5xkzZh8KgbLCCPWprz4Tr9Ra0jLLJsiVPKzoUTdOn
lWWamL62Y9xsIc/A2K4/Ad9/O8YfdyhR5nWWjqfT5CamnsmT1mH4rjCRNII3ZQTZ
VUuBRFtN2DLSJaog7o0puGLxgZ3POyl6ZjSv2iXxB+QnO0PabRN+Y/3AWugg3TEb
XhFPxEnThnYRx3neTNI8xWy2WgUp4QqS96vzSbHU+Jqk8JRMQnkLkWveJyfI7LK1
zkA882iUa/rxitB3I0P46/z09zBVxvtJbVIZD1prDMn7A5MKX0HgZkUrSN1Ql8sY
4x3R/xwfCt2pY5+r8tn0WfHI9RwCtaxBxqbM+jv0WMd9eCDptI80y57zORq653iF
RUytVK4Iz53CiIyBILMTgZLllJtkNscXHPEETrIdsW9nYwoCwbU3641kAbnHIBKh
w+QiXMat2saL2Ghl6aqAnrfRoT94deQX221TH5Bgxk+frJAS8+xgRdd0wpCaSaMP
XhlQiyluG0sQRpGZlj91rfPR4TYF3Hm9LysmYgemHyxmL8Qmx2K8aTXWG5HX1COs
aPp4gu+cdsPAVTUXfKbHU8EoTtqGOEPIawHOhiYv96D0ZkyJ2N2mjUiKmOf+EYkE
ox4rI3W3mZRKPRaRIrTeHuhnuaoamy8JZ+5rb8qvcPoJrbs9S2sKE0O9kAmHTg5t
RQoWhT0arzcRypNLRkuAjnuLydDDjeRi3Aa7IpWM9obPotwgncRg/AjUYpflIdYy
FUZLF7M1WgHIGNFQmzYxhbFaa/c3jMicYmBG1k5tGIv8F6j3jAiZN4XSzp+Ujz+A
Lg7hT2zQcpTLmTmQu/Fn0GgTOzXIBRBoOtU+52mr8qurU/5fcqdvBowZQ4hby+wY
Tb60CkhOnfMyTaGkequrLs9h8nIKhhwJ5hmgxfwt8TgxtW+WUOHKlAA+oXmpk/nh
3dB56QjFsKFLYPClPZ5W3dVuD35XoNoBuvzZZHk114yVKemBpzBS50ugbe5ngB5T
gUNgUFyrUzDNv4tbaV2YYKp1WsqmzhmwjDMRmFO0P8gYsLQztCcurmrbFnjdnHGH
O+tokZiihEfMbA1GUefuOauTwMSRpHHrGnL5nUWeiu14i/pSHcy6tF2hVX7EWi/0
TmDcOYj2QWKOiJ+XkZAGp2wPEhiYPqb1kPbUoGPOMklFtlz83FDZ8vIdFfpJuloh
ESwg/1Zpc/obuMg0R4Kzdojzn+1ELIiN4m2EOLVvpmFK2RsGI07nAn6zcpAO7DZm
ntXrgCLqUKziJd2qGAf4s+I350elALV7H3xj+dkyjRETiWgUORsy74HZFPZlY8WK
T0HYoraoArKyhOihPKLXT/IUHWTQdauXSZXweTlT7HO/yfYyvuHKeYpAB2hnT4wo
63o4hHjdYVaXlQCJBPnxK4QJFRGEZvGPqsN3+9zdYIIp8kWqFOesWMChNF8+/crM
l6tdUbHb8P6j/qWoqjJCXwT+5ywKtqWPg1K071WZzONMkVofk8IZGc20WqNI64a4
+vKlFEvy/QViLSBpiU9gg+WxV13tFqJwq2OH2rfpLzx5VFzoq+gjPhHXc5sjZOTq
g7xD1fFcglXayr1JvkBxuYBFmHJBlL2NZFIFOoouXYCYj/iCaDMw309hc6fxveeL
U0PkT9+tajhdzbi70NDcSFihTPGG1aK3fMVd18t25VWZgP12BTHTCdL0c4HjAFGf
ZGDCIrM/a/TpetGnAdBcGOdPTqzEeD/Z78A/o2dgfCD3LFlJlIvwN3kOa2Li0RXl
l4t1NJRu3T9h5eiuUstOtG7j+2u05FrdnXNQBraBQxQYQqJ42Ipau2QHFfWYF4+D
gQPdSTg33B8mVbwyHKfDTDXZCmSGSpdmi6GQBKHJfPVLhsUAJWaFjM6GIkDMRmSw
iOLX8MIcLQ8LjhVMXTT0xxGHbophOGX6EUeDoRPeaJkwIKazR85t64BnMcoq3RT9
5iH5A7Tr0z0NpuZH+E2kXFHpZ6njYjB3vWNoZyEp8VrOmjJR0swCYNKB6ZNQ84ZO
wU4rNGsVJzlqQK6fSeIC8MgBAo7Io9LpMR2owbczudvX8ZvGxGHtIXj3wO6adzhv
6mG3jy3H98Qa+YZNTAxOXbA8q2yylAWSzjhAlzu4IqS62j0/sc1pdFcJkqNhsYMf
zod3XEoI3g2+RodgiFINK6ap963w75DGXAyX2hwujk4F2khdex3UIdxz70T0ckgk
Smpmx9g3bFp7SL3UdXli825yXwtzq7BqQRmRPtttAAb5yyoTZ8m7bcBtgQi0f3KD
Vf9HPgpFByns35DY3iDqY+8kvHHxgbJkaXu2kw8NJuInqhiciH5zOuvtk1z5/BRA
cGDVdIDnlr6MwpKoS0TPfDWaDHA8pnmmYRT3iFVXmmcuZyVBWsbHjdlqYjy+5oyC
UaGgAiRI7HtjfeYxtubB9bj7XuETtyLFd2s8nnOCSb4PdaLDABbCmoDPeavZjOpo
9/h4zjN/5J1r38rEf4jhh/7TXtMLITTgNwCzPaIGlAXQsvyoxomIGUp1Zj2WAMNo
p6lfktG8ZClMJCpgg5B+eWfFZZo82SmLYcNDZF7CvLO+ZJu5bpVMlH7Etp+8dU4j
0YyX/RDi+EQ3PETg21YHhGWkqFWGSkyU/duLa4BGigomm7frLxfbYjeQOGuQ+X3D
a1rEpN0DOBynLYKEZZjVqCMVp8K2+vABgq49hyHoSygukNXIdHOBDZwfM7B8Wytx
QoY7c3iKLWuKD5INa5Z+tmTovkCpzlj7JP9Jf/8hEXFTj7NYmyCPB209gW2iI/Vp
wQ7Eb60JWo10ENauLfkGpL+q9LzX7BSNaa4Nn1JNcbgAro9w3ucOlaGhlonf4ZFG
HUidKVtnTtVLm3pEuXjoYFVSUwRW1pRbZIGKS0EGx4+9SqHCPXiaeJ7AJKLe9+Rw
W1HcJhl9LlOJB9VCbCyCYFvpRZDav4+smg+jZS8RtiFeBBg+DxtdENI37OYB6dSd
LcD9QXUlJRd1O8KSU/maIKPJppWDXMYIcOYoO6FRJWWdROpg1SMgGzYL4AEB9BmW
ZRDpDB90XYhjwkMvLRri7gsgmIccX3Qv89AvpS3TAFF2L8eoG5FyO+wTMNxapp29
UtLL1HA0rcNJBQLcAwjIVpTTWmorNRENo3t6roQTXk/QVGhLt8nTVlNterLeTfB5
DFgzTmXs9kjpqYuHs3p51/O/g+rQtQrwscVjpJsdFtvxvUgsbbZdoOYrWVr4HJIx
dJiFFDg4M3BeuvFHKiGs/DU6ZB5bfFuq1rcA/sdbjLF50bZRH4V5BEONw5WLH9Zv
W0sB81G9TBpGlmW21/Kx+IJn829sSgcyKHRRXK4uZWe1YepaBZtxr7xcAV/BI6/i
nfVCaWOJRr3y9c3sPba+TN8CdGwgTu0RGgWgcnP+8BwhPcTBdhBN8wQEotFwdJBk
HfLW0WsxUZUiuEZn2f1CE9Frw1ejVmRIKySbnyIZxrpEeWCnZO7zN4+Gl3vDIzJl
QhHRjTcCvlXfDE+fEkuq1gh0Tt/CKh/30rorV7YhrTVgkcJTjLsRxio8XiEGdTIt
Ya0gsQZkyrxN3aHuzjak6jwoGFsDClvIwbv6tFCZBgytvx2dQBep+c3jK/GA7uqi
r7Kswha1stiSWUcOwJ1U++9phV12EzwAPOp5GsoG0Kvi/nXkSx87kutBAU8rU2IY
EvU7fvYf2o3/r/1h8T57GJ2JBWFH2pDM23h5Mz/2IhfrWpQAlxi8mxOaNSkVFXfW
R0bPWIMTK5+nIKFmPC5EhVkFohoa8dFtM05CtymCKOObh6Yfb9v1N9aKwSeuLlbD
nNTIFeyPVhIstVTtGXpvnvkwz6gwuAljFoV4rET+u5yRU+OsPAlZn2lDwsaSFb++
k1dRFjkEUzrMNp9Bwewtr/Esi4ICN+Zu1eXUghp6Lo1lWJ83TjMKZVrST1fqHfGS
lwF9tiSX3/n7TM8K2ZZkSQ8VpxmXdS9zphxPBnvlJBRAGbe9dEuF5gfhobrwPA4v
fedBmfFmin2jedlvY5gKIoibW1VkzeYeexDgr30vGD7lsBFtDmBVIb1HraTcP1uG
gBh2LsSI6MCQQZrY6aOfi61RM3Tc/WjqijcGVUp71Wb25b6gzEgIVvG9RBlE/tS/
NP5xzsIxjdXB39Q6YvKotaZPn6BaVpHoLFjHp61x7huJz4a7yrMhze3GgPf4DtoY
IF/aur7F+5onNV6XJn02nTKaWZUZzrefjhBOQ7Lp0WAw4l7UdkLcQ+t6KrklPNHL
oicMLvTgsbVrvzyqoPr6qtC2sccg4Vgg4SwObdVms7AUgy+13V9DmSFYf6Hc2tGd
o7OyPBAg0QfyENtT6A5SPezAGiLIIis1ExPJ8YIC3ZmTLp1hMtimw6m6MxVvlGB6
ZI/kL/ziJg//B3oTJeiwYiVBMQeIF67Rk49k/cWkubHH8U9kolUUMsy7aVBedSTx
U4lO2AjmhI+etEQVIFu9ue4C27e0wuwPKa/riwl48IP/Tk54l3mninsT5HRcueeE
sLbcbkRnt/9pl0xgVLefcU4RCsklDWjfQ+DY+jUnJGdNzqCl0TK+hTxgVqQq+MLw
DxzHVDaxnlLy3fLDI+zqjdlB6CVe5+EknbuxJ0csqtSZ0ri2TTN6HqlhGkos2PqC
0ab7BtbpGdPt14lIOHcn4Hk2259kQ/ECOJqfpYYlNyi6GhJnvPIni9XQy4Xc6F9T
zqdN8DW97rFYJSN2nveG0Y2Gp62NAwqYQaLodavD2m9Kc2yiY4/5xUY/V3+HHFMM
6CmjFbVSdHGqPSPLzB9rnfKNTGC8W7UnNdCvy+Q7yb+j9ZxZGtNZcXVagBVzoy4n
eo/wYpEfBibEyaqryV7SU6XTpSubJCKnAlywTkZD8csErDK3LOSW+63p5FzRU6HP
FCrDvdVSTkmHrPUpuLr1FY7hXA5kpXWwnOzFhBjB9zRGBnM5Vtf9WzVnb8v36EWA
KtgZAmhmnmFjJIVEBXio7eHyT1v3LDPcj58t0lRABmSWgDDREzz4GtkHwCK3fQoQ
IQF5av5Vo4+MVbM6HRo7BPjpizusF60bsSfyLSa4LWIk7PREvM6UuvsGp+X6+ej7
4yHgRLvg8tSBIakkD/3y9kDP0M52aRv+Ic0ahDKdNdA1PGC2kMTvR8bUxxtiLC+7
aRFx4smtiVxioNOZvvbvNPRN8qAwTlXJhFXZpOzxUM2P5PGvN2t6WryfUt6TTmkb
hpjywPdR2Mwr6iaQ4NuMHfEAjsLzeL67REQ1tu/NcdpegpRTJPxaImqnFHUAwDAs
HqmjGaxXNhGUV5EYHpW0iFf1Ew74Zpkb2UokuZGJrX8WN0oWAQU7P93xLgqaUaCt
Y0GgRaPSsVqgj01+Arj8jynz2+8swRazKIEHKv7rpkJmXYCpGqBYpFoLUjkR/hHB
i5DMYXcIjzLGBtB+YDnfIos1HTct7+W+zS7p7mEkE2NJH641PtJjD/T5udYEtZVe
EEygAE/Zg0A46Dpl7V3JZZ8WcPuvQ6fQkZNZjayrGjyrdHRK8317wMyzfgpsHc9o
ZaddSvoW+YFK9umiUtgxX9DZjqtDzVT4cRMQE6ddPqHUwn6fu4oFpIhL2iDTJfPL
paQgtxTMHQ/bTt1HAttY7uj6LHV//67C7VRzNxtIX+e1Mt6NDr0KBJ+bGvRRIfWn
JbHOmEiXpwRgRkls2NsApf7LtmkHj9PI4Psd0MchMkp5+8WxDOCoVOG9CUjw2Pbe
FbbK3+VxPe5Wu/Yw49dhqiCJNpehozYIiL/+fgSa2GUgTwqdbySVQZ4ObR2LPcih
FwCXVCj1WzK9lQfcd/cDTmFt9ID9pf9IBKG8MqIi0uWMdEKzUYbvqgSvsNtHo9en
ySMvEp0pCoPv2njJSa7bULnyjyv1y4re6OnXTeYA27VrqzQMc/Xir/ciWLRvLnFu
6sLz2ikWRGzX02u8FDJhJSw4FRIZdVkKHb/fYHUDgd3+0zf8JCYeHtOevCqb4KIP
z14egK8pbzTcV6QB6qnxDZOJcrPh2plaujZz8CebaTSOTBUlfBI8Ft1ldNqAj8Rr
fiVTAB7GSCeCf1CLTZKRMuFBoEeD/VHSCg6Gb19RJhry1f8ca+GG1CC7OGfkdgLY
rdTnumhlwOvW5vsIvNZ/6BxTnsuUQLDw/hqDCjcvYHhf6MJFPoXcomDx40CVnxo7
wuZ6PCpuOZaACJarmVi2NL+odDEa3yi9hxnt3+BCBQWdG3lHCpSJSGoYHnHkdggY
/LtXHQ1D3k31GQ7EXFVGF7dMteeQDF89lDI6TdjGxQauAeNlf5sU0hpDPNE1bA21
MF+pOMppSaU0eQcHvbsrKuRLM6QJGg8ZZjFCLuS5WxvMOyBj4Piz5N8TCPeEZCsH
5yUjfqbgPzsUtSuMynd8xQfLGVzi3w0QZaIsEBEMtOL/y0UpwoEaXrD1E1JMVq4L
ijKug34mGUm+b4xTJQSaHJWr1U4tflH1vg84erMBnNmsTRkYSFU1TCaC88ghwv5o
245ZNEBC1t58Z5QPduOaKo9Sr7fGTL4yxDZPA6zHak3UK3NXO32dDpQ3MUHObqhZ
7SFLrWo/6i3J7Jd5waN0Nl8ZuXJMbp4Ca3gf3o8z3SSKZ3/rwEV+z/sG7HiB1lo+
sZAvy1CgIASt6NjU/SdcjGaubwO2KX633Flb2GGG6bkl4fMnV9qCpl8hOuJ3jJKl
Upb6wNI92mH6p5v9s0RzqRIRfCQL+UpTMY0j2/NkgghbykbmtTxXtgbqzYLY4VoA
j7SJ7sXgVcRIs9EDBKL710jIOmUrXZQYxmXi8ZQJ+J2V0BnRLwE9dMISzCkDV7Zo
Bje6lBailVkucByHAiizQm7AvLpcF1Bn040sA3eEwmsT9HnVo7Q8mo/FlnYVgtLV
aB5AVUi7s0CHRp+bIZ1BEp5xChucOo+bmYRz3uGzgaXbvIH3anx2HLSqChubPkJ1
m45LUx7Qj+5Qz4qWKkPdIJCLK1UskioN7kdxUDw9YDdPH9Hx7KUm6n+Bc7k+eMB1
SAHJVIDWRXh3bx/hLDUebX3N0tuNVW5BygKqxsfL70z5XqjZPeiDe1XsaHt5zj8f
JK5rrWBUPfwpNWX19juLFbkcGleXJhpwUdyFEjnOoen3oQe8tl9U+vcPyqiFvSX/
9zZnCJwsCNr/N9kC4qeMw+WBsfOvRW5pRuyX3qP5tDsl2fTLhSYcRGGiVMW3oEmL
6yhHzNr6nyb9Q68lP45uuR8lw/r7ZjNeJJdUN2lDw7kxQ6MyBgGeKhbRjgD3ixul
tP6lWuFxiJdugQnkEbMeQ07LKZNY9ROgALap8QKsnRb9+GJFBzm2I9IFF9xXhiYN
nOlPp670OBY5dutGPJhcoxq5ZC4cDYCEZF1IzTPsmvadEDJX227swvZRTa0OS13X
46RtFCk6AsBQ5IVNlP+Z3d1tQ6p3lvVuI6bP4IVtrqtimYkNbDEteesF+sJMzgf8
9CoshdES7ksNvF+gT+7iOhisvrZk5vka89mCoYsdyGLa7wx/KoF2/jMPZTlVFCSY
pFQ4puvxNClKTWmDDZo45KgNl03tWyI6XnvX/5hQWyOeo58dhGJtvsWgTBhc93xn
/n+425YrXqVUpbCdZbcFGuh3BEcqPkKZi38R5OACZfu7NPDK+V8lixm9YJNT5RLL
fhOjxriViVw6FU20gTFoq6Fn0KouE7d+td9mfYTl/Y+BPHSzuuiO7JUmUnsnaqnK
K8mixC8T1GJnwQbXgIdj1l0Qw6U8dWMx3uQKHW1F7QAulOssD4s/GaU0vewflQkb
aYpAv36WNILjOfhAOAzTm60ZEIzVPLaDcYXSQzPlWZap3gS895btzfJ433kQpnO+
qJUBPxJN3VsO9APp/l5BRHtYWYZxZd+2mE/kCC9pD3u8/MW2SntfDh6DkY0Kz1c1
u662UXUWKXN9cYTXPfphtRP04kIiiAEjQ4EQ455EBRwBfPFoVl53IaQYv4YygJ6V
z4793payEwXmVG8DJRGRWy8PubmYfLM51LAdDPJMV4RYX5EYHYjuwtfuvwFw6rlI
XFemy8GaNQtqaABWAgXebI7mnYRppB3T0wdBxNnzZEPEzg7P14C93kNfyDyvTwH1
G9nHANBdgy0cyLk5fJsQO06KfahoPW6Z5FUc94HICxTasALmkVLRUfedktvTsddW
ERZMwdTyfoc4CHW/GcnLlCcENlNiWZ5/xJwVYTSgkZZzQHvLigC8geBdyT2sShkZ
j4dDO9V6dVVMr+mmSQhTYbpea7woiez3fIbGS8hg8uLjAk6hIWEWIYJYzg3F4Un5
K9VtfMd940Lv0Tw0XUogSc/Nsz3wnNp7+mziMyDU5tC7UnTeAywo+HIK3kcC7fAw
qn9m3cxyNGla7I5tzTWiZ2WH0Z4X3gdRSVdn5swe+lzsVlIqMcWloJ5TYrZaV5tE
2bUdwFu8TWBEMqyP0mcRZszwt4NFmA7MsNxcAO4XDdaAp63e19y0fD9jiNMW1uFy
1rAip1TBbyzlYAkRYt1x3aa/y4pfnxR527FfFcy8ourXuUjEIFZ0FZLg6jNegiUo
nKJwZa1cTLdpYBbOzRtiDJMD20/RXniLCEYmBhWdUZR+8PdfxGNZQMIkCMUMXl7m
bAIfuvIdPHI+XZ988/n+BMT3ob/tMkyGCnwxVTWETenQEEeqhUxntsqkKVoWTCI3
WtS0dRHy8/PBInUg6595n8wxg8alqz4plpokm5TR//mq+IvBWUwn6aW5xhHqz+SF
UqV+1YblTxJc+cfuHObtCInvQre5wDnDOXUd9GUj+Eu/TC9YfY+pWgpTuZwzgKGk
IzPRB/ouPFuk2Ms/9xP9VlOao7APRNKi3s0RJwzDvgFJzAzKRTFin1amzsEHVOYE
PoGEOH5OkYFFVeh9eUsGM/arix9tDf9EWm2QF1RN25oLT2aIyvJwFp89Cg/k/vUX
6leNp22mBN5orWiYhWanK2TT3hZ1acII5H/bib7vnj/m2KLkdrXYqDNPhckX5bT2
/eVsTHJsBpctpBmYVVwpCdjgkDLKYLiaGAOYg75rKagxgPZ0ImNpYm3al0eYaDVa
gxlLcU3TnCqsYz7tyekpgnLCpLdgCaXIO8x2pkgrkpoYbuM9JKGSltX2OhmaFkCl
xgjFcgLTtcFXKgq0qpoJcvnEfk0ywUZ7O/SmYpQeinFYvIlh/vomv3/5ACURfs3U
V/fC+z3FZ0Eo3rjgkHDTl9ZlK/H7DkbOWLel4/kiS/HR3jKqTxIxbPbQ4yYUQhwD
znzdWeyStQ/qt0gGfkE/6h13r+wbLLE8mmFw9P8b4kTUO2sKrMUR9vXLmxjoPk/H
CVLxlCEauNdS7GGbMoy7c433s6tysr14aORp6kJcVIKYpzyackS0yhLfuHI67cQy
0P9STkE2nx7Gcj5QclmgGd5ObS+R26v/VljAJUpo4EjDk2EZsU/Iv9D9Jp4Z/ES+
Exc06wGKuLbwfcCmv7/9yJUMeVQYER40B+9GsQ8odKgRMztQj8Zy0VqeXOovWEgG
S2Cw7zH4nUJMjTheBBvk6lqdaAxRbJycZM8SeNMGyb2MQIdh023Ofq/wV74s0zlZ
riotnDIBN3DL5BNDGmw1+8M+BTLLsdq81sLjkySfehW8J+uaHWhSqIMEamHkO6K/
YBx332MmqqpB+mCut2iZT+8LxH7r4WqljgBWEc+kPUtzWSaDkIDmWM4DFufF4d19
YLzprPpZb/ATSFTXzcmmbMLoYv+/h6Euc3hki2tDoLIGpGbZ6LVq3QnUNUoG0ugy
couUZJOubhh/H0PfJHMsFSUkrKAEh7nqoJq6hag6VjY09A4CDRvNThkZ8ms8s1yZ
kN0vkL8qpFyojxzRfyEnG1lSYj1siO2LmY2Kn7rAZ62Grlfci3ovuI9cKy57p5vb
FASf+KglqwfITMy+glT3UOmbLB31rr5kYBRku9E7B4epWTvRUEQlxxTCG+hEfyCc
cVirztPnLsVKrivhiOzt8zbkoXlzYZFtluZvR/KC/sPMcMZbQtNrMeOsCpsUWbMs
2SJzRYTnL7J8FUAEZIg2wYUWeYvjBDGfycoMQLopL1VizyEIgkeg6Esb68huxz2P
g1W6MSN4sOsy9y49XSkFgm2ejptP1Y1BlsophZVZzAZwTvURYhIm747qPDM3T5r+
arUR9mrbwrY4WKnJ1gcej/Jx6oESmSNI83WxIgSKimAm3jaUbe7lSHgektRZvKzK
EePEwyhdlqNKy+NbSyhBaClJelKLxNrdb9HOmwrJvgWYdmA4hKOAckzcpCM/Mwa3
pn3NSxowescPBwHNvVJj7kQb6/POXmoqbhv4kw2IdxKARGnPJczFoCKtq1n2306T
ugcM4lca+9OSXQIaXr32SceNl3o2ZXf0W1AhRoC29uEPdP4WCeUpVbzbcTxGZ7Us
CoTKUwRCbskgYGv9e8Nrzy/H90kxuY1l4/92/KcdaJT9D/NxKFVs1PK8j6AJAH1v
pN91ejHZLFql95Hi+SZPgE/AjGWgyOF92L4OUV9+2rJU+TkVh4hnHvi6B2IIXYrn
VcMhqLIPugAwO92zryNdENHbQt0ZO01DhsiI4TVzGLMECnZjpXL9ZS/2OcCkNy1o
2NPGT/ooP78VAlv5xtqquXU7pnTOUyyPMSXjY3aWk+LSKbY7Qw867LSLisLfNAQg
n+3VDpUccFiCY9ZIeRYbA8k6KuFvxJr9DKm2h94/PqVypNwLAu1LnxyACFW6W5G9
CyMJcF7AzVtIivCQIkwa1LkPTVIpYpnFqk6WAGvA/EnRedS62ClazH/s5r1kBTQp
KD5g6CtqZT0wCiqc9OaYqjLj51jITiRemGzQ9HZclVCcMDeo/sQXtba72NApTZ/J
c/ulOkLE477h+b8HLBMikrJVF6o7edzi513oVNVzNzWdoOle1OZHrJQ7vP5JsN4b
9rshNh9B+pigNXtSRRtFYyAuVTatFCDFcUNQEMb6gciK3d4PGURvGOG0KiadGE6f
TZkvJAYu0Yx/e8/Vbk6ww7P0Yw5P1BR4JF+MunLdn4UEBVUAtrmaOSGfmQiAoxvr
hwtdeDmedMyi91wSbYNJSQAWUaBYuf8T0tPxVce+wpg9aLRzf5+IiODveHzxygnh
JKgeB1cMa8osv3jqjVWJICebmOSUvRf6OsIRon/HThBlYKhcyjBh/YiBYg+QMQYQ
akqTwNYVND00VCbwfyud4s/bTLRAGR/XjIziSRbIEk68MIG9y1KjCPuBVu8ePHks
oZTQaVaGRBJIHT18Z81fhq5xwM3FaR8/+7QMrRKAsZKDSCFfwBOhDKBYDTsaUF41
vz7TabHUkRxPk9lWYFDZzBowSVEtR6X7MKj99fy69kdtizKiGk8sUD8jEZbCvIaQ
IQdwBLs907yUxXPzAbexnF5ST3eqxz1tjZrN2o24a+kNSXs24cKwJTqpLL1e0Z9L
D76GIGiEwtyE2JkoEqsblYZ349Ghx7L2m9Ve8ZC99hxzEdTusAn/YzKxCCRoJW+b
4i36F+yOWhfT8FvPKAH+6rhPEwIqByWceJubffQJLbE3h/Rru3A1qNBeOifl3jdC
9riB/l6zF0v7mDLrzW2pPQq2DcPstZMzrHgU5TbXTXhYcg0sR0EqxTQpWwajtwwA
/sKZ+FUslHgawBkfRZ0p7MkEYmUgCsLFdaCXk4c9DdeACdZ4N7/9UjVI9WBu6Ckk
6jr354E8l+CPZ71qgQb5lK/KDc03gy4666lp9E+mONaZtUHK2Cszvjaj65omLGYq
bcdbgBecd/snEJ1OX80/zTF+J+KAxyXc6qbsMaxubwVhYSWrbBPEele+AM/ww+Vz
swoIi9V3LJsB92CGR7PCakEYD/03mVfc9dknirjj0x2phx/IZfeoL2zdUlsU63IO
XCjko8EaSutjx8hn4EU6uaNh0YtqmFucIsdE9I4cTq+2y/kRlu0RA6wB+KmPdw1D
2D+XbjNCU0Pbtd+M2d6WPcxjh1iVOhupO6hXYg6QzIQWegeK9em7jWSD0giUDEvd
PM8rpyCn8bxymRpk+VkTp0DLTBHsqD3401Dp6Xlfd24mCxgjDzX6dyDMIGF99dRx
SjhsY13gvBIRaf3SiYJwFsqKe+dEiSklZ8hs6R65sGXRt3+j8v8dk8HZDtKBHx06
ea7WeMN5JWxUMCR/Fwdyn/D8b/J1kZtwnQe/5lPhKlaQNJYoJuRjwX2qIJ4cwJsL
jGf/wanhtIX9qlCkmh2skxQ3a/XswPut6Hfl12TwS3xeKQKv/x2b+SuEwR/kw5tc
w2ZQpiapapQn/q0At2UFbVSnEB6AImuT82WlAAsMfi22tFYyJTQoIRly424eikR8
PruJr3epZWrdlt6C7T1mP0SdlseGCJZDiQCryw7h9U9wQ49AHLCAYDYH9cMgSEyi
48TfRyo5bVaO4KcfiiUtjNqwEB01BiBQCF5llviIYuisDqRVQa95xSPZcfEGdfbR
lZji2wPO9PmJcikWch15JV6Yq4ZiG14oPcTWyuMy6eJ57avKfqCoZPeRA+OuE7se
g9K59fAuVAlqG9UrsdPGHhJhZ4RzrDzLOQCxLZ2pj9x7egj4ifZXGAXIQpg+JS/a
aNSOf+TOyLkmFIeD9v7EL35D47aP3DFyYJR29XaaucEAW4wXuGSt/z9rgJUf58q7
OA9oSfvglv0fps3jgVFhak20adB+rTb/8dn91YgL5EBh1qk0fJXMhO49Pqvfy5C7
6iOZSW/cMaV1L/fwy8XowsrsSHdCniZRaExWjHaaXl8+WJ5NlcU8qdiPc5H/hZUm
4SXAN6kVAvoqSyWQqtxuHHqRsZrXbJjG25DFiygwzUFiwJnv8ouwKgOduRIJU8ci
ohqoGz9Gq5zEUoUEQBMJUccxD+yAxnwAlYZYmmBKi8jko/ByB9ZR1AHlzMfQvXi8
Buf+N/bwkLcwCjFs/8i/n2l5uVLiH6/YBcdaexGP8lJGQ0oBANDGXe1AEYNVITsP
npFc5/9QvZqkpzImwtJgB8CaE5aafhSIV4T2/UIvaZdKY5dOVhqkOFXP3hPaEF5s
IdW7RaXHGK4pufXxhx05XEyOq6fOssO9oAZyS+QnPn51BN+IToIRch4gmHFCS+KI
T7PUBKEjv3HH/MUwUgb/UT1EY5K7lTnGcM9aszHD53OKXghKqvMDdWHXLNAMIw0e
/duJP3Jgb4LTBdvaTQZz/ajZn6Su52inrdx/7R1ueEfadF/gUNWUUk0n3DHP+WgV
NZtDKBepB1vXtWogGmscVnPd8PveR3QKkV14JE6EZKf2emPKAjq14290379HzUk+
Z1Na0EF6lrn8kv5dmH2Z6CPCUmy9oTSP1bOS1mB+bhUXvRt1CdChYpOHrS+gLct/
EDmrTERS7qTk6nuO5MTIeflBJ8+064JNKNYvwqI5rr29v3ozHIknX2S5DT4Mqfg5
7zOkk5RZmnr3gtNhOfhGtu/YoKSeuww2ai6LVE/EL0jihxwEiMfqRfyduD0gfkIF
EG5GqkAv6lLmvSG7KrC69V32tTo0QuqpV/Yj2txbJKUh/sFrO8ccdWOviG1GZ0A4
px7aoTkwUJM7rQvz4urOt0SPbsDSPGdAhCkXGKpOIFhNwE+Yc/teATx+gwy+g/VT
76JPDRYInIxMw4fC5TvlgkVcZrpQ55CsDYs5wSA/OnNr50t70PR6dK7P9c5d6CNb
mOw2sFSLs7h756R/APt/oMKBSDPW8TpL7sZyzxbgjS9YjaZiTkp1Qo2RpZ/f4qqH
XeAo7FEt1C1PDyWk7zM99iSAhfRMETcZIsdgR8/UqD4TkggeXmUjr1PsGXHsP8TE
5wLgqmxVq/AOtJbP1R4wDEFsYZEpvB91+WU5CtHI85qex8fpkat9Cme/gaKXjueo
FdQIRVdSNF2MzcGYadDBa7ePycXNxkl5rOqUB/Hl2bLS7C3GOaeSyp9Ho+/YS6FT
ejFKIOZZO7fRIIOuIL9vJ69v/kiEPRuJz9xsTk0PVpeDhDHhce6NlyY7bb8xeYJs
cuWd94BL/dyVjhspfE4WtXO7KxcrtNkYGRVzzEUYqjXlyndaNpGGnOgTWJX+DwLb
C8mezjpymfaNecSo13MvYCCtT8U819bpX8A+jWsbAMdpaQ7ZWTitqo14b3raOGpD
WBYYs4z4WkxEiQSQNzj0Oo9G7VN7xvZYXBBkI9c38f9JC20r8DuAIjy4ZQOjBnKr
7fSAU5TddXx9rlRuKqXYeTwTKnT12UX/4WMb2i7nKasa3vDxmIdHPbn0BiIQF6pE
MNaJoLbE8FOT8GH4J0/Clewy4zG6h41TaZZAuLOObxUl4b97+Jhy0cjznghtQpm/
/cUF5/vxpw5/WtXVFk2WIevz7qeSuSbmNbhR4jDpyGuo9V/MpgZBJBDssuu+BaAn
qkCjdJVIGX+4oDPKLajKLh0IpeV4aPlu1YUZWeEKvrOvICfhdIpI6JinYLdxdsSn
+CGPm/A7dayd7fgoBZF7IGKQAUTQD76oby59MdbNIVmQZUeThavIxTcKPwwpTLoZ
JOE5VrAXQ+BQrz0UAvKP70xcOiS6iVIQcpaN/hKasb8o8ZllHS9ZZK/i98vNTkfu
jE4Zm7fMzk3zZh4rp0qb5rRUDT1ayjXaq7+XHDVuKpsxZvfa4M8Yzztt4X4j9fN1
vpafAE4nDJF07YE2FfIoa1PFC8brXO2vBaUf41pEt//HGkDWzN/YGb4WZXUQGefP
EvSClaa8k8McyUW+oq9lx0AszKcnf8EN4YYvjeHt+2lCfrTzTIakMXI+yZclcmzQ
4l8p2a4Jg/F8V2EqqyNoMZA+k7/bQZHq0sUiHYvNrU/Rd4O4EDkNcqIWvWt1p0LG
gDsnM/ko/eXFXCUvuh2aH0VLAoxigxlhWMrzUYmqvMap1R5GGEY1/TzJswrsawfa
r5pkg33+9D6b9q0i7ZgjzBTIvqkdIu7qi1YGHTmiT3Dh8sLuqhrCcK9V0WfK//Mm
O5lbMMGn4z1itkOEeH1OzDtVZT4a279wNoTs6b/ZAWTkt4ExOeb8Q090HR0RSeBv
xtJO01FJll8Xq4JLQsRVyXIj4fQCFXD1GUICgNTCiZgmp+uJMiTR7bXwGQOOzYwt
6lJ66GzCX2ndrqPSewQmnGh2sXPoVg1buaEx7dqUBTVfievBqUKKeyu4uPLYz0tU
xHBgPw6ip3ix3Iccq4EDm8k1i8yI9SbyIcuSg+hpliPKbAa99ETXMyiAQfIFrBxi
68AADoBEw+ueXhkCqx8Zue58KCcg5Ueh2KxX4lovmHL1oDuLxb1SqaO5gGXxwQI4
tOhGF3oqNeGkvkkuPs8O7erbbaH78RG7+o4HV8Vbp/MSlY5U+C4zvrexNr7X9hqq
IBC2a4b8Tw7IQnivl3ydD+djkDH/dngnfg6Nafpo4t9SioJVW/qKqqMa0ld4Mvb8
o/JdgkC8b6WbFIklalOI1hO5YI3DIUtaICg41RSlc+xQaSDITmPqhwW80DolTCxv
jDRy+VZ4Rbsb6bjuhBQQEJWF3+wHpBqqgZgYt4JC0yf1RWXx0Ox11VYUS1Wqm38H
ScHEbcoyrItlwIB4R/v8shKA3Oki/z2mqJqlMK+K1NFV3AkvEy6YOyGxZvOzvXdQ
AbGGriQuupPijavW5pDESNpevczAIYXIFB122NZEdwrfLMkCZfpvsx3haxiKt5Bz
rOMvAHjfHezGCiyR7Qo+Swq4Kjb4Et3DnG9A8HPclBO2B4hJF0hbnDSVjbg6pf6r
LgkyoHiGGS7C8zvMFw3D+ylJJOpiSc7t1GgwOnB/SiHS9GmzaAYmQ1gunD/RQN+E
B+LJ9f2MkmlPDzXGzsy+7wsqyLyKnmag8L82/tOgKSAdRsKHElQFDCmVqnxL1ECK
vEcZvFebDcnJOYbrT9QsRcv1mPzeKdJY6wpJ/SYvrH5L76BDyVirji+G+qHtSYJ2
es8SETB+RgwSDf7pUEjqfx5c22BSW6lT+4DCuDk71nW8AqgG4WxmkcL6Gi69Rg5c
SJP1zcAnaHgmv4vubVfkWDexSaJXQutga0hFTaYYggAHFph7rlD+yfiRIn9ixra6
SnFWMKpkvEaXBFg0wsMnobKtrzG+krh5v7EKj/1JrRu9d1e/Ew5c/mtrpJ9JCLYG
68eXx+xbU0D9JnMtHvfiLZIMzVKVF9LrKzxylbAMW6EHa2N19OLm6s38CrAqIiKo
pCTBq/iOnlIVdEJSLlWghGodfjRUzPzjWLhkotYhC1ykUxrRBTvkLBRHaQgrOWHQ
KzcrJSnC1JJeOejfxSz35sE0SmlQoTyE9xptj5Wue+liyJCzwoW0iuIGRlvbnK7M
BmeR9sFGdZNpdBI5dy2EzH148P3OrWipDuk5rFjHk5n0iNHTF2ctCNK98dB0bzhV
8ePagpdHe6sSz+lJnrPlnAqyklRuC6u/qtbbYmZVfHh79p+nFYPe31ehpqP5PQQI
73HV0teVasGntarfOXOBoU3tpz/xlirucMhsJ0IFBiJG/ZEAMNYK93Hixu1y16uz
A5LWdrXx3fhdxfc4zjPAMl06Wyw3u3au0Y/ZUED41AIpQIb9r9/LlTgtB7Y/FntF
XGD7/t3ViJwK48DaPNEsnmtkMerVfZmPoPb+0R+ZDXRepthxoPq8aWOZpihnd1k8
6tdBXJNXB/TDYiDU3YZzNhq/6whHLhwkw2iX5r2ZBnzXQ4NcKAWEdQ8CKYZtwBLm
Lkfs4um8C3bxDbULeQGgnhN1gtWFopvirIhhWQNtGq89RXGMuQBS+FpECTnwuomO
8Ol3EN+zGi5SJMNPqxEZ0VD89AdHvQAifvm12R1kw3xWYM+0679CB3yLMKXrcfMF
+/psE4LklYWGvgPwPyptTGYuvEIZ25cgYPjK1Ff89UiYtNg0pgFgg6NUsc5AD62W
nfetsClIz/ikDRZ1YKr285s/driJrdWLrqoXfGLzecD77Onk94KYij92/3v6GDoH
mnNZ2ILPoCSMMQ2YvB0IwmBllNbl6tHMZJpptLEKjvq7yxrgYz2B0xehtVMW9EDy
muOLSdQQzJfj5356YNNBvQ3gVKgCsZcGGopRVS5uDZP1+Bzgdq1WvakmLOKE3MM7
2qKwtJ7t4/UD3ZuhgQ3rEqO/xigXQpcv8CnT73WTNlQpqjG2FZwGyPImwIc2xBxD
zXCmJW3tMJjOTnvavywnrUPzxmBH9MXiH5W05vgSdgVV03Uo6SubMsK8B3WUh2W1
aEnHnUiEY27A5K1ASZUIG/NpAzE0ENKR/vvhiP74g/1gKSQ5LqSWjRV37df9TlN1
/eXHzotL55oKPdgvsgb5KUZT/meV4qZAPmboEjWaumEdlVOVBP3hPPGaphOQreoo
l/3AL/4jtE0pVM6r34LJ1/WXHq4SxhNJS5Zex8xhTiKt57FHEdaN8Q4yyDAPRTiU
HKlJ7lXWgZTyuVK98fMfeLWoqYo0DouGP6IPl6Hz3y5avR5g2psMPYX2Lc64A/XY
CujRA3aB9eP66AZNLSic3oKwmrqcXkJzsUb/dQNb15WbjCDsH8/Sjrv/7EqlYQOD
git20JNpR0T83KGbVyVgdIgYpvZWsbgkLkubMXH3pQNKl/2idXjMhwxDatWw9uIf
8FIo+Yq85i7QIDmzm6NfZfuC2ZTY3AWLsQ2igrokhdUkR0iBvpKLwJVBnIPS0lkO
+g3HhNANDexRLIijnVCLWcRd4KbxrrK6jMCs0aYkrhAX69iGjj/49B6PFoFdhCxC
FhK/TduvKvpOA1csSdy4drTYrIwYh97fcUn+Dh55BOY+evVOuTBaz0UnCCljNPvF
oU9k//sHZ3yeH+lEh7iswe93M9eBVp72P00NOnuoeWpW9PiZp+FKxKCrXfGiGt7R
2NvBY6IpLIwdf9unZT7Z6MibGX0hN9rAKtEGdziOBZ5iAtQkFP38ZsdPQJ+vENsJ
gkCIV4QT0I3LuWtpLzg2RALxzxC90IyfXMW/Y8RaqXMDHfOhb4Tv3R7rQGVKexZr
v+Poi4phVXUwK4lktwQ57czCy7b+LEZXeUd/g/rPD6cwjZReqfjWNusRWuPG7KDp
zIyrCHs+9DmCvmqDshzHkFD8JYFbbJkv451P5QxVx3MU+ivdcoNZ/V1Ha8fRuXbb
1LqIUp882+Mwm6wlffBQc7Mh6ZSpEryYoWaC9H/9/XoI8bAlAfX9ee5GZpPocS3M
I4rvEMLj8s2SDOiYIbVNkX0Pd062anoD7kwfbvMcwh6ejovp4EAX/ZTPv9OlvyCa
242d9IHSrjgWjzzS97PNR1wluqdaVNWUUe9y3O5np8J7t5OBue50UFrxE5BwfbG6
PP8pEpuJWmLyc9cr+fC0TlDMCeI0bSRtkzmFZSRgzBkcVHrrlgE2bf8NVZWk67n6
yeyfxDAcECpHlBTiM+o1dmYl2U1Q9oDY9BVZamxuAsiYtAZsA7NEfErkB9MiU7Zy
78K9xQ8EwI08KEVEICdk5Bs0m2NvqERNsZ5K79wYdiiCpGzvBY72c3vMPfj+aUuZ
8FAzXdu9qpc6y56RM9ZjqBfAO9s5vSlTeWQaqurlMkCUGF7eIv3Bownihz53EFxh
fG9dC/HKeGWfP6o+syExFiseW/tBjvBqoIYjZvjE/pYRXuiCjPCZr/8gw9Xb3yZc
Z0UMYuycu99otsxUxPxqvmTb9ytSe9SgHH286cw8IDFApe3FDfwIg8Ee6mvBo58v
rdkpT07D1HfcHPynZ50L9fhnhNYu4rmcHHplfLBO8ZbrfN1PIMu5boBRWyP5EJb6
mAi2RjX6PdtzKvRpLczCgee8O2pSEAkn08sR15OLFDPft4rrH4G2Li6VJ62Gxkry
xXhXfl1T1tlyyLKXc5yd8D50SFn/tVcS0pvoxpnijdCmhCPr7xYx6MCSQNEJ6nIZ
3gZgNVGrJC5ad2+3UkU29EU6XvDirykF6+077PLkt/KJXEjQer0Awv2TKKUYdXmF
o/yDDXtDxeQAvkUrSytNkTZbZtABZUwHgNWAcmJkM/MxUMKxmiy1dCDI/oa+bpKG
s1JTTbdVfQJOcAB56gyQxzKtxX3vSxmCwCo/cbCjCk4nPeisYwNxAZUDg9cj20zd
JFfMBamIkdAVuziZogQaEWIdtJqsQ+eTtn5vh5GHl20b63BTb+XwvLJhD+85myAT
4v9IXmsfUzQ5f3FlTuScWHojCPLGfUmVkz6TQby7NEcTdezVSsc5d6E8jS8TGl93
ZIhyKjo72u/Ua1nPOzkv5qMVWoEizI2R4XeliVK3R7Y+wEpXZc1TbcFDgRnYWaG6
0R7wiYGTYR3PDFQJV1dsWB1fMjw1yAKdQ/C3KVjdHynTfFsga25iGwF9rxKXGqh6
netdY1YXK5uvKbOTpTY2+9UjcT7Qq2bnnp0pqD4S2FDGd6HI7AfTrIV58/5orW53
y9x1eV7mkf71pcMsPvGeOIo5gHxrmS9gTnTL4xI2XtgLWmwCE2RluGgqapPVNDfV
Ij0RN0Q1HYIDrCVxBBjZnjo5qMIb5huo5kMimVymvGqpQZQ5IbMyNs4VGFZR07X5
jcih9M1ziQYuA/IIa1HPV5sp9Vy8ULcV3gqpc/kt1bQbP+shUOMnHin9SXLwdVNc
rc3RI4vtkYnYMo3ms71EvdDN5w/7IsLRtLLm+NEep/USKKaXiFQs8Khe0iuNGGpT
WGhDBoZ2vQ61Pd9T+q7KiuhxEvjAKWEaBehI18ozPSlL4WkPh72rqTsaESyu5cJj
slxRIZJgIQcrq9PmCF+5xClZXc+wE+MqAP3HitBw8/uRlXtfEL2pYlJGuwAoOW9G
1UbK/5zCKA4C8BL6Vhpif4h6H+6FjgtxPodbBzlBU3yLtgtGTUAHbdns9QgGX3La
+xsypqACkhFmM2Uhmij0dMygetVQ09g4odLMZAxsc75XemwWF9yJQYmrNEf7Ff4c
njLYXJSpMCaCMPTW9cJLXO25tNMDwi2qaE/3NKKv92g29HURftoWJTAbV3JLTOXN
vSVsDyQPxXGKT19B/SCFPGPUvLseMSY50d0OVCMUB8EtGPFrAk50Ya/dWPGJuiSe
Qez8pwrJGunD4rORsyNChuW2ayaB2M2ZLyBYubrk9Wam1+ok/cty31ho2irOzc79
Qjj7q3BE+7Z0JQu2iDOfJtul6Cij4FZpIpvgnPO8NJYQomolaG9wNoTvm6dDmDvI
SlM+tc5zaxQaKag9ZKpamiV6no+C0wPOf+8MrKYHGNdIHv2SkjjXF4ydO2SJF3dN
4ioAcqZMVvll0dY0hF/9WfRutEZVTilzdkkPB03xxmz3Su4dMyzDmT9WWe2RUy5U
qcln3kGYNT6K2p5zCNg5Nm5DDOEOuebTMRRQJyN18RCnD4/XEvnnbJ3GlbdWaYWw
UwDLqnWbnej1qdAw4/DKHLcyBfuAkPoLDnslrmMRUYH0qqBTMasj/bKxUrJ6Kd0G
OzEEa+d4Xtm2My9b3DK8NwhhaCyfzAcs3he4INRNlE7jLFc9ErXJc7qD3ZiCx/tW
KPdTxcrzc9PKLHrKa2w9q3/1FYXZYi2G8OFKKLz263iJxwoPsWtgb2nCDsgQnKna
Zi1jtK31yvMDyOaSdZaoowXBC2Xdb+c0vYMMd5GXowtJrSOzysEb/H2zVOe4E9e3
xBCXkVGT3nUB9beqR166/wPnlIe5pnvlmJn4YlTyqLzFOF066bpgEvorP70MPzOR
Z+CxFDAhtOSQQvLzKxgs6gRSUWPUXAgmx/1bXYqgXMvac1EU5aK3NDPcB02jYKjp
De+mLyytRFzOTEWIaty6pOj0AM+UnMRYVmvhbsCecjVxATQZl/SQSh2QrzkoS7RU
/z280WpziNFhRgI3VDdw+8kRIhtzVwvhN2knVkcqxPV9T/X9UN0gbfcsjqXHXPGv
k332wTU5gWtd54EREW5Gi2sndecltmIplMc+vbH0WL2zxkFdpZDP9CeXqssQT+51
k7YL3sHPugkaR/a6nNboGh/k4A6otkh9GDsLHdcq6/Ex+/sinXnjUxNRCSble05O
SU3RKp+LN9uH/BODyeOXt7fPBWmrKMz5y/oz1y238zwB2QxYO7x4dGZW322GOgYp
U1fn+B8iSWqimSLghnUuhefhkG20shDFPx6YvAxcHRBSo2JrK8QuOm1u+mTW+w2V
mEzMPGy6YbjhX2kUUSjPEexTt8Htz6yJw9VWOcY4S2AT/hQwKH3lM/dKy83eZflS
FXYSnWfCrgZyHjbfdu0QHSJXf4TLHh2FBqQuYSsCyFsBQ5U+V3Hy0zKUB6oazJRG
Zyz5UJDNZRK4+zT0V//kAT1Azan124ALsUkx0C8pU/JitFZMeytFLBA77fQbjH71
haf9eooA7U0PJfnHibQxzA2HZU4CJoUaOZmrHJ14eLP2yDY8rWwQV7q2lbGC40Ve
a9rxS0W3EoIl7ZfwmA5szyGn4TINcBv/5QLKHwz8oiSglfySZMozM9Wd28tYrd0E
z+LVFCfvj5xZtmCHBGHHF9XknqMCmSztACZMup3WDMogA29CEpupOk6N+JfTRxLN
jgNmeTxluVnSt5HgqHVgrgEhNcUXpBH47R6iC9Tkdj1XWkhFhwBA2Lg2CYKl4D7O
Ps72crPPp+Q1d5wtQzDtnXF4EsVZYG0TGhv2iErX9+5Xy+deuO4CcD1/+wFA6N4e
slbv+Xs7npNgYuLxxBsoz9dEZY2cRcMrvSUEWy6Q3krEzGn9dV7TU6LZWLp7ymM/
GL4ZxTeMgM7dzPgYEnHWLz/8lJCPiwN4Eq+aQWKsiNqQRxO/BzFmuaYKer7sadLr
elgVT3gTR5+DNU0vY0AbazdX7xqqwDwKPTiP5gU9ye+kWnE0djKIBf6j0uT7+OrP
dPVl56nGvBnFRJB+bDcDzfo6H9GqqVsENauuv3/rFaihyKvLXITPuIlyulZlngKb
2E8Hr0GVcMD42j23VM6f9k31ELwD0xv5pziiimYFf9IuN6hOiuqqpAUA79axLI8t
KZ+wPM/tyJJ5gQNMFG7BdkiGU0mMY4sz68V+EsBOffrkr0czXyldAgY2hspwl4jC
yesObWOF4VEDYddOqrxJXerkmUlhxrlODBLdgY5yAQvs3FDnZy/AMTMnW4aqZXcm
6Gq+JIPX2z3hM29pInDjR1v9fSOVLDXqSontmvHs2xUZvwxZI9otE2ODsv4yaqka
Qd5xiMvRRgrVm9KNK0n+sij3MGfE2G9CEO2mZr/AmzHyHsleT8IwC+jWSYcdRDbs
SHsXHvBo4mGNKltdssl8+W2ior1VHYXs3ZU9QEckBhtgaDUGn1IKLIrpE7qSWHuQ
cIZz6xAgmZmfN0DMx/BHMGRgLC5s0uSclJeThL62UhqVPwpo0qXhSST7m2LxiJhp
Tg5yMlXA0MOsBzKuDcJc0X2RhR/0yDKHS6FLUUX521Y7hW2nTqOnn1RjL+i7kF/Z
d4yerke7w9Bfmo30KGiPbfRbuaBGhIic4PWREP32rp+0VO70jeI1cnjd1KtPK2qV
D0uwmJ1mMrb2abDWhTQKAYpZ6eW0uzR4KGWVvRwf5LXuvguG7Qx4PG3nrAJWEj1q
7Rag/9vQL3ixmaduMTSbW76WsvmGH/1KdMX7qNipzN0ahFvcBO0kSJTPVxLYVcem
8+/l0VlpCPm/fl8w0Cy9PG2YMAeYk7ZSMFGJNHzVlEDfkBCulXpSwbgkBuNerWvt
F13lDshA2q8UAtQ6gu5+hB/HNNYDY5sdB4dJd2B7y1MA4/YhIsfE9B+l3rLDqiT2
MedxeWcgAfo7wyItI5xZ6lptkIxIVT1g5eSWlmDEyOH+6VsxZr9Sw7qyGL68wfOj
V3U7jtQ7g1NQHevbsGWCIKJs5eMx3pCrbXj6qxJeWw4AZdgzKW5o1EwuSsOm9mk2
dPQC1m6QoNkYIOn6g9EMsOM4UCkiGhrxnBNaByV2Hlo8kjuc05+45zZ6lPaYV6Tg
S7XH19tmZMVBqF3zv5IRMySFcFBtTsFwuwLCvkVV5+QaGtBOz6NUXx0We1Pc3luU
AzopaCwrYP76aqbPWCYc9a8QQ2WQiZpYO9lsATvIq3X/uj/AAHMbybTOcUzpSBC5
DfVxz4sS4dgLHNL4TSlqDOrWJ26yPDsDx6oSiW2dwOq6Nk6RRpCGZSxgVeccD5Nt
VR598u61a4y77A0DfWJGlhiaseKxZxAWiNA9gNUVDyJKKIecK6H4q+DGs5RCvHkk
Juupwnm8nohsL2cLqKBVOdaUFlu52QT7DGOUDOEBDfxMVsN5oQUCgzApjaWpRwIj
ILdmSJ6b8pAvPy137I1i8NfD9xo+phLfW/KRy5YMjkKv2TXmSkNhYXg67GDXP5ZV
HEaBrtD5qb3qK13fcTWjePzB/B4kd0/t8bUiqw0GY7jytZ7XUTVk5nmoUcb7O5lu
qu8vzQzZoptMcZpCthT5gb8lM5JMXXuzoEupIZnzzjlPhUJC24G1ejwhmXj6m4eJ
yGOWeNOaNYyRlJVGJ/nGf6L4OOfuspfpgiU78XBtQHbD8zwzg8+xA+5gM9fcxDMj
XdtTw2AUEtTg5SJUvQgxerwkAyc7MczR+ZUBVNNAokMtkNOguEaWb5gIRkINLVNQ
PWlwlCU+veSaFAXuYxcyUxvw4EMvgv15BJDAo8oIbp6T+EXPa1qIRYfEHRjqENyz
blcmAt3iQAORQM2yPebJ2KEUN2ptPy8IbBKktIkpsN0CLOI1b+80rW9FUJnm8Ohz
V/pdyj5+8KcA3cvyII3TX+gTvyWt8cje7sBFj2xLIUgqG1BvmIED55HCJQBTyEfB
ougX0kggf7tpXXRngvwAzeqUZI8JhHmc3pPyQniGbWTVMzrGZtuEUhu+ybCejc1V
kTdSwwXqcIoBeYFkw7bgXBDcZyeezkwsXffvP4cg7sVslhnMAcGD3e5gaLU2onys
BaQ/c3NyZL1CgJR1aUCcL5MPOpdGnGb1xECu5nJV1S4E4Cn0fqgvwAvecccvAgtf
tLPDle5Cv9ifI2l3z3utl2gzZTJ40LRFgtyfN9XacTYqW5BstdTlhYBzAfrhoBC0
j/xjP50W2vnIZRQwBtrFeAUbQmRrlM/7EeRZznglpFJheTN7mit4pH3bqZTGV9SE
pxbNYFyddQgD9wX1myknVIyb8UeI6+0mypo+N7AKiPCB5SvDvEBNW4vIlNcpM/0E
CDGUc/pq9Hr25ZaY0Ou/zLBiib1lej93BQ5PXXirngnGX0/kRwi8PpjnfxFYZbwS
TH30qNByu/OTcCMqeJ6QY/X5+CBHiFuGg/lU6hGD/FjBM5KVo7TQgNxlbVaotg6w
LUYIzoDjgXwTtmG0V2VgYpVIsF6GkKFWf5Dvg2ztZ2x+CYCrLAEEl1nJELusuEKq
Wgh/1x4MeepN/qNTZI6T85KpAoTycQJ5tQeEzgQhzrlMmmKfMKg5n6UMqsFARQnR
0vsJl/P0gMOR9c6AuGPzisETk99QSQLNBYKMT/H1ph4bHtOfoHoXIiR/WKsHkLec
4JFQ2LczhLG4+0GbmNZvVcQhARRX7E/2Bb5uSeNOoe8XuSMCdJSU+6SI81pL1sm3
vdv+o7Z1B81UlA2KxYN/aWVefIpi5HWgCT7+PbBz72gkgbLD7Ob0sH2+iLDmpB82
Xjb6L8kFyd7ee1y70nnchjdD08olkyCe6/1bC+5UrQuzJOtoUVBlt78bg+Ad4Npv
dBbriwZxrNtF+wl5+4zn5hxog7gjdC5fhUe5Lg4UtMcyCvC1HNikjpCIG68nR2JT
5LvZFPcDzkXIEsHw052YEQR/8V0XijmaU6SEUDM/ot+nfaYnzs9h+SuFIKMXk2IW
ijbDQbG9FLx9rJirGviGUQTYiJ4Jmwyrgshzb9IBv5py6M2T3C3qP/tRaMLeKmBX
n482nmXaqsDFR//HWis9JSL+a322A5l7XtzwS6GnzOt0Xivkeevaq8azp/3Q9rp0
orLdgAoXs3BfvgnGeK2dwGb0XKq10xGmXpEvKNvYKEL5/Qx5VCTP0n1AvSlTEqRy
J6xR+dRhJ3d31QMNltVVGjlDk09nvJZXFHpT7Gc+0TX6+nrDhKHV/URd+fEyhgK/
0rKFs8Qjl4sDwN3eX7oreeM9UN/6p75vstkemOhxjgC3IRR0OxV+9n8HaG8qawhu
VJdkt/JwjXAy70z010YQ2FAXK85j+jPs5smRe6l01xu4T4VA5CteIbwz3qLHyj17
3+ITCjejoU37lmDTpcI/KSi2D1tu9p8YgnZadUBHhYaT+rjs8LEvytiExoAWg3Ru
Z4mWqUBoYUUMkGJJBfyX3JJZ6yyK+kETXPtYFbb4kwfZ7ihnYVh9Qqu0lMTrvxYC
H7TUpNffMbwj384ohXputjIOs6M02xTojp70eJwGYSZjfKVzB6FNF9o1cCrf/FSn
DhdY6bjdMvCkgXTMrQItXcGN4n+PD/YKSd6duuVV/mCAE3mhh0JU0I2aWLMaPmzl
rhzim7a2ob40RAZnBI6yGicD9fv3q2o1NlHCg2rM4DIkwxwFiZQJP7/jnObUR4X0
DDUWafoLurbEz/52qc3fdIMF/OKA8KWD80rl/qGf6ERKQ4q6+Fl//AKNoHhXAEho
bGOshus+ImrfI6QuxY3uIdmW9uwL3/yka3ZevWQ+B49gfxq5pslDkEJcPcEadY7F
PXQLl01Az2bZoZQxblIzVr/gNE7+O/lB2ivhdNWPIkClXF+QpVkFDL4Mbipeg6v/
Exs/lzBVHoR2T3e2n1iXHtSfOwP/bZpzX73XEqpT1ewayJWXvrq+KPCdb8NZ5qeQ
LqAa7s/oNu/ko/teIlDqDDMHPezwK3CRyh//7YYJoGqnXHtaU1CxcR4L4W0Pvmv4
xF+MpltIRAon4NS/pMDpjvbZOwtH70A2F1iwv4Y+4MJYmyaUqb9t4mAYSnEErCqo
SWQQWbb2btqWcnECfQmuZKp4h55H2Szk/Y7Qo5wyNhEQ76v5L2QRHtVeAp5vgO6K
3L08xJSBCBZFu3CzkuRy0ALExLVpnUMw1wSHWA5zwj0abkfLMCh9UOtbTyk+xl4x
Iz+P7FWEuxa3/s7h61r+SCuV1+zsNiGiCmse9Y7WXEbZSXNnR4nVGahkcdxq97GN
HftvcFOYLhenxVKhHOvWo4pNk/pUxk1GMmgtsA3ZEyAzlZqxY68SR/apH6B6VPZc
oQ/Dwdc3j70Nw1jvRSWzWMoRLhNnQe9CG4aL4/S0ai7UNRS/SsfOIQF6cJ8vuGrK
iMojebNQQEpj76a2aqNd7//3EUL/rFmbNYQTsPngcfV44Tap12MOFyAFgvy39+RL
WbPQtlQ1+WAm0hq09SvBrGSFHYrJ2HaG/BFKRuTVVEZZ+XkySViinqFO1azCaayy
LAduc+/ABDuALhUywWjoYdyY+McXAiC3jWyf6DsaiZMf3KMiHLioG2qOdr6dZOva
OXLmxXRTKQHbSf9Yl+0NWe6SdqJFC3DdiRrbu4RyZfQhKoHxwajKqKza5UhaAwGE
FXJaz22U61oeo0QQSin2ecvbkZvjnXo5uUdIbozQ5NEBN8PvIb+13UlLxB/xDSjv
OMqrXGQYoVfQ5bE9D5cylU0EV8KOf1APk2n/YhwkfpfrZwIAdStgnE2vMlM3xFPq
ilQ2/lqSww4DQP6khjmNQYiz7+Y5KGh2lWlavyFgse7UOYMVm6caodnAewJpxmJO
5LBc6hJ9HHZBW5gzNuhfW0yPv86SktfTPcQcmUPpMqv2+75YXZmDb6s9R22UgYd8
das39Ck9MB2U/xE+KXGSUoq+8gN3LkUtUgBEY2/QY/VMcmB4XtMtDFsVTkVgGGtJ
jX00VFLhPJ30HCk6ib9/asXUsoBYtFl1UZk8DtHSd5MG8iFBojX+/fdIjZ46YPvf
6wtpdL+L8h0zlcL4Vt6Sg7D1EbjJnrZISULJTjZmGI5nVrmn3PUX6RwF5MgPx1Hp
E2YYwxKn126WW/flMNDLAG9NSL20qHG7JdWe+UCU8HaylaOnnXEx5ADT/ElIf6D/
4nhl8K2H0NvgRgJibwa6GTfnCKeTDXje+kIXaKz5X7VMvUCYsyF5Grm+apXKUGh3
n8REVMfTWd0c4bsgsbETJU7IWHm3xmRB2M0rvORTQb5KvV3q0UqOK19lDAmmXAZT
VpBez3bDkeLKErA5zCRI3lRASGK1tvqIqOOiyl0qrKcW4ixN+ghui4b+Q2MSLWj6
o+y4V2pbSAFf0GzNiD+T2Y/mA/XKvgM7ubGHi2o16T73pgCzfQcv7sBt1t/CX8hX
dhLWuyNWGjHtre+bMLeX7ycrdn7s/fD2auNkH4t7ETBQraz63V2CJxalup5DcJSm
69kjqtLkuB97dx2DsY7Va38d6h4QGlGgvUqf7UekLxp+cdW3Tr5nsO1wtbIo0a4h
DdhqPgGG2OhFHjJNWy0gJRv+GAZoByKf1rAVxi9mFeAVzXQdyxQu1ctva2TOGGey
Scgw9smFcMWhZS6KWFhCzkHjbzg/sBdraN0p3YuKP+0+RBjL3MS4iRjolgHuqTTt
iV1VDY6pc1yqQ6Ug/UDaBmI/YSysRczslBmGKTNnBZn2gGFtai54pJSbf6VFV04L
kAGlv7c47XEUTMqa3KoQoWhufd85lfdai3EkXKvMPgwH76aFw2vMCqguCuhJ8tgn
j7z9LSoSjKS9vgYa3pWYBHFTDGMleNO098SConF58B32u5EaGa0uIO1277329GFd
Lfx0dWBacW83UhXp2M6/gqAOWt6x2bOo1ONJCZWoochraqnFUY3x6gAKZPfKaP2S
EbQ78io7QztbOzeLI81zXaQmdDCZIo7A4J84Kh9os0dqe3cvP9xJ9Y4iA4RTNU0Q
cMb5yOcx4zVAS20ypHEAF2iC/2G97F8kBHdAXfu1xI4SK5u4v9AYs/y7ixOgOVbK
MSWtFjjDpfd0J6CNecX8wyR21hX266OQD/rJcubWr5YWM+eSaPcO13Xu6vwmPivb
fY+eMy0T9CQ62eUhkp4hKulAiib9gSkGHG3nftRv3nYpuIRVTYXeG+hly/XwTVvc
0v2/YtlEUSojNdZkiN/XY4BP2Wfx3MxOfohG50zARJtzjUbb0QJp0r10HZZIHN2s
MpFKBeLB8lNG75fSronAyP2EE/Af41kShjOr9VlVVD3EPhXscSXX1LchumgFwv26
ABJMHH0+LfEjVDMm2kLlsUA8KQ6Qh480Y9OIVUiWlZRJMu9P62M+n8cJtRc7S3Ia
JpQ1R8flMNOLiPaK1dalpJeesV2CsVzqLWBtkTC/My8huUK4R513XZ4GzmVnAdGB
Woi2DRj9iqieHP2pO7DxG8+Ips3doxr5fQVuJShwIgG4DIfvb3L/IxMfOOdr5X24
WpgDl5EzElQSI0FdPSZLSvRzciax+zKu0vE7N5xPPm2ZlA5mg9dW24iUD8AMbZ8l
EDTAQOfWIF8JAOc87/RqTv7ZnmFc2xx8o1sr8gXcgGTL58Gox4KsZLGMX+J8Erch
fEIY6G0UmVVYG1FixuCEOJV2rnhWSjEkoXO+IuscnmxdN8zHRkxW+FJ91oV92ECg
ULA+/ZnWmZjln1HYtvqKIt8PptMcFa+5xd5/PsWGEJ28fWywRYOPKVEsqYUHciWV
p1Wlh7dtfjIOMLclj64NnHKbRP60oivHmtKJMcguQiaxsQVCXTSTDW4TY/+9vcuW
pHZZHmXQx7LOBqP090AdHLCmqDfo+dH8tmWE29J2TrrP/C8afxmag45a44ERjr9s
ojRVvPI+n3HHuNJ4Hzr71Yf7L8nmpcP6JOZE1LBetjGdxhZFjgT8IILyGe6UVvmv
X2A68iJAlF2N53EsR0SzGcPbIuCNJtajPPKI8aNuO8Y5ghrA6UmZvhO+9DGxPPid
BFzXsGwAAcSjZ/Gwnq2Bkj3ZXmevpS9mFNIptoyVOe+R8sDK64/p+bq5ug/7hsYV
n2xSD7MEC6x8uIZPy4b5efnlM0NuE9dUe5HFk+6b+VRleSCKicmejZ3z+qQOHZfE
Z0z40zJivC93KXvuuAtrDfKJG1KB4vnyOWuNBvXkEojDmCevZW0ZcxP+m1gVCHKn
GYqIpi7krClN4oTiV7971uHvFpdypSQ6dWJbZAKAfa4lW8Ij2qvv6KYtd8P0Wp8m
2sj5TQvcDMbgtl0rEttN/7o4UJyiBCFO8QLfXbBNS6iAREUDBkh6QxikQL86zcl3
1G9NdajGYetlpYG87Jjsi2wrTL003//CpDYBLPnJNNL7VQ18mzgyo3THcOkd+qgd
z1UTudnZEz5ZEknmQ9ifD7p3CSwJzD05oUjQc1l+Zg1OL95vpPHqLGJZI6d9mhAj
Qx3AlN0yNA/GnIJ+X/1KUhbY9X8/pMiaPf6P2gN9VbZxL5Xi4Pl5RmAHTkfEb2RT
WCO2uu2f+z3z9ydh706r0uAQZILtQyYk+dCwfof+qFFP/Zp1atJNuboU0i6zY31Z
hAIIP9LTWwQn4vRoMTFWdUvGOLKi3OxAIMXQGaG07OxmcSEwx9GuaNLcwLKyoT+v
gUiqJ4nUa0GvGuvj/vp1tOlQoEzvFJYWs2MVBeR+jlPyu5T4HV4DjdrzGGXM6PN0
PwcgAJ5a7Q5MsjlIwWCuYp4OFDtytCqz2hZ8sPXu7fRvdo0PaTYgbwtYrqrEfSVT
E0jc8m2FhFXgtVHVRO+SKrlNUybtj6KRkOJSv/7Cnp5SSpWeCOVh2xtUxN9ksI3h
nELp3Nf1fU3jtP9bh3xnEsBbNlZbQ8JeAG7XLsx6QbK5MjuvTZQaGJusbOIxQ+W3
vPzkP43Mqpo8Hou4bjox4yvBwnvZmfNN8gJw8Olw2TmV/deGIAmMV+0Ia8xpMFG3
kq4oiDl5vlshtiVQOpv6txPrK4UoNTAUQZXzHoYNu7U7Gb7aqs9H9TKGHbpohKZ8
jgCGZj826BEGSOPhd6a7Vp27nCA4YMC2eEO/t554zqVwmUWcYP+gvGQLkYZqNAgf
opbRfVKej7HBr5sk+zMBPWPJTLB3Z1YB6cggPpyDK50eONtoF0KHuhDmCEyme5vK
cM8hBBHwC/shZTGxP/je7q/bJgHSvfW2dNUjCEBolrHpadznCv9VSPuE9rC15Axe
ozUR0VdDT3JAwaAoXsB+dZLAdrZMLt6QSomyd3slBzQmL7/Lt060gp3DgLONlg/5
TFtBDDw/MvFK2IiUmuErrtC1Io7INcXral5dukecp2N2NZU3f2rVyBJNN17pFDqt
5wVVhI/5+wARW6ba417DhFAbijTa058BYnr5GW2hUzV9CoBw3kP7fAlnSD4bb6Cc
CPE48QwTECr/hrd7OcdeK/5F4MTF+V3UrAHWDLnCqzAygyCCcp5DI4HXs00ZXAUD
0FpkXxj7WYSj78Ohj4UkHUr5uwWLhOdzkYjmdud0QRS2FRlj2wXYVTNmVoCRXIBs
9hmgyylsXIi3KDgbmQ4F8u5saklfVDWIXmCf/tIYkwIAnCFCwinzy/yRDp7BnapF
V9aFUFlraeDFNMzfOBjLLQ4c3Hinw7uZ+x/dLnOE0xI5vHANYcD6nwJyb1qMNqoq
ICNflXp43+vUlIab4omvn07+6igpS/WZQd8vAS5109bdRA8kawwF8KePvEJR7efm
dJsds87ao4/bI31pCdablhM7FZXwckU8GTqecUDATNPItGtQqiFns4IzwbofQCuO
N5KkjDqLD214Z1GsRQeK7ZL46C294eICRkpmVs9g8bneqZ/yo+YNCLxBmcOF98ue
4t409cE5onr/ztnLoNtcRNElfN3w0FOV+vzI1S9dkZgfPAJR2/wEPoD3MAC7+ImN
+hqgpAUFIoM4Aiy6GGsvgKjUShXe9U1v7zQ0VUUQvoOE+EY2hoe61BSemElmqYaw
gh7L7io/d2PVy4TvGmads3rQ3qrryJ1gp6ZbfPxSJnM5NC9IQFw8Ob3LjHjV+yZk
BgKtJgVX7MbRRW/q/79SYn+0Cz3hB8S8h5g7zFsA6unK3zo0mjz5nXuckJpx8osh
kbkTwOJ5SFKDFTeUBAXKgJrAxPNAVO+EDC8UzcKVBHLYEav6OSEB5Sv8TyhQ1w8C
6JXIAM2KWHLRNKqAftBCjI9qKGm638c2I5AqrbDmDLyC8fg0kmKN8RFxFci76jtJ
J2HKn4SJWGes7A9RzxLi3WrIczaQjBQWBKuIbpClWc5+YUt1/BNe4hDnpq5Ss8xB
fJ5Jcs0TRHruo13lvfpUv88gc4Gi+cGOBjBPYRErmQ68DAR0a1kVTDvOLxtUe5/f
QvmhPNnTtrJEnHMau8ok9DMXV1Qzjq8NmABDetxtXkvsK8Jftfp/eilzwarQz0YO
1/48zsgjP+GsyiP6aCNmdZ6fUBkaI2DWa5iZaZrQAZZOPdIEq8U8XFBRtNwVKajg
h6nXPl/xpHHgCD2ddNxpfBlS2juaRr+rD1PU1m1l4STVj0n0Pt5a9NfcPtwZvx1r
nbXeSMdSvJbCiKDLGrv5P3VWFbqF1x5bVjENB0FX8OQPdUswN3wuKN6/MhUbS+Oz
6gdH/BM/V+z8QMPY0jPosNA1d6wxlbgwL6qQKKHqt9Fg/XqSZyy/haiaoezjbroz
2V+WDrELcHc7j61FxA6OwSqoMPfQhN4/OntE1mljpyfJyUN07OipSDk9iB0uxkAs
DN+kwS2LXW2maPiGRzMUKitbyYqZ37tBpCxph3nyaXKip/O52sI2zg/3g12s5BAj
RuR38u0kPCPJRV3/LAYCaekK2Y1AzQfX4Oa3Vmn8ZTn5RH3s9tiLPC3PXKmDl5yl
xn7cwtjQxdyMNz4kWiIT82YCeDJurXdrgCCeK318HD6WBPJQSK200K/zCyoK6+Zi
RrBVtaBnYJmea5Yj1ZJ8D5YwnTJVIhOfkVvHbvsOA5deMWauBmKBtEkVYClkwcK5
la9EG2rE6sbh8+A0Mp5kiCVZd/tNjCH1pDtgxQH0Z+pdcUZGbCoA4pNbJFScD2/e
oqcRecPjVRqkWK3FJAbauDfOZn8vIW2Ak8+9B8xF1Xm+3xBKgS3tsvUzosnM+UQN
lu3THDrGohHAMjBSq520+XDtWx8923zY/LldrfE44ZCFjqOQSX+lyvFxHO4IEwmD
Wfae5QBqJQTjP9oLyQ+lit3bXJXKWLjVEW1rkbm7ayoAM13GQLgoDcyCRUGd8VBE
gqRRJBuMKNdFxtuw4BKg3NLZ5UwADBOU9BybaX/f/1xt0m0W7+VwAzSVAYwH96tE
vtyR2RwIgAuczIUU5smUKVRVk/qwU3NvTrfnU4q0371ZZffvLJqxovsDsBmjQ0XA
bJJkvYbS0OIxzsCcOPDw5iBjTMebuLwkYdTHxEa3leRc5W6rTuZfsu5o+KaBaAOJ
oMCJfJxE6rMh6iqEIdC/xbMGVq1R9sAkVABnDHh/5iVK2sk0DTaxFFJxUhrzMIck
tSA31M/oIHFBhc/zrTDlYPQFvOVlL+HKc0B4tfwX3ib/udpWbTYjwrAtdnBW5jFR
GHmMDRk8H8TfrGE4ID0S62gAWl6TiPMywfD9nuRHzG53RMCr3DfBdpul1pm5/kHU
RustkrXsSR6sCR0F2ciLII2AFkTS8cJM6LPd2jOjSNQJmcoLYTJR2z3QG48XKCFS
0+G9rVj+3KeLa8Z9rm9m8IlFDxj10Q+z2l8b97KaXFu45Yx/gnrfFxJDR7+sDlLN
1CWx4iLoO/kz2DQbGvGCOXehNfG2ztI4a7dZkYVPomCptE8DSea7kgg2trA8C2bj
fuEH79nTD98/B2zNG+3ZOYJXvNPgADZK8e9up7/z6fUDi7OLbDxZ7rJqPV+Ffdcl
eYV8RcVU4qNTxbWasEoMp/Fishqbcx/R8bP4RTAuXoMi/IJIfR0wv47ZPjFIwkHI
q6ghcfSc1F8bBNLqOM7UNrV4sS+yute9atmG+dBpStSo/GQg6keo9XC0K3fyHSoG
3ur2V0QdeE69FS1UJMEnaPZUVuay9Jso3EzRnC3mOKgWsIbm3B03XQ50irUD2B5w
5HRU0SxIgvrmP5U52Gk4fz97qVgPYfeNzbanDK7CUpC+eremqrpU7cwNsVXeBE7s
Jb1s7h4I9ub4Xo4lWPjJIsyNHv+dsmD5Zo5iIPzM8LnCw6rYQPIUA54yLdG/gcSM
Pqnw6UQfpquJfkIuWZnQ1zWzrDVXakcbDcqNMlXR9RBvkoUdeCmmLUWb0QQeMe1H
YyG9LfIUWmm3G9stQHlfgSc0gfyerIKwI3yldVH4DONAtd7JI69H22Tth1svqGuV
4KS7wbLM5uZob/LpkYXPdfoZZ+HP7QucT9f0XficbMYKr4FvsuVuAJRG5+57c97g
jHP2gVqcbsSafcJlR2RmMAo7tTc5pD4kVfN/hbRB1OlewhcnvWbh9s87CikF2Ebt
ronFFCK0z4MfLGfhUdOWsGYPMcHKepxeeL+u+RhEiLKAhg3ayPGXp1PfOX838viT
Lu/x2Dk50HOi6PMYFZmBOoEJ3ofSLSEco6EbPMC4RmnKJjEqaYn3g4yx7bvlfTjg
zAbO+OX/SszpGyKkTf3Or9HJwTujRR7PikS4zGofDHPXKi+KFiCx8ELCIScvCvXX
EdwMbSlQez/eXRavihv3vC9UhwKx+46raZ/ox5+0+snPLmN9azruZ4Nn0K3V7lgU
W+ovKZSfu7x/Axezx1OaYubL8dlmiEBTlLPBBVIApSuuNjbfrWpGqQLjgL2icNfv
x0i63fheXhV5OdgYEOaoU1zoFzlX9mslYd4sRQPoL10zFBByfCjHDkkATwfz2XT6
o7Xyq/am3ZzHG7XGNlhc7KeJf3pjAaoUsuVwMmlpOpAryo6kkyLFBGRFT9hs2ZFJ
NOpWPBaPQsvloKd+wr9Nl3jnj86KcI4v9bVZwGqMuk07G695D6/3446LtO02g9VJ
mLWQ2kUzxrIX0ka2aN0iIfq2c6PdFPibeLGRBX9LUGqaQK7OArt59hxfHymjgKDS
6Q1yQvZfdyI8OGf63rEOoVpGlu3eTzJT8+4oNZ90id2poMM8jj9oqUjzxO2O8OBw
t4Tm+Eq+rl7mmZ6O/HNwNsafM9SHINe/pmMroVCxTjrydOqRDYlh38Fb+4oteAKA
oKGLD0NETsMF3QT7E6t5U8Otbi0/JPztgJjjKGvZlL8PNW406+WWkSgTJIpDbicq
ES9ha+dobZU7+AsL4ASBIUKzLQChxGtoP3yYxd8YAoATCXMk7hFetFZEDkzjeX2S
4aEVmm3eWra8Uz2SWUsgeUL5RPyasXgRYuS9hU8060VZ9/Z9pgv4dH0uRdv8TaNJ
A73Hwv0LL6zVMXgbQCfvOxZ8JxBE0cUREo2SwUtvyHfL+6chxfZXp43kmmLg+gs7
vf7SMEFZTj7vMpN4SL/FuC8GzptApuPf/UIoBDcSNHtsO/f9VUMUCtjbAnnIBOyF
D4dm5wodAHoJmszgBWJyiMtmlrtNNME1i8JA/5dqprtvgy/l+PhT9ljSj4xmw/gD
lG8mnR4ubbPncdAFrne8XyclZUefZNGvuZ2CIxJ0OZLHHEdbNIyYwtbqywNH6Z7i
UHdHyRlP8AA/FPET7sK7SE0pYHJwHtRi3vMcgwQRJEA49AqUYBRdhN0IYoh3z8un
BSRp6p0kuoAxp6yL4jt7zU3EzjNMgEqmLNfVoOHOCBCYCs0fWrDfHdEpEG316vQE
aq5SapaxyIIvH+XbOmx4a533mn6ul17rAsZ1wBJgd35jsrgLPpzyVh8M/2dVr9Cb
7V25nYx70ycuu0oOzrgLb5ixkqumHOMTRV0r5OsDk3EZITiIsgBZ7wDxuBO1z0Kl
Iayr3Gxj8laknoECTgiZhynz5kQazglQ5RnLReIhY2ASfqdcOxxULKbz6GLvl65o
wvmDMWwJ79PPJa8ZN6SDZ8hIfKa2Fu5EWPDOMVltrL2b54swSXdE16hTb5gXeAfi
hcmpnGxMjix2FtY5gFjO/d3ZtmQiozjtDVuBtpOmF6qLjpaKPYLbE6sxqfdAjHax
9x4pqGKfOrTr9Dso+0uwip7hLjqq2+yv70dykqlR5BtHamQQnuGUGDKpY1jsrdRq
0utb5fvYkV8gcLAJ6roKXqJ0P0uV5hURgsjKRMNxJDHyW/FekCGcoaefBoZOmh32
L90f8U+OrQbSBe0y8CmR7Ce5qsJ3tKSOnaBfdKFBjTOvQAH/9KiGXoIoJJklN7ym
r2hVunRiwwiTl4qLiTk57qCxHFHMe8rEhTnyBqCc1BY9lwvDE0IDTcCW8r6lbIvQ
otsAeLSXHdOhtKESIc1NUQBwYPdEJbG77C0+7JcFgbUxqdrvdT3Szc9bowWisfTV
3oTM1XinUeD+ubnuEgZsH5itJ+CxUemqZvhAyJrIUvQp6/QFbMM/X7IZZfzxKFw8
v679FlfcmAkaOi9684G4/9dX1lVpcOLFXG3bQICtBigfIIWCyw2KyzwOH2ydXEzi
3BCg8dWxJgBy6qjc63d/yIZbH+wpwvkGHw4Vf9FS2wUb2+SXfD4Lc/5Kk64quCTV
HmSsDCPVd/ZluS7dHjroaxkDRDK1gaT2qcWtGwXOtaSgXab64D2ZCIjUuSP7ld/4
ScPXWBbNWL1X1EPmaVI4o1+Ok31y45CqxO6DGA5fzQe4e0E4wzIClEe6FZ39DRai
F27ULTL0Ajtdgqh+rPMiJQmg/Ey5jRZMlBh5S+YTuwnjimG4PCfMVAZjPclPYhhx
EjHKTX3uF7S075XWF3SLL1NWBj89ff/EpzuuZxb0K+RlsuOmNJSY8ufl98j7uNu0
lYIwAdYO/oESWysuPT8PpvnOE9yBnyKZ8bCmeCIiriC2dXKBuDZxeD2dJDc6Z/CJ
CI1ONvlYeRsEyto8VqGmMloa64OSVQ/b/iGeVBI6COBnovE//2iPsCzGJ/OlpL6s
kxXMBZbFc/yrIHe3g/F+D1RrGqYcmoYD6xcs3fqu/x6lAI3BMzQPVhlLHpesqXER
5tYRwVpwujwgMhFY8D4rA4DdPCOpez0gheRJXw8uUnNTiJ7hOo/AUS/thCnaL9zs
efRAIiIZsovzl1xFbkTDzD692scLPbFnVgATFTY2jzDXRdhN1YiaB3HQps9yjuI8
ryUFLManzaES4KXMdY+OYfNrlM8veYA+VwizpJrewTnn9iyr0Dc5HZr97Y7Y5cG9
3iDCzf533k2bMTImSEaMd9zg66+UCPGmmqab2ynUKiyVG3KhLldosGZ3S+b8eNiZ
FqAfdQzs3DfQIsbhygT+OJuothicb/1MEBG+gNjhiDaxxBVnVv6OZ6zpSOIvutAz
L/8xGW281P/OxaVsBZDilqtIpQFLrDEnMAZgW7qkh4rTikJ+JVozpu13WT082Puf
GJRd5Ox9juRwDWk4nRkL4Bp6+8E8kyd9eLuVVgm7llaA2ds1pGsvXnCZkXQl0tvz
bPPhDkOphTiMJOa7+jk5BcVYl65uBw9iK4fSReFkmzMzezju/coe9fl8aYuFQE0o
0pFJs06hvLCS2GpfDmY/PtOSNQZC01IdPvhltS8nyvcTvf//RD2G97I2pfrIZZZ2
QvoQUNqtg1FH2KGOCiGraAyQt/mXEx/SitCsJTiNVwY5zQFikK1Z6eX6ImISQMck
06lFKgmC4trS8SLKTYSGu3c8AR7NWm4cUnlS4YmgV3izsGnMI5j/CTfTZn3DxYwk
1OMS3w6/fkXysKcGIIwlaWpv4t6GjuRRNDraaiwYq0Sj+6BGVrMES+rUXUw2inIY
mmAzBfHiuj+cjWuun+/P3TPBkg8r06BjblBCc9VISylS7xPv4+BtDip3Y39yRvk4
2tIjafpHrJk0OJvpq41vi4+3iWA/OV3+aSfCXHQZnMIa5b6Ykhuh0s9KE0Wbi/WB
5fYsM7+a1FA0KN0qPTEqHDmt2UUIW5fNnOFACa0VL9OHZj6fyWukDVkpJ/UGu9/2
L81kVwllHZJVJ5AAFDjxXdcJii0npclxFwwsvYm+TCEwBkHdeuVdliOVAAZc47Ob
iHnUS4FBcMGrb8e734AezueNTWElPmbwkcR//7qLkjXLe3tY3IWZ1Hwe035C3JGa
h8G4ipL+7JVdZbZzVywvJXK7/ho/Is96qwikvXye67Xx71+4qZ12OhuO7vsCyQYg
rOWbIxT0IUR9vTERBLRIDfN22YNTZBLmMDHXpkSjyrWlPsTMsOOMkIGmBYowRpvu
uFE9ZxH++Z74Qvse7kop9X8K1DsAAmhBjfXCce8bX68xly5orpJiczjEgwoQBfs2
obvfisYQ8SIqEdjeuF6cs4ihmtmoyjv7QVkFA6GHqfhaPUizlEgCa0DPgfhVkyM7
cOndXoTETEP0yMPZ4xSA55P3pMtICBknHa77DG8z/0XenRTLvF5sjSaYr6u4wnX/
LPFZX6NN1ydUUHWoPga3J7HeC/5iQJep/ANjERt3/5qLgshzi4oEWlVO1Dfwtwqb
YYMYznX0oeIl1yTeu3lnhf1ZhPW0z3kFGrpWId7uHJR5TZaJW1+KcckOQmlTyaET
993yxWo8Neip/X++ZqV3JCMTiEdM7dx2mjg11ES5IyRz/omTLmNw5qlD4ejVZKny
8Mfzpg3zpgn6r+5fYPUbLAUrFQtPWUPGjI+5JBP5Qy6r+5ENRtajGwWoaTKDN8mY
0MVfgwSC5hGCfDJChVDepJjcZg9P7CirXc7UzTvViF4VNDA24GMAvnIrU0aoS21r
1t5SGry/GHh19jDlg/Nn5zyNrrRjIyVdbr4tT4q1/DswsREyNv6sgaa28xitxLmW
gRJypb+ly5LhXEynIxr8LPmB9iNgQydt0vv4EWlWCOiPyGBn4j6IWub222FeLEPg
wlWqjnUuRwqGSlZBzkQlmZJ8ACNc+0mJB3snKc6iwaFSoMHGsgiRFLHLjJFC3YDQ
vFoupYdL4bMEzmX8TyyE8pICcDaKLCTvXAi5Sv0YIaKSf09MMGSI92lTWrZ6FocO
jZ04fqlk2N8VOhDZyhVJUtzlYLj9d3WbA3dJc6e3vr47cHKNQEWcjSbOWRilgRYW
MiZZQUxCYsCh3gcsUb8N7wL3XA/bs6bLzom9odEbA+znoVfx8qTOGtLi+ro92/gd
jYePhKTF35gc3vmuNLHbDv8lql0HyELVfwQBw8qTvCUlfASa8k/QA+EwV7/b50kf
+pPb2P8qGmaJ4GmW/PDKYqBb/uX9C+jT4KWtIs7ykQhu5//IThf31MKd2Xqv+EGe
3XagttRs+YZAQ32XOhO86v0McnU34B6jrIU3W2JAJyjC3iEnS6SM3mLezmeFnQT7
l9s1hr0K15C2wY5hEbp3WrHI34SE09C0KjMy5BSjInIEQfGuUJgzOU1jylxlFPpL
gTmqfOubSG5cgwTVoDpOuJmY+Jl2KVKgZA1YnYxSR9e490lYL/wQZXNeCfnCgWCE
5Ozrv6wnLzz7PIjrCtB0uNbfhJ+D/tKegdegLetsUUYkO+6cym60+sej1ykGsbBd
ebId5n4GJCeVo7z4vvYVfVl9tINx7PAaQ3s6S1bBZGTpCUQjJ5xhIPGfFILC6aOs
2XcM4Oi2XOS88XRdY0zEZbiuQdeGveqThe1rNpp9hweTCLRugjGaXhqGnCk0eYbc
mW+b2FPPD0hvbKtSlT6N9kWvZQtuTulPZiPfY/OdBYu+Qj1/T/OEaDj21DV1HrQa
xSPXlyX9hDcev/y6jb7GKLCCTq/bHVlV2AJ8URxvb7q7qIoREeyX0D3m/rry1EKU
OoytUZKuRDzelihbauW9oUy9JcryQiVUj8nYdsYGa694GC4cAjHLPhr9O+LaVXxS
v1ixnI08ZNCYpbGxYTBabRqB3YCh1KPRmDh1wCauOoTU1k7PXM7dTamlEDYkkrb6
rEbhGhj/RgbpVincGdo8tR5D4qDvTjYFQRy4PpJymts/yumScow6O8EGB5Xpnxdc
THmXiINMp5+CXsUZwRsitv+NTVTE1kEtU3gQus0SgbK4g0mA6THoBZBTYHnQGZrw
CrQdG2XLg8WZACZDGOFLQ6Zdt3+7KvTKqXVlz1WKgpT0WF5YVAgQqpIibFY8Zeh7
pZTNA+fZPaYIzUCDuQxY7t/vow58K2WUA4SF1YeK1urxZlw46dBSLQ+Mc7V9ia2P
A02BZiyBL9+X8XbYQ1wVQc8rGbHV1HPxEg0TTbIY08KaKAqvCaobRecFKCNXE5ah
8xglsWsFtmb9OEt5VpkpTbKkZ6K9EmArJVrt5EilTivxSXLu008xJncmTS7gad5r
l1DiGw+nZ2IAHIeGmyMY3hO0FMrcVYz2LU6Ak+sRC6MlMU8B3nBN5GbvjoIZoayI
wzUEJDb0NDj2Grg2Z1wkyBoAi+Whjyo1yDAr5V4CZb8F34tLexynOvKSue+zoT72
dXtFF7gDvbOtVGw0Nv1pNx2BC6i+dZkQXTCSV9km+nA8eG1P+hTSGdVuaYr+Er/y
qqg7akL0qkAYPcTMCrRzON3Fv+ZdFKiVCDsP9P+MymZft8muW8ER7sn7o6D01uZA
4I+R9dgKRkNpPzkCJIA6mld6sEd0U/jpOFVbbUXXf0Ey5dx/gRSi6RFo8+2e35Dv
StjP7vWkxU80HV5PF7coVtxPJuNEZLh2Mz0Ofk/F2lgoPvZCVgFeyf0K30s5X1sS
/GE6JhcqgQMMHhdIl2CAbZTV+egmzPeTXP/9cW7CVbfEYX7i82hytAjsb4WlT2p4
Muz/cf3OvtcOrQsw+UfOlqODbJL7XSZOH61nqDL+Mn1VZhCz9NkQfhfJ1xbgcLWN
PP9pW+R9BE+grExlN6k7F+dB2Kzlt0xgD2hJexGkSb4XAQJbUcTRg67ePOLjAjeS
KRayXpuaZfN2fx8Nt1WRTZG5YeDGw/lTyCPiqRk2JgeYHEXXVnXmnTwiuePMJabD
U4ba7Qs5PBzWj/CbxIQczP+hgHGJoBHIueRNsLRP0yPciHvI9pCBqLAO4Y/5C2PN
FguiIUAMU2rgoGGp62wfmENrX+HH2wO6ZT8zdm6mVWHWSj1be4ndjCRtwA8QpZhe
makbOUNMRePqnJnmDbYflCu3TXkmKgp6J/eMbEaKkLHP0GhzdWoHAiPRoXRuqnFR
amt9xkPIbpu1BI0BP28yH2+c+x/jye7RZdehxpoknPuOeNe7V6vkiKH9WIgDlZCk
1reaZ6WOJaiuj5Hq+KZrCD7Au5xDlk3ABLDX5kfXF3MXXqdoRFGY1YKGK+g4dlA0
+r7/a5W+0mNSGOUxpCDlGkkbf7Bg+1Pozf3v5+RZnlqQI8Gbq4Vqq0/kgDDrTSbl
PVYPAHKf+xc/DSHFNuVnqVvUcnLnWqLqT2mSexYZtAOg9tAOj5QIo2cnzKGV0I5N
hbxJajYe9vtIVEv9inXvMwqch2T3x9pDRQxPnqDXL9A3WUJqZlolX+lkRy5H1/Hl
+FEBUVChbztRCpuNKmQHVH9oNVKzZWO4svDAHKl8mmS/o60yMXx+bzDi0xTgDNY9
PuA9iI14XKL0QxTjB/gg5lHqbC74vpyYEZQSIXpLStK/iQeCc1DBF9ymOjz6hugZ
gj5js2Jy+OASxPnVbQluSWzXwQa6cqY5ZWVijwMmCXSZ/fmI2xOLlpuemzN4Oq0S
3fP61m4fqjRs+87Zu7W4g1HnoaRNjwW3hbV15SP5oxoQZqBcIN+zT2OG9lvjiPif
5Iz6phniprWfdY+sa1EhH+y/erUqRGLDIHppnADJ9Wu3KLhIXyHVuzN2silWT0AF
E9M8UXycNqQXAuVZCNmY2z1oV6Q0d35wQg9/Ol7VfJFJsIWrUqFv/2wFx3NqRy5A
yP1VG99s//uw3QAzFnFWulMC0htB0x8epjAFvBN5YULMF+BNzKPLDXJJ63k3DycG
ek2EfYsBkAk8oCQZ6EAhqUsxomk397tHbzYQrTSuSTQWFaQT22/gabG6Jit52LM/
+SAMJ9zxEvdRdaK9cynfLJk3dHxfMZdN5oATkQcz1aopWcL2dHOkgvohZ6RRz8Ds
+NKSdtAp99+IVsSty4McsGwGz5OoRTJ2CJ6mio8yO7HZPxcp7UYUwnSnhM0JWy9P
vOoaa6xxgE0y/TZlYtQEr/LAwdZeOId1LT+8ZDWeaTDYjeVcx2VAnCB+cgRBsJWh
ddhNAujin1Utp4CZBtQJ5iXnxhx+qpePTlcQzXgMFhPJ3yM/lsX4xz4/T2GYerZb
7cpJbkhyEaV2gD2Y276D6Mk7jBKv07OpA0Rb0LXxhbN2s5oDPbtQqA/XyD5RnKL0
LKI4QFkNz3JnrxCJ8FXhCXSWKJF9QmNlIx2DCgEnl9VtYfj5OrrmEhK8EhGcdIXj
fwmBYVmnmyhDzboBaDGZRW9WBUwUuKFN7NyvxYopr982kj79xFDxLCeqpUS/tyZN
D2mICuT5ivJkZYnayTKWfAxb0CCnBeaIWdzMPQzNqo46p1mi96lOT0jeGtgt9RST
GlrQ4OzxTyiiRLvVRn4Az8NemOUyZel/vFKfW8szMOpmya8sgKdAgBB9ZOhn6cb3
4JH4/VnpzNYE6DolK7LYbauQSZuCybKZ29becbCzV808O51WFpwBDtYU5hvJMwd8
E9wTCgQh4NqXEZf68i26Y0drFSOVxWtlNRWgfTCGTk1BUUEhLnZuwsyHG+aUc3mn
PyrztI6TCxoh7mKI6auG9A0JsgFip/TuM0kUmGW8X8K7zOwHlBfT0mjRVWhIqhog
PZcvisoM+jMqjsNnxZ/p4HoKE+HfSTOwEsZAc4bbXkEc5+Qnsg5+wLn+lSoyiAkq
5C3Esxuo3uSzjVoCJCuOMq+WE+Nc+hZ3PX9hjdy/nByVtKaKcvTRTZZP/yJ/y+Pm
RmX3nYRFR5dvE1V3NoZw62jGPN5elR2bUkcluiNgLOza3+6mcyMPMVkY6Uf9Ko9y
euNfh46forNZ3jdMkx7JgDYsQMv2T84LB8lDOc8hxpKQtN3fCuNu9HkjFjowd2LR
MUhDcjURZX4ZtjnltwpFIKZAzdCV00THIfIzlOaVSijH6fxuNWe5W8xpnkraX1pZ
vFbWuB8yag1RZpsoQU/7HLj3qicTM0UnFRfFUhKlM1Xmw3oc6okIKW2z6kfuW76x
ADANJoENVRu2UZ9zAB8gqG9MmcZPHfhaIfkZBQg7+ZRBTlZMnc4XkpXViB+N5NPi
5RhPMOxbzjnJipAgBTcuT1sK+GdwbiY6TzgBtnmMAzm7h7+1SEinA9Yd8SX0Cr+M
SSldpiC4lTfXm2aLHSyZfJ03SCA1CWocnsl4hW+ZgiacagN5TdI5/mEdQb579/pd
zJxAUGVQY6Cz4egWBMaEkPjw+8JwYkdRqHFrVWLJbKvZ3lY/5qldzeTnvquz0wQy
oLp6Oq+WFtyvH4bOYrO6utqLyc/LiQTx38cXjliLsxv3UCIsZ9lwUwNlZE831TbK
/S6Aqqm/ED+78bB+v6WfpxrwFyMuCsYBo2BTsaBOHrRTmK/XQC0hMeSo5qqigBcQ
AcNF/J+4S4KT5qRPEF54ssPj55lqA9j0VwLMF9dv+ub5RANTKblENEdP+tjizNzy
ibAv+1iJBavf40BTjafuRostgYY+VekBoLdXb90+pomG60ioIcM8IVUkxbrc3eQc
nVOKtNrW5pMuhsUhXT8RpG9k4Qxv459+T1i5g72rO6daYHlf4eJRJpPAmKK8YiuE
NLWdCg/1D5eyoRn7xgovQ39IyRQrmnHfqpRNAM8UsA67u+YpX4c3g1fu6qM3qV1A
C4v3go7kva0k1LJKWq3eEjRBrGgigeE4bKJhiThgvFxx7R/gDdCboZs4zphUHjAB
PFsP5wRw2omCpimhcjJXGZNGnP6litfVgvOsIdNV16NV4OdJpBeLtlIsUFC1lJ2M
hxkuCxr/BXRVnF6Nm3mfRoEoKuyOgWz9DSVzqjrYwNs4xemQiNo/N0RHm5O4DSrF
7l2BqgGdnphyRp8RPk1ok9ULLpHY9HhyUdCmdsTcxd8Gy2MhrPh4tLnkIKuz4IMS
6U7b02P9toEGlJ6l3JXzU0j+bz00WM7I6ZsRG8g/2Y2CHUvOvcMUxmMHNbB4Tbjd
ipf1OFMDgoU44XFnvkeJnj9lgeEOrSPtCAYEcP7wQ29cLc65x0t3cIA2cxW2ubIm
IKV5Doq8b20IoUCgXQGUYXuwzUII634v03vkyjzqImORk+TCQmm6hsRDMQ/cWs1s
SXvJ3rbhYu25IfDsMoOue6N/TBRvK+IXvyY7c4uNdZFgAqdBP2+oU1MbmsNUpYBb
3MaNYMW8+wmQR8cvR8in0vYDnhu4GoNw1II5+2nDN+qc+m+rzsJYWQoPdX3U+iTf
uQLgb+c9nb0dt+SY0Yl3T5uj0UhLF1cF5lrAIlssOqIbTlyMQxOmlKPtffcqHwaj
oY41tdiuHOfclL9XYjs2UfUwXPU0llNvey59KYkGbLxa4/d+oGzpNFJLbucqeObN
lBgVOIwydYogDH/eVAFJAZqpi76io1Ds5BRYEunlMWbxCDiCohwNRCunGCaeHsD5
GKNyeD6wWPIkehzabjF1+IyJB5DGv+KFoo33U04HtOjP4fepMyTAPzEEYhf+DQyb
kgsqJfLW5qXejSTrsHSPZhjdZEPqLyP3R8ldr7aFpxPWlUQ+if6Q2JTHlrkVjdd8
64shCKhJAueaeNwRemhL83rrqFJKch+ErHwhQPphxVF1k1ChdxKW0p2tmYhBrgqu
oiZC/EPHwXd4RDuslDKIUZ7X6SNsvoFZaoNxHr4COMbiS6kjxmBS9H+1kuCNeJsS
gNJ6JfaQbhu+M0C7acdRx0jTlDeB5avCB5K73POeVQvPf/fBDT93DI0ciL38c4Aj
NsUtr9n57rvp/frKuaWJQ6ME3WU8jUcvImBiRJdG71pU8H0nUPsupg0eoV0IemmT
8gusg1nYiAiMOkyIiJ9APtA0ps1XgQN6MJHIfWzA5FKNoSpbnAhuSEtG/ae+ihzc
E/eoiwA3JbNEoVD6W0r/80frPjMajn7ubZNH2/qyJOozRjPIVi5fk8BDNIfh0AKI
ryT8hQY7No3YnhwvHcg7M+yBNBm6KaDKsawxTVBFGB/7jCDxAjew0pF+lu5FAaq0
tVvq/wcpTqwr3aIlbnp2BLrzYDDxbmbeB8E5vrYU3RtdkYMpK+sYjq6pX/zhaJt4
ZLOCs4UBWCC4Adagt2t45GcL3A+vT0lb9opCAa1gGEYj0p7+Z+SsELcNwvw+f/X1
TVzPcFGB6iRrDK8MNlwJS2Yq7RBMiouaoTyynDn5qNdpawMwK5VHvk7jNf37n3+D
MjpoLVAV2NoyAa9Z4NzBoFvR2gXlHkJ0mEk6jPtv+n6PCWfI1YcAeQdmioSApkie
34+2i+0Mwoll54+IHdsw2iDcptbid5eLF615qT+6rOUJ/s9adOkjTqI+56JR8hE4
DBUdNoK42QjYx/NQQX1FLYMgyohHn7VlMIVZ9qVVQD2Ll16UxPCLtNeaHKuwFA1O
Pgev9vnHELiQdxtd8aHohqB+goiKOxyYikSNNYXKftkDpJbOWSBQWR+ZXyjK4BLI
N/xYO0AV+r/xmFSzRpvtL0hlrIqdt3MROHi763kGT+ZsLkgX2/scaNOpsJ8Xw6Gg
7UyEi7sSyMx6iVEi5e2AqxX5dEcsLXjYQKd0buclGr1YFLvFUOVJ3D+Myrf+Dz4N
g7yGFr+Sk0pPa4eNJ16yWVP0Z2VrEe5j+TZ73Hmcmq44EUA62WjX+2odKnn3UU8H
BZz3Aq7ZpIqpgl0AxyC7Gqn6vQ2cWkh3VXhobdssJ4LB9XEsE0xWFe0LaYsVfSrI
lyUXiN3z0FVgGCUPA6iD5k+loHaAPMCxpAfXm1ekFiVpkwukdPJCInofJWMXQ3QK
/3UU5Xl3tCsaxfFkSN1kP3ZE/4B7ZdnGS91Jsm6q80g5ZDbR/AMQkhu/A7P6ijcW
NRYm8N0mrIGlUVDH7sZT69nZlrXiDNAKRAFVqrmr2MwM2yO/tofctr/8Wf2HKd/m
DdomhRDMlDYDyT1vp+94vm1Ivb2swujDxjNlx6tNhSu4kf+QLeaqpKB0ysthlvxY
D9/lMXQnGYsuae9++uP2xFIJnuafGsUddJhNZkyKktcI96Lo7AhltLzD1INf4EBq
pac9NxFVKpOpZ5fUfxT4CzCWN6NfRupXizEsweTd52I/tMXFFOKg56k6TfBd3PlV
BmOGWOgeEm0JzaLGVlOlcca4uLGAVNVxx+7jUHfZvGSzs0YozD6oNSLLivnPFLSz
91sGfsXq2azXw2a9Ad+WMB1C7UFpaBBGsrfcoRAiSCc2j33IPQtLTzgsBdSfPw2q
GVevmkexhD3Kkeo5hso0Ep77kGeENUhK97PxLFe6KDcX32lojOAMTZl3AsGsAylE
+lZ6Zp5CefppYeRM7fky55mH7qSi/2YuZPJT0F6euFa4QicMHW8wA7Z5PQF9GtyM
ERCoAoOBXbFSkDu/VA29ZDIO1wE+jP/cCTskuznwqUQ8PnlJixZ6ny3ijea55sej
X2KuOA6CdJzkEvv41LooR+qM0yb+OSVGvOmOF0npxcfoEDZFRlf6a3c9EoifH04H
WYme1/+9S2Da6GYGdFhgMpSbF4vXrQ8uJMz608Wyg5V5tf1kgyuipjw45BLMcxmm
LZi+Z/2BWuO8X+6nCOrJ4xjY1tg2uBa24s7Edxop5xgNawHCULi9znDY89S+xXfi
8PvvXoVywd0f+uMaPdCKYpNcflx8LFSHiHYAKOMSUwoDlw/SeQxG+69gPGbk0oNc
A205LIP1q6Jfnnmn94SiX+PAa9lzlygJEBP4L+fkbi+tzOBif6K+QPypfWYR9qUN
BeJqGndt9SKymIF8uu3m6xrFZh5tYOoIpNKk1XFWcqnvHvu48zGBKHRA4v95nDmn
0yA7KKDvgib9ayXqv/KRbvsLw8f137ha0JbZlJ2wbgND+CBsI9KiBPn6oveOrIEG
q8V45QqWD3KiSVnwbVXz+PB24udDGXHPyryUDcNshB92+r+llrrb4f3Cg/Tbix0J
av/VGoWtML3j1n2DuGGJGhhB5i+W/tMDgATw5dX1wL42xJleLqj6qXOwKMltMCUC
JE85hFSN+sfyEbgR/pOwbdhFbc3DKUQGoh0KTmN2zuAbYe+TTUqESu9Y+KFgHglI
uW/pcART4g9GCzSmA3fNV0tNG8iQJW1D9bC3k6xN1SbUPVy4mo0WpeSUM49/qxTs
UzhQpcREsC7EcajAWZNihifUMZC+7u7CbprZUqF1mjIoXL3Ijw5xHLkODvnuyqal
CtW8pVDQfNLUzuOTYxO1hG1vXuzk50/NUwfVb/z6ZuyMrqh7foMnvNKaS+WnyCyM
YdPAoqbxbLc4oXmRenKsWaeMKZRy8fZIX/umGLTYA2Naoy0K/R3jtf4d2GTj+PD+
KxnWPxhUl33JbLoHRwhjFnzicrixfQe/Arwjf/jok2XDTAnQot/kb99HLIrjos62
dM8U7Gj2FoyRkQ0+sQ9RtYaYJSfmUVs0GKaNdbhYD6IwMnPcMHy5/uIn4sLstxwl
H1C7Xfh+8bqrm+pb3KH4lFda5WIoy7qNbEf9aRaMaVzYNJBxOS72qRbYXhuVcoZV
Z5v54jlx8wffwwZk0C0FC7pikHB8Vz2FsqP0xlmCWd7O/6B3EXcENHu9t4qXZ9wz
t2k2fw7lIBj9YB/Z+PNIuo4EFExmKlV+5Gb1Tz4ERL+fYPNppW2+8ZlLvzQngKq6
kb3+kXdi+w9eeCQ8SwopRzPkya8WF9xZX6/8aOcduXaZXwS2FWtL/cUr9UuDuAaW
4ZFYtgNFB/ig7ZbjV78xDekHBz78TAdy0G+uoG4vp4zSApnBc8ql2S83BYsNabOH
gS3aRRlO5jK8uyxDYQ7dOuAxmSaqWzxLPqQN18H4OTTxcqeeZtfX/87x71vRDjmC
VAnAonWFOE45Qo5j2M3rPxOqREke8cYrwXhnCRpu21vtAKU9Qm1pYPT3iOlIKbES
pi+F6qUbk2BWkVjtrfyuEQ12NChq3dteeA/Mz2E6aurMsVygEkIR9/7CXStSvelL
wnyGBB0N/E66lg+RGj2A+4KJVOCzOZekkGbYUFGzis4HN0VqHKlBx7gjcdj5blNH
uAkmfNBXJVVub4Ccati6nyngHY6MCe+EQXKEUx+ImgS+zGyOQ4V9NG1On1FJF/V2
gcjKeDu3Wrt2Ynxs0aq8NrQWamYQE2rfrOP/29syDMjYJBFQlxmkCaNFR0fU/FyS
pVKQ8QKfrXbJeaM8dZJLm7REtuYMt0juA61vVFgZ4vtdFfr09gZB1T2eabF1TiaB
V0cImSwISIfEvWxvn3N5tzW5D0lhK8eN0RIUd4ec51No/ob9/DC7wVEgXRiDXvR2
C0EvyxlnY3a+mP6py8E+4nqM3BXPgbtjTl9QzBlFrL24NtYe47kKXzca8z9OXne/
89eIQZIzobyQESANms9IQzv3DuUGc57HXvH1u7QUUcFnCtgN57ERgr6G/czuocXa
LVuDxI27zAmBMzGAbApPd4GJXVOmtK9FSBcBUz7Lw743gnshbwKCFte4W6KXbhDN
w1dcopEaVf48NppxbLnhCBQVGd2xhMHVu9HdCXRd2LAPTBIJTcWZ+4xQIIjjx2DE
+H47E73qnsLO6C9OXeSnI2p3D55wtxiusQEIi4PmNgwT8Wzn4TiDsMUm65K0+POD
3qPZFYWMJVCfQt4qOp+QnvsYZz/gyo0H5gDIGeffo+vprxd7tXkqkRb7WiFMXtuG
BdzupRQqEFqePyBI8ExnLCayc8DHa9qI+UOmJE+a1tDCrHbHy3WIfWDBPlQKw6Y3
qUGGsqKS2cVKhzEUm+lmDpwoIOxK14M72cxCPT8cXPrQCyAzhQuUnNkmAUm8i4gs
XuKfDKfq6QHohNkik/+yhq13oAURF/luTNe98LJB2GEW2/tL085CJ+cmq0Isw2xQ
JeS1qfrYXl45+WN9oT5M0XCO41Fax9lAAw3T3KfWuHlTiJFeMwkVU004SjefMmQb
YVjdFyTP8N8YsCnUyv+tk9jYD1dr1c9FuYjHXquHSrTx8hmFP069yKnjcMVxUqPk
rmZvZ/7V66n61Uvz5x/hWuPPj0gJH+UsK064HvbB+QuHvgHu0Glg09LyjIsohf3t
4aom0Q3cR/VOdd+wnONTFgaN2WxaQogDEbF2B7tEUgs0sbbJhDstlkAbP2HQkT/I
VeLnBsLQPZaVlCn9X1E1DQP3M6fLLYjimQf0uRf0QhKVZhF8eNTil3SuISyZyvZe
fIBNjqkAPwqmdyfc7D07GrxzndtHEyQYqAhBVnuw7hqmOqx6GiAItcGV1w6U0yRg
ecLU5n3rrPb49RNRLysBGMiTn//3Xnu+y9CepBfCUUUlwRgxgye8t3p7J0ruWcPU
anrhLM/XMmTrZhEifhIOI3rfcAW+EFs8iSrI22rXXVFaxtckwN/N1c9V8kdKAjQy
8INoyBRszemWOT43NYN49GPouX0rZ7jIhLWliiRtlwFLcMVya8B/w0qZ1cOqZJDx
O1ecuATKDnAIP3LHLyRKa8ZkocBxkGgy9/YBp7L6YRix38JcwGY9V2SEwThMiu7R
v5qGfv+CjSITx1CGA+zxnH1fSTlqwBF7oBpAOBb5J9a3fP9/kn7OldX8gkz6k24y
ffF9TVRAat46i51XZQYcKbTgEmZLFEz1jPoHNRYaa0Gmx40X7EFIOgTS+vJYzv8K
jIzzcBRBzFXcAMqrOvDnamv/2Wz74VKvoesbMGTk2wKCSHioRqARSirZ0vGStUXi
eleLWHr6Zu2sLueaKWYl6z0XQSKdK03hRJJcOzt+L093TSjwVlEKMh9g1bU/Rwbg
9zRNCUZFiSlulRhn9LydZ3cqhtDcGosvLNEKFNa3HaetN4T94yFAwW1XiZrJEHP2
MIbekpmDUBDaPRz1N3NQ5osCWAufQsozhJXlYufT1+9GSFhhRAVlfslEe8I7KSSB
zWsDcgrr5koMrv++spFxaCV3J0jMBYYlH3PICb40+HnSdsOZWuitct/lJvRlNHf6
wBkC7Jzu2PYBw3/b+eIpFnn5EJ6bF/qATgWIPP/o/eihTSWKHUdDizjHqZkqeSFd
JabhTrITAysErEDA+m2GJR8Mkgrjc2UUUnMn2ze+8BkEZ0tppdNHTCHhjCgkNZ+W
ghO9YpWbV/aXmjLxiIl4+jz8dg1WHJ/DakiuqIgRx2ixDP4wx/AEyaCnk3nOGZkv
JZyLkHx169kKNlWxXcCNop8BuXWUeRJSddBDkk32bKpe+t2/9lvDmaRbhnZDs9c9
h+eLe8B36E8wDjwIj1jDHG4poqPCTqjGNTZxMepPkNYC6Ny4QN+4l7wvhZl1MrHT
I3F5K4hXGKhscCghIqoa7syHj2J2pfOLjkhfNMXBk/Sial4f+8lkO8XBtdrWuneU
WjafexBzRt3aRqztSJbbheXOrFAIghrtH86UH4IJOHMe4ihTzkRcTm9YHkIo8NCr
OUByMg1dDsb+UOVN8ll2Dk2I/pnp2pxwuDNShJKdvEd1Ngfi7RFA7FZ4C28USRbW
UdkYDUABMyOC9kET76HU4h6uE5bqfpgcr+ghvDK9zSAtiGzr+tp/wT5fszrjVS+m
EZ1Bpw5f9/CnQCyMUxYLlNWokrbLehbZmXJnszumXdtR4h5J4j+gsaD5x69owgKZ
3EUQWcLDRIIhlIxlzHpRS3xnPlQAzOz6zSPSPs5XVECYRo5AF6EwJk78yXWIBgR5
5tjqsAwRw1pVB9CilqBdKake0mx7B9TgO+vA/xSeZtaf4TQlE5fdywncIoP8NV6h
S9qQmFod0blI7qCLeD1mQi50nM6Dfb3l9uefNqREeRiE19uMxHmyMy1zBGnLPRxl
lz0vzqdDQlKpI+cUju76XEFf2cjEQyz1w5yRmujTMCO8GBslDxQwBL2H4p8sXOVM
CB2ampR5KppSmQQfl05PqgLHY5mtbckajZD8kkqQdmT+P+lOcHF9cmJBIkb0s6LO
fi9j1h2XMGwGxjIXzfzQ3A3T7I4Qp3X6cmLrAzjlUtsQ0KRJiPInvupetBFM5Yxi
S+DycmWHkSl+Fa432tXh+gNBKK9B0ASGOqn4q3ieOAQSdtvyJ6tcr6r6YI4GZ4Qb
DvzXpuwc79DCYVDOw2+RoxU/RigG+B6dnSV6afRUIPe0/if06HtZAbWvCGw6dCbO
ed5qypHr91jYWx01DZzeeRbELyFGwrwRa5YZouMa8z6nZMQvl6D3Z8f3RYY7aXw7
Km5IsoHi2FSYslnKdM7Mas4O0EHfJkDkqD1I5w/F2FV7UA2x5g5ktZiFl+/aM169
k7wcOMJzRejp1V908RZ46/QTbUFGaoHlrgGaGB6MaP7JE660yex3U5RQ6y+wlDpd
fCUZyUer1icoKqhhuBmjGBqJ/mS8WNbid28oLus4rkaCk9mxa2dMol9L+X0aR0lz
HIhfV5+qaDO9RQtssjyBMYYGoko9BAAymkaknoTjoUP0PzmMlP3hhEXRX0F+As1c
tmlWyyPsV8X9kNkm65N19ZT6FJ1U+P/h54rncoMAwqeQ9R1Y1Bi+WAs24I7tegEP
uviC/VqdQd1dkeKOa2Y/F9xchddO9Yhr1RY0hjkDzbvjFznYpdV2LKHBXiieH3kH
02j0r3i7GPiG6blMiYqk1q7RjiePhLmwYYpFVT3SlDh5OOLIzIo2fsT2pt5j97aE
swrZejozmCY6NHD6wI03J2mf1Y1//wFuZEFXf1KGzzBX4qRhunGI5Wn/WTT7xldZ
YeRsapHYvAXjdhy68JKpvberUVd3H+UGWxh7T/LzU8/126Edh2y0tXFxl6a1bFvP
09E2LUqcovh/9KgAVaWJm5G/9edeD78wrbABpO8EzMlOLZuCUKgHBdDehkQ38DGT
UU1JQvJ1NFzzSeimf8sQb+SmrXam9KvJgtZaTNOzDUU1DVazTF+Dx+R1MDldU5jo
Krvf4yGLmw+C1iJlPIHUY1adlC79Fc2yyP1nY9QRBvD9DKcZ/11l3qD277MfLgJp
dOtDq22IFVMzt0FD/gwETh18jZhPG6tcbb0mgd/SH0h1Rp9KZnSoyqyU9V+57YHz
uUmvEOUojN54R12X/s6wrYUjVQ0pcuck/awj1ljvg45cF+uGHUj0zH+PREcShzxp
zP0zi2YMPB0AtJ1re7EdGkwxR+j8qNhcNq+14sAavzgrES68Lr11vZFMhoqQTjYv
s1lWB0dgkM4LPP1LHwZBfAjklI4TXDgKYiIfBXA45fPRybyeQ5U74UTM61IBmBcp
MuSoD3/boLCfWWMQgTXkR6PKpxtWuTaOK1/8aP9mIXNIQxUwdx/jltCfGalZznZf
Vh3VXlm3B7kzNMM+H09vAjjkNhn74V/YKdFCBoqta6b2/H+urlVw5efbCCl9RG8B
ZFh88/xE8//qshCiuRdk2U9Ds3nBKWLdfX9YP/zShxO4DGTvXYFQ0yidIk94GemW
QZ56SuU7o3Q+XKmuBXCiyzWLhZYYSVUM35h78akAWQiuRrQo197/76mJ2TjLHWKp
+uc/o9tsHn9SC2u7LIpRbe5p/iZYzWdFHHaCIEgQNMJSfDJUwc5buMG9EQjALZ5d
yzeBlvAyTT9pL9pf67BnjlZKg2ml6+y8rnucLWQ9a7nh767/qSphSgBe6FPayDuv
s3hmLV2P5As7WMMMQbr1hATPRkZSFcpGHmdnAnHYoDwlRMiYQ4xQehJNQzM/V5Ua
Z5lv+5Ndpqwlq2P+Gyp2WPaqdgP3/B7EvX53T7xw5AuRZr2zx/Ezd0xnANXnx9JW
8idmRrypqhZDlvFojt8YZ4l1pkF5Am+rH8xpPnSDYShSerVIS5o+zy7KhlIDoiiw
9xr5HrhjqL5/+YHRf+V9aDEYbJ2lFhZttGwNae0cY6+ce9jqAYmwGe0ln/n3SYo2
LPt5wUHzspmKkgLp8+1px3FNV/UkaqM7UxYHMqPQzLI6C9nJQEEaD7cksgz08yph
a7tbbwpNXEhiERECxRjQpK1ao+H5d3wyCTtceMLeSecLiJTwCwEMAB4/LMeTk6Qt
L4tPDCFzHCWRC6hsCVyI1TcpQMmtpQ7zmOSa5FW2tcCuRn+AtPYPJDCQ87ti0iVs
qKmG1ikzyuZ38MPEfeTNUc+TpStImbXs0SVsYznKviL7aCX017HheLcFBHAbHCjp
9eB/l7jYTdaSsumkb7ndFRnVwcxIRkGCaFj44oRPUr6O3axAAQGkMXfNzAlPErxK
mV8WEq+FvxQEbdAyj9nhgYViyLmbEK9cTIBQFXLppIpWFCZcg9KD1FT9BkH9VAMh
zpFIBO/0pKvCv2mjvCT43yKsttk6ymI2UpWWuW/0AgmytCjd7Lijt7spR6Q0PfnQ
TlbvxVEmQX5tMjgUz27EY4dU0t8qE09xtrfsuepCZPYkikMgfW2L95etH5cMYS8F
hdf5NkOto0oLXxdhNSfUxYi4KMe7Qw9SIxquPRzN/FoqF60IiHJIvhtnSLRWsnxI
xbTmvYIVGrrLeRimjofLHpWGlAxbCWmU9sbvjiYJSWyePiCRU3V3XGTOvnQaTKJb
7SvKogxaBh2U5zZYiYXdE4lG1xNsARweXXZ1GES91pabNGc0oex+ltunklKgK33n
bp23cfCNrsnfsFe01bvMNbidsdfrqjaVebpQk14bY+64jn2s6AWcFT/R1udAyG1m
iLUWPKuH7GE/lqLoAWLEmhhi5ium8LZVqPKlycgyZ5E4FT8z2ST3wCuas7ln+BDu
M6NHnEn4EIro+cASWCLurCP+CRDGSffKkFskpg8vX8wLXV56R7E4bhOysmviQUR8
OWCKt5ytcneeUH2a1iFWjCyZ+DC7xWL5FO2SP/HtzmB635BsqQjOPu8j1Nw/sm9Z
mex9waoL5p/89LF/Y+0fisx1+x3Y3xJnjyM5FbMtq1YIbvuGkQ+wnmXmzP/tooHV
ul+v/eSpfxNT+OOUV1ZZtKydCPO6PgFlwM1LYLmdwo8mbGNod1gXFJ0nRTOvh69j
HZPz5/zOfzS8/7ruipVKFyVM4hhfTvx5+r5AarS5xgPnVaEDshtvVXHJ90lXw5Cy
8R6W2aEvjM6Zs+VGHHrh5yFpnRBCqRChJTkLGYjTsELDqn6GRP5LLuRFBh4Tn620
RgPD9mNS7KCkeZ3eEgcIXg56+YZFfapBCDES4lut5fR8j5bXq+4iFIqEd0OMVq46
Dz3Nf9x3UCeLA7iuBiDoGUhpNUgy2TbcllatcW4nTL5RP3okFsTHNG9PW1x0GJQD
ij3b6I6pwjtnBLUbGsA7RZqvmguiKZW0zykTk6Kkpr7lPhexqoILa7JpZcgwtuth
UaNYzLyQsqjkmSb77XKd/ROdl/meBBpWA1MqCesBlVb5huIU9VrGgWSLSdPKBwwl
4KxaJ03XMHAKsdwi67RGUPF4PO5fy+KMaDhERKX9xorKvmCW77i5Pdx4i2loro6E
Ecvddd0htcYKuKI47UPXhOlPCF154qOveXbToHB5/G9idVSfu9KXiLNv8722nA/v
iW9nG2OeMkP057l/jeSJ3AysxQmhKFFu1ZMZmCfi0zyG7gFbaFYzU+LActKc7FRF
OnjF7MYgXONPRL6wguP1xzvACMttGMgNm27MMBeWKJhUqRGYXViJWR692QBYNoxe
YZNGJ2fgD71gd1RO9Nb2X9jDHLi6ACOmTrpMagmOeSDA5gm3E3a8qpSJJw6iz0KO
lS32KQ3EOdgRLAHdNli6eHq0+A33OXmZPu8JVxiDNaNUZWznt7kDKxZvWsqOCpvQ
lOYTIjgSTok4dWSdWGAHC9QlOBK3YYkodK96MQcoVnZT3ozebkwPDZ5j8OsesaTp
N24NOh7Y3BBDkjEhBgTVxJeWC+p+shiEzTcPdC6BxpnXgdhgGiXmfrT0pgJAmdop
VeqjVh79JkDXS5uAzqb+3K4Ctq4Hn7IwvCDEjd2AIJk+PW+uuK0mxXhvBfRWmrJb
Gw04Oy6PDEBAe1etOLO0E0TwldHigCLJsJe+WL3T+IC/rm3fwM2rx7FXVhRJlSa2
lX0k2qWTwJKdrG5rbpTfTBdcpYYKqg3ttaHKtguzPKXp/cFUV/bY3CiqBTjl1Fay
AwmGN5rEHUgzRJITdn1pcgFzC3NhJ/fnWbiSZw/B5UApg/Aj+ztl5ViyBLRu847E
RgdVpBjg3fSjpzlpCag7mlLprx1Onk1ufu0xBro/Aa0xEXthUw1n8X27feBYHIJV
FCQafXnPuL7Zk0G5gZOJk9DuhxgCr942lzT0luOR23NipVUf5xlIZf+wRLwNdu2P
OQsKeMNQ9WwY4185/BvhNGWQwZ7siRKm91Oz9+aBEkLQMLgQXEcYP34TWmn7/GMj
PLWqD9Zy5xzHF0r/aUz74CXOvmnFBQagfTgIplF9sP6SMye7pDlQ+7COzw72J85o
QxjhoHTtwl6DsUjroik+tUcv4o77ljzfK76uuBvDCJxxWJBOjcCdOJo/ucAzFNki
PcT+LaXdQ9ffCnQn2H1VzIuneQ3bQmNVywBNizQNbTGlTL3ce8W5E+plLabCzK1P
lr5k4gTDfwHPtNg/SzXMqVnOzz5HlQv21XOODHxkpjtVVzHR6ERbjn4At0Ss61Xx
QzQmM5LJRmNGa8vavoc9PkDd+aWPBeHms6se+uDVDF6cDcGqfXxLk9hZe0viKAfu
O6ix0wFBWtAWnmlahdkRpSeMdq8cq4xu94uiXltILzBuQy8cCXBeY1nKEKE9C9g2
oX3XvNVgu6Y6a39bkcR2Xu+NYfJjNVqL06aWQoxtWmR8C8YyosKdS1M29hRWVZEX
dBVJT/0TZlX/LKlPGFA7lN0aM5+6fnAq4dvbGAL3FkRtxtxuyD3fmCoemszNeLEC
uNN0RThd4ftBLD7CDBMTc0YgLgkPjJgFCWF3hqLk8/KEz9Wy4oOYjAy8S1hUbg0W
PWTgJ/79YRxa5qGMsSR3iQXAsw4TeKUhIJp4ASjuCCULh00+/zrjwb/U1ZkCZNAy
7Uc5Cdx+WsdUft4LsfDnX0pWGONmKJAeNirDLDiaXFyIYgEAUxezua/0Xu09Rdh4
hh6FaqUGO7Abk7pb+RP/Mt2zCa5ILBcuGVqKLNuoURAf2zjMV4gkZuMbIh5UYnkE
Ozg67mI7iOOHRDqu+WjazgB9gTmdzyuCJsoTMdnbRPWz4r6XGnJ03dxQKjjnFbOS
2NwZN3d2A11GzkXLhopA5sMCGS6xuISMr61IpCc1WYclC+opG80IopMJzUVbDHYP
Po/VigagmAHEr5qjBr8Y7whpulXL1z6q0xTb3gZFPrDsoXiNYvY7aFCbRfGYH/cq
USWTjY32VSNCaeSdihrthIBxeVp6XyuO7Fw0/or4uYtsNXI33fmgDH3JT3p3mN7p
bkaXvCT2n6Mj23h8Y0sZMJ50pAO3tbYmuW9Vm6jMsIS4KWeaJlKYnz2I64QrXA2n
jUa7b2VrmXvxEcqUNMA4HJw/4nCThOWESyVRlFkcrm9zIoz4x+DuzENZuKnC3Hi7
u3g2OgtPQVtSSOWZ/wE1zpYESzkKubDkLd4PZx15aMQo7QGh+qg5huEyF4g7Gyhk
q5JzkPBbYNMoPDc8NmXA2Q1+CG9AbHc+UUk6qbqOhNQkgIzOwYQiypD1LaKN94Mb
CPxDJvo1EMgrBK9Sp/bCJlF/+AGpa6ZVOzaFajsDDSQh/jxIZwI41do4dGEeCrZH
Q+i68gjwZeZxkgMPWtE2xNVw8ZSqU8DWFZPIFIZ7/GJkzZALxsLFUY1uXYphu5a8
mD3tiunUsidAd3iKc79xFRzsMn65I4IbTShgO0AgSZoG19GgN+tJWF1VfRlM1BJ+
nfl94elzsNDI2uHSO+QYNHX+H4cUQ9iyrc08jpvmMQ6BFSmYomc+RUVIBQw2NmDJ
Xo8sMyojw51pdMilsdBthhB6ce+zOLPQFtZF20E8vsqk97Wm+/KM11HPCiqDKEjJ
87JzDywfFxeCFQbyjEYq/Pr4Q774WMmNJbNls4PRHaU8idB4rS7TM1LGHfNgWLbp
Gum2YZXY8BKMo/nNjjQg39PsB1KIGEogSplvsfVXVbaGS/xD6vsxM0Zfpjs3ZcCh
63U50KP4XTxxg9op4E00eeRFiXxxZSLXeegpAkrJXXW6PZ0Mx9trZaj4umztq610
r9tfWoznbYbuhMxM/04K+cOMeAR8+LblQkgv5ICRIvMCCHLFiKTAyb5YQ3RdeR4M
KUhMzXYYYnHeTrvDh19x2rHrnXP1a2ecNCYyKkKtONdz6tbjn1HgGADBew7l0+D1
Y2OTYFGe0AGuEB+G6Pet3PGWW8Gmts8tg2dL0kxPvaTpvOBK6QHU7SVRPSLfdpMa
7vrCb61AMlDMxfPzmAOvS/fh+iEDzwrNxXCuPbROk7B+oK/2tx5tG4U6Qi00YRLw
5WIKigBHxYgRnJhzeY7prVbijVTTIb4B3gw+0FPE5hkIUZ92B6KMG1jRTLkaNhep
LnQU27Amqw4cKsyVJR11WvuUWlaAANXz7/9ecBdBEFwrHTaXLJt/VKvb/YlTbGaf
72piWzuHHOXp1hm+YbrPFF9HYsY6lystoQoF1sqqd3SsC6/UK+tpdk7Z5xNzKryQ
Y4TQ52b0BVlo2QwaXTgRWP5LHF/8SUJ1GB9OxfM1rWQfoB/ABR9di4izD3tUOZR3
p8sheB9u9T38RLchadV891WIfEbCt3Ty15+0sQ7UdVI6ShfbtqDQjjCxoxI38bPo
+znYue/EE5ufaQ6ppfyTvpfaTmBFz3zUwRTKWHc9ns8VL3CBGUWbnSQXY49r9aTA
SxTeiKcOEjFtVGPMhpCoDqBjSNuaC7CCsHkDrYoY8UQPyyij8WkXAsm1SCnhc9pk
TgemMOZS1lmkjFtjT2hazbUrb08osCVjP6j02PITt271VQJM2OI8AwXRjgvAvdeo
ttHIbiaozjJatOlWU46Bnsie1WNDAyDkZySBtvUQ9khqj5vAflx0sUIyMyMhB7No
UyQMVEJ+nA2ANXtprumGXctKw4+bMT24vJIILlw589G6CIInTf20YsS5cIkSq6Ju
1dilRA/dexStp9Vgc84KpDfZWj0wlSjW5G4h6AaV3jmzoNIyIeG4SMbrgOxIcaOj
aLAG0yXHTcN49+hwd7yhiC00lARryiAKBlAW0n7WhoeTTKGEwvNZAastLs9qVNJu
8qKkWDKo5AR1Ary9Ba2WQsqyFfa9TcaAYd8pCCyUK0+jhUPQPclSo++lYYFI9kGb
nNrZvyyVSCqf/uj0WlV8LibgNF+PXPVnoKT5US1FMZi0tVOXh0OHWTSSL216K3BJ
nTkm6sKHedOyNzPfdlDQm9i0WypSQu2R4PQYJDlK3OC9POPL3JRI2PB0W4+fT2Bx
V/ZNMDA6IX4m6JHRLzccm6/5Aua/a5ajVVJJubiWsrP4BGJKpHeqk018aglyCxFN
d7Y2YhpDLxAeQfVWI1aPoai5SLq4w8Zety8KCnVTvcy4EdUau8sg09sfphBrJnmF
dOB03LZqa2xaS+AcUoemNt36Uv1NQVUaNJuB7odZ6Ae9edDPWo2WMJhaFtId2xys
liQmxwX68GEC1RJ8sUwU9MojI/lBdnUpNz8g2t/qJrpnLYPlQ9c/4dM3UQdQ8mQr
wCCLnQDvgu3doZGTQN8HTNVlkWsqYJgAnztahcgejTbo9ukGlwPcE5ptpQr+wQbA
CvJL4lcuygAAZl5ZD3LWlK3edClI1UEk+ax6Idi4jRUZsL9fO1mJwBqzWxQUHf8R
CwQauipVKMJKwsM5RS5Rc7ZOBrO6EwxehPovkOxyKapOrSYR5D9qPv74gmUvWp/c
5gZdM4P5E38JDHeQrn0GpPobV6w0PGJ0CtSelvhjUvGLUO756EKNOQoJIRnmQHo5
1BakwYlKdt/b/RQwymcvjYRd/DXcvS2kGZ2QQ9KWSVRJs7dA0+BoEGMRWOk+HY+F
EJMGiTR9HBAQx4qSlOIrL1YRzdLffpIAwROK2bEXNNqRonp1CGu6zdvKSTVJYT7I
vk1GsFiliru4kESZJn1XhVc88W5T65EdiQcjp/5i90ttj3Cn54fAC4fO/woLhveB
rxBhN0itRY1mdAJfFDx/tug2RSAEXh4GEdoJ0m9RH0yE8JnTYYB8sZm9spfQIfTf
fDj9n+K79FRr1MqpRwXZkE1wtL6o0UXfpzdah8Xj793tZoiBUVCY7VO4jL6d2yIM
MoRKRGU09yZyBpGzXX2YIfuP4vYmjkfh18MsQsMMZxUaKVbgCMrkVeMHIHw6sRxz
rifvRtxnteSD8GxBOqnEofssEwIwgN1mwyhund2CaIHjKZRdKXsaTb3uLYfiRIhn
eA9jVWT6HoGnHzD0BR8ldJhoNGqmxDwYY55Zv9QAxoI0RfjprXTmtW/6PGjurqqv
aFYfi2Jk56pce28chhnnerqhNR6vYvyqXfescPaeH5ygsaG6V8sZWY5tC+GWP1jX
5ON/n8y+MPJJEWMRCUfgdP0fb7RxMgU/oKJeXj/BvKTw7cQnX2lo+Zbh5go8sx5J
VoSMkWFjKoJvRCfmm+2SzjTQnhrU5d6AMvewvpEZDcFi1/IFpWqCMoJdJv+UArH2
7YIVorfxW747cQZFe+SAkrkvHkrpTlh5Lm7ZvGeB7CasSCPIUxEnZly9CHDFtSAM
4xeDvPXI0+8xK2S71o+3v34uDVnsLMDEnI3x6L3jX0aZsFLsC0d3EEa4iskTgzhc
wMXJ/owExwIVasQM/VUdB43JmrzvqWK8trxNHmZ2C0hd/I3SxLQ6QZyqmYq4dp2m
0q3jXEhvHhsnhCnMLV9pSrpWf7c96hyOkVmzfDwZDH9YFjw9pA3HbeFWAHGtP6Y1
E7HqkUDmM31LBl+0Ts4GQ8RfXmTwmcgFPxvAFXmxybLERZmpMTCkPLrsMImUMmcz
RE0o4a11qkh0XjvvJ9aHz+6Sd451KOcla0OsrleZt4MuFVA4XMTqoU3RpWdPQKeN
2PxH4l6I2etcf4MnS3UulfrZP4XOqgybZC5fQTqbcqOjR6qAIQOPsm0NNXmY51LV
6jc3mZg4qV4v5ZUqTuBodcl6g24UcoH4OrSF8OCJoDGUsjeH1aqiSJb43gq+2k+N
npV5gn4QPVduP2roSIEIG4N5xvIVo65mR17tG3Lgphho6urJyMY6avgOLWApXGL/
Lvm7I7oqbCKFOYlVtZgSSDets9rH1fEL0ryRlZUnEvnUMHrwnWWOvcARd5UMer2B
rmaO/kXz6l9BQ5iz8j38smYZLKAGWF1kCg4lMut7x8q6S5A2hhA3IWwpHxU6s2Fg
2avTIrJS6IVEUrRzwd9FC4gg+bicsUjy6yoMpUMQIPt922KK/2zRVAopZGwrjSpF
OxQYtUYxixcMCN7HHpFo+asC5smZZgX6+JOz7V7OXSKWhU70yDd8Js1JTwYRPchW
UJsCM2v7gbmOJU80jhDfDgF8N5vVrFjNl0B/tZeYXDOeMb0Puj6SByJdVGmeODMV
jPqtQREI/y9yzmBtQhCDz7LNJca85nlRQeOeJvGETBefwAK4eaIQekywzEmjb8rS
/4+ZCPrrE6H5GT4LK1rYiG1EkcoN8VLBlVw53BPny/Tm1Py/rqDVYzn+vFZGJLLW
GApdk0vh+6R2bj/4MFAp2dDzGGH89IwQAp6W57vLro/vesz+qvPYxsp0nzK7Mhg+
Eyij1qZ4f1gJuY3U12anXVxjb4YvV5vwos7ruQ53Hh851TEqZWkQHAL1GUIyh6pG
AIQr8kpyOTmG445+2g7Joj+yei/JByMm5n3hD1FSwY/qa0fF58w2IrdxBG0AnoTa
YRltshlFG5s1Fp6rxtbkIf0RpEgDMPXByjpV+nesFNl2HSynS4rloGavi1HtHerC
GZRHuCra3yqnaxG+IuQNc9k2mc7TVwOOxxCTmGpzwCoLDuO1wpt+HDAh1FcRqgcj
A7D/rshSHoF2WfzrDlwhyQnBBYcfyQd+ivzJCFk+icJOcrzTBDXnExqWBKPw+byG
bVN4QwH2LTdvzQUSvKoWXblArVT0SN5yF/qtPca0wAmF2YsrMnWXqzUFhAcqlYf2
H1sG/Esy358U+X7juK+2/qdZ+rABx85f32jttpUX8tlI9LCd67nVgjgLAiqhy9TV
3msx4EVm2yaNxxZM9vn7I3kN7T0IeVfDSdjz0WUablXpxHisV/PBSeBMK0D+WRIM
8kp1HYIHjW2NKHUkO6ngSqASZzEhExmu6Zk0MqACNB1atw1POUeFUC94n0MvjD96
ITS102ZUngQLKwJCaSHwtwrArPYihQHwNaZbJPrZspJ10k94gALLWZHzRB2DbYQz
DPeqt2+6+/2IR9csjyGYefU80SR/rp3GTL8zaZ2sz/jxzxAgw7c2MxotzVreps2i
JXECdFL256XYTAN/fRynIynylazXPqgk8JHDX3uKTk8cwMzNXE/YO6S7fe1xDxKv
m5Fnt9Qz1gQ/OuagtP+Gp5V2xNowhCCjT3cqWUZhOpLz/AdMCJDtROUolREtMSon
fZ1qiLZei1FQgoz+okojViUntFvn6huBWaHFYiU8o3oNG8fXuhqNbnNRgVI5d3HP
HiWNlKjXK4xG/V7Mvfes0gC0BNTvSRUWP+HaA+6ccJPJAGMHZxr5PsDvEw/aKvgo
iqowHPQyGDTDcZSMIo2AuEbTX58iq2ml7dgMwC4s/XIJptOXYnHGGDqc+LjxNSNm
BmXVqzpL0kt2Jsz6xCPoPtzMVvndryoArsFSLMFTeA4HjIIWujDnviLJ4cuCOoLO
S5mQ6FuLFzTVUVJxpHy02avxeW0Q2UADpv5TJc+uckYIwBMjFCbvaSke8ZsZfRkn
3wid/ruTB3+7baeLamo75m9wRLyo5aF5GkAwJiL/Jn8ZprTvxzOmzeD7vca+KkdS
THey/g+DmAlIQ3h+wkAJtt5ejdkcRMwEz95p3+Z6p4HUHIKM2s0H5hW8lH01H/9t
aLST6+BO5ZGwLSuhZ4tk8FHIYqz71aUrQkzLfF7GPakMQbdRwKab45Y8c40deB+S
ykZRWy5ZOgBjjwTL4tLi3nM/Wu4SLptV3pOn++NnfSZlCOn9KAji9xEex0xYbOzL
KSVHJEc6FLzoEWiP/14X5LqTtnUdcf7PuCxhU9B2YD4bq6t0eVSRMThvQIuJqp5o
HNg5vYLOTw+bUmKwzDGCzgy2AeMDlno60Dh8LGskqu922qc+26+ck2U8gSIGc4aj
vddz/CzOZrExNNruXRfn1F4ISEjjfgrl/6nOE8Gs/k9NTapcBB1GhJ6si+DRHik+
fbxwmjIQTcR9xmrrvONccuR6CWsT1W7UjBy8Szhp+hT+eWb/DfgS+yvvQWu1LBrz
x11jNNKbC1jaI5YEaeMYAl+CEUA4z4E6uz4P/F9LHPaJsFIUqvP24se3gcb9nJNW
Vm9fE2Gk25U21sfJiIMDpWuy43IJkzDaTI7lDfNqQT8aChcH6PweHLWFlgOMNevT
JEiiWmLluAqoKvvbHqw+hh4Ql7y6qFUJ3esmWQs2dgDDFKPX1mUXiHbeQmk4ex6Q
O9JFjgNFfCXY7KIZjni06dW8ssVrwXVPxwHZr1FETf8600yG3cO/K85DKG7rFEge
osmC3UxmmrZ5qeguyYmVvJbE2cWvyj/2U3eimmgWN4ZpXQcNtC+bdrJT3m/2VsqA
u9qU8UUOY1Vx+7kRnDkj4izBJvuQIKQSguCG+MTinaAisNSPhqM2OInh9GFDuW0z
qtoX1PeZKPmJRR9DdyWg3lR9qfLw2VZalh9KfKN+SYNRHpZdEaGCe2fo16KGD7Pw
8YShPQ6nlWld1hB8JL/Tiz1uOkrIBs068/CH/KJxtmvtNmG5M0Er8TJLA9L08zql
Wg4y5RutIgm+DujCmWRwX9Ku2LwXaNwHBpBfD79yEiQkcGk/s0lt3JboX8Gu+Nlj
T5IgQWA81IEMH3er/Ph9I0d9zKUafJmHZzKzm4E0c+5wtqFCzFBZc7JLGKpgEZmv
M6nQZzUDrjE5C603LJrICWGzRTx0jNf2nqmAN/m5uT2SY4vNfS7os8LRzBjNCwVp
zhDFeIcmxqN2g2YUul+oUVm1vQTT6TqWTaS+9evwnPPoe+uBVIf1Kd9G0+/ww8Z6
+ayGwMjEne0kZQo3Fbbv8JSkgqzdASqJcFuu36UDuBKdBKbIyXRaDNupQ7P/phfa
MSqSRZCMNltBLJ1wYR9Fkzl5AuoCfS5AjEuCOajAzTGRAZsUhd62NFkuoHQqH/1R
7N3Aex0kULuFb3CNxjJI4uyq5ntkL9mA1Qo0Vo9cfGg=
`pragma protect end_protected
