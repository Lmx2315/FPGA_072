// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:32:40 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
VSKnfDYrL0bmCyFusZ3tbjmI47MwPDCYMYw3CJtksuqBgx7wI0tPVYrlPrq6QCBg
Tyy1r7pqHIFgx7tTAw9PqMUZopwTUBSLFOKjNVETQAubxOmxwRjAMEBr4mEQtWsA
DPhkl5o4Jl7oJQcPYNAjk9p/hDXkITJDLDmTCoKZJyY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 4784)
mfErQWa2kOste57+N+lF2nb7nyVo7sTjf+E0sWuPetmjCZEgvSZxViYzlwRvNReq
B7HDZO0YmJHsKPR/KmkTnwP+74ho70HIDedJDZI/TNeUuaBuRvPuZ8IR+HgL4oaR
sVmICLAeW6ijvNsRKDHcBrUphZJIRmQuHhvVOpl3TGq7b6fNTJF1qfS8d9Rl8vkZ
Tl2HAep3VNQJYo8nzHqPaLSNV5fScTpG6CTOWsSNnDIgl1lbpOt41vJfXbZesOmu
KsfCh4Rws1Aw/nFBLQbXmRMvgjxCMgHxPb2xK+vpjTwukr55M2Lmedy5dboLv2Uc
RK69X5+xkDOK5zPDqaK9yuxQVyrXLLpJTNyvbF5v8BTvTdwOOx1kJZRAB5pXA+/W
A9cEqmqwPKg7SmYE7Oxcfohw+0BshD+RJ7OCjB9ikbl5OFPyXoENXRtnPMIukJUl
Y9xUWmUHxwS18zHSIP9snhBIlCcWIPno/F8FM3ViwA/MiQRaRQ+JweMU2apUs99Y
ug3KnQk5Yy6HTd8H6GoVbubiXX2jmCL8ihJZ+SzGPRzLEfD/SfwJPn/sng5kGtM1
iuqP+xU7pK1hvME/rpIB81ub2XTHXKazHRLM+DcxR/rY1OOD9w5BMhFA0prpu2zz
4kH8ZVfWZE/zDrmE0K+D9tG4xM1jBTZqTg1TaWTU/Bdy30lB3ipeVZUiC5Sa0/sm
Vw+bbo+ZTXeEvoWVtcNCgcpZJy7qMUw6u3njE+d4Ddhd24duyMjjDBGHL3b/iqdW
oLuyT/G9QqL5lNgnMeouzOVYut5+7UN7+2F6R5c310Ogv7bntf18lLELlZqTjoVF
hq1WkE5U9QcNRqygoE1C9T316Dt6IUmOvrLQZJc5fzoNTRZiBmOto+j5/xQ5y3ch
amMSX7f/IY0msGrtwv9d5FUBgEbybOD0qoNVeQsy27FMH5Kbx3YLWgBLAi1z0J/L
x/DGtUz6W0ye9e2GPikgdlNuKox9ACkuI6EehtMt/fQP/becS8zSKY605zJnysfK
BwdhphtN3xLF6sCJSU7tVTyJ8mVhgAowTYO0g1WEWB2GbDgOjI7oEu49FS8lcFIE
qe/gPGqsLuucb3A2atLcuZ/FJBlx2qiX0OSbiY4lJ8WyQauXErnyw6YaDMmZHsUD
vUrNgP1/T4Uqh3opuHYcL3GmRhNbLygnH8bAnTZz6agcmHvwmtxkbncRalA0mdcg
Cf+j7RoXQh6IiTmTTFAPOQ9Tiof+nJjvs6XRyOV4z/K4UDkorYM8bX+sOUc2YyXg
bZkyG72fBxk7VQOS80FoBKBCFMRrPsr+9BpJpSH6wBrtq866mWO0CNva0DorfS+Z
AAWH1uXNP3OuK04eHdAdzccjspvRGQ28Eyy8f0KWUgXTPcL7GoAWGGN+LopXD6xo
Im50hAuEUA+QzCJpdRaSpmB9IFlga4oQdc5LJVxPwpUL5RQy9mZAECvcb7f8IOSK
hy+inDvoKsRZEwTAjPOeNizQgK6YkbCEtTxdL93QcNOglqJLlng6tDuAe7epbMdq
svog/YW86jzBkhrilJLgtDAAsw4WRhgr/QAcC3qaO5wYJKTl5uc5XHFOs0WFOehu
HforT8CivnqGJzDXLP4wcCkMekcbK79seui/EDgclN0Beb+GoMcVi+noLJuAs1FH
Fj4e6vaX2CtGmmRWI/C22QYd8JfsrwIlAiP/RN/0vMka0OCyRzpiY1mrWsaxbu1Q
y5KzTrQkQZOr02zyHIXaM8nQzdyWRZnYbbSHw4jH/NwcVfm3Xn3FnmBtRmE85cHu
6Djxdp2+t/G7CHWUvO2eIAH4TWG/Kh4Rc/S3IwOVfKNxdcjck1AtW0PvFgT73A+s
mZQGGoN4P9ztJCOUYZ9TpMWXOr5L3aJifhjdlIWJu0ZlasAMQoav0qHy5nLfuRee
AZ0ADEe2dsYFYENqSAgyx6JKwNNpg4FN6RZAFofXxOU+JCNp/PUNg1+yP57KrVtO
ujg6Y/i5ka2081WGGjA4IMfLepSMgWFjvn3NdepUxwgFQlkE0Xgq1gxLMG3lcwKo
DvtmDugisGfwlH60u5IJrNHaONeu+CvDvi2bBVqWU+QJyuvHdsfX+5AHsBj+rxsx
zNhFkyR4PI3iY3g7/2FPUVJMplmyWYuoeQfuy4Q126ZbJ6BsTGoA8j/0JWlxMrmB
DZohy+KGB+yi/s2xLIADdtkWsqSokduV15ZXZZL7mRf/OIb1gjkaicsCpicKhnE0
miSiTbVodRY6/kxCpLnPhphU+ccwfas6jwq3WPkZFkPtMHOSNG7y0JY0yHDvdbK5
IJ2lLK+71FFrn6XqouBdwXK1SiGcTa4Z4SApk5kte1vmphju/iU/RIew6dFnf8v5
V0JSX5C48lk17BXNK1uYrAeGvXNJZ8gTgyDG4EM67BvDObpxBRpd0zDKupvJPsdu
D3FfROO7Qc5w3ytg6pio14kFyr8102/Kaa7ctZyFRbfLQmYQ9adZRKlMOYogATWB
aDWjKPnfC2P3Bw0m5YUM7VVv2oU6bpw2GXsRKe9dIu+7lJHvRNbTccdL+JpEXAFi
gAbDR6A3BRa0MxmRqHd5QZlVIYhmZSeoGhJxxKF5At/Fa1rv/N+M0bcoX67aIS3u
G1Tp8CufU3z4ANKE69Fh+ZYlzm6TYRsKTPAacrENCYBzOTehPgrdF59MxoAPLIr8
QuqcRmP0CPgQd9hNu72dAsCtqf4pHKdvKVebqbq6cDiYPQv4z0jwtISoBjwTfMBI
19Y7madr4yQ/nWkCBQ0+3jvcGmxjwitwVE5oFUumRsE6qGA4vTa2w3RTZejwNgvq
o3aaSqFRi7Tg/TEwVfNgWua3mcsZ/pV8ide3YLcExPNuflXCQ6yC5dkkGT/Bs7Vo
yYeT9Dzt4u6OgaTDJoF/SXpeFVuGqGDpvSBQGDGntlG3WsjkDx6MTOd2zD/AYakN
2EtRg05Qla//iMi9OxeK0yXaHf1kBVl8wE6ZQ9FIqE2F72ZAo1L0SnQjOlZW+mYX
SQaUcKBo8yIf0aY6/Q0R+G3pW6n6r9j9GMSR0NIYiR0UJwpIxug8lodDcGxKPZf7
B3LEJD/Sxi2gWjnWdPw7TzhfL84sSqL/RzWujFHfBzWHeaVdubXErXBINMRnDpJE
wjp96ZGclaKqOjhHF1SHgBY3ZGvTkFdMu3vLl8+mN48O2+eslhkWP8COfXST+lJG
iiG4tUBfAdgHlK08g5YZ3RokTao77LfqLdDjZtFoPcp9oKerjPcXlgIzLXl6zTXd
m1BO7XC2C1Gv+wWtofCRgezY/De5zHtmKhA4P10M8qwDMFhivFz4j/98cQqIaRIY
F/HNltsp6XUFbvLXU5ZhRk4gX6Bq5EgUHfcNIb0/co0HRy/tvmKsQqsaKq6jBJvb
WhRadxlPjlDFdAFPzwisn7AMIJoVehgCxbyT2guH/65MKSPEKXMS2zANdaN1LFBC
yISi6qv0K5hV7F7BvZMMHVMdqdtN/X5NkMkrFCnjBkbCmv0DyPYIwXCM/MEBcuGN
B7k8FqN909DhMAXxR96RHu6Yjnvs4mAcc/hWcRzW62S126V2OaV6Kua3yHS4O6RS
WSfNiDwFtDa9NhneojMYjpAAcA+q4/MZYn8KiBaC/xyKBkPFszCpQM5jX56bUCgX
q6C7JjQ0G26ZTWf6nbIZb55/Y1w0fMqCBKaXEDKOCCLkrc4Zn0J+96uioOXlySab
z/6LTrPQEFmkoVIvlr+/nZvZuRZIqZbEWs+YHVHuoGOmIp1u0PFxLU/lGFYne5UQ
CiIYUNNRtbDll0Ko1+BXn4nIJ4GyL3Nwq26573Zscc1udT4NLAyasdl0vdcVO2KQ
sgFLVOUvTx5inj6FS7u3zLB+f5C9M+kyJRjYk+xCNGYAE1oZmSFCev0meD2THvuV
mV0H3v2zjKbeVZTFv2BoU5aQcEprJP7/XmBpSg3LF386yyexy/s7VOSqBnjqn/DW
kU1KlMvRz0De02q/OQDLsLmI9N4xCmmaErT9jQrUdrvkz7HCiJKKlBZYmv8ULgLz
U4kEr5enOmzA7zY6WuZ/K8oM0PxVFTY5eGnk7vC2IZ6QNR2e55vz26S6hxdJtAd/
sn0DP+h43jWmvXXu8fnRBYgvQ0SSF+I+In+q256okJDFDJVQ6BBZC8nLLad6RL1k
BI6InTwYVWR4acQC0pME9tQKeN5DjS7L/aqTzp+yq1b0Bqf6dXGos10ZtmxnmcPH
JZK6tu/cwyQwR0hA6yQ+F711bwmvVQFm7yt4epWzrrIAGcR+DXNrmF1vnL+Ws9os
anA3SMUjqRKn9RZ43X6yQAmqBtm8jFEYfZbg4fmpkWUDNhpiH5ygfPm1+OguC5bz
pfFVpnNoriRFpKBXCk6RTlWjrBgBrUCuxD1+5STnhKMilA4kPRbCND7W478T7J1I
iiQh7j/CAuXMFUnixMXpFOgYi2DKTWkqEiiLIcolhkuCdd36mJrUkGiXN/nxypft
FkT/qWNT/wB1OLLwLXLxIm7leiqLMypEL5eWdGkrWq4qeoj5UtumvV+GMD1+omv+
4vkEW+INNUKAbxsAictREQS5ZdCLTz/iHzqoxHpe1EudXj7UI8Ldq7dtO5es9080
EWzBo/hHwuC311+V/j2eHY7xe6pD/X7hCgwudoVlW6h53KT/WBFdBZloSHy/fXjK
ijnWOggLhvB7n6zU0dkf+1pEocaQdFz9BV2wXjrKAd6RFcogHnVfX/Lyq6q63bE9
Gnc9eT6FgS03/EBQv5EsgnEicC91xLTLgvHPTSn6CcE4tQl5x0w1axtF4GOKEQrA
Ptz5CyM8lVLQ1I12SZl1yd03bGYxRkSCXlk3ev7ozbTjKK9jOWY28LW+RwyFZPP/
xzaOtb6+35HoEMQL6JPmnOg1MKinAAIDLNlEtgzjT+9AZtooPM3zcoUAfxM9TaTg
zUt8m93UKiQNbRbCPBNDyKIK2cQlHqIKb54eOFsjih8LLSH/nreBmWtXWtMdqElJ
hOikoYbY24CEfAnbrLNNahpktMHg+dCK95UALYINGjkLM93qLfiSGWrHa1usy3Hz
C/k5gIK3y+i16ehKEHo2lE3nfiVesQxqPUNxDdp6jKtPrzUSNmZ8IxmOavE9LA8v
gv1gf8bmyH9vjCNH+ISJsLQ934o5AdOhZBGJNnPaQeBBzz63E5nm6TPaSp8Z+7vs
Ns+UIPFRU6yfm/V9D00eBvKQ20ebhra3XWOzsKd0oheiuwyvFkC9w2Az61ueF/9R
MTH8EMZfxxuTxVfNvy8pCMTZlKbpAmaiKnDKhO72Kvdz03IYSrW29jGsM9ygONvM
mt7EMK/uDLucyzMeAkOQIK+5WRDcjk8PhzX5/CiD8mu7sZ5z14/gAoGdh43HtH5Q
80gE+WqMVntH4KztiBBrWSqkdZG6zGTyBqL6M3kW0WQzvbRoaHlshvfjg+DYZPWM
u1F41FDcmPLVCNKAZXDWFhLLYj8LzwDdUbS67PT+3Xtl0hwkMDUl5lE1SvjiEnJU
ddTvmQxTqK3hFzyK3VqKrN3WMMojjAYIn4WFLnn5cDZfx6slzr5hkAmAB60scfn3
mxS1YYyyVsGdJ7CbHS9zGidKQOpaUa6MDYD7wKzKuYbVWnv5EtZT+XAbPgIzaJ/v
G4wQB4DVNB0TMDQB4V4ZTkYAmS2lsYCP1m0yui76r3/JiUW/OFeloZyQmxuU5kz9
wMTzCDxI1kT6qanc23XU7wRvP03AuD6qZo2C/4/FE96w87ImWkqdpD5Xs8dwIJ4m
fWZIIF16ShwZeRokoaZ2Nz8YBBvduZU4xRt9wlPzYEspJzijndRWFrAHsGqNn/Ki
qvvvtRSrWK0MvuDSDLgwCCPrNNRkVm0wK5sfebARTSVqXQxlmYUgVR2AbgqyPY8j
53HpRmFPfvxNuo27vpioaFiQ0wBFU96Hx65s6dsMzVkbPHK9lVT3i9Lzo6SJvIS9
VYboXYAq4LyIicmyKZ8fskJJVrCAEHC4kKwfLQw9gggei9eSBBmzXRMDvWnJvIsL
HXjKG44PBZufZtCOew+0YrJWFemXZnJfBh8x3WwdmBnr9+wy/l6Hpp0fFWiaspfx
RHfclTl1omYMPpvJrWMTA2TjpY7myNKBDVuHcF6HccIdsgxpJVsTXYplQbuXpJRN
+/3dsgfLEMLBXi3VFIrqkM8sfi0xkYNzvKgCAw7DNDodPwQy0aWljG0WgF45fMdB
jz8LxchtFUBN0NYEcVBN7KH+FzimPBfWByLvj/e7AbSmVwMOoHwQHgnPr315hNuK
OrezlfbsvS5lBeXVI9QbXHRXzx6NiIu4XarKSOZ1lPvoOn6rPc+V2Kz8SrrISo3f
C7tGeB0xqSniOwE7cw8/7bizzs2xxjN3XvUCeI2Y8zE=
`pragma protect end_protected
