// (C) 2001-2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
B7tZJMObsGf5USvgOdj92B+7xrIAVLe1oaoHMFiQ5zwYGLczBtx7yQfdQ8vDaPtt6AcNDYwZ+ZQ9
R/mq9lH5AmjXEohVUrUBKEDJ/Mt3uho0usTWsAHY4UpkZvUvgPjcfuKTzgauz4k7UA2Sdu3fd7Oj
z3rNeuPYQVCRezhmWU7gHPk33kfaKWxKO+nK7BfqZK47D+fMFl2IFVbsyQpjvqg/bwGAHGH2bw4Y
+vlKt3gDAzH7DhvDdLLmM31rOy+EKG0jco+ZIxBYIeToIO0xUkYAyl/i1BqjubKAeuVEH6IVE/OK
/EUqgwEWsatiudcFcUm1GHkYFpBswtIAjUPhSw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 24432)
q2X/nqCd+zI4xu4duevCWfkBs7ju86ryJYWwmc3+XllmgejT8jgf3TR+ENzSn9gYZjWLXrkre8Fl
WL6v5VzOHBvyS5DlZNLoqI57Nx2bjyNH0oV45icfNmtmKH5RTViB7mveHRDSoxnQJnzPcRZQAX5H
cAcin/R6QVXQsNOY8jO7OYrIkTW3MnH4q1rL2h1YCn4RZUZkauNcpQ6ZZBW8SoAEHo44aMGK4EpM
WNGepXPj29ROGe9oD9MszXY+a6V5bxHwpI++qHj1kKt9fLSEpiEXKGsy48g9A4txjnv5RRG9Pk0S
n/eVj3FGZZ8jCRvm4lg3elwOPxmgatP0HxGXzgrKiShufJ53K/3LtitnTaB2wtNJM3ScsVQG8HTV
R8MnieALn28ue5a+qtFMoJe97PbWhlLc+ZLgz3SVlXdKnsykNdjXqMLOomjW9NBOxa+CAVStsFh5
Djs70GG0IO7gN4WYYK+nMO7/V0mcNAKKh2ZecZaHIBPUltIXMUe9jNMOnIuone6vORpNs1GkSK3b
uln+GhnnUb4vEHAbUIf1t1XfO19D5s56hDtphWPJJUL6xkw1zRCab/2gak5cuXRYYCj4BxtDpz4m
7b7kmm2ElHI8eY5kkDu/kR+xl7VYtid2QycT4+UikcWDNqksVXaHm7+ImA38VwLFBK3s/IqHnKKu
aQHa1zEq8W1wlzX9xBY6GlPbeXRvp3T+efDFkIXSGlA9+zflGxD1s3NNkOBmWz4i5WwqjxrY0aDU
r7dds2W4x3pV/aME1rrdnvOUStSVk9oAauG5kDA7BNaw3zIM4hn8EmhJ/k2QtE9FotT7YuO9RFQ7
taOETuGalPGMYgvwBw9q/vihWQGWcOY+ywZmzMu1tJbp7pa/lIDetAWNN+tyivq/pnvd/kv1VTxQ
5rSKyVzuu8zCNQT4wrjyxor/p+WkY1dxxJZ28Zo1eLU8eOZDI1/3/DL6oCaMuGkwJjIS0wg3fN6+
VBH3xnnTHtHJv9pDUTc3ws1V+mo2f6QsNPMJMkMAXcA16giPqpn9EqFNHj4d6CghwE8vP1prDLlE
jRZ1yZ31Y78KvVMU1XsOY5yS0RidPFOcMuMTbNUptGT4NFyQQQUxhD/vZRDwkR/8sHHUb1aLqyoo
ljP9VG92ymye7VUTXgUHwiE5k3OEpZLJ+DZ5og7OzGJ6sbp5ZVyQCiO71K79qnBdhKlzvYQqgBpD
eEXcHfWRnMePZaxCO8zQ5xCRr7c61ihDRjRgFNJa6M1b03HTKLn1JmxqjvqyMj8BNOnDa6ivMGOs
dVROPQrC/fqaJ8AfpSm5UqTeoruB3DFJ7gVVr2IG3DMhZYASS/c76zZljgjMVJHT4NuwSQ5UQd5L
+ZAIsq5gyI+6dotCSSS+2ymx5oXc6/1450wyzcpor5E1OXquAYmjJMQwf1iqZ8Ke8ERtiKV4PH/B
Za+T+fi8hLu2JkjT4+mOmCfmp++erckIQ4hOf5yZy/dLlEBZ0OpfgndhFJz2yiOunZlG+MaI/qST
vWfIOQpb2rKtpV4d0JU+AAn+YW8pBtwZsx2iW4aI9zAhrpd5V0o1CtADoRH9VPdlahZTVipcPqvq
XNhRCjaTjoy6Cu/lLbZTFMK/ZfYUXqYxNasBO7nnwmX1SIgYG51YjPzArVB6Vt7tOPj8p7ze/UUt
Ob56KjN5ykoq39JztpPs6f5vnRxxQf7XMi3ar8pT3UzGGg6/EJUNdsToipBVDQB0qZUJ7qyWZyAi
7anktSdldwpRLKVmeLCGaqcPCzLMxzrmi4YAOT4OPMuCXidAdb4bcjtDoFJ1/xk7WGVkrEEAnIDR
aZdG+/c2eMDrxPJVZrrNYZyDGGIvyo7PKk9w0FgupD36GclObi0Q5T81uGgieQ3JtnTbzHeqVA3p
HIJOk0MI1ydELKwB3G1imPk015MMn8pDHDJ74SqPxe+4rWtVgqSU70+9C8rbJ8YE91imYZE+hODS
22g4J6IB2V0l8Q0cGtJQuXjNKL72RVxD7109TeGYIBLqzgANS04Lynt2UhHBhqB6ClVYZ61E5Euy
nx1nKJQak+HKf33doFdV6nrwiP0K2n8cYtBdrwYqXa8Nj2hm06OlIyhSpGSiFItYxFApcNjq5OUn
HgWo1xcrbA+rIskvIIhiXr0ZukLW+nauDthjn1XZW5ONPQuzxmVTtcXuJYVrf0MMBVFd2nXnS3us
ziLPiOq1RGFjiioTL8p+tpn4nryLPlzcAheOm1VbYSh4rTpobs8i1p5flsVsCWBzx1wGQpX/Y9wL
Ob3QKkGZxSDNkiIc0hWGkUxAa05cKDRD2S5LZq/u4+nSV6Oqwo0H/cMFz4YCJx89VaNafSCVWlJ9
E3u9zhuo4fd6aNdHtM3OtdWa1tsAnr09cwaBwN9dKsB8ZvvTEGy8Pqj6ZlK+edRA5gGI1oVgWToh
gQe5ZFGizENGvqtevdApXrZJx7lZuW5M167S6+JZqpBoUivv5c3CmF2614ltbQ55B1Wc4QGEED88
rY7FBjlB4+7LCD8Uca31zmjWfQDUEQNaa832W0LwctJWuym5kK9EFOhF7/TuXQijzg4FzFMVFA9+
j2k+xd68tUqoei/t/F6s3bo+Fmv54NOGuvgI/uk7lSNXoiaKXgqfPW1gTU6BIBsxUSxiujJyZTHk
u86zQnQM3uW8WfP2cw/di8mIrz6ewC4tcK3Slw3reOdetMMXqnGbSfl6h0dxJh/l/+f88er0WSrv
0QePmt7JAs7K2zTTJrVODicdHWejN07D56PW2a/wczay9KyDw5gVcqQ7H3hcdAoOVrzW4+LuI6Vo
otCFHMA7R0Q7lNI5Stnel/JuBh7DFY3bpTylWJzHhqlLPaJy/0t8QJyyRlip4j9DjbsHovCvKNPy
dDvkoznexDL7IYlLYcoCuggciwx3ItuN8cQbshOFVUESVuIa6Gwv3xSnWWlOCpoIfe1WBs9GCUdX
Fw8EUxp6S54IGjM3hvoWDh7H+K8/V1DSDKlUKfoU7TQ8GHAza5CNVjlNsrP1f447y4QBrhoE4cbe
CZ+USAdQcb3V8T1varO/gdou4UerJ5IptM0SD8XRuT4hVvJsS3gzh4yJMscz/n/9YzYxmxQ3qkLa
Ovwd1Mx41wS5XLfeHyHdfQTsGscsezSmVMqFgt0kGLEW9YJcCHiqPAWD/zmvrnH5Wndud4en8+Xy
wX+dAXxlJEqChp2s3Ui+VK/YLKXQKUGFPq/Fk8WqqIF56U5nP2zLfPfU+euiShbk06H2JnCmxSwq
O0uOMIg4pLgbcWD/Vi+gFyVExAxYjK/5sNhSu/oh1NpISxqHtaTT83VQsSL4P1IRLbtHVYTDtJHL
lEdW4DcZdg0zCd2xUfXIVMAP1iFOsFfqsSeU4M5iSK/0Mk6VTj2GGfDnHLtWnjkWKrdknrsYg5VN
QJtRY5V//ZaSfcnigw3sluezASpkFVIOdbjJeo4+oiBKHRgNaYMlSYkzxC/yqC2NcBN/HR1gfVpn
jGkNJe0mBj4AmGM/M4aGAaOH9U32xJ/jDwz/LozsCcjYLUQv3ohzmG2L31wxCNGsfWg7W6ZOaw3A
jNn3QZCTzj4Blo7UGIUhuulQBXsWos3BACRl81WsrJURsDywgHwF56pHJ4i1El/CHGE6ywwz3KCW
uSSYLHhq44MA91zQX4CdPhRWqjDUO+4x3298njK/J81uz8V9bh0LJv0yOrSLuiBlgYsnjWmZHZ+W
e7WD3nERFQEnaSbByyvLSp3Mxkuhue0+x7OERZ3+YnRbITdDHKS7+sEFC857IbUitbitm+bF2dRv
zM3c6e7bT+Udg10HYh2GF2YscKZAmfI9fNUEfqhavRfTcKU+qGQooqKPAbRFMCmqwwgCBhfBB5vT
0F8J0WUzL5eH7bSapOXiKFRCglrX5HEiRlT5MT9FYf1dQrKll4Js7TMASr27wOz0TTg80KDXFqTe
BQeqlehkErl6S48xKjlrI5EOoHG5d7sQAGDBy70jC4gJq/vXvjV9FBJR6jn0x0Ra7bD8Xh+zge0X
4GBNx2TUUqYXAFrAtaly0nO05N67yeWeaN+QpppSHandMECNP3exfhEeuV0RpgFRFKNk+1xli9Jq
Yes8CrKL4KfOmUz1FRc5nLmrd1lWS0FUCkz40KZLx81AMJx5ZhQPsPzs/uJxDkY8P7hlp8okZjX0
IUeDJSe4HLdqp7iJBXBYPn7VkEWPjr1oSumWLFTcpaj9ORD4OgxMk/NaRgeFXc+bENs9EkTpzgX6
yfbB8uigTJrWNw2NBi8HSnN85wd4LwjqfiiSMJzDTkiqulz2V2ieZerrEXIVuK+0Aud3KN01GN4Y
9x0cdXg6MjKaVZKFYZW/Tq9lXIgUcW1322cfnkiwKvtoEGEaKYF2hVdC48WpclvS0fwp/9JrlLDz
N31odSca0JHMlJqvDWVbRSEv1jWtaPPPOcJ9CtodTabFazMc1/sI1lxcPNqT5NqkxymB7sVXMQ0l
z6OA2z5vn/W4ZjKbzlMBO95dqk9jEJwci60RRTDAJqvbxgPA1tLdEcNH0kiCXxKAxTXE4ywPw7rf
haUPOQnIOrIJmf4coDcWO9evGeqw+aTlQaPHMHRUz7wGSETL8CeTSpD+SyV6YVM5uVrIZa2s2JWK
P3dCUlyZgkqaozVv7lwFk0Y9/JxEhQm1JsMj/ZjsNctXgKb/VrM+2QjBZGbzP4zpqhhFY+nq11F/
Yqy7/r6dlNE4nB1ODaut08twX80ydQ1YktfERxFKwgUXsZSghwsyjaJcjsJlXZglLc52Ip7P2uH1
2l5vu6Vt/yjWsnG0WKD16dx/qjcZfLGJ1qswdfwIljzhykcFyv0qR047uU0hz+vMFNqZt5W7HdmR
hiPC0CcjGmKt3faeSmnYkkqdmXKu6I6oicobOnYEr2Fcw3Pb9vnKkJMnqTyAEneV2bDfcu2sWSz/
A0qXwMuFQtZr0vzbkIy5l3qyBr+3SPfX3TaKyzlIqUikFh/Stlo0sKdt/RtItiNDQfvdDvOvlhrL
zPDZoFsyid6FiMJ+B+lGcfz41zp1h/KzhLQo2Tm3UtiGglXdyiDLH1Kgza5cQpw7QRDxjtg/PLj0
ju97bJXHjOGKI4AX1qfb48MffxgdyzhztkYeYz3fPvm0wtG6XwiiDMhr76QcUAlHl066zBevwCoi
4mnn4Zhh2pkSxPROZpqE8gEawUmJLJZ82+2jPnntEah3jZxjo1YfrTGRgE/hnGe5942RiGWsAEt0
z7lG3NMAY35IizUf4FI/5Hb57M/QgBfB0vM6k3PcymeXr79UQVZuaz2F0TWJecoU9mT3mfEto8Ra
VxkPYf2//LgbrANuflOtmoCDoQTgMoy3zTYpCyu6S93VFbJvBrFLLjzMOPTnnccPOwFWgSH7/6rF
pwKstbOh06IKi3FUeSfcDdwb/gIS+ZpRsdo6SzTzf7j6LslCv/6ZZXktAnoC0JgzkxQLgi8OY1lX
d4toJzalKl45uznZeok2gbQw2iXRYV+qH9GxPFRq+Yas0z6Df1wCIyyJLCRXvLH5ypdxDJeJyH3f
KPA73upcU4URQ2lCa/bstZOHVxrSxNfxhHdu2erizqBT72RfbZiiLvudrKEWwEljgpycklBo/CrY
iBP7DHURJmphlM/xNTO/McK5VPCH1qYkXYmR9nd8rMXhceKAWrP5jGBzpWNT3GFIkTKqlXjiEZtY
qqXavhIzxnVChiTyBYMRRDc0in2oV8IvzoEqGYIdQBeQL9uXPrTpcAlVtWs3H8v9Z15L89rsiGOy
wOnJMg1tWMGlNoiT4UUkEXxMhL4mc5F9de2u/erIf0aQsubl8oOHG2UYCW2bmZIXYpq5QlJWqf+J
GcO7NvstnVOubKJbo7EoJu4MaTJGV0XJGWZeY2ZFA4gSlU1pPaU6HTbSkFwUWKvS/agRTZTaJQQb
kUEAau3YX/sKiAhKeH7wNs/Cmxb1NsXOBLKMZMjh4BOkb64vd/hox4+Ln6OxrFiVY0IalbCiJaJR
2BcHeq3KNj7mr8nzXBltHKjIz+NtYAUnDBbNai8FNpkpatqGzb4AxbZm/UH2kyQ+Xci4uokukHRi
8If7PeYIQaEwAx9Z4dEbwbRHi7b3dgPZdscpGuLIGx8l9uPz6th72fRGzqDRJ5IInSgElX+o7Iav
vaovieqeIPMnHfmFtDIWQv3lFmcNj5eeYasdMXQOJqAh2XXKJ5coPTXF3OR9uD1g02KOt5pAvS3R
EwOH6ifRZnSngb5dVGMcBZMkbnOJWVGM0cJyEWVHfPf4M9f5WbydBQxfznZMHFhytzjI/CLJHw7e
gltKV8KiYpTL2P0G0ARFSS2FxTuSBKyiCjCe0+PXIa8SfSTBrStuCVtkWo8JeWztlzzTlzPMrD/k
/MXolLYkMd/68JSI8XI6PSs2ppoYj4SEaqTOgQ7kVkDemhm2C5aYL8CPcbrwwSsg5GEfUFDy0z8L
2mjppc3J9ry2ni/sjeBFJccDvwEnqUsu58JC0pnbresiCXwzDV+P2q7D+JLmZj9O/MCVVd0KGoUZ
jfyAEzhdJqxEyr/yh4v4iQbUcA7MpWNy74ILjQqo6P5ROFdKlfANpHPBzlRgPTXgbUkDuHsQT5Kx
PqTaQxHRaX7jEd0hn0V3PLpytpyKksJDs8LSo6Sf01rEyJ3IKbHc0LOdyGXMyKHn0P7ZkYYvnHe9
7JvwQR4nYlbxGKPnWGboA3Ar+xB3t8CX2Z5AtOUalomEqXlr5U4kpgbcMt9KxolnDr03YIJxTLrk
+qINhIZavYfsKu9pGYraKBGZbxkG7HEzrHUamstj/i1sYU9UueXwLOAmDi4JrDjZEd6RN+ju22L7
3ZC+YNbTD9n/J9nsK/Yszgyqg84voAgdEEPQaA8N+5KwG5vt+rORbFWDKHhQVIWl2e4pCERhmzqh
axVz8lv6Uzvbos5mw9YAW9viDJJV/OGGo/33rvb3AuuOKcRvRxdQTf9+SYNEdpCC3AVUqsUWGCx1
KIky/EL0Q9R7sBNVHZlKdT2EYFeJMcnpNfBiToYD4N41taAMFmo6mndEEuh8ZMVzjrcykBcxBclM
Xs3p71/bDRSWVZDKSeJXsNa8/yikF7QSyRZz79uNWW7sL/iqHjo7IBlHq7wP4ySm2FkLQ4GZm3fR
4Ahchme4Rf1i7CQ63l6ONxhy1AstbxM/CS4URtSwnhgTNcW2/mGR+9JOgvqataHIPtS+ZYOsVauz
TmyahkzYJiQRHNlA4j3Dvu51UYMCM2rZjXAo6/woQV+GwHq7QqGRXZRfdQssme5aKxUYFFj6PvNe
vrsVRAEbaD9q2c3cY4V994YlrV+LvIbKLJ1nRFFVYD4QtekQOlMevZL7HOBAzWTmTsNb173umXQ4
Vzibuhjnns2DhMCwKQcIdgobUgLQPJfB92xZrTE1Lb8o3JEahcDGoutBGnnVAVeL1cuAPBVg1MVH
9xjswKQCr91+0FWbv31URxade8JTXPesWCVy5elNcffhIsrAAqhKXpxLlFpXoHtHxTDB31WbEmAT
THYmNF5eQ+BCMREX3GIJh9KJHV0JXWBvABKSgv3k66C1lLJakDPvPPVKgHt/5vLDWGC8jrA7I/lT
BDLYEcBS8n0W7mAf+uiMf8+qAyaC0WQ/tg6/gNmnN9oV1UN4Khea3sqHKlwHzNS3NFlMh4KXAe+r
CT0E7tfYWNh7oZbpRi5ucNKTVGN0ruoPqAAUuqw696RWTE7F7kLUn++VgHsEX8ltjaOJn2fHZvmz
GTRg01VRv4Qf774IFAOARz1l4WlUlKU/ztDULUZcZ3E7kSps3Rk3BSCk/CUcJmUyV0Hvx2iKN/KO
de1A5OdoU35N4T+zVOL8XlLa8jpU4RYPXlJ76g/g27xYhiSm3LC7WWJR7HCpSWFi0uOEETLnqRNe
LkpJzhLyjiAh7xNLmKBpJdqkD4g98OYBucGlGoNvxmfLuSu5bEiNuLJF8VsxidxSOW5FMkyh74G+
K2nZcU/px1aMBbpHjQYw+Vc7fLT32BnlI5BZX+qExFK+1tiWJmjn4JwFOUa2SOwmp/nTzVzDX1qK
9Fqe6FWTSRmiWch9AesRrdy/BeH+aN1NPBmU5KoML3C0Ojx6crNDS6RlrY6z/MKOU8he1iORdLY9
mxPNvN/27+RTZ3tgAv7L0VlpDoIrQkbXwvOVwa8Fck/QAmtAdKF/EGoAFaAJEIaRpnZcmwERhYV3
rgCRSRTQka7ycbWbSQdr2UFNmPmuyF7Kxe64gse91wj+W4JVxneCXWtMEEqTimLKCdugD1DBZ0xc
hF/7vOs3+KMhQFhSRXU1urT0KLKaZ9EnrNIJi+zK7nCsCuyMevQGbM3wYha6yW7cJVEEBZyrDhgg
R+lEBlFg/6CT3553iHjgu/aWNCZUCqW1acuz8RMbfYFhe7oLOW2OHH0SV1hf9IAobiYVjwleUhx4
PvADOZqqnnQxrsxEnR7AonDMUIlL7DF1rKNa9Tvyr2z+6S9uB9t/cXshNUfSNoSU/Q/gnyMqHDzu
hxqEwaBJv83PlJGnA1adERgXHSvHotxh+306g7b9RKgxHHrcsfWoV/lv49in2bOCo4zrz7zX6g59
xh7kagssJTlNqg7b67gp7g2F7fS5U4YwN+mVweIDF6NLzHmW0Kew/UmC4qJl3wxBe4hHdb3qihY3
pvAoCRgMWv8ZQzbouMheXS/4DpqfSlRaPj0IkpCybUn1650o8LEwPM4SNwLy6QQhqPjYLQX/FZ1m
lVRPAOmL2Juke2N4kPDP0rTvSr3i71GAxcfOgXL0TMD9qJCoqXz5BBDJ1AM+GAlSQMJcAzI0Kjfz
HZHA2Wy/wBb9MOFg/0SR9eKeqxOTbjGkJO0T6PNv9oEmfrZG9ojv6V6HsowUBosryAWRJvS38JO6
WrTwB+AYCQxhAFq6h7wWsGAFXdESJQrTHMQGjxlJ0GwBMnf2JM3UD+hOhgtVmH3uS/JzWJaO4tqM
ZBDErYD5NY/paqng5Gso7icGDdnrN3WQ5AU/sQi3GMQWiWwWnM3igc0x1McCO7iG9SA/f/E3qhVQ
l1JrTkQqaOUCChG+9Eptj8fGgC3ro3uWcePWdmKK7wVIe9h1UxvTjDl7y5/Dh8p3vKeeDy1QRdYh
MGG3fCl7LLheJoSkWCGQY33DvXo0by/Br/gnRt4GKk7MYCg0Ts5bB842v+myYJABi/wgZvIk7CVS
xpSosiHJfY41BWxAjjfAvGzbcKlD1w6mTW1hQj13zeiwY4jbvzmaRzomdebPdc/s8XAVhSKccsHK
ucfmIV0M8+MZPIspzPGOh5qhvmwrdyh3KNZw/6xsWe/4yuIVddONJcAR9uyssv/i3dSPjc4kciyy
vqVcGxgpoL/FKHic+Q5pyPcAvKteZNSWYbQz3Mv7wXGtf3EKrx2GlAuLxyTMwNMS0yVEtkKg/f0R
evYhcAWHBcPaMTKwRzECNn4Sm4YIyyauy9WD+h1lJtRsy/fhmJ3ONB8HOTqmaVyICVb2xLCrecwx
FS+k2IktSc8567Xi80GuzVNnqqbVPrOwkXVhjDlj50s06N3gRq4Oj/KIDnMm65Tk58ih++du3+YA
rPEAknEOVmWFn9YKZJHqzqdOUhssY2YGh9E24Qu2C0PQFHxhfjYb9/CFLWhG/G93H3GZEFt/9ep+
mE/wCGX/nk62YKzM7Qe+MKt42r+0GFjzrppGyZzc23YoKejuXABKRVq+/MWHx4oWJI9AFa7wIjWL
tjtJzTtzJV5mleASBBX3QsV+lpfBnmAY57D9fspmMgj/b4L/tzFmugaXjdAb24Wlq5sXFATfKoKX
iuKq+lmSnvUIPM9MiLnIIsEkoW966jt33Ygl/9eXeU0srcQIwlYXDjdPpW6gDxjAFVydHVqIGre/
rjERrLVKIm7ZAsTy3SmsfRi4fvWToxKEuBfoBijC6mCB4LG5RsMg7Sg9MipE4i2Wlyxlj12CPV1e
sSMw3EeuZipVW359mDVe3u7xlD0aPkSwI0ZwrOJjDQ1CC+9j+aEPgTsNZcQVb8+DjBOIclujkRVF
t0ofivasEf7txRgT8QNPtP4lLfJVIh+1mj4pCDbjqU+kHkjtZA8zJTztuywdF74xKP1O2o4qGOc4
Fp3jo21u2JGwwTdN5FYlC6oDHbiSNbkTH+TknBjga+Ow7F3pyhQOxsGTTsVVsrLyPSHgdDCSKK2s
yFpzDLTahNWirFqfg2DoRcJnahgMi9p1ld+Ofs2A1ZoX3Suwnk1baI08Xdt9PY7iH4XsGzt8jyzl
FoXk12I9AErL1/n8qFZNH5xvYm8timS+gFN6lqtOhqlIrzEm6jvtpvtbRbJcVAAFLw55n4IF5ISw
6GkY4+DzHCOb1Qhh1C9sLrXUejEMUh1heWVaJ+F6A7+aOMQZRRNg7OF/vN5ybg35wY9QCevkizCc
Hc8Nj45S1/8xsfTev4lyQ/igx12vQX2cwDISjUUc+TTK+ilEjKHmd4RJ5cBD4QCn4rv7l/L+8Kc6
jVoDBzQx8+LIxDf4nG8BC72UYtUC6JIiIvGFcj/5JW8y6VESzo+ErFmOjW/kWV1OHepAUGC/auto
Jj5vtEeW1p1j9wVEDJNlcilKTeAFsW40wlZeINMaoMEIKnxjyHYM8tLuBKiLVGo9rAvqVy/qfT1D
btW4HeAe56qp0l8mVM/KG0ZC7de7To6y8FRP0C9Wo9zK5hXII1JEQITpHkcwAa6v4BzgBLnYqMgz
OcCWsgtmhOfPPI2qEhOLAs7OGVRxw5dFZpApC6icCH66M0LhwNhipZ5b/tXrfGCpfNYsAPBh22js
jlGC+ESVfLFLPSeQc+XMhmsH/0bi/fmdwCsF+BBfcSNOUgkL+9ovro2xCSEl6qARUeH/m9Peoo5j
8I9NztaMgpF9NyqxX6Gk9/TFn0f0i0Ur3cPLrlMDeaN8+C1x7CNhUwxfYblHpYwmhbcuaCpctTMu
oFBs86BwVMepx7LBDBv0c1Qy1o5Xb6wlR7UpYC7pj9Za1UjILvoA00Xgb/ma5YSGbYqfqIoMDclb
OPdz8NghHT8ECcBkJxDZIqauj18bL5cg6OYUHrKMG7urd1k8DwO+xwzZ7RmfQD4WL3cHL60UUVvQ
Td7sPij9Lw7uTp/HiTNZG5ncPfLs62VH/y7WDbcZivyNM51KZaxQ3fmplSYXBC4DLeztdQNx5pxx
oPVUtPAZXl/38x11JvR4XPvO94dv+2/CxjUChP2oVw5qWnYuT5tRz9y+n/rhxQ5H64EDXNc9bt4C
AhBbg4zz6eYL/YDb2azZPqjPc0RgiEBbI/VIrmYc8aUe7o9X3VThkm8LiA75nNkylIZA5Yg/4F5D
/kSPvp79dABpk7FMjszLC396Zo8f1JdgZ4XN8eiOE5XH/zopfZixJnStdcDa+M+iiKKR/gwp3mPa
WdIG2343/T6G9OAHJOjHwe3bfX3fQGs+q0NFsZuT6W5OnLd/K5pIIhZ9SUF/rlFZ7s8rvK40Ejzo
998yVafTdC5uvNo/Kc70FtgcU2DW5O/ONZYQspnhfJ64WtZ+0QYhNeZf4NZ6EpP/sFRlySp7gWj7
oceEsiCt48zyNkStutVAWHvecwpvImbs8GljSY5rld27EWXxF1NqVUNkbU3yKqi10c2htYTvFPmA
WB2FA6C/0GwN41I52hbv7M4Kiz6SlnTfr1xj/tQ86m5REiPb2NNjMV3oJG8RYH2+dsstZIYGFq9I
JsQAIUwboFrD2ZUX5JtMhRjAzV4xKtEN0jJhYtuORpXcBq2PBOonhmO7m2Kjgq/sZAYfVHt74Dut
uZ8yovcdioyOwVdQmYX6nyBd+8aln1ceUrHZX3WeILFm5+kilavaUxH4wtb+i/ZGKAJ5xQVkjwXH
KkLsUKl42wPv1mC79YdYOLyG0HTHxYBneTzcMqSoUZKQz3zTFj1TvzMlWAT2ENRvfocEUkIbIncl
O4MVgJH5LkZx5B8hnCzx3ls4IFvzKIcd+8f6HusJc6AxvdOOX25Tmn2bYPg9hl8X8FDpibXO7xvz
q5HEedIN8oTR37DZlt+ywqiqz8blTznxPn84w8u8+zOCx08VwibxzmdE+4+qa8NTYkuD9GboLBC7
l8Y8NxsvvQXUnZtShrIaT6MG8girJpejukMjLcp101+gVTQwP3rI821xsx7DZtGpl8IVpOAryhoG
+c5u/OXcJgUAv6Blhn6D/2Sv0QKMSTYqDrj/IBIX3Rl6VJkD/7ZMhWmLjR31hTlaWPWon4+UggxO
q3e7vCNVKq5e0j//DxOWYc0Pt3l9qrPzZMVv9+rwytugELgcFyQpE0bdQDAV/hCavA5FGaX3s5Xj
p3ulxd491qh9MpvuBk4N/Dx1VbWoPkaQzSFI17P6WlysYzv5QPy/XNyTswGWuk13mSNVAN9i3SBj
yZvOekr38uKAUL9o0pAcLL5qqaZVZROjnISS026bH9Wkvnu45oW1pK1vneSl000sVfU12o9li0zn
07v3aMuodVdzRkJ/6y0FEPQmB4wHXivG+2TzrgSXQCHreZaM5uGaR/ljfqTSahX1kOuBwfPmp2GS
TGXKFJEJCYrXjzxnY7Aq8/sbYOoUsxs82dksxxEoajsWXOZbORHhCs1nTtEJrkfs7ZG7BoI/V8e2
gLWj6iKghZkWBAtT4Tilu0tZS5otkk8TaZAJwETgb+LEsoR9VF4V5Q5XF7yRQoZe7IMPszSiEl22
xeiAVj3ceBlhiLsosDxgYOBEML0L2RUgQp5dlCwcFhdPseYwY5WIhzClT6uNqClK/lC62m5ZUoc7
9ITHdHYOhyM58CCn5mNPA43MxopYNz4BiLiKNs+xRNnXE0ImgoWghMZlzBbjw+doOrRZC/XLF/VC
CrD0y2knYbN0g30gfK1E3Tk4xCdoXgLnL0WhWhkAio9k5X2pkox48o9R1OgwpBUnQbHEpcEVv25h
6Q6u4rVxNp23h48RH220AYH9Hc7F93y1GK1wUxl1pscd651/3KALU13GQjeWkFOOn1nmRq0gRnyL
dR7ZYgMcajNG+jhbwicv5nhkP49qVNoV00B6hi5K715oxkIFUMrWALq5sJC9Q9iNkFeQivd0v2OV
hYbsI+1pgXkiZNfWvpYowul5aS1Yh/8JL2y5WaU1b6BMtJr3Yo4Py+9rSPkDDqiBHgIt9k5pNEvE
ADQGMkMMtP+Jxzt5zvehGubd5Fpvz6dKBNDfVpmRj8QEtj83TTTyPKNd/MFGG4Er3LqNLSMM49xm
E7oie1icvyzTf1XHVxvb+NFOrXHtbbXoJ9Fw7QiwcuaOsHqf7DzXi/hjzKYo4kED1SKKTRq/ZanX
QR6Ppp+1g4h0zK3q0LalK4/aYa8bTvCzXhlny6DAhlH0CX8AdSxgnC/LF0TIrBPyLeNk3QWo0A0j
hvfiOksPqWxnG1RLMtf4ge81ToHamzcf2Aa4Ainpwvn8QSucs3YE51eEvqgh57eXTJzFzUeTHRVm
EuUwyiA8dEh2NrEoJ7ipG1HtyiNY5O4svBbXDRGMZi1UF2DgnxhDyYoVP3mYlwV+MVhDx4thMake
cDsztA/u3yEqY1ikmvP7Bl4jIYvuVDGBhfAZxGdRLHNPfGrO7hHSsvDewhi/wE5J3NNPFHdskdx5
IkLVruVRDieHUt1X6KCXMdYI1qtgTb3KdRofoLO7uv1KnMOo3kAJMalC6D4/PF4xNpsrHmIpCcT6
N7YNTxRy3EDrq29o5GW/olJ4Bw0BxCn5tmLziEiO7reSKsKNf15RSZGfluq5hnb/TjgW9l7eeT2y
vxAtQ6OZ4Sml8RukJJzoZjShySZnOhhv7YGE7lAoMcJBuXviUD+NCkrzidj8tQvDY5cO4nsxyUg9
qiTLW5Mlu6JeVTDOiqnx62LWGeu0EhQLpsv15v81u4bXqp1e3iZDGNwJgcDFGJ1r5lsJ+frYSoG3
6JK7yfsEKzJgQkAjxFmb2L0oUKifao9aZ3eqPnsIVraKDRM/fleZ739i886IUWTOBPPh6ikV5cmN
cZIbpJ6VAa5HL/OP39pepCBcu/PukPAGIkYEHIxECVCMvdXo/a0WtiBHyzNN9iMCF80scVtj1TQq
E68Azez5q/Tjcf9y7YeiQRDscP0g9YtB4Bwx4RDlxYYUJVtfGYd6oRuqxcXvXkc/hDaCysWQj4DJ
JlPLzrbcow/FbZz1l7LFrOscrAI4UUtSKSaELN7RuRBop2RQbwHYTGVkLbib2ZpJ2WPTyZvgGCJc
7GtCwfhGReRYL4crdl6Yx3dDYCgJFKe0mc/S9Jl5dUqHFNq0joPDlFbvGTLO0SDQvwluuhlV0QLX
nFAkxQ91ShTXzEFpXhNofp9hHGwS4QFnvjt+fOZFueS0f9MY5WrTyogUoyLt6fRu1qX0f6R6kZOI
Pg6cTx72SI8j3ZIpdA1gMp47OUFXS5n+hljt3KZLqof3HXKwZHUV8BCThY3o17lCwvvLPalg149v
1U4r466TrwZorPwLYDUpz8UNmQ8Vxg0rEpU55bFGzFlybiAeAzZnvkKElbKS2wfspYYi8hMFU12s
cbFlnVm45Dt3d61Dqe4B+z/9j2VCf08K/0aMpyknNBD6Zded3HRnHrTpn7fhKIyw0HPosaGuQps6
jErt2Vw5omCrIZg+D6BpJX591yeHZlDJoX/gptbYm2PC4YgEiH8Q2W4zeeA8IGKbzDvvtoAcgIJv
dxfiasIG5nmYxGIg6ReGhRaKfgKqUHBLr+KORafwGOJocLGB6vFt+x1wavPqRryOthkhHFCCRQvX
dUbCnGG1qfr3f7VMf+i6InkCGuta0uL0OrzWQByHKLEyq0peYorIgZRufJ+OBZXaO1H7vnxrv9Zb
skvjtMwV/ktOaHq/CQL39pqXbTrXmKfw0ckmsUxJwcPcAGiRn/meFL70ns8KLk9sR9E3dBEM7Ryj
poh/gJnBIcj5HhWWKC2m85OtDwcM7a5agVi83XP+len8ioe7r/PgK47YdmZCWnTu4lxUOW9E8qw5
YiB4BO0yjjrUpxpi+J8iB6SiYYqY1Avfou4s6bFoOmrdA1gk12AV0APkVNNIfwA461rBlXaEC+35
hvI0F34UvBL4F4a61kaq5/tSrMdGwiwjvLQJv25zLOn4Z00eu3l1P9ePqKyWviEYc0x4mJ04vv3H
Sv0eVpGX2nR8FChQgnruTbiwvBNSPFF8sQUCOvGvoTZT9Gn6/k7p6lUwh0oO06cDnmZHDohFY+bN
sO0XM1qP88YI9+G5Y+dEsPSkJoFD4CybebgfnGGlCKbdmY+thVbolUH1idzeCWb6poSu5s4KRy1F
4MNF9SkmFqm7bxWzQYxbU/Lk+841GT+IykKXmG95Lo22iPDoUqsy5eLWdOohJozFDK95TnMKcY6Z
03Ack5Mc7LCGYoFbpJUSfsCAKHiPsQz396O/5FbH1lgeA+14VSvsUWd7iAgSNFcv9CekCdsLBueS
8TgVaXmIzds4j8qWEbu3PIs4JXfvVuNnord6kq0GC25Fkw/7ICSh77MuWWdMnfbu/E9a2gh1f/eX
Qh+3S0KRqtgZU3vzI558WCWDZoHTf6RevI1bInGb0ajQrY3ctekZ5t+eCBGCy4expB2zITJY8L9W
cJber9O8k7A/jBaD9ohtBXh5wm+p1KfnQWTwh2JyVUqLyxYm7QPxlSGdbN8SyotVVTQzFbnYWcOZ
IF0BIRLi5e+RrbdkxRbc6DyyyvEQ8oipR7ibXekKd6Bgphx8BAC9GqWZHMbRlkhTQNN6ZNcW9+Fi
DS4m+AuuCktl7Qfw+miLHN+NajLuBk1SqptBZka8UdbQb6zXedU4Xwyagpnc/Ztz4zbCocY3wBs9
vYp9Zd1wte3xa+vbyM3AM41ljk2rZwSHgTHAiPnbfEVTXjDiEQyGnlFAGeFyvM7/QZ4hVXUDYxU+
b/TAhOzQ5qBsqSfzAVzzZVs1x6WXHqWLO1vTZyXtALBuxJYKf5ktSfmfU06D21nHEV7dFq6aYHXP
O2zFI2zEuarmg8eGb4Dnq6BuNL1awWTq3ejqRWqKkSebv5gSuQhm+Zoe//vuXrmA5h1p15cO5HSG
b9IFmK4g+vihBemTuNOFYf3kk+Btg6BxU9LI6wHY+CegoD36boPWGpjqfS/OFfV0Fqe8b4P6VB46
GKySBoL1qByKwzkPOXuhUZilPlg1CL/q7dhprY0mJlUf1Gi3x3PFqOXXXMf61ai2pVKoQ2y8qVHX
CbpB/IptXXIqAEVCg+O1q5CVaRR4HBhDjZ+f1x+ZutwLWCqMbjsCRkWcIETB2n4oLTUranOy9an9
CiAvHmCWPe/ieCaQlprA35o0sC0XECHnviXj7R9M+vR61v+Ms224IGUSxxxzweBn1rhNNM4ch/CC
af66ETVmKqEAaNcwtTy0rDwGZPPr6sYzQbX2QhtfyHggkcakx/UfJlvKRyKy6trb56v/2qFpsnWD
aA6t1/rgPxycc2HW6/t3uf2rFxOboxnNXU/nY33qZRtG8vP8YZ+HuEt9oI8N0G0WBIzZ/7V/pkNT
zXtAPDYT422lW7EKIX8Qmk2L56f8TSOG9yyxKBYIJs+p/OMJbogtI6w7rPPptRhGSTGZw/44VOs8
2jddDCgN9aeRDyrLmaFKK/Tx82TGpe+OOk2pQLowB2iy3FI3bQy6Qbe+jjAHBaZVFbT4ElVCKx/s
EjwUde4+m5UINvhDC4QM7Y8f72Q8CWSnFQjGQY/bUHxqCODcO2yMbj52pKUvEnMiTpgAD9q51Lsk
1blKpGHpq6oJRrB7708X4JIp5kSH2+sykdCR79BFccbe+nU0kj0+hHToToZW6UP/2MJtgJjxRn64
U4WHcE/ZR1vJLXthrV8ray6GCV5BUj6a0NpY/GrsGH+OVjEsqVwVkEFg01P3cbjdoNOuLt2xyt4k
IZhUobphtopgUFj2m9beCndsYXhM6gHqXnuJhF8dV7QudIAxpWZ5kY0E19FIHJYeJWy5T5r1NftR
7n59/o2nXiipas4OQUH4DqdA53DkUQoxAdV2n4W+eX+XZK1a8QQs+exMbvGIVnYvECfJgz/dL4pa
hxbw+n89WoH6RpWa/mDA8FhlKBKW+LLiIRVBombvn99fwp/aKs+CQh09W4zwHU181s1H/l5/wB3B
ax3bKmW3R4sYK0unT3cAa/9P+AIKsmarERzbF/T32fMo8O/pQLRIK3w7MYpTuhgEmSG5ww3eFRsG
lL6vSIGs6zvVveSqHBWK3EZOEtKvlIf7o2P/FwiY5sDBeqbcdUwUyF/v88G5Dnbk78wrBpIeu00o
tUvU6dBy1Y7V9+ZA0hPOkajFStgNKwHeXgQkAHlsSnd86QIzB9YJ/+tIu8Cw7Z7qcfLSjjZ+HEE/
e4+pQYNMAhqKR9UwuDwXqjC5dhe4qzaCeNR29l75rNKRi0p5eRInJmLGAlMnH1L58Lb3tGObTw8p
Y93FtbJ71VLosOwdk8GnDzhi5ppGrNUqH6cvNcJbNG11g37TfrLJKV49wZzPpP9vppz9zGKQkLKO
c+POr3tvnKNQBknaOxKDYdjSgzXNoogxiIRA2xiUf3qvZgmcftKd3Uz5zkaVH3olCe+dNco60yzH
J3PQ/hdVkRO5HGEY2nM5Q1taEqzvZXTdUAWqfK1E20oBsFCg3mGc5L+RVLWrz0bsZjuxrZ0qGjVX
n1fEAm5435O9cieeqYA90G6vo9h/bic4fnRtu7FS3DY/c2opr9Klj+9UEv8YFLPn2ptK0tx8Ua6T
Ljq721MMOEJeqMrbMqJqZ+Ua0cb45tWPA0AiJfaKsQfilHEzs3TO429Jfx6/Us7fUDkJ0Sl8CN0n
HTM/v/x5nmhy9xZHZ7EzQVwCgevr9SeeWMySe9EVfPEqmDEwnZEUoo067NUc9bPFHh7RI/wl0tN4
YNIhwDlXibovnl6gbadsUPcxXOmH6SXAQVcn6qdPjMVeDaqoDmRHh7b+7rYFhunxkD8z99gUe6bf
JlIFN2OMsVLn8n5mkT6ewxoo64+VN9jTW1n5HC/ylJEWw8J8smOlfKYzpPY8x5cJKyfBHWqvS3Nb
pQKAFY34Raiio0v4J27U0Avt4s51IGOnNhfgHA8bzhy/z+lJ3LWc8WI5A37nrhF+q9mCfexTjo7i
BVUANzalo7l2ZrtJE1FJ0ki3tGTVSaehZJYm7kE+t5U799GzZfFDjY8FuGtB/giyc3c1thohpmCa
JR2thJfwb2iat8rK3GF+x944SDzCBq8Fk6C90Umhmz0kAUAQGW8YkjM85TQX8ODB/krs8gRm2WQ6
gpJFD14dtI+kbSE4/YgHPfcQdaj19chlBT4flqmSdUDg1uf1APF7nGkSxCV6OgErfsrHAPDZcXsj
7FfQeJJpinZhuqbM8h0986rRKnUdQX5HPnz16HiMNVNs97eaT79SM/MQt7u742yPTYHmfPn3s6NF
aJ/u0eyLEqQ5BHEHNf2p5/o5C3Ep/iJW5UL/dsZ7fb0Nb5CV925TTHzsQpjdXHowYo9z1zpFqQ3I
ITSrWa+Wvtibhn7k6WnTVFFtEX7I606xdHCvw0pucLsTyYAYRjlMYr2s0/IZXYmfN7cGZGWuWe+D
fBixgbEAR79hoRmGSlNdmVkyq89RCv6IL+3yuT6T1FNlGB2g5S0mT7dSFdS4aIj+WxZkjzITUZYc
zcZ1bAQxlWoRdNrKzy3C9diSKniyjt0eH/2gU1xhzKiT7V4KbZWQHfbhdgSQULC5b0RZORteTYgf
6bpiCX6WAGFJSJgdOoacGvqoGNnguq1IyIksgYWDa2Bt+4qqcz8R/LGXqYIu3eqvB6VYYtNQoGPl
KBEW8D321YP6BMXxgoXdyKpXHOdnBjT854aQJXwLgVufjAHF5SJL1ULc7WoOMVKpABGrkSy2mNug
sV27BDiEyDsufKMfA9Q1UUrGSBrL0VPhUlVqIzk08PfvZWB6ba9G+xa4cP0upbR7JnZT+JMHUU2H
xqCxvLazUjp+u3jt2PIsv/wdeQm15pZ3vjRHAR8OrAXktmgBz2mrFdgRRIvqG26ISn5+/UJGsvLA
VBk8POEvhhF0pAFEaYumaeKlbzuAQcR895vfGvqGrqQbzpEMHTX3Ob1wlMt4DHcQqlE3fpGB6Yy8
H9iTtI+mBAr05Ic+M0XK26/59w+ZdspygJGT+fy/+ELrD7c2JerXUkAojr1y37dKRymHjy5hE5lA
00wseeCQ5/hCJ9o/09Q/dzgeWszYcajgfmj0jbalEklITjW+v9p0BzOMb7NG3Gfdy4TakEq9bAWl
aAYagNYSJN6lpDg3EBBsRn4VhKRjkoQDVzaSCpxWgNOkfF0DAScLw1l7kSkFZqCEavpabYE0OG/g
m11ASDIpFgqquhHb3YZdkFvGnLK5DluQto9CLjGGcCrfsZi7IN9b5GagOyMXi5FuOwfx5afh2MB2
891B0bq3VooH2F2wwOgaHmJISJDjBL2k1Lmk46vZzEzq8GTqeVki8mvp+MEmQMVvXi30vpAw8x7L
GcxZDarKV6v8px6Hrae6EhlXKf3Mj5wpn4gA3dXiXAi1MSoa3R8PjghFkx1ntFMKocI2SQYgtnv4
XFeSvucKVENC6LOD3rtD/kRUhcNTsYGXy7LZhV2gq6IIkCHyFQ2DbaDMniwmJTgkZpd9W++c7Otx
5vL0eZ4Ar5ekMNoJKETAIfSw2L3+yqcPmWHq/DmcW8CG+PPUq+AHqtbN/oclqhhxjlGGb44T9nxb
7XjTwccBA836DGfTn1nq+igfw5LLn4XXeL7cCdcQsRt+ZrPpf6m1WentbLkP5ZHdwfrhND8wUb5h
FqFkbsy4df5pdMGbI6UMUpSEW/yl+V1596stointP84Z/aLIRn6lY5MqWGGa6dvBhVWRLuFyvCQJ
cuhLh8+Aw8MWag9cdXBvoGPDIkKW4e9Z49h8XLZGn98rNSrla//wuks5Qqb6fo3q7U3GfWMvTqnt
UE5PVnwKUB3rCm0CxU1W2EwRpkb/8ADRzM9XHsdDD12/XjugdX8fJ493zpME9fs0mlpgdBoud8+h
JETi4vmuw2cbnY6PpCUZarSeBwB9F/gDXB8qbJHzAvh7w+kUwq+kyHOZsYxNZLKX0w9UiT+zMpHB
l0gaY8H4MKMyv+wkU0k+7LVmpqBoVJE9OYfEOBpFf5yhzHcMliWrUkaFSSvx3Ot+QsQ1SCRwITWL
cCkxJvrNZU5wa2v5kYPhK/sRq57wxNwLGits80aPnCyyYl1DtBLjVMitL+JXmNy2bbVC5dOFpnqU
JCSaslEoGZ09Bs/7qsQZwXus0EhjD+Ic57vSK+L5Fvlc9LmHNwjfd5m/Cwpokx7/1vJiMFK8zBt0
UiS/qbz+9jnvXRV3+VrgWHgYGwXPMO9812NmximAGy0BiWYrplhqDYpnxJE7qqvNZp9AQyG2odN5
fUwcLPkVY29EGOF8Nmia0hXAeQAvKq/S8JOgTLCqosfE5XNylEwscg5y6RBm8FqfQXrgKEWiavTQ
T7IFRgStecojYUDva+w+gXX2O9UdqtcqqrmeKGG/PHT/dUINQTDieXIxr50m0zHobhMbJSaEGvwb
DdYNtzf5segV5l+FFyFO5XS1jdVg/a988/iBrtxDNTn4tH/IW5HRwoav+Cq3dI4+QM2ivFhdonw1
kVJTT8t/uO2bPTYp6kUA3cBMxwyRD+DDwbJA0R6pzrFgWjNVEstseOHKTTmH2sUE3bMEbWRFPr3c
W6ZZtHqKWgdQz4ERDvrx1vY+oJYsyJfpbFlKWdkaoEBsLSVRhEoZDGU/CwaTGnHfZkW9AJVNxFss
cHNuaf+ZMkXQXK9E2jXYC14q/5QFAdo0HNTC9dczVPzf7brDLMD8qWnbtMhDTNGzY4iFMuvcYfuu
c2ttXivYX9dgMe+FchhigEdE7HM/0SW8fyL99P3QrXfq9Nuo6945UccI8UxihZHA4NmdbmtPJQfR
RnmbcvFGYi9PbykP/YEaA6P2O9z3I+ddcL6REG9eu+MMsflNEZTpjlmmMpO2iQckyy8l8jPEqCws
P0cV2Jrw+2SpBvitZ+dizbRivtUCz5PMyd5qRvf1W0esqy3rdvHTXyOfUqqerqWiEtzApniQxGgb
DwM8mSnSfqcNnjzRjXOHq1Oi9vW8liZ6/DqC02vZ5TPFwid7RB/XZ/OGHkiO7TU0GstrDZyJa+ec
G/ejncDTB7+nogx41b9srNQewAhX9x6Bq5eVCXhzTdbzUl94tMBYX9Ld01D3mXHU5wbIO7ymXDTm
gUqwu3J7GRGHE29dqKlX+DwvLvXpikovMsEqqDEe0nWL4AZJ7XRbcZV7U/dAz1XjECrL3BQDxRfP
M5dnWlwQYiSK8AjuEoJ+YQiYQMM2V0IIHI4s6n9kBiOqS6hNqZE/IIjZWNqEZWFE02Bc05B9bnOZ
ShjDiptCqxhUxdSKqwXRt+tHg7h7xQ0R1IyvxuWE2gWw+3jNJIM1aTZJcTBvTxy5IV1VLPmXeA0o
kZoPvZ7y2m1oq7/JbmJU1KOsH82Fm1uCNfPkeHUDIfafyqBP9pA6M8jGCE70c5HlONPKkCFHBnZk
BiwIRsns/4BbE0FKcSgX7rIUeLBu0fdwmymv7rLIixyml0vb6i1LMfXmgtw52kHl3e0uApDWhQMZ
xbm2stvNONHZES+0TvuC3QOmkSHpHFVzAeJlTamr40PHLRy6YW/7jl9VvYnzrDzZ7BHeim5iX7rU
5VGUwot/DjfOAGAgFu03bh3GOey7/Mopt7EGLM+1FeOLv3KblLJRyuI5gsSA+73sMasqtQ/0HQ5k
x551zA41MZt0dhO3i7apfziKlLgO9EWGIhjZaYF+yNySSCXpp9ZOLNBGvTIi8xnVYBNRxdjqP98O
N1ZoV45fUQYR5Lan+KXHqGCwygtFlRqKPLEvxT27FaToMvXkzaydtZppFpVgMVZFc+74dhKjro4+
0sY49Lhh/LRSG6HhGw3fbZJV9i0vU/b0HF2D6B1Fnv7+XR/55t9TNxQkdIvtAuYIkM0+vkHVauag
3Uy3lpkPNqGjbUHczWRwwK1me2YV05vqeb78WiIbexan3vqpwikuWNu/DIosiTSurlRLcP1+GP/Y
FOrQn4QGlcJBVOkUHzzYu5TRO4iHLgjgAP4/T+JwUhZ0NLt6q2cJnIrmE7+Z3fisyfobB2TdTcxk
YuuMZEU68DtmGaClcVyJor5HS5ypDIsyT5uR/+E8gRaq3QZNxhsw2UHkH48FIkLKloEUuYAALqRj
dXvuVNmb8VY5YKUkgNMKoX/SdvLSgP1guLSfQgmeF23eMDtRtl6goRJytPiPbNNNuGrvyFhzYZYl
hVfwbbX7wohEVYskYE3YuCxNifpDHWwpDhTdKmMYpWlIdCtA5vY1pP8cTwpeR3roh1hCriZFurTD
3/3C/2LZOVcplFJU55Br7H9z6SdK6wRyunVa6aGj+pWujkQdnTOzRUX7Rxv/iK2/FH68XyAlVTQ3
Wh8m+5hHLcv9zrvGDdAWHN9OeIv6yfqxo1t7cbFI2R2OnirTWmWftrLcsuXpok35y5GVVb9K4jRg
rrzJ1F5fngE0a77xiYbTtTMiAAWQsuH2qtFqL4f0GmktAWfjmvDoAax8OhOJpDyBe84p1d2AqFyC
/Ue1FXMgLSFzPJDqcEKHkKPi1ANRHQVErh6iGQjJRiGN96PuTKcXcrgRuEf5nd5h3qoAdeQrC51x
ZUh0Y3aIT0bUdZ6yxo3vIMGTzl6lVr3jl70R6UgeTGO0wKFhwCMgw3VJJT/aiwjbMzOInBoeOeov
RU0jyzSFiYeW1zHgtYw4Iz0jmkYOhRejLcYnQaSgo5c7VJw6AhO5wNdkQyrMXygS+cLqbRsLqiJZ
ZX2sL1pHNzF0vcZ1zPiVUsDPm4jJxm47olgU837UnJgmyBCbxiE+lcQrzUHMp03yUGCwAV+o+fun
3n72g5xtciQCmYWTgw7hJNb9nF7MeThVUxMm+5Ar9lUobyy7cev8vuGjmpnX4dMJpxmc6yxmGHhj
EiJpkyUmvcStN6cj+tnJdxV0QayQTYk2gQ+iGQxuIEs8P4FJG7z5Bmpegha28Ir6LELenB/PevqE
IzaU6GJy+w42keapkC1GCskf+gaHK4GQN9sCVJf5AVFnzTpD+CF0SXDD5LcFfDozzrm3eSIQNew7
CEcJq1hBrKTeN27qseOjQaYKl6uyYqixJmp6MGYbQvO9jgwbOaBcF5xks09txMb9l4bKM5qG6zoa
KyAuvIU0gWqIx6uy42DPd7bMQVJh+/u9EXY/PPg2lO+snI6bQycspfZJHlUqLMtgAkDqcoFoFSRK
JqOBxphPyrZdP2UHp3vRrX7JRK9JPAf2y9V4SaXVgcn84xFqUNw/fO84F+yzByZW0GFEDKBQDVt7
f1xiRIDd5CAs0u5r77+6KbuTuuiNsT9H60b5TiDSjuPxXgjdixoD+N8zostF4DpWUoakAwENbiYU
2vO8jwxRDwCzzVGF4IYpl7XHpg7vhklmr+a6a7zMSkK+2fCllzlxG/sZbn71V6MEuOjlNaYe3SzO
HwbMGieDrJ2ZmTDGmZ1jczIF4IovkiucksHmy8I5AEJZsrnTOcKcyqZBZS0gu2MFYR8jThc3n7CM
b1RtobV2pu3NeGK4ohrgpodYdKYNiIdYendL9NVe51yCTFOevl95a0OLoQhvuKJRqH8SO3BXMhLe
kZwhdjNKHJ1UcjsdPzM2Oc2aWaS8Sfe0pmsaiRRwuu/P+m7VaDgV1anGtUXdv8+PA4IToRDLGx3D
3SAOibq0PZOsL5FPTFetos61QRQwAUgmOhL20uLSFfg4XQ5gHAfPUDFoVc/gD/f/bQr+vrFgJVRR
qzJ7EBew05P4DTfQ2kXUAAD/sVpgbi2nhaOoBJaRYck3/FvRpvVl0cTd0r/7YkyP4Zjo1pQUd3+w
9lUUHcBQZ84snzMPwWNoXKLElnn36DXbBGA9IU6gHEJ9cCiEnWu2k8WpER2/2wU3pRBTlrCKZvld
nn04dMEXU7Zt5Hr1E7JQErKUHCtYKzcBLyBaus9MvuouP2HzCVfLU9ohcKX6Un95zIMrLim2/16o
wCdtHTcApGmz7eWRQ6a8IQjyTiYyVtNBAL1RpW3bsJiOFvjsyXkKRbbHivUvH9JcflYAfpxQB2SL
NMBzPjwVUelqkxwBrLXkGBKEoFmUD9zP/u0FrVHWyDS+a+wjnquwUwrvCavRvtTiLmmxYGHnGHcu
VqvLG+b1HPZcKOViaqKbD4h+ohgznIW12kkiu/Qf8rYPIUjL78gfVy5SnXaaPXscmAF9JAxdo3iR
fs2UzUGwvMtjWGJqTd582QTebkFDGaJofnaG1W2p0y2lzzVgafTnqpvVJssNxVZuNvO7jdR2wx2e
lMTsTeueRqV16s1QkvhRBgilmV5DXsnI3EyzHA6JMQw+LiPTdNEWid0Qn51T/I93pfVmRJngF3kl
twYq2tlb2i6V2rcoMDZsLAs9D7wx38WkH/y3YU9hjTMv+SPLNXoxfLH/IyKFbQa1b5RCHZ9eFJHU
a/6VXTeiT/zLox8+O5z1CCaam+Iu4t/k4PLKcG2EyoPR3yjNKJifCYGRAqzsHxP/D+yXUaleIP9S
bo50wjOxVHVKahRsa7aELbVaN9Dq/b5Os3GEoo5WMaBEHNHExZEHVvEOQKT/+TDaRmee4Vq1lrCK
9VViA7fqJZPbfrhxXIOh6px6ndyw5b9kdinR+ywRRDdZKBr9T+3pRGdTqv8yzWxUH57eIIruTFmr
MsvKPwVEeSWmlW1XogyOf+RRcEp9z8MRoYbrfj9r16s8B7pZgoOKwuys/8fyPnH6YsI4BT0I+Bqw
PR3aseG38fH74seO6bW7Zw8Z2jNRI9GOFU3gh9GTE1Lcx9L1UcuC3QXzHIGxlWEXbygXxVtl/TY/
KoMX0PB5HNnb7qIr+ji11GjUtqSv1cIFYPkyGKseB2DXT+LMOWktsFbeJxKPjzL2ZqtoIYZMsJuo
7KX3LHF3wMN/McFWEUPVXuIuMI0bdOy5lTqBTUyB/CZIHAIv2PlUHmyKus9O6k0W/kLn/aYX5h2M
1QccuB4gJxQ6M5MZSSuh+eRreSb8GpG3h4itHBjv3cfaVskqLTwcrReXvgp5vQI0oq4giI8yYbB/
EfqQh/xAq3BbS9fS5Fxl12gsvjL0JiFuXl+jMjHjRISch99Ts9YP/Bv96yRbIcuOijVg5axuUaDX
pysHNtj7rdPh301nl/ann2J7rVPns6j8CqiUnN0WJS9URict6AoF6TtSnhYf/sGdb+2wKhM6JPn6
1ALLfuCKTpOTOA6neDls1XXi7aOkokxfH2dS8RxXgH2UBI2fKAIw/UH9tpNdJc9bBiohf/D63M1s
cpic62+X82ZVRUXyTRMoUlU1OaUfmX5uanSnUHhQmLregLaUPCXvZAQhKsNsXMRlrrupmtRGd+4y
0abB2R4s7ezL4+Wyf5PE9cFpGtzqpVJyusS0POIx7K9hqFMI31HFFQaIlqTqzHvm16yUTg8qZDAw
kbYaqp0IrqBzZ6PamBWQH8D7qdN6RNcjReelWfe6oDcD6m53i8C1S5vcnQE4vj4NozCJD39mmzOs
LHe9v4QlrcVxs1yIDL4CFPABiioMdYdUoECuSUqY371bZzGZWZ8TFbYgpnjRcz+Rf8HqIo1oLqc4
qPzHAkacl2eTv+vH+I13mDnPG722FF4Grtz2982aK11kI4U6P2lyLXjMpRn1Q0mWB4U/2MCK9XjK
6hIJQ0/KWRs9tA8D0+JpuYjY1mERac/G2A5De2Q2ufue7hrxYLyIwhAfRoZsdBlNkHCWJ2GoXAWU
yxIbJROcHrPxSRH8Nhvb9y6jIJhj/axYFzd6a77Fv1aYDCe0C4F/LIq7yk+5m2eZXf+AYCxEl2Xx
eqn3JP2fK/obZmLKs4aiEV6joU4jOWOnWwPJDXcNqBf8NOj30pROJVVNq8IjyRO0WQJMcMSWpO20
3rjHzUZB1//QTpgkUVsFZn56LfKxadgH2lLvhsfXX5iLBj1yaCNIoz5OGarSjUAHXfQDiaLZNWiT
Jigl5ZOV9E/wG6Bj9bo0hLxnYLn94pejp9NLWGY8mIeqgs8lzHSsMvAK82L63rq1lP1ePoTl4XLo
YXVX/0DmblC+oVpcNBlkfvpFjQWj1lgYRDDPIVr9i7pom11GSs3yMEbihPKuJ10XpO+uBpJl88mC
YBkaWYPTB5cRNfuv7UQUwZrut1spPjqKkYCj0zSmyJ7wP36UetKLnVkP4KIqLlicDVIG5h3HB7gV
tUIDoJsUmwXySuUuBogS4SV+Wv8oHu21NzRQgqRVpqWYBJBTI9fSCDZrNnz0itK6xd8Hjdg5hFAO
hWpDybImI/7h55OmBPeAc7KtV4ykSeys6TdEWrPuMOUIGpCXE9HtCegadAe/gdG05hjRmwvuAhXH
3nrBXWkxqwRL7iedaui0V9fkpPCc/y5p4tzc6i/uKjJmu0WhVwmngAqWT7Moqe6Ql2DKRx9V7VQ3
DiXYX+QCZceJbGU/rv7KyBcj+yJWeSrfpZp6YuLOzxaxjVJ+rIIz+CgqJ+ehTrWmX0p0RB4EUCFq
gfPbJQ2PXJllOZn//17A6Bb8RXduVTdRQkf0OyE5RMgxF3gdFvL7lQwfUV0cFVLtM1Uqa4i7ArG7
Rw2bfb3qyjoPyGgWq/rLd6biGR0PMm6R2C7b12oPrZe+rAu9x8vSlBzlCXjaYDToqlAk8M1HKGTL
JNv+JxlazYDG5Psvli3uQPk3+OjSSPLulx2r9RZZIZjlIfzEuWcY4Zj/zlVXGIVsD/7paoco2LVV
0d0GClfBRKql3osy8TJOibZPXbvczgCzp+bTp0G2fX9OFr6bPkboU/vD4eTY4kstyq/kr20PXBPv
NxtamGQxGZ+MVbblD0qA7R07m5ZTPS7E3sXNnrYlIctskXQhLn0blBK7ZMdDi2174Ot0isyOXgd2
TzDoDUpGRgHXN6UWtvVvM7SxmnFrc8c824t17DuZna5E0zEsNCK9Bmak5ceywkXX7MSK/j0BFxNb
JpeZQc037Qve5ERhX+JWDGGjdvmd+4VSzShksQsBdI3sxuYCc4Kb8thwjN2M0LwVp1nOYE4/MPNv
j9KavnKBNmjbcBkauBXX9YUbCGOC8gWxLTZbKp0u2PwCHfhy4xXNHcXU1tkm8NoXnukwd4OJdLVA
KSFpIv/he4HN2rljHoX+pF0kkM5ocxD7Br08L9ZGvRMUfCw3vbxZDHzj7q2gp+3tfgz51C550EQz
lYa6WEukIOzXNKptyIBbVQs8PqkZN/Y+KAUT1yImmfvIe68hzZdwXsWE+PnEDuNmElDntJ8vmZ9W
ItrUwh+AN509LwFFCu0B++95Jl6oUCoH5Lxujn1ONDtOoESmmuWNilni0uiUcKBe+vfHHLRG/E4X
UnH0zKkzrKiZP9NbR9ptY+Nbd5UvI+Fz1uAhyXFRuBmabyHuxSjee2+Yi313hoyiuyslKdM4+rsv
88Do6tGWxi5/4BGJPhunTVN0/z5rSZTQBn38/GKpLXx9waD8d5D62SXZUKtnBrXAgrEDeFNlGoDG
GCjhSy9nrrVIpb4VutWGu3g72F9IWhjAFRIj20Ms9sLrpzsUPpw9wn2n2U1M5Y8w5wqupGpxHNp3
wCQjR2bg8ZqQKaRZaCsjcswGfWq+b+pfU9hNUknCw4X8HNet3siYy4w+1j+slQ8oa29l2cQzrSPP
MEgA/9k7mTWtAM7mNFNKRtA2VDqVnIEfjiYiBggTIKzyEjdPg+iqy+kWDS56as5xbLmWEjLPYQTS
Ra91s2dXge3zoLS2OQ7XsEw/3GcVe4+wKXNMf6o134eXyVIA/KdlHQ66mCou6s9T+VDWWgy9vWl+
yvOx7rKrSCZyYc1FPl5jTjY4nSF+7xtcHXE6AuVSqwRSQm+b0jKm0AIXlKeNY/dq1DedmuUDjhER
Z/DyHfar8aiX2dBt6JwqD9QeBAsTnXwFGkg2GgXMoPlMjKkk0SsfrwVq7H0gQQ5Swd+eWQs699Sl
XyIqp2Xkdx3SvoYOKyCADhzhOveupNgpnOmHUQomcxcbzhSz3t7RwGIJsF5LPWgMQvOfQqkmQ5t3
t0a+ExISdEFTHaQZ4JpCWgDlSwfaxfTm09jBm7a81pKpcjvlhVlOut/1KH/GvzeH3HfezGTLsJaB
Pj3S5EK1w2AhaBL3Qs7SJ6h3rsJEo4VVG+l7dIQtg0ITqQM/x53KAcgBFli9v/Bb+ush3IueYkUh
LinphKyGn8BbqoCYYXHZkgTm5oMSPlliRbogRwJdFCI6XLW121ep1wXOx3yWgAjYL1vSws0AsQva
ti1avjkVXkh+7N0K3bTzgmiLeEUVVbq1BZekHFkIiVs/NkHtI9g7vvnDm+KjRaC0wlj8lTWBwRs1
LJNEDKyhozR9UxHbaIS8im2ePewgUUdqqQNoehcWBRC2rBUiu6Va6rOocgStcWsiGzWTGB238c3W
zTHuzv70d7L0LX/xUwKI+Rq4Sa5UmGwMCNrAMYrTlmedHJPBHIomfUAamqQ88Gg4V+oudgH3XKP3
x4sB+qwW98tyiWR9kuy93lraKzADGmDBbzeAwRYJ/Hh25DSvCYW82U/fr+3rwLimXfhQhFnnegep
nnV4bDS8REjndC+h2E6tw8W8hlFUUddbGZ0UFGFW5Y8iIhvARnsW/PDSuEhcer2DFf8D5cxn5336
Y6Y9P1IgNI9deekrcKqImgEv0GNOaMtiJCO4K9qeGa+6kpnp9NF4wqvcaMAKW146nt2uXW9RjwEP
TX3Qe9reifGf6kzP4oCtXnTrgcH0MYFvX4QbYA6QxCOSRq/RL8VfzmA3u9iUkZj3561uLXqDchgU
YHSHjla18Lrfsm086ItMPongcygQN10Cz9Yb/rhICXdG9rWR73pLjoYRIytWakozvNW/phsyR/ZO
jaxUOvVEYSB7up1zYjvI+22QCGJXFtmiB6TDQVVYs70G0SRQ2fYiLzgU3kJazUqvtDiKZbAkkj66
qOr9hVBN1l9VLdOfRX0VASWdts3AlrMYx/YLinnkKV2xkMAv4mlV+TBOu7ug9RDV1n1DOMsvX9wG
qGO3Aj9BiF6dSxdvmWSZqfa2KPBymMoxWqzj7o7qAaOyV5bu5lzfX9DMMxNgQr38g2in8iEMm8EB
XUp1/rw81kq2LHOejkbcPgwDPfGP6OuE+OA+1IVaeRorL+TPKt9S4dKW28pr/2XHt6taLBr/h9Ir
Ln+seQJoErv24EXOHCxuPALM1XaZY01DZPRRJUIfQ2tUSE3dKV+PFKxAPkYUHtlgP5Y2JSX59GuK
/NjhJmC4fui3qTR3r1UB7bpHcIzsBmbu9zyc3Rhqp8eBnAcSSzUR4OY2btNeXL0Av2DPgoct77xt
FTByD11ALckYyIwEjjT5Sb5k3uj8kx0Ri59vUTqsnUCcbsCHn0OnC39yYadIf2nXw5jK+bIVX5I1
PKpuC1P9tx7GKhIbWQjAIky1+V51V+0nJTZpPXJ37L0zRhf/gpRNfiIH5i7Y1VVxQM/rGc12edyT
wSp0fiKLFoKVk+ZHDzAZmQauJCbRrDZMQP5I5rG5DhxR9WJeSfSC43t+W9wKFvPmUmSIZIfY2FAs
WXtVimCuMgMd32r0BTTQiREhtEjLFqwKhENJFlIQJri1Qy0nYtkaG1n0Uqh1zJzh3veuvy1HdQLy
NHwcRKtRVdE4wzJz1t4+EBILoII5IKoZO9PL7YnqLt9f4xUaf+iTuMphjXWrlnixT46WCBv82b8d
hIPVB9etwL6BRxCNEB1txT4evlzjxE+4EL36xmyWwpOwUaQZabWbeORylKw3S+gFhd8khyshjNm1
GzgjBWK+l6UaClJnXHX68cgzxYV+0AGi0o4NWqfR2pUhainGjxc1XGWP91YPAIrSWXMJxHLobaDt
8x/8cnVy9Ksm1wfgkZDLs4DXAKq4oblQJOt0ofnxQEvRsf1HljK6pD26g/MW+Y5q5kY/pVoGu7BX
jdJCuCeuT3/YMizFhRacX3R2pAK59IYireDb7NO/0rfihWh3HT+YqF0UL2O3womm+SjeHk0j0nBN
8OtPiFjeu7vLWAuqGNUUobD1Wfg/vdiciAvzH/tAJTVm4WfFiGXC9iOjqoLQa3nirc3l6sWGl3dA
ATiZSBMOfg3FON+/Wm0seWIUWtvxCDitTGP8HhFydVvlwVADwyD8mq+/6MY5liDbP8J9OoVk/EdU
b6e08eNLLbnQa6tWy/TPizUeKa/lzM7XwCO5nVQyVNsrci3uhOWhGSyu5bvyl6mSxnqixCrCTa36
vX3yVMk9k4V1bqcZf18tgqxX2TmHPcHB63xNZOsr5HOXbU6pClw7FXFiWbtVxE382p/R5fJSGsH+
87l9Qt0I7LVUY50M1kHWOQp5Yuzn6iMg4u6ElTpvhcFxHX1H4q784hgeXdbFDmDsCCOdc3mkkMY6
+T454lL7JY8Jy6Oi9hrAxxFWWVDizvbCZleNBjebxd9yNAjH3T6j+oIbGW9S+YyuK55lMcrG6d3v
gecM5RTQWG1jZe4fBiAAtX508ahMOZuszIZkmCsjcALu1DDw1gGCj48j0xsn6z2V9hYO2sqyT/mx
o5+Aw3suiC8AyX5celO3xg9ScbZ0zhcSeZ9xMM7aqF+e4oDg1AY48my6s5ThFKt5epE1xgvWWR9z
eggor/xFGIJj4hsth/o5ezvQByozDHMwkndEe8WC95waHpeKc3GV2Wj6WVcwbAwb3sqjNC2Zlclz
MuTQ1GbESOYSNtNkP9CWt/T0oDWLFyVgse3vN3xtCWjA7VIOHADSn8ZTziFsgzL55r7AqSKOv6Na
1nWIyovH28fDrexmPSCqJB6txyfzehTgV86s4GKa3+VKvF83DQMBrUftm1EmLvrQI3/T2aaQbtgv
UiJr+FMbWlHyUofnQ6aBA8UTxRWEpcNZ+bwL2SNfVUeCeu9dX5RU1whN//L4k/ZE0hnbXKiUs36J
TKg4CwuFde5ordzOUltkNc0PYxWBjABq07aiJIw0GDVDs4jnazLimL3yxDlCNWevu4x+lK/KT5OO
E1YzsWnzFwAoUxCx3VNVCO7zojBzvhSwYwBLVAKyRmtenCaSPfzkdscQgduMwmEVPTe+VUS9SPtI
JHhQKz7rPaKYnTSzC2rn3m3S8TCIRV75AeDhe7XReXcQaBxnad59ZDlz3k6V70fD5ItZsFqc5bh7
RY31V+cLX7R0j0CXE3FJ8AhAB1D468bYid/LPsLFNsZ3VyS3XusdHvQ4x7X123yxKM3/NCFmQbz0
InrcPGOI78QZWe1CVie2a59//cHO1TFzA+SVUu98A43h1MA07Boitt88X6U9XdoSkPDJoiYAEDLq
p346pAPE6uWcC/5Rl3wEdBpGPQGhobvgxxgRYXZB007XMLrx/oEdilcdZhyC9wBjQqtk9Mz7gb5j
GGgcsWrJcqgchT17nRaDs3/MP8EFlg0WC9uX2TDiabimyA7A9Ca013Bx4TYxlM+JT9PiZnbO6Nff
F/BfpnAGdgMf4NIiEtFOkrTJolrnDqvi9PlbQMYKWOddd+MHVBGNJDEojH0Y0pm5WoknFpDw4peY
0165oiczHdgiDZI7NRNpVjf7GPOc6WirJQr4y1cJGNiEgn3PJOWwfOpGBUSC4V2aTySvqFFfqimB
gpwd5ce+NGoL4gHFKCtJW0oICGzxsAd46RZpmW6UerwABrmpAzxUYHIMkj9R4UqANbQlYj426hB8
ilvbHX+Xk0uqrhPxjenBbV77kV6609WMUrQrcM0Z5797nec+xM7TTYKvfNYTug5r75t2l8eg/Ygu
pDOrMbaZcfp9WptRdtpMA+SJSLbhSXssTKtq3XR5oHcAJpaACda3ZnUFP3+Q9AB4HiOQStdXbohN
1hnceBzNEzn+pF/9YwnhUExBVWgRJIAfk1wLSKnno8XNsGuCKB4+kFSST52UoPT6IeMJCBopdJwv
o4wEfhXnJ/CzBmAokErNjRhYQQCB0EfDjjs3hIvhVrKtf0PYhblt/3c2Detbat366yWIzMdXtQaI
PPGFrLKhQyigtv/V/M28X0Ro1voLSAqZdetDsKDy+TWoW+/M7i/p213PQCv4zRaq79Kh2KrjPh8o
zQsmU8KAgs5rFwgtL4pGrXFXoCARCZBJjh83VaGWscNcg9ntPth1BldSB/HZEMg9VpHCRWU7V84S
LoGL0QfinZo8OOw8UGjI+DTCsMEaoFrrW6LgEMoYGGyDM31XHQ7OxaoZseYI97dmqKHVLEDAzh+z
A91p1b1DtI4BxWECirbWeiqM40M0LfBoGyMMIk3S9FzQBAeNHs50FY7vfMHuMRNha1PC53KAzqGs
ZFfTmF0Jfctk4SXfq7ozOXcZvphpKKdhzBZFtdoysvckRDhWOcRiBpHRCOfe/sAa8TUwCk3pagco
K7/SNDeyD2L/ACY8SAiRnUTkCDnoFiF9vhc1YQ0TLux7Y+j+7AG5BdK724fx0VY5DyMlhLLtX28a
U6QNGT9hq9o9xk8/liGKvmHBkeqiM8/gx30BYvIS4wjobe5gIKanDn+nNFLSC2LvLJ7pe457vgsV
zvdKGSA4I8WEz9Y7gF3f+3TqUt+WN/cb3D2DhfVu3AYSrakv
`pragma protect end_protected
