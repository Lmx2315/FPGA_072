// (C) 2001-2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
LY82cj35C1f9ogrxoM6OhASh5/NhyOwpIJnYBkGwZWUHBO89cssVUKuNO7dWWAPDWmQGEgnQUtB5
j3zn5uVj5YQqGFIHXnyYLdNLBslTRQdGeyxlRQJRTFPKlPPOdNPRmIc+BfJgiPHkEXZlW+GqMen6
ZMRRC8cEBBFB+MOGsnXUtuWdYMyhAG3wR+Fnp5BEyEk5PGfFeJTKWsCeS3uk82acwkZPoRdbFsTi
o/wBT96nvlxYI8Q/gLBoYXilNO9s6Me+E6KCmfMlIK87bVef9kYPOlb8LgmUv1eIdwbypo298RfR
rSCmQzVKxy/0JEvREeMwh8m4XBc26w8wUwQXcQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 10944)
mfATxf/hgHnF0in6YFFRW14gg6fFphfS0ucoPYi3n/Ap7KYh1pEa66PAC6y4AlT2N3yaC3Z3uwOp
Zm9inKvu/216kZUXrjEF01jeA/1GUVZ57/LLdIvx9ibV2scLuprxAaa9Q3BDfADYoczCDHNHFcDx
bJGZ+84RiK4536v3M5vO3umuY1cxjiNF+ZhXaVjGm5Z6Vgndbn6gSooioGKAzpyTtcgHhJEBTkEG
fvog71bmi/p7vpSHB9x1UlU3+fNwSy6TtsHPrhYfp8LZrRr1EULV0xfB6pxyPmcaLzs9f7J7MYst
IDgUCxT8zlJIkpSR9fsXxmb72BdblLXPxH4/1CpxTFHAkWIy4IsR4qhQ5goD3sIwC7LxlUO37xUR
gUYOLYhBW1q1jKmhjLyU0uri+p+DJzpxOJczKXFTd5DdTAZxRp21ASQGB9zkkNSVLYWeccXURAoc
d3E5B/Khwr0gQhQ4z0xcFK1jCgHz+J9K7ok4w/OjtyXcIdZhrEXFNrFFqP4ZyZ1Z4Q9Hwi259S2g
qT6KbDIYES+DKUAG57g1BvbOo+SAMjZHlE+dnsF1mr/nrEllj3qUFN9Rj7sBIUGhex9ajJNealDA
8GL3fuTlDLCL/W9shxU1UiErhvUaH77V0NnYVHeKZs6CBhlm0s9IbLdAI5dTT4UMZf/RqLZ97jym
WeF1XpNR0SjLuefZNl4oOB13v3iSlu2i+kB/VBQtPwwfZvmQ06dzBYZsK1LoMh49XDNrm0FmVYVC
6qPN7OGL45Db7vH7gQo9N9VEpIy0ayz6dHRxIXt5cuHEqHUZn5JQtWXHv8J3i1ICiPGC4Axu92o1
2qPKV142CQBeVJ7TclkIG5EX0X7+PFItYVSKpshtLGTmGE+ynBBscTWZpvDSZiuIXcc3SC8OZmRs
D4rwnlUDZgO5H1HTC9129AiXbVWS80midj0AVyXWd7pboFL3bWY0M1r/5IGhQs14cwjliBHyR0y2
f6ekazrON6y3S2Nc6vbVxMAy+HEgljn5QGI+8XcqraQSyZIewIHc5Z1z/r/yYTWj4L/m+Ye+uGb2
nLDA8JVFr7uESaaw0D+WwLYhUDhmF4BiOIj0nHhx5c8v2aDNPNMguyhMYgvQYSPpZVNdTTjokG/z
HhvG0AR7xaDh70lqHdR0bkwmVTLb+YT1gv7Ro84uNpuCNC1evHE5cYEFOViU+azhn3fm/0nqwcgY
283BuxOlI3SknMlWDN5Eu39DxHb7g73shkMkFmy+S5MwlLUtb/IYMAXb+MgMdTkghZt3wNi/6LVW
H3Z9LsSMdba/iH+KbyDc+4HO2202Ro9c56URa6AI/O82JedOdhlTjtmdkKbY5HR9MY4WPn7dGWmA
nf1smGZlFWKeFrehY6/cwJu3qrCKvUwIKuU7rVO659XK0pp9MqPN7kIrOfulTIy5RBcICWEbJppH
P6fufJcnqEVTbnHY2nALFF+7OQhPmCCJJ78prNRZ8a0DHzHV+zst8VH85m9jqLHkcA00urgX+4MC
SpG4z+BBkEQQoA7CvQq+ns19XQF3albeXj42cUCMLyqruWMFgutGKDm3c9sq6/0Yu9omn6rTDVfH
ssSd4Lx/t4ER6j4ELlrsVB8UyQvf/tgUoEj+DqDrdrJpPknv8uHkpDAHUvRg0vGvyg49A/ZFN5QU
8IIfVQXY2f3y83K1BaImVIQp+fn4OkEnxxkOPS8NNHpYPFCwfUwFkOAo5nJIzi+PwdFh/a3kouBG
2TFR62zMFLX1nMC4O4khrkNN0R9qo4HEhAoYgHkR7RpzPmuCcwTwJUY5QWcu8z5UKBLWVWxOL5fV
7B2Oz6XqYHUDwtTKOd3GUvjTkBQCvkrsWNw3af291SzOF7cWleNTtuxlJmYe5ygarlEPwBKmtlNX
MeC2PmEHAVExSLbasAieJQI4qNkiDUeAigds2aO1f8SA6ilYBt7LP/Ccmf1t9eE50XY3icEMOS+/
zDAg/f/DhomLwasNlV2GVFwk0gHZgqv2D5S2GYZdtIGEibnM0dUMq6mLyIpnlZ1ArNuZpLGqe867
eYq3N3zp6ZuS/tqN1nc3CJlhK2mYNPvO9PJuuA345QJspjt6Pbg6jhY6r05Uej4e+ulRo5H/Sn2K
7W08a3myBI+4dMgr12E+bqYFF0ss/aNA98Ux404v6KdZ+hnqQLbwBwV/Fb03j9toX2BxbMVNUmm+
MFKnbMaWRmWab8fy85WAqiqL+Kyk4OeDuDW7riLUELK6hafiw3DUhbrYZetjDVAxU/hQpXGGDk3M
qZrW2JhX+tvZbXxnCb6Z0MeMZt/n+Sm8QEL6evSAGnPSHK9V8Mnzw7k05+VlPdyl1VsGDScVEUXD
zSNIGM91pKuKj8FHQLcIBH+gJsD2GoNA/d4MfeUSCR8AYN0UyZjyCLQxMKd81MfKOxEb2ZsWR7CO
TX0FiftcBtoZ61qFHYQj21eEFCt7YUCjtxGCbEEUZ/tCz1s6gMHY8VgXpNzOf86GLDK0tlTgdxMW
ukIGCWNcmJIZ2vHr2tTiZ2OAhT6cvJAVEqbfWXLHKzTCkcHCNZiY4rbZYmc7J5+OkUJm34Y85iF/
W7uMyQrHJ3CBF5TKiiT5E/1T5Q8t/Ri2BsmY9vFpBxhmOvWJDg+omQGkhIhlBmp1Y754qRJ51GSj
kNEsJGYXE0/GPjWLFraaRGaN8aRc4B7x/Df5mZeTk4QYULUDTuGCDqxXiNVRcoj//xdQtuL7gcXd
4y5kd/iENv1yA9t6nr14v1b7x2bqEQbytn3q2OgBBQN97iEai0cjeW/T9F1bzRUKhRDiLqywz8J0
zOVTTcKic70ifnW0DcADte8f4xELb5Na0fPS+usSE2Hsu4HNBuEJEF77BHRjVmQHgzSdUEIoRNfX
gwJE3Hq/v8CtVPj71ffs7dG/IZ1YtfpMc3XoqzmAAEHlKEO161HrCT05dkdKKBbXP7mTwFem4pdz
YMvTg7c8Wkwc+wil/hC3h9nHGOWTKmAla7XqFjHlf9fCplYg8WcHIqodvgZZZAHMWaoHOeUY1jWs
/h+Vs0HG8UTzE3qaWcqqqpSkeO4BK3oR+TgoHN2EDXVYmOPjoLr8hpmAkRV6YTS5UH34JrDk7iXh
xowPn8rweE7kNB3sAz1ENEaNiRM+5ZjqH3u5531+4lRhZoAdcBB3DAYm6h3y3wg2bup50+fbLdbA
erj6ym3GLJk13aynCDcq3mn4IJJiEVn+DLbQKZUcVVOz1ckPMKqeXk/ycsezHz+uZQ+CD8v06KMO
5ZjCltspD0ghVFqcaNGEvpzjeDuy7pC02qrUh47u/yO1YZl4Hhsy/EuPC5RUyFjoGI/gFdIIBkxz
JaEvIi/ZvcAKWOpy5FRONsadd6TWDKbeuSMQTB+5/9hJ0vx3bp1gUBuEoTOvD+fo7cG3rLKlWrO5
+lFzr2EWPszEp/XkoabhsdMQewAFjq1WgVtwtHP1kGkq8EVUjPPLk+Ps4lOCemT43SnpScb4tCUM
z9Lo5C4HP42cAyF5uZo4w9s1B7Qt0mrEONUt8uA6/MZrNUL3++vxLEGy4muGO6NtS3gMjTTrnBHl
okPQE4DbGGU4X9lPqyCnIisL+1KDhS6B7rz5sBuGzOBxDhxQNis5803NVU5fTYXTRAr6SlWVVqls
ITqLABdnSySU6uWJR0HwYeN9917PMoEAT09F5Ab45aRqsb/h1DgrpkKefxJPciPZUcLpkVQTqVWi
uTVy0BNkkszNb0698J6NTWg8cx4iJTVmVsc6WCED+OWN490zr6n+ndn5zsAvabgR0lN4CcNOZZzs
1hzLVIXDZLYjNFCUIIuRawTG4FmyUAoHZCY8avhKPvH+n+DLvu+h4qrpTCbIJAW4ZstSgwQ0GBrz
jkY08B8jZr8G1CZPOOPO85GyntY2J/NXk+I2TwRaTv0uWViLviw5k1yOwLMvJ6eLk1Cu3+OuHjZj
cAdZs2a08xxBAqiOJ5Q6ooPOob2zKWpnLiPdhnm2LcpMvIAe3qzObr41V2v5PiBEIR+rYDoSyctW
+ceyeOzAnycEu9y/0TABkqxSw2yYXvCJ6bXs7714SHWkJR7LtXTtRmfwrQe2jg7L1bI2xbPxeEha
2s/ZFLco2WNtAfBe7/lIOv2mOT4Y3/dbUB9bwkY2s6IU6P2a5AgzHyzuGGQ9j5gzHHHRNZH+Cz3y
fND6KeH6RTcKq32FO1xZT/NGD793ji3aBGbLDGiijTHLwI7y2oahI76FXl9xkWbG86NzTaXS6zWt
HzFMauMr+Ubsq3s2Pclv2l+DVHvIolWbc6oGI63SO7pSqfU52o+TM21dhIlMnfOwHuA6+6KQdhi7
HkMp/RcEeX7Uza1xBhLg48tVOaIszDW2H5r9hsLO0hxC+fyuGwlLS/IxUc+gBBLsSsOP6QUV/bYq
qRbBbkIzyU7UBVVpb5DtSD6GfBL1rfktq4ZjDJkgb3t8PaHbj20hgiUaRLF0oioK8QtDF/mcguiL
tKGRkB/Dw1kYcz+jlK2w/CVMcoPE2N3Trf2J8OWTSEsdAIDoJBM5HXM6TXoJg+gA1qWP0A+e3EkT
x+R3EgFObzVqjs/cNHwyy0nFKxWfhH9C3Q0BZDF/7QmbGG2s4DAR6cxqzXImmVPytId+l7EPhl2o
PotSYLG88jJtBlayO5AJeHhEgtBjMCK7gb4qBYk9zfFWwapl7Z/nQ586sq3RBwEC6Rk3r5gqK+xm
mW2gaFiYn8Wr6IwFOnXpsgx7w7ZaYnKWoHt3SqhXtGTDSPy3C5gnGT9afSatjOuzF2Z4iwtqxc/P
W3W/N3yPugmM9FOzNIvfuIpZQLpVlsCuK8ezngczFI3LlLJ0iOKjsR9jy65aswBg7nL1jynxAHbT
XpjtDAwd7mxFWfTu4WMpvqHofb9KSAeWXkTgiHtuwNrZYuBnYF5a3p+l+P4eXBHku37eOqg74nQT
KXKJBpe8BGJDXqHEmq9uRBIUABslZHz0ERCtahWkE+LP05WWzklBZxii7qsHMG9xetH++xXBIf8F
ZuapLLIAi+YNifJH0y2AeOM/2eHYtKl/JmPKE2/36jqXq1/NuPHFyzvAJ2jdgELXIbv5OUOpOD8M
BctF909j6WMdYIaz23+6x/uLOLhm3Hi7tb+LFm1R3AAbuFcUIQO9VADLapZVnK1vpQePnF3+5mSZ
EO9MiqZSM/eU5MuafPDdodIpgrgKCgHmy3gE/ZPj+S41Kva1VDGb/7PcUh1NrUXoXwyYJR0rPosM
hrKC91LnsOSCiZ4YWdNefeIc9JZf6FbmEi5LTR2zWlGKDfTGC8mZ/WGnORTfmyEjTCOOhBIiY+/c
suLWlMRqAjJqyel0Ve3xJsPy75wTuKFOPCCiAlIB4AziaxoVZ66Ayjs+Re6HUlp+NYWK40MtMELF
s5XgDAQSQRctkoKDQN2Z9JjZb8/Mt/QPSTukR+fFP67OGkZoxBYbO4tmo6F3kvJ+CqqQG+YH1VaX
AKwVYltS41dm4FKpitOObNqN5bTHHZj31HNq3yd1Sc6P7Fdm30MiURi3R1N5sgpjUxzwm2zUXhPg
JT4VdWNPCDCSOvPy3aUHvyq2zcTv6DzGXUpXz+UbHaqlNcBEqi55xrDh0SCtLHkrOpeOd8uY9spP
JRd8I6/C7wTaA26dxlF6eWXaya/wOGZVztejssiP/tpT5yFWxcvemA2B6QHjVrwuDOm8mJ6lYG+0
IuLudEOoM+HHytOkP/8iiODDgeKR7YCMzNt+OHUzfD+M9q17iQYOsdmGli2j7wp821L2XedIKeu5
aJzVSzto3mfqAXEM1U5FI9uGBGizRCHwC8kayNt20+yTn2oz4MakrCh4oiZVZ20UAl9BjDw+X26V
4MM7L8aCCly4Gywte/nklP1fClg5DVuY2AdYU9amuu8ejU0HWO7PROqHWImyTbn4SIarWE1J7a5e
g0Y08WtfaDi7akQ+6rZzr4C+syGdPJ48vTqxARfWuJsrwMj0rkYRACRa6ELyyQPh6GUNCOtLP1GP
lV8QTo9HJOAzvRnBdWs/uMm3KadYrMQXlGDngqcUPTkqBLW6KGGrcK/Og1yQCDaCanYGPbRYkTVV
dnyrgcbYGGBMXCS6KqcVppa1PUR6JQb0CPlcA2sADb+zFxabcLw14gnlO6FQIhbrhxwNJAoagJYB
YK6fiIVQtvtcmzk/X2jS4xB8O0sI1napN0HbuUlWTq3NjuoP9Jei9tWm7mqYzNsEsOET18BhSnf8
8SsbORjJgClDJEbDOWM5Ljf8Wlf28GPQ1jW6wtSd5bJIwNi8Q4Hibnp1vevDtL6xsZzYjlMxgZCQ
Pbo//WLRvJhwyLT8ACUGn7E3z+tO9yQPGQ75DzFodBsGl39JYk768klxZpY4AEeOze4n6LMfMFor
C4I9T59q5BmQ5hzamst4LFVMBStYHAtP1f5zdODhwUQgO/SEEa052JrWELVN7B5qPVRBZxE/YZOV
kYqybRsNqSSkVJMe2OCJNBqqKuPSndGNLBVgPuvVdnH1iO8iTRYYjTFKFyKv+KsxBVFHamVwKST8
+GUcaeUsIWBCO5nmxC56mnu/OMkBlnlXrdJ7oBtOj/IBm4arkxutVBLWCT/INgIW2BxS8trFQCmj
S6okqm8cCvrU9ZPxb/Z7C1lLW01AGiwnZV0EFSHDppd/ujbpB6MmJ8JMKu9e9acBGfvgJcYojUoG
IIPQD87q4AjawKHTEHWcZiNRsSEXcACW9Hm/lbsx8pLbru/otyvV0N4/zUhJJ1Z+ITWyWPfhRuE+
4dtf933wzWpiewUD6zeTV7TpZK2ffqUnD55A2UNToBeRh8KTEruhWKZcsEAaSyLNaGyhv7bT05yQ
Xms9dHMouPD+8GtLrn+Cc8zJPpZbrydZZBuzyoi0nNL0w0tquzs0IQcjZ2cZ39RLdpqfrEH/XY7g
y5Z47iXTp5dQh9ixAvo4t2d1CmFSxrrrCRWbx9nyCnb+47W0zp0n/54VU3itrHvQFX6pXyua4MDM
80WS+QkraQRe3k+jDK8gyngBhWWGm1/ELovA7DOcEyfD1458Mg2Ycm69ijt54MkiN+xVdnBDpc8P
tO4iQtkRo8Buyq3BTdUNOaspYrTo13deOBBvsyVDE5So8sXVMTp7PJrOWojGM1bdADPsY0CHSUzp
wPIYyZvXlxCKyVPSzF2RajYOB7jgVWSzYyYKBh7TA0A6X+aqLqWmi3N1jO7fWdmihYwz1j/y7+Vy
TP8jK/2oHKrLwy3+uacMH8msOo25ahmyw3QO8nvdxa3hJhDKJrKLzs9bTRecQi7+/gQYF7xmhHBX
UaUY1eBbXnluDtoCOzPj7k3v84oyujTJCUpVU32yMjrQ6k8aPR0O133h2I670lWiW6K82uo61ebB
eTT3b6qgm6+2PuPr6daj4yoDppIw1zBHj92RiaDRGkZuA9Hv5AY9+audFj7WK1GCDEZ1SVHffAAa
7uFjD+rcGLrGyN5iHC5mK0T+/ZBf3V7SAhj7jv2vMe3oXPpJv48YvUWFRvZRLnytS4m1lhFzCeWn
/LMBcVIqDiq/LTjgHEVYFEDRkYQ86weduIjOEWJdOT/1nskEwHylR3KEDV0vGznyznhisfd/LaB+
rwACPhrNvcZG3L/gsrLZQ70MKOwrrjkWWrsDY/vWGpS+uL8ffbIgtcm8Y0SZLXFUEIS3XB9aAAdr
+C0FPjAzyXC1WfoU/23j7G3PttkRrh/MGAFeXX64YBLKA20uTjE8R75ByaaBWPyEWtljywhKIkh9
OVjX15qrRQkCHmxLtsDph+x6gDQ543vqujLUFyEjBYtirAAS5gZmjLGlZaA7Gyt5bqcDUJlO/bbX
bLy4wy5j9HTZOnkVORUrim21nH8bpV0BYzDji//QYC5hrBa6joGppURG9crbfEBAV2N9bguawjoG
ekrbjTO7cXBnOCXF7dfkaMfnzuv2rQVZnTdTPxZQa7kRK2q9Pw9Wsphno1zklYToQngS8esVSWzz
Hup2JbEgX+acoejJMHq8A3lD6nv+A+9aVWzx2DmW87v0ZL71FFvxgJNZfER/OwSwIMbQxlZCCd/A
9lNSYyD/U4KDNzZmcqJ1lEMRm2xFbe0dn82/DCdkn3TtyOF0+UXqhKusBZLyr8NMONxsBQscVI22
SlYTrcC8igYppFzApYcezSjGyDBfZxN2QUnClQbfYyXSyLsjzCWnTSRj8PT+Q+gJ28DlkLI7RgRx
xxgHFzVKNmgKr4XjK3ujLk3eoM7AU01Xsofw9sc3lEl+umgJHUFFBTrWZVR6+slnUA25jYqdEJBD
Mz8Rlf3SJDkC5N3i43v09x83iXzNpthqPhSNkBJ8JhHkUNNQtCox6P4k3Og/VB3nJvclkWOSkWaJ
uP9bIHWk9Q7w1+BRZ2UKgDlVZsmyt+dbppfIQiTYOiAuQloP7hK29RHIZQ2QUzPUhNWK/CBhKgNZ
PS81poiDamL1LmYyjjW5ooy6rGdYZC+bkH44ekdhBx52xLXpV2MD10dst8/v2lmWD+5Gm6gOQhmM
i1F1K8bcYhWn8dOmN7MaoZ+ZrdqhJQtTWjGoitLg23X+40f+JEt1UxnaFpM0rFqJgVJH2jAVUmPf
VBA2MEJSFygPZWnMDvUgFPJ/AAxe7jA0UY5VBfJGwvHNg1M3N3mjlsxPKuHh6yaG/9j3S/YD8ftT
r2aRzY4WhF2iTT30UDmTOkWe8AMG2sy8rqQjae5/+JUDkPiEywITGvr3pMi6LrMlZAIvN8XiJnzT
3x0+O+kIwXxVNXp3+HanQ8FwD125u59tKe0+LFciVl9sYiS4JHO1zXZMv2sWpLGfKYSOOqQeRyAY
lh9jKRa4azPRsYorFTwNngtMvQFemt3FZScPMO+bNgyzt//4OdFCJy7a+SN0Fn5+aAUJPH08EdyP
FCZAE6qmzlDDS+epDyl/fMpzg9oyGbz4DWKVLBqvrjrwg4xBcGoDHCYsOYKpwrJaGy3/oV24j5y8
dOGqJkiODr5gFP5qFNkU/JBr4jYwcGo+Bu3gXotn2EtRwd65Sq5pq+2M3R4+BLk9ZAVRiXgcS+AU
UktDePXNk4rEdLbU39wPdUCpiKEatsN/e1IcmTImwH8IptO+FVSJGIdLO6PHud8zxeRZl0Jfmmic
RwWPKwZQLrRaRxooNYpjcfipblVQQjuJw4oG2x3HJihF8hj4hQFAhkfYJZH1S/0BU/LX8M6lZwMv
ACJfhOrY0zchl8HRZbgKjkodYq8ynBlpdw5nIFqCk9gI370nThHD0LEJWstkbB1dUMgJVDB8eYif
9grsBcCjxeY4UIDf5Fp931A0fuHUA64rDOvi/pYjN2ECIy5I1/sa50veM2OGZEs8FUfB4fvRAJ9K
CCd9rD8gKic6isPI+AsylEpZmK3+caBzEnVYWyTRpgb5/my/unaK2M0LtOB1NScH4ABmj7gCdp3C
jllCCZDOBgJWSCUBaQusEuWMvxjSXrCauDgBRFQI7H7o8I9jSiUF1lWdCFrMEkTsQbblgaeZu6GI
PtlnDPH1zEqRcQxhkL04k2Ze5R2EFsPa195+YdsXu3O5vr6gI6NclpmMiiKOeyF6S6IT0ewOI/9g
QwEohDczZRP+O3d7T404y2CYY1Zq4GeX2DepbGDiFZjiv3xjSGk6cRulJnR+POWZqpLQLkebLLzT
GCi97pXguoiR7UH2DkpFeRMIzmTzkkUhZcZNhq9/pWguN13e1NeSW2+gIVoocI9LWvA/mE4ypLMn
J4gIZ8pIVFIjZf4pyGnuAoGp3pxUES56ct8G/pxSboVHMgELcX2cx4nQElaHikUYECkqMPZ/gfIx
E4hsXGVPYkwpReTwfHFDVrk01K/HdWdy+lkunTh0VVS8CzB/Lo5d1MmtTwwbKAal9peif5NPDT6x
5WxPZP6CU79f8WcURFQtws5pVk66NC6xw5eQFei49gfvFkE0Jqu356biRKezpBxlGeHiGkbRf2wU
bBdKYB1sKMqixDeSrHXs/MO6lnmqf1Yhi77hqEf/8CIqy6p3mvnrJrh22PVFhpei/vQdn/LESPTY
xiDILE6lhtkJY7YRFI7lSMUanYFND4ug+gIiLx9b7P1X4FayqHhMv8A5scknpU+endZifvoh1AgH
kaL2Ei8teLTVmx3fy5+KKiuUibaeG9mGHIL2m4O2wjbqsZ6U9Ya9MVhvIt/hkZC/StOBAlbhT1Ac
UIDGEzQw1XtxpTUJJh4F75EEf/b5uMSWgnYg4pgllQJEbOakDioAhE6VGwiOrkgUnMs91qgpovG7
KqJ9N+frtKE/Rkbteql249D4yud158+Jb9U5IEX3sPcLLlGwiyKVq8uzpm+LWaCwwgwDPGR8G82u
SBsa+xV3779NR5Jw2ESxRHITc+2nHL2WD8eplXTADLn0vN0GYZ+ZGYYnsrxsKlvAM0aCYitsuD6/
By26lZX4NSVQFiKja7WinJUQH4ULFM74miVWOrt6JQHZbswgJ+jY4HBMP4hr2RhhesOu0XcTDjej
/i1Ai2+cngTvqZd9+fylh/kq+IIluNlSxWBllNcURUJXuYuMrpV4eruE5oiTAd+iyNtI8vClzSzn
2PwbQZ7BNnFSASMbMOiYqZONt1xObdAdnFQrdhNeQv6AtlibntPU0lR/VwE5c44otdmW/VmBxV6y
HBgR77DCgB2xXnPEsRd0O+ikbTnWnLdxCn842+P8XDWr9IMIzBaW4QLkcv7Sl05TDGrJqrQttt6G
gZviye4rxcNa8AfXJiSJa94nUCG79aQD9a42VkS4h4/EP+pxzFXBaWPRtS+ixFs8hYcSkew12ycM
jClzOTgY6OTSGkg9KhTdudm69PRgKRu27GLYKw81w3Bgk8QH6Dku8mtXHPXRAG4GayTyrzfbw1KJ
hxDWrMlHMyW8qLyhVC/m+Vu18N1VYhcDOfRXYSC2MZxXug848zopcFM+6sfcgud6Mz4v5roID/Uo
n0TDFS0om9h/0Y5eAkJqZlHudF7yd5l4HgA7GSBC4iqd2YIclpSjJMsHh6BB2P3yVccy/LrOKyHh
UIwZErG//eWJR+0E0RUx0zqrTs+53nakXmSUcupq1f1V2647g2bYfBEuzPmHB8v9Zz9+BgEnfxda
IDHwMgIYmBGLsZNwgLNL3ZYv8/wUgUwy/ruY33Ze9+N1y2F4APIDV8vmdKdCnyB6DzhGlUtczceN
vkJjU1ebVrCmYWkNF9R6P1b8ZVrS83/C3EtZRYS681DmAPZoEZIpuXNiWaXOlzcMJq5jExW/OVof
HODPr35GEVTl4r8qbip54hTjJTJt2lv1eP5lAmE0RxOl8/Sym4xTQvCmX3EjqoBLq8nFk1+rF4iv
3MBfEHi8/ItjoZ+BcFqAJsoqfwy1z//zhqPktZzjda5JAiS2aQYyqNa5yAc787SyDuDMetzmdSYK
jMkOfpN9Ti57zu2rn/RQ5/bZ173X8/FA/jtg4yacZh/dte32ZSV5KaorEJ7EFvwguIfFlqYLrFpw
00qi0u3RV2bHiHsnqXM2gJ/Oq986E80EnCAjp3D7D7PlrjMAvdxVpv4uEiLli3zIMB4ctlMHuV3G
wH2HQKh/QkbSUGDGB1xkfdOqdnNnPSyrq0EaDvVWxIFt9b9Xvor8xH3e7Bc8WnbXDeY3LZktfz4o
1CmCPki6URk/78WRkgTuizwnWaPpLnIjGnghR5/ICWRwrTGhX5DYfkCwVf3Upjt6pJu5WU5A2iDk
5YZERGnY16LEYJ8WA3EwNpgAUXWgAo4+DqU19FO5ZpebLm2sTd0qJ2s3xVsB9HdljoMRp6UU+H9Y
HVxzPKuBcuJNOEbHmcKm/47akc7e8VzMMvc/0UDMmhKua0KsSgZs56eOTuJ6fBF0Xxwpym3fQhOg
CbsgeKe1WqB3XIZ+zRDlSX/DKrOI4j5LqSOk96jNhH47ya0MomNluv9NsFrph+UDkNjRIcDNqQux
ADPJkelUlWfFkM+a+C+K8F/3P+SuaLlE3+jCEpR2VxZqL4dYv62/F3pmf9L0Oz2VZL1MjHlPVros
FkjqTlP5ahiK0VF7OAIt26chiqLufEetdb+Uc+VmSvAikQdLgSXCbkrsrkDArONe+JyxhjD+NV8h
i0hRP0EmYJsHJxpjJbw/rtjYgShTErPvTn2YCLN4VE8Ci6ovr0Klpnr9wuyFwiyW3BpOMtUXzqtd
VkIg3A3zXEguhRWMYPyOy+3bnUXjb0gK33XPBzgFVRcjiEM2Y6L0dSTqsn3UsP7RbwcWTPzdCS2k
BciFKw89iFB2EMuQJESSOAXHghbZsysDHS6kiEu7+IhFM5PLchN3jypzbBTCWbSPSejAXqpLGxZi
yov0n3r00I8iQ4VbQjhiGfQt+WJ7h2rw4gf9WeYmGFXqHuSq1QXrdT8DlaNoXXEoqzSTczB5178I
YjLpqib3BKQjYx7W1g1yvZ0DJbG6+EeEXZynZXfqY3nmhD6rHdltJREKQJpZzitdJOe51Y6mpAbx
a52Xy1zVSZHzwqU6jnU0KhAEgNPWfngLIPSoGBGMbVO4RQ5s6KE3PTdBgnyVvRdxdMSJWxB13Xf4
LLBJcS6agW6tCXs2y5WQoR3SHUuVv+ehR0vpFMwb6w/d1LghfovoOBKt5DKc0yeYXZcCXu/c/P88
nABVxLMNOihMxrjiwzE9TsrnRmM98po30ZMTwraYobqHJ/GCt+3yZAFbECF/UvmirMPWvs61Q56x
jjLIQ5TNh/mc5ukErqXY01eSaQzkxbvRM4V9lO6cRDhDfpH16PR2Sdhrs5MYmECLJmo3A2OVf6db
GfjLwUhdgmCrrgtL9QfkrT+69fYJd4QHY+aSJdvaSt/hQ5DmOCAM5dSECCmUch422RtsGYTGHJyn
vZI2iUPASBirDVV2EOuhUI/4w+/4FkbvaP4dxikpbYyi3Z9lVUNPGraQvDPuroYr/TX88eFBkGqr
+HWUHoa8bVY8zB9xRO+MQXZJkZNeqcXZRqj9FCz5/3Ojbao/CnKrTvkjIMATTBLY+NXtgSoo47Z+
5EXoRrgE4wd8JkW7WSXWii1k3K2/nK47v7Wj8PzJBIGWXH6Z1hora1svouLbT6MXW4745bBWLXLt
CcrHPFgQpP8aVJbQd8z79x+hhFyMrgS6X511Pu2+bOa7dexak20v1e/g3i75drxHUQJDwWS9k6ua
hfHGngx/lLRwy3czKLBfZb9q3SfxAmkBRm06WcN2unF/cceOQHPznlqlzG2944mb/Em8fD1efYbw
YP3cRFl93RTkb6art6AEoYEcu8aHjcDsWjA3VRZV7YePeed+Jyj0BX1C9fZNflmkgm45W/rYqF0R
63qyaGgjUh74l53Sthgaq+hnYVKYTCPXZwiYFBSCXqoVUqxDUKxqMeerbwAiwH10Th9yL3Fzgs1N
+pIQx152XUWYUhqYsY5UF47mt00lkx/3DVjtwbXUwLQCaFB9LB4LisZD1EoWdus3CQ06bt35AbTC
euSGl9WEI7qiNJVXk+qn4fGzKV0amZ7Y9tNMjlb3WkRNsTwqCAcuQDWmX6obK4hlP3Ty+1rt9ioL
Jzhwx1XDTKNrnDNlTnkXZL+cnzLzsdQsyhwVwM2kmIdNeayDUouwL3NT19bhl/oYMo3TQ9X16zEQ
gzcLHoHH5zkgET3GVeHOTWeiNDri84t1DUX0q3+w9+tDbgj1NtS14h0W8nQRD3S2obtusCEelaxV
yrKzvp6zUsIURQHKK85vU+fNEAtiTA8LpD79ok/+06bIAoRmgS3rsJVm9y19olELDDtVxeqDKTN/
dspdOTyizjG441fsKX1SgrlKptdewGDnO/8ory2cUBSSkwVaniZLqhnZevMEHLO2f3uQXuNcfZjZ
BqVx/ly2ONZLhHbNE3CvElDSh3wtgt3OJm3Hym482bviFdS7fXTA6vVp0Ec9WEdeF2uM7k8XuItw
1boykohnLTbcTZylEV4FZvCzC++/9YB/H1qo40gjrO6Wc64hxgX07XNiV1yNG9VtfpyFGhIeM1XP
MOPWEKiO8INIEymVRVVeDas/3oxVC3A7SRziQQcjx4Ftlp9u8IR1THvvtVQx6FhdcwdDEZnRcpnx
Iu+dNjgmkd+JAWKCd0odbSOJhV3SPax+HvnXyzsyYhX9lsuKLGIKx6xka1jpTy2PyhZ8fUBshRzN
JykzyUm4apihToOWMHbRjA90K9fQEADC98hauMh3twzBgU3ltnSrNl8GFwQ/goWk587AKVmr/5nv
QmfWxR7QR2BS+pIQXspF5n3vKanASPGwNHQpmf8RDZIBPwA/WkZudS2F2j3yiQfBgl+MEEtmjdkJ
OZUMtC1aKSj7rEuugz0cnepuHTo8JEx9Et8z48cyiNeu/Opg1eWBVP5v7nUNBBb2OPrgAwIGmSkq
QkiCC5H59jF3s3+EXpcFNCq5gtOCSBG0TF6+N67+fByfuI1WyHZLYDRU/cmMpTEmQOzJhmq3YqeZ
JpQf9YUa6ca7pvs6tlxWby+dIBqkmPRlee9FgWAdEdvVHCgcZLevgUp1DP36ATnM7PNNpxJhKEgC
dckine2GvLMoutPelFkq92pgT11OAn7L62+9lvF1CpMM5fosRgAcwQ/NXc6jiTHA4GDrddTBEAmz
`pragma protect end_protected
