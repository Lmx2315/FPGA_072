// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:32:39 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
sG8jOPFtVunTPPBruvL6NDwUKqZwyeZRCm7rf9/wnRQAVtEb/kFDa78v44egYiA6
SjCYKPsQjBHohEc6gt99ran6pIkQ63GOVGaY0q+AJSpXyy1sg19QBI9DwKR1AG0w
W2Rx6H+Cesg1TZ10yKa0CPhJ5LDHPmdAt/rzuTxH7bM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 28016)
0BJNb8U4jZtJWuZ1fyB/333cZaq7vYXd78EBjizh+fevbaMPTSsV7yS9xVnaOxJH
s8r1XXlCCXkQbGt2b6rawS1EQSmqZk2Jtid0ZOnYvuAS8mQnXhTpXKyV9FcFoPDp
XnzZYV9qwoU2pdpGD8eVPxRVcXqVE6aRIjDs7xqZeFkDz3IFLYXuWwtRD+jSVoJ0
nRhzvQQEK9wIQ/yEdmfm06qvc+SU8N13xoGBPsU+gSfjsB1nfnmJenhnic2A2NhQ
dswF+Ha+5KaBDIoVPAmMGMkcHgpDBQJk3mq7xgmTWLrfDfnKqyJu+htn8AraZ5qj
g8cjW9kdDT8OFC6VxaoDuTDTE/9QAhDGO6HV/NUVlE6wa/WJOiwezXrBQESnhahe
IbVWjB0U5Ie/FFMYS+ZXjXGJKkCxrm8SNwe8jpES6R9zScS7QTwliqo48d5snJBU
l3AQZTNJrP1NFn6/ubzXtrwLPru34ODeyOHjeGJKRLDlL3L0Ftqq4p6j/NCyCLO/
AbhNUBN/yMJiJOm/4+aADLbTQUe/381ZZpgDIGwDvOvCRGJy1DteTEQazqiuUhqZ
lz932AJOB3E0N78s1U4rv8AtL0h44SfQ2vuxmOzbT3mqxwTI3fdyp2txNo+pkuIJ
XDT8MM5H0QknBdzmeg0ldjRMFYNIo1S9GxXo6JQADX+U/T9/9MVRDl1Jf8puFwOV
yQW8RI3Us/Psm3fpNaFjiSg4dZKNBMZYZ/l7jQhdGIGzm+PBXMLIHTf0G1uXnLkf
YyG3YPO0M9juSLlbQ3j0TXW76rmcW8rvayBQRgN3xhGL2cYV3bJOSHZ1G83BGa/r
X4zE5IPyu21JJixbQja3gXOsczWkZCsDGOAIioaqzqxg32+Bfs1L/eg2FA99lBT4
/EgDjyQHUJOrhBkMnU4TjjpTWVCMm0xEAaXxlJVHiRBk7Uxo9jpy5xXJf0dBZtuA
Te/lVYfiGzEIO1VFS4xo5HqujVsGGQNhJIy0rAbCTK3ld8Hk4H9o3malnbRKtxUW
yEffN5XTDYurso8+Y1sXUta9VW2AGpZpjoIL8OsJ53aAi6vOGhT5ysTxtFjiOtWV
KXYVk7+NwEUQnXPXIWek+d/2zU1dp/dTXffS/Fc8fC72TQH5LFfxo95YjmMBJVkV
2N4cUL63j/8cZG2iI0xk3/8sFCg7UY13ptOO/QMfKSP/NYtLiP/V+ZkZ0z2jLgMh
E5/InzXvylOcxnJcNj3zdsclArAqYznUpLfodNCe7mYTccBAr0B5hlcaNHVYiiSI
nuI3T1okMKB+a56taMn1sYT86KMJlflNJmSZJlQXVVu1Htiso/8XOtyNGakR6A+3
GtGO2fvYShJa3gMk4fxuQFlczGoih4U3x9jwiY/ItCbyoMl2tgn1elr4TmE4V7xs
SNLrinntrbhdAcKFQuK0AmLY0w66nC/eSTThvboxTisOEs/XX1pW4K+W6Scd0ckr
MVTLgptA642mizzlYENqyhj5hpIJ7nRT6V8pR/8L5UMiNDnaCS9MQpZgVGancV16
5kDfQo05dw+wyL6goXAi9TUAkcFw+mivhSQg+bUc2fHqF4NkGHs8MB01hc35VzDJ
+t/SxGlPLeAOsNPEPWpuYnPvTOm2QNpkhYzr3GTN3g+puMJxzKYaG0qMnQczYw5/
OLJc2EzP9brxxSvFhhI561sGtFwnbQ6QWkrY2uakIvxs3jQ3NnBJG8yREr/XAxD4
LpJQxHyxxTxPm47KfNaDk3gI4fAtAR4wjxWqw9hdwu44d81rzNJUKkRuYuBRpg5d
FJfQ0nrJcFHrq0RJfk3u+/1kln+cLjDPh0skFqKttsL9HB09/uydPDygorvjp++0
8cD8R+9UO+Z6Y8E20klmYx1JNfSlfuD+dUSj4leochGEfKdItHVwcVhy2LTEZ5y6
TmrKoLOzDkFiX3B0tTmxaMenkYTfEwm0hMvKfgnDK3T7CoK5bixyjV5pAzHpMDhR
+ebmoG6y0SAbm0Nqb+ny395nzxrljsJwz7Pw3lrNBHFyS4nundgsa3fhGJfr6ULi
4MQRDS839f6jWO8ds3NDcQFAx+KHScXX+eLe2iLW/Bmc/t+s/9F54dkai6/tCsvg
EfY57FJr2Qh1g/xmLJtkp3x6ga8DRgcGSLDUeS/da/9H7ROh1RL6Nps3saU6o/un
ym+lgdlD42RC/WqA4fGaA7MIS18M7GScWKDR9TsAtO9b6LcjAw6xiA1+sDKc8F5L
83Mmx7mkASVjUQu36lD1BUFwwCqSD0As6Ij78+8lcl6oiqlXfL5b6a1+K4TWTWkN
5iQkZmnB6wQErxyFh7AiRKCkuw6O1H58x6aIzwRKZ5FPi/dcKcBJwb21/qt8bSxB
40v0elXHsvtUDPyg0n1ubXxs1c1+3UKT1dCYHpWt/Z9cmtHRExsre66VTn535Vq8
v5oBSSPABFWoV/CQiWMiuXGLRW9YF0NIVyJTaRaYtRiQiqBjWEG5k+2aiyl/Lsqv
hq4Z+LFDRCqb5LIRfjjZ4qgHyrytusQSbP3XswHur6sK+Xl8oql6rcVmqH5uBOCl
ZxhoVOODV3YGrEMpWpPjaRtkItxF7jFchtJBoGbMr1QWxXvwZXP2azSkEdufXYrm
rk4CjY3haEAdvWmze/LA2VVO+VXdWwI1iXDs9AEPAVzQsLgmqMzduOH5z8IMo6H/
Zmy2LEYS8BS7cmJXmLYeKx2KyZklQ64owgK7ldiBgjtrzom+rMmgyPJrdBcpcBSp
QVjHA2EWClJns6eauL3Sjs9RcSa6GY2tivhvGQ6Q8QDWU+PySEjKrHQqLCP9pGBS
IHT7TqahQBD1F7437KZd0KP3uDS10j+z3wBD5gnT/liNrcy7J30Gxow4tW9yDDFM
cuudWLvVpCJisVYq++rOuu19Zrm9d3i3SGWU5CwAUxurEgf84dyp9Gij6bmeSgIi
A9JimEuGjxBeq5St6pgkre3zHRpMUZrM5g9zXelFz6m2MwYfDsTNvJ0gsewFXX+S
Up4RIfa4fnVMuGC7gXxWswtoMmHmNmkhoDwuJpcGvdXnmAwpll0GSp1ysFIZ0ySc
v9MgopRgWG7d64PVZpwTKYyaT1LrLqsSMluwLk6jDyrMwnXbDrPHFvQx5nS0DTLy
gMIHAxpF5M7pDeAuZS7S4tG2sz717+/oSGFF1vUhVXMJkzkY7tb7eI78A9PjMFpp
j8nWgsBsvPGy4BXIlac9BkSzqa1ayKIdf3ka3ptLx60V/NwI2AglIxtXqoabhl4S
o3SmLNtbj3oQasLbOHcw8MulQKJtkKsKzue0YGFi+eBWCfAgPW0unvldWvcSosti
7qe12y4+Jf0dowFB7JAcclQyHkNw/XF/S/cXoAUz8JQS11cfN2w1iZNO9ICEsf2f
diGMtnPULwkjH829C4C0m4NTjx6a4sp+8NgP3t38G9ISefFWnrWxDK4/fveLFmx3
pLmtcwa8br8y+VAx0v56fzge/bL4yfJv+7KBRR2gjcJF/FAGwmtERGhT1EIQu0Nf
w11EAyp3POR4nOUlB3ibPm4y0ObaebvkZzeIuVnOTOd370x1gm/YyRg4K6ymCPuU
ImlW3SaMMZ5hzoeoHq4Tiep2nP8lxB5wdE1ePCmTnWCui9jTPMeaw41sDtQCMQW1
U+P4jp/ceeY1HPeLsn6FqYJIkijrNU/p6WwcMXlpwixnK2UMcWy7sazk7cAyhy2v
hgsWo+16lUYqMLfAqpdiED9Ff4s6fBgwawYX+hfK9/Od9H4dYw1u62iho6ofG0A3
E+sHy3gmw1f2ofsocuUicLGcImTpMx/JlWTC8IyP5ovXvRMIIZ2hE1TvQMcMBNZX
2em8jn8hUhgpad+i2OFdtm+4xveu4eais4H+gXN9AciOZMLzGXIg4tEoF8YicMaV
0VAX/UhOcFImdL/j3jhVyOjSbNqI8zLtrP7klIVqu2eFXGRHUGz33a66E08/wnXG
jJEhlzPl/WA5fcOH2iXhZxkTTME1P8oc4O6J74q7Dwej6R5y8JdLhIB/vk0MU0SN
OHo1dUTHJvqVKPgaB8EkWQK+vMKC3M0I7NifR7jwVbtUUgYLnZMVZDGVRqFLiDpr
IES5bq3a1VGQ2JWEjBmlQv/PHo5Q4Gu97DxsMz1Dbh7Sa7/+JxndAyKKukn9gcF5
MKEsjIrTH9RuQwYji1Ws4RjHYEhhMGDd1Q2CmmeXX0/GS01AeuMRaZv6pU/msDmY
3Ww+E8Jty7iM+zeY0F0EQkDUTIXHbvrcDNfCWQEcZqQoFt0tgKt0A0AaxONW0sQi
Qndyff3nMu452HlxKMQrdCP+jfu6bwr2T5epGO8/GVb3D4WRDOBhD8BogHlBvuis
tjamFagMjwqUbVar/NHwQlqm89XF9185wJELsl+/U6hWaP8YF/JBToS7+0QrwxHz
3WNZYplMaxVd3/b9bveO52hiSoIrkffEEYcRdnWSUCscTqgcUPd3co+Sri9YrQup
q3z66P925MV/I1OsVg7fgWkX8Y3QxtY64RYSPHnj8mlWhQL1ub3PRf/C956tBncf
hIXbt85MEZg13BLsgl8rGIInFHMbqRlLT5eICJxzux5aRL7s0DbzgFM+++e3Kf/B
yWqxrYsMfDJXJ9RNkCSwf3S/WVm5V+a3m9NJFP4ajYOx3KMI3IUM9S2bAHO18D9U
5rwXZWe7jn8GT6VilANvfNYS9lQAWfT/c2glN28xHGyU+xVLJ3LimZjcJegISgX5
s2jElGpF9AsLZiU6zlhdYOdCYJS95K6z5OGBj4KHoNfITrzXmeax6EXSe2hnrmPx
f64YRuE+LuJQK4heglZ19XalgO6jrcPckAcLPe7wlLTLE7BmwNNYrHjCZcvB+IIO
9DMylAG9gTsIAU+UKxjQhaw8O78YUZNuHz0HQZqdV29U+Y/LHTyZU0aTeW/P6WFy
aa8zLAw5UDY+OnTzwdM1EWRAtfR5IAO7WATckFys+2IwUq+nW0Z1TxdYzt2oN3ab
WjbXG7k3fGdW+PjdcrnaDAjwR7xqlKFkSl5eLEpRjpFRJm291iz/b+NuJ+zCy6sD
47Ju7LB2FOo6l56K8wdzC8AThUMLM2kBsXxqJd9vXffkAqkSdCdewBIm5uk3aUH4
LDhy3gbxyaqb9yu/BLlOv+/fjK1Smwt2/rlA9bsyb0KRlp63WTv0IVN42orqPyX4
XgSTj69Zs6oKALPB8mjHo+VrUHKSY6Vkw6LexGIZBLQux6hx+d/kZS9snA9e5MAv
9Mx/+TgYNCP7Pb+VY89j+sWQvTdM4YGYY/Wfu1uxJMMylsGRAR5ozB0MwSQkxXGr
fdF7vJIWoKbQGGVeE0dC5J/drxCN/iBRlwySY3FAw4v4LXnzcNKk4R42++f5mS5l
ijoV+ips2B9OlrCV29qgAHTAlnDhaY/nTO/o723VXgK67zas3B6ne9r3Mq0TCa6x
l45YgNzk54d5tPKZi9ToiOTKgmvPbUKiWlIZlXSlO4rYYZ/sKHBZrotZPeihIo7B
M6gfai77iQAj5T2+Arhw+6kD3mn52PJnF8qpopb05P1guN5auDQ9iO8Sdfp1k2Sh
I1357vkpsJ7rTD776/0FdA6O0P4+VSCAOXQ2vtDOvDKEb4za6z1uiesPNxInDFZ5
HjAEfX3lkqj7wlcFX4Oa1ZYPzH7utOGpoisFdfPuAW7BImBlgZ+Yi3zrfnUWssE1
iJfY2D49xB9jHDzdMw6zpHXpcUT7PjtW2Yw4h/Ncfwn1NXdCsiWIbz/Rey5Kx31J
b8hvS8d1IhLuX9RpkiTnW3jiNZRWQ5H5GY/WcsBQwQiK5yNUwWP5KgdyBkM8QLul
Vy1Q6uoSTtCNsWYBKZ7cizjUUYP40WUjtSilwx+hDhVnyzcpUZSoX7IqT3IApVdR
Texx/szUHjol4areMSUzgScCZcgRvpqjOa6YOBtRSzshn8fD6Q4EF28f8394K4RJ
+uiOOJh6dOKIphWjtOF2AYAuKUX4Jj+i4mx8kByNYCNpiiuekevf0VGzaOK4LtYr
6ux7c5pXTrXUcq3lfwdRRHUlKakQ0QmkDRest9WMZHqu0T2ZvZ/XG8VV0k3iWnyq
V+rr3Apmcoj1e8LLCarMTvy3ygBx9Ln+VsdOwFbFYV3z/f4/AtF1ZOsHj/QbotoQ
D9fgSQJ3iAU9f9czsPqWlqHTVwiRXTVT0XLyS2fBF5Ietj3GLcgfUlMkkiC8/7I/
LL9NsNdlzfS61ZRHXVi7epYvNpjErXHwhdeHtNw6NeRIqhmmPcNvkMWcBEeMEKr8
gIHr2IJrC9/QiDbAlU0CPKJO7HZ58ODZh4Y3cMJqazf17wWqIgyUsJU3DR4znyWa
EOR8szqtg9Kd2yMWnA2UgFohwEFZIfHsJfgoEOYExNmWtssMD8p6Ykxn6b7MvPJp
XLM+N9AYxZjX1rlzFK3af44K+9Rm3gVetbyhByHMl4bD3tFkhTZHVSC8kfXuu/t8
z2Q0qVPVJEjxn1wVvwShEqPAG36zEeCVBwfxtp754yMdz2mB3QdlOofY1t8WNReC
DLKSJqGU5FJ591UtGplLk2cz+HxEDrc7rzXaxLh83ecr/DhlgJ1QtEfUYNiymA04
2WhEtMoPBys1t+NcVb5LjZrxr4/EwF6qciLg57w/4/Oa2tOJre0eJxncUnefoxGs
9JO66HyryoYCfPt7q/OL2vUpev5gVsf0dOd/EtbJNwHOopOgUlc0qXsPSan2iJn+
bvDCaXn9gFmJyxvBVMym3J2Tm36cg7Kx5T8xsEtzdcnBqRllnTOcSa4P5LiK8ROd
TOlVnxl8S9h5aszvJFCyI5dj/EOkbQZVwWbtczgiNhs9m4q9C62DmBGuu8L1jYvB
+qCGlLYFylg+h0UXJz3Cc+GKs7Fw9JihWgIjZkw8joifTGIysMV7lqxJGeaVSACQ
zUv8aSODlkfqz57PyMJUN0X3rFoFG1ab4KidLpWdT+3Y0ynhjrLJ4/Ubl4EYMWiN
qDJrq2IUA22tM5sTk4qUHUhwYPT2E5c9i2SkufQ2uqssBsSC4ut2hvFH+kDzSMVB
brRVC5Dexe3r4J2BVl0l0jCc3CAG1Y5+x7PnyTlLeEfGGVd7aaAFpoNzgy1zbNDb
apQFMGw78PE6Mj7LL7llxOiIpp0omCu7FpXepH+qeGRvlW0Wbs22vYpVm5XRZlGZ
4IhkO1PLE6cb9ahDDrpU/CE434wkiLXLZta8lC1iS02/qsReeb2u73UaGUURPf3a
MX/OkUygvw2ZYWDbCd9OxFyv0z87Qrw3eIubF+fspMZ3aBQhhXB/8xA0U4y4uUtu
CFchDEfVYI40wSIy5SCSS0zrMJslOj6WWoACWETY2OXyIbsAnxd23Mj7GB7jA3O/
HrN87wA9Wlbfzx9nSkhnJxGgegtI1MZA6zwVXLeNN7rDGmfASofkUpBsE+fecAFJ
IHPzSODmu9gP7imN9Gw74bxMmZqJyhxS3NQxAzv+iSreuaPoUYaU8aWBqgxXBOiA
TA30PEKHnci2RKmmnoPMzPNogF8TVjjQviVBi+8Dams1TLfq3hvmRY3EypPpgyW7
4RnxX2uOLWfNuMdO5gJiZRj0nua1v9UdU0acsX9u63CSrZmU2VACzvZWnjxB2QgC
p/cv4tWXIwAoYFdIseecWaQWVG43xRfOwgJJgICsGBY8quf2j/s9wFij6pk8Fimv
RwTz7AO2yp9YYatXQmtXwQy9tQj7/cFbMGpqxZhp/ikqN3WGujBOhAuhhQwf0k76
AqEKq3rfxuIL2kr2sBWQpgPBv+r4/C0EoRUrwT4zgtajgsb24XoymAC/BReFsYRJ
7n0fUX85ptqHam2Kn/Tv4jY+p44lJeqbuRN3x8T/URBdSVLdVPeflmT12GUiekRo
I5DfraxVIlZKNEH6CZykweupJSsAkcEJpEymnH7MYIHNw7A3TMqG97OSf0pl0WMG
t/pRphpOCFuzJ+o81T7boifIYy2DLQlPZ6N45Gh3GBuldPlaO3FllQY+Hvtv3qva
De4HKhGqAb7PFY8JCbAs/MHnNy9HEVm3uWmg2sAQ/qz3uBDXIRIlVGVY8q8Q2OeS
F3mqT4aWJVncnqpBVuphNj9R1wk0pzo51UVLc31PpqHQLOx4jxqot5N9cmIY7kye
KKS+ARiVrf4R3Gdx0nyyjDkdAqb4w/DCtr+1aqUwju550+8ioo3QbSC9scxNvQXC
qB+zL1r0/jUInAIswcF0nWrmiKqzAxiZXFr9IA4UD+RE3Iw8PZKqKz0COEZqcxb0
kHLWXXEH/tmei1uEg7MYh913OMbYNp2/uUbgaAen5CGGDwSuLUw3NjHEh2rTbsC6
oycluFORHhjBI+KJHQ/qoP7mribH/zzm1DbQc3y52JjgB9llBlusy43+ur9CvTAs
91uHx2GLwLpt2GBD9FuSQV8w/CD30m+/qcAHMfSLDRoQW35ldLnmSV7oFFAPURYB
SnxQELO9ANUQfJxCfpgu/xIJMZ8/tE5SDYpiBQzAwwlKRrqAUntFhM7/6AfpcF9o
8vBf22hTZGV3TGH0vE+vYr2RLC+eg7axl2aUKdl0TYEp7LwXpJ88uPwTdpoI1Zzn
7OdR/H+rTFUms+9R3CzZHZLBP46sU/T6Q8cnxompOU74uEHmRqcIEyPsOEI562sR
BygjJjeOSW+lizNu0PTAwFDStaHy3YQzyPqXpYFWDbrnLDV7EpLr6DAgHyixoUK1
x6qPrkYrpHogKnZGvYmGtJGhSkxOnAVqPrTg0yLSkBTLwrXbE9I2QaeaVhb9Qx3U
mKh4O+yqnpmWhvRC3lY46GUipkkj1MxbM8zqhX7ZUU5XyxViBD251Ianf8SNTarn
UqXxdJviWeBjQV0pfmE4BMv8eWEV1NHi8r9Zlstg2v/XdhQuWrXb54HKGyKdtqgK
wXqgF/mNFWfFH21qUu4UK9IpU4wPy7gVa34hgrKvA5mXT5dCI+tuCOHovgRp//Bq
jnZcqZCsgcfjjT21sBG5GvgKwiDMTpADUAkLUK89+O7A4f/zXgk+LLkH7YWTL2Ub
355W2X5C6DN+9z4+ZI0TuDnJpVOXmpA03GVtCHRg8+lEOVXBB/ieBi1zyhygNidp
0O9eE0fyzZFXLFVJ3wQ4YWavMsI6PDyCXbdlwLm+17DQp3rwxjdHF6jLTkcpaJe2
B5bPYPS0INaPx5HbPP1D6wijmr1jc9LNIpp7eH5ymk8oBpzptycNueN2lELN2PNm
q18oNm3Z0nBGSFy+Y6yr1x4TdW9+OgdrZWhfUzXuifkdqsgX2DwNuHI/jPz8vRrl
7bi6q+middroDQ1u7iaPD1eLh8yk7iIOs9kSaHyrRcnoUzLiBjiOyrwHR7qa9bfk
8g3AlrBiYUmIRL54qgNWnELqSTXJ1TD3YuNx6BYfyG5QSPNPCOLyP5VXpc1zGbCz
j4+HlOq2TiunJX6sWRcgG7mfBi1jqfty00AzEibaOf54qKnYSvUKLvhyCKUlaAjh
q3fFnbB53ZbWOz7tIcGZmI+FCfU6aCIfn6A09IS95+cT009Tqyi+VB2thT172TEc
bQQJaDEUUtGQDFPQ8ikz1iE5sYB4rgU2LDDCI/WHejEB0YRoU4kbXPLRQYciqG8x
T4atme4WAZTGnX3sTk1dgSW5NZriYCETylhm793CWYJHeXqxMPKt2dGqjCULjMaP
Punr79ZUMWQAiGa5ZHGiVDy4OJKncL6KvLCy4Yp6tDQP8Yr4H/tiV/Wog4nYv6Og
oYObBRcRqDSgj+sNa5HrN2b6DEJv2u9ttDUXi1glTQdxTY7rjoO4tMKhaaluwJji
YnYqxzTLPHFWW/q4my/sDmdoynJiWpUZcGw7NgLsBa4TP8IAnB/N2QNa2YgeaUlk
ZA3vyTQ/VM1NtuD9SZVp1QYv6Mc9i7niEwG/O9OOv9Tm3tWW47b+116BWbFfNdZO
qkJ33MffUv46LcZ0FChwlGaPg5Ps7TEUdmBtADOSX5lrlJHGqkAkgmplvWL6oBiD
bdfpp/thTcMRNf5ybcQ16RdpmaJfknXj6ZeRnqJskq1mmMpDa6oDmwfjZnVn2R2h
9kDZJ4kHBhs+f60pEIhDrM2PVhK96EcgqrJdvAgx0uzBAFg/K5awK7+R8k4UqnA4
d0flvp88V/rOQfFZvARqPla9QLQhPvO3qXMtLVxJYcuRgZ1Hc/2Uzoarm7V+2lBC
MEw7S+OrkhNG5kDQN9N3iyjh0nSz7gIb2ZCEP1ClR8tSNOIOfxjm137wCNShwlhk
lZyrfITLxjt1EM069bPmLmUThK8QfdsqzWwfEaDUr/ak/xU7kZpl/VdYdcZBq0ys
4rc2cYWzVEWvzJhutVzT0EUWvi6Tm+wwrCD4+qZdwWJRD3BfQ2RA7nd/TC+vIEAK
+i6bRzplwsSYgRylRePgJZUQQGWn1jgikiSf/10PTDJIyMPA5lP5oEj648n8HE3s
uEtBhAR+85WZwxmDcX60YKtAzbjWldNHkCOY2XStoQzEDPJbTG4xdC04iGvYRAzk
hgXgh0LS9b+Y+qkRETaAl911v/uowxD9pBBQMH2S2jHyFLnNMn8dLXMMpDWr1UbT
mxuSpfEvVUWi6JjB8sKh0EGo/vsok+hsgbaugU6VJopg+8UWS4VchCV0501PRdsB
ZWEajp1BBKpj9jf4GaVWHVrynGXnF4+YAluqqeFdPc8nDpJef3xDjmT0RaDQxC0x
BNEf0Y9NIcRq91g5DiNZ3kdKbRhRxzS0L5bEI0cm+BtJ6BNOVo2gqxYOkMaKFa9j
Ad9dUhEI3j3vVo+Bx+nR/SE2BxRSgZqpPOXjWdBNXjM83i31jf5I/9n4rXeHaUsS
2GmRCRyMmNi0YbvarSWhK3xCJhOdWS6ywdmraEeoYD0BaNywO2bthG5QxTV9hKxz
2Xb1V8paj3r7B3bhrugoVbV1xhtKIQz45rjXQyRcLA9CY0l3BIKkTb76DM3ki8uI
XrnZCOw6AG+yGJn94rxHkL72UuIsKIcD6gwzPCFyQtoCPzxCOY3Yclybm+51+6lK
wqb3V3L3PaHe4bppneeG7Ipos47ARlkkuKK0QyLCpB/vjoER3wPSu0u/3E4vJ8QE
1Njx7WdtCVimv7fBgr348JZKNOgwtqL+lklfwlbOZV1qa0zKecJVEWNmWUSfEH7M
YGOB5iFFPH3D8ZWTBd4Wp8BvC8U20lIlEp2UCCj0mZ2bUAi3oSzrC5D4boMEYS+z
koBSYmvXoFLYWPXcwk/8Z2xQN9iMxJmMum/H20uItasYVEFOWLw2cHE90suYTukx
dtRgfdU7v28Yy4C10AqHjqLu8psqeMsxbla358obGlVsdEAMet/+g5VqBzc7LF4c
MHwDZkVRzAwhD1rDAe1Jh2qTYK4+95WQyIr/OKr3fVvPIrPPjXSpaiArL/5nNy2/
HNDczK04hNJx8mi6X03datAMyuzaZxlIGs4DyVtlo49zvCylhwQpqmttRfhq1sWN
YnyUk6QEcv1E1uKYuXbJpnWf47Y5NODEAkXSgsvi1Kldp7eHAf7YBGtf2Wnv5yYW
Mu4kbZFSOUq3uGXFfNxyaRhtHwdAR2RdOgfyHJ0U59M+JEz/RxbKcymYix98hlVb
rStYzbiLIZWjAluQ7OBZb/IXZWrKERzyPP1VAKUjJsznyzx8A8+z8DqB8mvOZgaQ
tp3Wj2CxN7pHB3b+8epMl7GXaGi4lgP5WFsohU6Y2SGs5Hjg6JO8QPCW38FSQFSt
H+nPSkZi/eS7ghDPE9ksyd5MmJiNxrQxwvv605wfmaa3OrrOregc2BW90jeWH1Pk
LVD5o4Pv9qBRG1bzs/J+tw+H6mozPnOMvGblIXrhiDu6iRVtcOa1mpXrsqKtEf0p
M47A+KviKf2wH8d+JBSxB0zW57qNATtBYWLZZ3X3yAz5zBPqMmkIr9LFVQUDtzL+
bJ6W3+T8cPQxveX5fkPYD+Nbk3+DJC+1dqlC5vZWPIoyyvdajzPswMapbqQ7RBOu
WlPHCek6wVyrpw0Z1idCxMWuSSXbyxCATMEhuKHrv9H3cWBOxN/5IQwdYkLac3Hv
3TSrnuqgCP3NLx3KJRmX8rssKmXD/sQgsiqISnLkEIAkyDHW9/VXG0O/88+w+gd7
AtmHr7uemdIQ+ZhbwTlVmkEHMbxkB3hhaLDvbXtnnAvhhLOPoj43G0Rc2w9u/avj
gzZ3hBJFIGU17AMNeMYArGhaKWb3MjoKZKX/dhFl0Ylk2ZAZEwIoUPKIlbwQgDXe
sAvfiiGJmNNYLDkJqyspTxIqcW5icLf4YptXr//UZqOjhw3u6uUaaE/kKwNOn6FB
XVybVTpUtEar9e0GPM1Qjjfw2I9+q3KUpVRbYkRcOtFMWaVKMiS6G6eQGTn7/d5s
9hClFv2v7KrLtWEXSoJ0uWYx4ogXL32Rst5eQIP5awu4hxD0vepO8MqkR4mm07JC
rTqilFY/R43ZTOsoD5hYY0A871TrN2PVKj8BnmtEQ11BPTwZuNUiLX6gdGHtlv9D
NtK4+9Oplhfkam+mbR3D5Hvjxyp7rcDsWp+jEL2FXmHhxPln02e+bHuBNmn/33ms
MEFYSmgv0WIVhdQGBFXlznROQIayYGzT5j5fdXejgWoyZvesVNhE2NJXnY6bSlMP
isGyIUVcsAZKc8ageghOrZ4vpxvfgC7onzVSwq0R4HTDlMrOLELCDi7wYKN57hMu
WL4+PF1r9BjwmCfDHWjtR0ZOWgszOG/Hq3NhcJX6temCpBwFgvgSoz1w4ovvx0+F
Lnd/gwSLOL0Qt9vcuM7JrrOWliCzYxaSo12OTxiIpq9jFXfGTA09+sQWbK2AHnQ/
FBLyuwOtLKb3srQ7R0H4TJKa3mYSYlKMN9/hclYVJf/WSILfoWzI4QBmJQy7RV3W
idK/i7b6oRBIZlSJUv1twG0lYGNgk4vbIJPinHhLS4zk1u0vWWMAy0WQ+95QysKF
vmm+4yO/XpODKUJf4nfPD9g5tI+c3nu8JTXzVyVEvWrMqVjds8gayZbO8kN1kdEX
+QiEwNBbNj/Nd5gwUXaiilcA1hff99y4Z2mdBdKlUEXSsxrKuNDhmP9bnBlbOoCd
BF7VEkIFYbboq4qYgkwml+Gk4pw0lSMEHMn1gfsb+3aQYhHQ3rnVrdDOAzliYm0f
rsMrb/jEJIlVjlH2GtVURjuhR/to/pA0rEXEWC7ImBarGDjI6pqmmKwxRXXzbPm7
W/p5yuADUIE76yHTULU77NIzNgCiDJFt2eHSacAbxnEE+i0qL6/7ZFf07KoZcwPL
uvHlZC+iVqZM2CcgHaAGFJzLMGh8zQ5VwT9+ByGmOC9ksfbWzY8Vr1db0/kdfs/r
hQ9UI6haFNqRr/54FbQ3UvF8fMiRKBODxUG794b1NOP1Ta+BKzxRP0wENH+LoH9q
wcZQbMZ2E7UShZ3dv/W8bUlz8NO3aLlFXSlSkw4K+bGBXJlQSzYAWvAS/8T5SU3d
jS1pu905sjZO8T6ac2TrybhsHR1tdsEHVK/b+ldoP+MUucQVF+jXolo43iSsJROF
6CCTKZXOQdFBvBRExe03mLCePHH4ygx/e1mn7x9V4Zqej1QHOrvFjH9FetLYkkbH
V4uZUxAZACUmm7RNEUrCgGmNaGl9qy66tgZcqF9xmQAGSzoaZKmZf1AGBeO1ERxB
y3wtyKMLYch+QL2lnRomfJRYgtKVVREAedABjNjeYMG5styQhf22kUFTWThgq4Dp
mj/hkYW0HE1XLqU+eAd90F6dQ2gJI73TpA2PiYdR3MxoZDsN0yisRajiP/D1jYCY
PcCHEMHx3J7b7Hv2Q6vquYlnykH00Jvg3+LQzYLoGGPG0z88AOp+MT3lSNmy3AWd
1xJMKxeQ4a9pZcQDsmJmuJxrjpX5QBgfiGG5NDGhODXCJs+dI6UYuUp3F6/XtYHv
zzPjKI41S4X9Ij0fp/bT5VoTGCcUa4bOI4x35/uhBroGYGvn2m3pDViJvPYkWFb0
U0ZrJytBs7kKxwDw339hQZ/HQFfrJYCw9QY9HPwgaaeE/eEO98yWBrcDk11EQ/er
YnJAlfeqCU/qIb2u8Ks2W64fiOPy2+nJeHYbYNSNRgVq7G1zj40J9be9X58E2Kgq
fnpPTjt12epZvsBAiQXcnpVXc0C4zn3cTYuPt3vNXe3TTQgfawOA8NOSOyTnQDc1
KkNqyCLF3+iwX59/Oohxh9ON3Cct3gymp6WUjoxAMGgt8lj2Fs9YlyHDpvsHDmcP
FmRVhCEm8wLyBMc4p7pF0d43hbIVwuYKCxHdfISkLW+VbDW+rUWnByWgHW1fL7sX
9frk2WvpDdMakvpYROZismRAdLWXZSnlY+hh7/fkicPq02NiZrpouPO9hu4i8wSx
M5n7DURMhoQT8uEUR6YCVSwxAFCHBsGF0hYS5RGQfOKSdlIYZM63xDAAkKzMvO8v
S9H80hB+kvwS4W5RNIR9E4lGPVX4Gck96baPjoFUEJ6eu4BW4oBMJ6krM7FzG9Kh
6yukT4PuoQFSuAxpTWlzhonumyZVV2VpN+yKCq0RBqcRgisKmVXsLEpL3wekLZsw
h3MdvVD+AVEZWZupJ2jZl/aVJKTfCiRR0p3qgYUfcwtvlRMBDABEZkYRH2xydtMW
4ohnNTDZ0KyYHNHuy1tETy4ubeMFU7PJMTNrPNZMpR3Wm6wJGAtvumEWAUfKjY/y
zdMwWWqyF3LLZkDvxsynQFO4S5rYJeUeGk0+6ck2AcyD5YR8oMnDANfXaRb6DBl1
wyxwl65vhy2jHWxeqSiQhHYg59rwiqwQd7LT1gINUidAvpaWHD9FNmS+U5whk9XF
vUUAsWus3KiFh9mKV4umf0I268nqW8tY64OVtpChK/WK4jFjnB+UphlNZkJU0t6o
U1mrKX3dIJbMKmY0p2IMNml5DEUYstuflckj8w8AhoTSxUixScLDQV2fW+Igt+Sq
IokB+N1K6arTGCETPesX2GVCwY8sF+6H6j+HRTtdsOo8YS7hjond2wEg+ce5oL7N
u26dxuVkey2zLgLYPLCWUlQFcCUO3bZmmaHsMmSBQ3Ugd+Mm+51jRudqnF7lYfC0
guZDwaeV33gn9T+445WAhMCzjP7QEOg+ZmSCpBpj9T7w/jtTc8DJYoDAlkGweUvh
Mm+LTcMYx3hk+PZ75pecQieCNdY9MUABgrCLjRjjfrSgcOw4dsI99Ac5zcoL0o/b
KmT2NrU1pfmh0MLDXjeo2QlFsc6+SKg6vUxF8RWugDQGFFo/L8ER0/OrD2z1AFcV
dtcjNNTrq/O/Phq4DEpTuKqlfimnX6JfPlBtdS/V3EoUcx3DAuJZIz3Bv8xNSkto
Jer3jOk3TBHAlr8cxhdYWwIgVrBTsKUMrejoTvDug5766EoON1a7FY4XfTj2/XWN
h8v55fPZK0aYMsqQU6JdFSFI13hnS/p03hX9Abn0sNNlRmmMIEgsaMGlOf1PlSg9
kHOt6nBG4/nLRYm/xzu3NqKzU5gE8Jo1Sgewg/W0CLMEiIS8tTDM1JH2MsIorHak
7sE+FWQJo5PosWPdQPicKNckLRrjbvlgOf7qWIpl2oHxe0Dk2jkWYlxTm1+koc3f
DOBBq4aiynBfEyysB2T+AC2E/T7L+hXjb/RvZpPCo0+8YdTz+baROO2hbj/D/DdY
23poWcxttb6DOBKrpQv2MVLFmCvzli3+omMl4IUZ558vAH4z5Ni/OGLJfO7h9wwe
l2xlCXtzzXJUnL4b4Dv7HgMg2Wiv+fHlbX5+9fit8AR1RP+jQ3mtQaf5dSecthki
E2AWlDl8jy/SY9gsAe7QUrOsLKyj2YI9Lo6/OoAbnnvPJbkIRw3nbint6U+HFidL
TZdzhRlZ6IjdJbVYAkN+6PP+B1Oa4oANyGVvffYyT3hUp6h79nSi0PXs5HUR9nVs
03sB3I7MLhWdmRC+Bdd0GoX1p2aUE+Zq+S6DawdG3DbNjCGhOt5cX+Uivth4c7xz
mtV3xv4YHpMpUwb8JwgSPCurPtfTy6xZCxov9jjWPnNd7mu8YDnhNj2hEGHYmGm/
vJxS+SVOah8pWwTuJ2SV+hSGzErwYgQ+jb1wZkD9xW4fzZLXXTo9GQ07qpjd+3av
C0kmIseomYaD3ralHcUFCBeO1Os9/9iyA9/ZwMYxBU7eYydecH1gmXQwTIrZkCsc
nUt1D5XiM3efCgxAhBCywsJuv2zAOWcvhNQlVVq/kyTdAeK8typoI4Y07ZNCGmBX
0txFeWb2ZspeSWFRN8z8bjI4O7zXDwYg788aIi2QZnB9PXB/fetoU2Wx45ggFmw/
3ka3/dGRuxaP7wC4jnAdgncwKbHpcRloCzm26NXae50RIETI0Q0T6OYy2yIaPCBj
zGFwkCbbh4Gu07jun6smhqh5PtsIlmetzrEh+OkQhkgSlpcCkklHjTpa1hZZa9O1
GCwJphOXp2lzCa60fzZ38V42knzFv6shpKHjJcaD4JHcukqmNdqHI3pYcB5BO6VA
fIsT9JEiUB7xXaRxCSNLfgvhJ2Db31gggFqMLvZHNWWUyAXH8JDSRZ1ge2JNIijB
Wi7qPPB+iam8KS0HPSVsn3Jh2c9fon614JhScT185ofcHPvrHuy9YSxY3gAZNLCj
dM+zT3OAPfgjwie2IFVw7bLStpqzcjWjTk7oxBIx4OESHMtrr4U7GisQJ8UWp2hE
kJEcR83w71pp1Plrir+/5zcFnWgOItZEKfcHDGE7vmeU2WpGVnRtUqHK2DvNKzii
O/L+6eq/Pze6n6DYqNk/ziERi02XetkRYF0p4yRIqzB/UYLli+T9bGxzt7cP6dr6
Yj5TCp6tVdKR88jbK+XOkw5GVrq0Kb0hOOcl09sQ/X+gkDNoho8JotRlF9KXmyjc
+W3BU/iI8JTharAuoHL8rdkUhil1K+R95I0HqmeWX8ad7krExZWS8V2+v3mEFp2u
r7KdOWeZLXvEVzMfwJKRiIHTgVQ2SsCo/iHsUBmB/YSKBGS13pALPLheGXwtH1VU
X3OBA5Jdja2PibDaMDwIXMJgY9XqHFn98BaP/hiT19w0d5vcbDFILMgZr7+vAVuv
bXJ5O5StqmXO9k/lpQTqyLT9MgvOErVtO51qdcJa/+TIu+hZ69JUUbLtS02DHS64
rFY00/FP+wdYaq/jI3mnwRTIQGcvOQx2DLUlvWN8ub6iEigP8tgwnEKkY7eFJQfi
JUBmJe4WrAo/mL1yQVGxT7Z51BN6m+r4fdLPagX3LzgCrhEcDhF30AYb0KcAU/5z
ih+3F9gicQcnt2A+hTqQarQitIbadYbCtKFfkSpRvxZ84Pf+wpRQ5+y0OJjNdj48
IWasdjG/iIgA6tWXg9ZAemacago33Y0OY4g9oAz456J392ubRXKHSBrpz6hqCWiF
EhKGQHLEc7LWUM4aH5E+j3fyyjiUdFBaP4hBDIYMqyQhB3JFj5fWgiJcZi90zG4q
TsaUwylwjCJ+o1Xc2nHHOPAqGkYy7GmtO7Cub36MT3UdYttxusP+UriQ2iqscqdV
4Mr88F3lwRX9Qu3FUa7gVQkST8WneIDqNjr+09E7mWprPUWacaPSx8wlS2VWewvG
9r0V3GWgM3HtycKWYO8Q/TWc0Oy5a4AGHJJ2SKMmOVXsexSV+Lr4vzhFqUCM+q+f
/YO0oQdarPv7fvCjiKLhIQeqaGklWzYEuePo4J5r4p30E+I8XoSV/hpVBVjJBeHn
FAPEOSqISpesfIg6bUQW2kIH857KbTf2SDa35PoxIhlQQF7z+wG6MWNZ771M+rJ/
VWxYSjqDo/ZTklkJoTFkPG1XQpw5LBLrqdbMjPNwPvRGhQfz+gY/2aBYke+sYUPs
yJmJAU0ivsdETcAPfYW/QADnkvXSfMf/tcD/jiickaEACCN9prdcAO4a9CS0l/hT
ANeXN/Wy13QZGh7gPvRgYZCfqSxGW+4zBzSXxHS/MK9tWtLZjw3utsOSxAnwSM6v
vuTORmXYI7JPPiQoim3J/AVgABvco7lkV8eS6+X6mBexVB2gjU/M6lR2CQo6YVhV
G3YZLEpjxbvqCjlpIZhN340eKs+KKjSq4AO/0Jfr9FUqYd3RWxMcnO58eMysBVOE
lBMipcVR1NelsHaWc4vb51ncYTHnPIW0WEvmfAg3yQNaj1E2wzaxi21qHNGR2jy9
CLgBfuiv4sQSxIgXcPsInlXQAs2fKj6CjUiew9xDNT85068RJjj0C1SUY9BvzqbH
zZ3wTFMQqw1oHZ7hnY/af+3xFqwH9h4Jcsg+CautZbSW5unl+HDkF8FpLdt8rdoW
FI11VfpAxr52avAb1+lY28mlylKqz8vl01OK8Bl0pH9aGpDZGu0w8MXfcERWKmFf
G7BzkZhjKYRGNL1vaYNm/rPIhBB1j4yx0algxUcy3fwgonc7eLG8txIfRQeLp1Kx
hjliFXnUNNudB41E+B6h8YxR8BLMo1fSGYFtJqqR5PT34q8AAo+1HNboQQkOv8Ba
wAXuj/WxRExQSu/s4lhiTDUvIgnuh8TMFhh8EtzQh4D1/vMZ/s0dEHhh200YTrbf
tanWFuLUhCvhgVeiOshqZrwvYs8VaYZnuZpjrKpznY/qZW9RRwbNneV4i5sYbjzR
ldZyrt3vhqlQ/2hF/wxsXiFNOKJZGEEA04DdMzz5ZApZDnMH/DZYevhOJeASbUjN
bp35vb++AabbTMCfSYaWQXWrwM6qOfQQEpv+mTGnMrjc+Q7s4mLmXzZA1/8a1jmt
+elea1wSYRHz9yey+hKYNUMhCvnE2Vybu+l6QNxks0Yr1Q+v+MZgu0wIP5E/LPkh
SXUzB+jZrnGh1nqeZz8MK91sg8vXQkGf4u1yUIiARvWu1GuXbybe6tAAold66S/L
W+N5ayoxyxMPAC3oNcSnJhPOcMJ6P8Mb321yLXqvPg1X7IfZf6Y5Qo4dnqTWMvMv
WaV4nl42vkz4Sj2rOs8pvV/v4FQU9yenNLlL+2dLbUlpL5okxggZeGwmrpJ1Gw6u
8hvvdIwcjVhFLA5flakCFN9Ihm2eUIE05F1+ORAaiDc675Y58z0DsJTuqnrbcmAM
1FHREiX1SGlZoantmYjQzpYLxdnurxrmm6RbW34AeU8SwnrDiWscN1nuuf21cthn
kOFuOihlcO+hsDek4/9TTU+RSeVDz4cxwUI0i7bxpdBudGHk7ROayExIF6hcPix3
HyQVO+ovQVq0C1vxmzNyi4v8K+A5hX13ihez2plZIVHlDlHqiCVvg20PUDAJUz+D
oTmANUKGrz2ryFKAnGYIWWSFk/4W9JAaPtvOrz3/FfQKfwtwled370oNgYWwx2+C
GnO27FzVkGoCM/q1wxGNHCbtB3v38gSoOFBrdq97xbsaWSd+FJrAxpEG1IOKnVoT
dEClQy7ZvWdqVyXrvwa0FK5nrKTQQAnkakQDEgs1gkBf//QBvKCFyp6KxcTgjERw
NblYCuAsrwyw3RZIljm7osuGQFtBIgUxdrzeIgvBegtTY29RDXylYPm17OdKEX2e
pVYqQdbHI6ucNN62BoZflmjqtSYucGzvkAnfNKsfJMDUNViWei/lnhGyUhAGj2pd
BfLRX0miev2PxuTdO1GHf1hOY/SvBtxblWqdbiTfzvP6DWyOGE+sqqSd/yZFI0d0
P/Xvw0hKYlHgkCqUyQZsb90pLUuBKeUyvM0anaW/Ha6XBUko+qituj/5az/5abGd
phXUOYICo+rkE5IqrKzbcAM45hyMpuQZLJoSkrdkT82CW0e+gwJZqAUMhZSXzjFu
iRxzCB5k82IHki8yJ7ZeGD3Bi8EBMwkcfa+pU4Uto0fgq6oPmM65EzzOQGAVU7fc
lxf84fqzUSu2TAsGVIPKJBQZOUBoMmeGuU3i2hT6/tqStdLsY2n4oHpuychnq859
8kQ0BpL2eXHl0u3cLgsCK4C/C3MqKset1nCFLVnbp6f9nsT3VjTpvXR+n2C8kVAc
ZE5nl5uYfBYq9oxzIh6ODCS7lp02XmlPvpUvQCrDZRffqDmf6tnYnosUHqU9cRlC
WPqE0GbcuhJ2vvo8wBaWnvH3RAkcGOzUj7/Y5JcydeO6eRxQ5TwQR0cVx0nozocd
z2+1wuCcmcUXQxpz0tioi7ZUFMoPACa84dVKKsdTdVOp0cN7lYjm7US7ByE34mRX
ufH6IQryQwaAqxV9MWNAh6sDiVBvewqh5iijyLYecIRdXAMdiw7uvwtP5ShoezN9
mjHA0nnTtH7X6BeP+JYzVgkjGUaz52CKZpKZor8GKBgK/B64HCxcAVGBdRAGFGic
4sKZZY0ZOrK32+1Cdd/l4mDe/YVMozYpd+lZv6MhCB415d1Ve9CtWLbAXSt8Lyqz
qHq797oGy4P9dkEsawKLFQiDN2WNX2GGmTXk5S7hWaxfs0O7/loKLE/wgKtI3ddP
LDA5l+iR7hv3znB1JDUnslB6Z7u79zYbd9i+ZHixCwn88VfhAAutWX9tUmIHpmHY
A5LnL5jW8YE2Ba7MtuRL3v/hBRocw38aQwVi88xOl78V4JtYVtqK6rU3lWx+A9qn
+En7L6RBfIdqCMVGKuy8fpAot7igewKZGKB2A54I2RIBGNptQvnMil9VEK/MPTQL
r43Q5k/S5iinYhT7KeaM2RcBlXxzMPy+xi9mG+r2dd1zJFrR1660N5FDqPrrJkxK
R3h8Bn2vmudDoNrMucoOVgPQvKffM/nv1SPGwqMArwStpxKKhexeTskIuc+GTEPU
qcDnrO5EvNSxVqAsOkDsLmO9+NFc51H1uPMbkB1ZRetVDddj+BRD9z555rQ92+ge
TpY7Q+aoUijrcAml4zne6Gj8Nm80jPYVbftmTnkZe5/pv7rFHPK1ipANWh9pEvvc
O2ZA119u/cC/wi8UcT8AoLR8gTD6v3KLDKEYGJKmkG9thHFUp0mKQuKcQfhFvMX/
BA5O51xWsySXAt5TZ84a0Zvx1SBDDIPQMiOAjSTsbgLisD6KoIVo2FBoNp/BKRdQ
EPV0hNSpxCar+/CmPbYXYpTMFO0jRlROh0XvJoK/DNdc05bhq5pdagqnxdYdAtkE
UuzgspOVMlT4PeOzT0OlvNSpU2dIwjvhLRwnwkO8TvwWZVbnIbHmK+HIYj+ua7s6
I/73UU5TwQttxR21dchj3Q5J+N7pQobfwxB7X7mWvzVj+W8LeaJH1LmtWZTsy01Q
s8HOaOht/OiQBVomKaPHXa5YwZz1H5DQVnmIP7wkXOp4JgZrMPo3Kxw1XD34jNle
5mn2lDG8X0vOuXE/WTSQTd84TaD3TN0WiO4XcNJ9pkr8NvQqx/omOzM2l7ynRS3f
7WuLRoXp72N2adoUjMmm6YifQ730kBKcoP7gWqHCWuN6rSaM6WeFaBYyYKP92Ho3
4fr5veEtFsX552g+SxSalmLLHpin/WRT2Ut8HObHyNZa5b00W0SiTNIF1wAIFzaj
ygV6h+ApLlCvyI6jajGu8ki4Jal3iT63YkJOh3Xbn7D+fcj9fbhd340OBAi/kazo
3Mn+dMMt6Yys71vsy14vcJyo5PoFd1dHTqwMHp9EzCizPQOvSNPhmMPXKJR1F9uK
w8fl5r4eR7SDhuYMpCMurVhGVwP7qu7yeA82MoywtGiZvlR2OPxJrJvn8VyCZnMM
TPLc+uNrh/KLYNu0aLRLfqUfvGV+qxN7S5g792nNyY1g6TCi9hJCZ8amFyXu3xR2
dbQn2bGr6NRrx4O1/jP0DAAtNBXgaAd3dHvFDCUg0a4Uv2IUjmyI/foYoCyRX4px
H5PuEUIS9N8VK69hwDz32tKW+fColeZwYD13e6Kt+YaPfhiud3qUzTGxwybUv+6r
zyq3G1Rjr0OPnLFeZzo+zM2m0vC4fF1xblODGxAY2ZgSROg+kRsl3jQHV0ph4nbx
oWpR0c+J0iMCJdbBY/EPkNf+N92Q8ootQ/7/PEjBRTmz9rc72jWO1DVvNrGJPDCf
qEn1+9RbL6k7x3gGTdR9FjcBF/Zd7v7r7YN/zU8IpQuRoRoZjEnaHgbTUW4TUV+P
XMzNDP2cQcf/E6oqwfBjb8SHUda5602Mv/iVeMlmWMbPxQGaNFBgk1piTP8YFdVo
ZoZEqlYZGkgneCOFy/F9dzl2fJYjoNWfn3E1Ddyb10sLpujSpk+WyG//pSn0r5+t
ZS7pMaVb0YfqCK5uSmSlAg3V0oOjPkyXiM+Gq5AIzq0uol5sEulGW2D49/2knVLa
R8FiCvwwMvjFTLOrrHnlS5EXKcG1cPUIivk54a2fOIvlPt9Utneh2XLx7UqYVK8w
/ECLkeFeiGYO0HSVcDmO+ocyVcR84XcFU50RjHqH/B0uc6Ux4+CVk8KezSXiPxeH
lrsALCnJv6yepYCoF+AUoA++nAc/KEE2OrDwWodFm9mPagpitqwOX2u7JMkd5DBe
cnOQ0EWoHaGheEI3knGkpnsD9HMOU95KwXKvhHjdVvHhjBgkzWYnmLzP5gRlFztf
zkYZ1JE8ZS7z8sibT/omk4eGW84QluxHSQkDeK35lsqZgPM8k98WPq35K3APhYSg
ZRNpORmlMpTxYGSZtxWwaIQwJchO5q99f6Fsb3jSNThLIjBMQbONkF+USsJ1zv85
W0qCiV3XMyme4XT7sb6ta+BdS8nlCHvVH5YveYcrjTwrD6+FYu6qVsxTdsowC7Xb
OuE2u0PTYFEf2yUiRLAsN3WcVB2QTvSzrv3I6e21Ar7sWxD6R6PCdHczNLSGCJu9
CbCFd/nOc3Pc3eCaOkfl8o5MPBdHd3XOoPTnNsVkaZ6aatI7V8ILobUS8QcPzU9E
vcQ6P87yk6wIcqj1tR5B1kEonfk/EOIYFKdQRtbkpy7U6MljxLTI7iF+URuyduYr
C6lK99JMHF4ZSABTLZ12jUXrpOfJm34qXUUC/6X96d9bBu9hw2omSV7rK3vHg/WP
6C5EXxNNYSKfyOqmJdP95autIUEA6vXDZcfULztK1n8HVdAhgguT6M8hz2ZRTUIv
iotBezuNZJj8Vlfc8J/KLbQIyAdHUoe/rOKGRmRKMk9tTTeP8TtBwcq+DY55Hhpo
ct77GMMen80R/CZS6OzTdg2HELopQU3xFgqFcHHd743f8sO8koaoxuIkasp2B0cI
c9RgWWJBKZg9erB+mxdKkU0eRb1Aq2PLTWzMEHYcNSTwJjwTw05f5urly8mwhDkX
VWUikydhjWHZWa3Ryn5TSgI7eKfP1Rwj2TjbGotb1Lshjju7ABTmIA3rizjt3CYw
xd4opMxaDFUcz8WX+dBS7VC28kT76V5wiUTrtkdGcyMucBpilcdsQ8N7sgrVqLG3
/iots9j4vP9+crN20JUTivaKt+4o5z1Meqhc3EKk/j8+ZUXBz/BAuQSk9lyjvZe2
kNV03AkffP63VKkcjtOedCJbBzu98Hd2k+EQjKDl0IvFT/YO2VS+9C8jUPX1N9jW
xjHa+fETh6GFTpZWsRaYIQ8EEI6Qn0K2D71c1EW1+W4ye6ey5qO1S1VmKeuDY4CJ
J2sO5c9an0TRlKejyGlJGAQpIG6S70Q0E+Vaqxy9Pg/5xcl396da6bc2ZbI7o+ic
isW3kh/CeMGHFeT47f84ckdx/0RbcMtqQR4ac9A87itHNZ37He07Tl5lTLtxFI76
eymTacQSszCJgLIUCn4SfGoEEvPZBT5HijovGnRBrDoETyEne2ByjEBufzChfUEM
8Y5oDa5ljhTWvJKK+mKmmWUb0i70a2Wde0helW5xMbLY/SW4pP0RiGAP2NhvgyFH
j4KuImuCcc1hRmmO2KfokvgcDlA0yFvgfkiAlKkUdR+nF7q+UkxdIAEIRuhLdkZd
Iv7F6o9wZeJIFHj71X8rELvEaD6foerd+SmLJi6amRZN090v7Dc0iiBIwxDal1ee
+2OGgGbtslsmDMte9YyTMp1PJh01cmxahpA3Vzn4xc0U4iwrNcbln/8Aa1ih7AjV
+mQCfrMwHVXZ6di+RUKN0PjxaK1YM2ULR5qco6qGmvCUWXjMhT6ZkbhWW7+8jYGj
leJzMGo6MaDCYHVc8wXPdGm0F/q6cxtEeA57eU452RZ2v9suaVIuYwHpVKN8uwzh
INlRYlEs/bcDjAUVTVlwr84617ILBVTDu12rPnoN6zI/NAuNTRN7J3mJsPSK2RDT
Wi4nfh6cp8fMwBrfhodoV/NthKs2HsCSYp4gex6UooHn/Sy8E+iMz0B9xaSJibYK
nptYzqijh2/veU7F2oziMA7+DqjHxqDEsGQeI9JsXZn48HsuoalnechE4cEmdHbF
VzR7mIfgGyFzeOhGqPYxAKHlJci+Dyxr/yEbCXSK3vK+jgUXtQPrrOcqFIoV0nMy
NJFiklRlsl8DD9OVHMGr+aZAwy378cgwxwfSUUxHURskwEywryo83KIY5Xz6okAR
OP6AzLxMafDpI+Wz04yFlDeLZV6lFpNeElN35fqkI9XRhYYFxOtqpxo2afoCW1bm
kg8WxN6x74yQOpUGdj2UBYbZJMtKCet56pf7u19TWC/BNxlxYCvH3ZbyWv8yd3zN
0gK0cwrqb93YbRv72jZ2ewvPH8kSUSGbkihxkfALXyQDBzbRkYZmHz3ZatVjK1yz
+B744g/sr5guWN1S9EI2JDfTOSuvCDZ/mXXJOWMJzdqNAtyRyWCBDLcFv+o6tpgE
VRRDV1gN3wb4FeT1wlQgTZK5iTzlQeaWSpYhoXQHvEJInx5yipPnfGdT7s2VHFVb
rp0iZRa7pqhoU/CFYneNUzaI8GW+4VqTCDPpv5ziKm6TJdWniZFSbEiRED9BJO3k
oDulvOnySYWNR2cIk18RHzeoiFeS4CWM9JP4j93FdjsOYFV4aV/Bu4GIfzC2RWCX
EkHWumTCWCuVw6ED5dBULOjWmivZGHOVjb09hD0H6yEQMW23WIS1CnCreF+PXJAN
OZJ/0s9NSTcx541IFbs5uoDhiHC1FGAjiCsVmL9ObFJFXEE9vnXk4DHSwCfO9Gyv
+EW8LTc5NAxjxBXOy8kucsV9iIDtSLRztMFYIEqjm2w++Fi0ne2LlNX+C4sDRl+d
AVAm+/F594TnJXj8zsz6vK8eJqONpvrirRG9ivFXPiLToShfvJMlB/WhxVpkNybK
HOVsuWU8CdGSu+sUcgVpqE6rsou9ubaFzCAdnraj5Py31uqYADFPxvUCrrBEky0L
GtQ7Xgweed4rILkPPSBdYe6JMhkgKKDZOEwEyV+W+0eFJsEfgBpobNksoSGjfFP+
g/b/DRg3ZSmCRVNCFPtmpSIbi2xwBJKU+Ff/G5/Sxga+/M2z1u0eMEGjdYPlMgwk
Y5VyC1HR1VFha95EcbT2DqZRctvDh91A+oheIPhrRR1AdYO0jzMrsppmFtnLtMcZ
oePA0+XZeFrCRqEOT19kSOxFmla1lK5OPWiWSqXJWeGhH+jv1ym6B1bzFIPU+wte
iG3fY1LJ+HJFz3Mc2joVKJA+mnfhKo6bBe2bX2z6Z92/qp1PS7f8mLYe5087AsnR
cyAkE5alIhmCWo3gBIBmUtTtPvwvGdtSHqgWehm4uWI2cd9EV7t2MKECcZx8/8eh
78kPjGb51/SDpDS+fQCh7t0iPWZNin7rGibsf5+HiLUbeBiAmPSkbMjSLOj2Sngj
oxK7jdABQa+dOAHKTg+oP4ZDhWqu3l34w2595kL1Ljy06t8u9h4OsD774El/Ubgu
YVmvitGX76MTNNMuEfw0B0dumTwkY8S/famqjd5p3z2saYrcGwNx02sGL7naEBBy
G1LR9oYBdCRTomzb3WiRxbZLBS1CRGmm1fgeLL3rEXZrvkB6J73cU+6oOqePnPl9
m1ZEY35lvHphXN5bS0pqLPOI/eMvtfEUEMPHZJSWMLAmBBDqfRjnfUDZgDG5cxz8
XT7G6Rts7G9jwCBaft0ePZIz6dFRrg7Le/MJIYrmrEccLGosd0L+c7Ya2YgRABa0
JNNpsPqHPFdJXF6gne9ahGeXb29+IhJsa2DRYR/VePeBM5B8k9PorQoQMuEEWPss
WI7W0E4jumVSf0b/o72bWlrLnYe/Wlfrzz42XmVoRdLPSOstS+4q1zQPQWc22kLR
EBdAtG0yFtyEQTx1P7+MUDmw9Wgsso61xgmWWqjrpg+cW0BlRnUeU023xLWkF/u9
YCIz0afRGDrBfzHWekhb7BDwkj3H/vLDA6bWq68NgMSaxz4hdqNuSrHNmC0xYV2c
C3BHD2TeKYvMqBq7j+xGaJ4tb0urFeEv0u1ThaYciL94ye6a4oGCR5JwAeLjaVFc
xVyrZC8TSX0gXCYlEVPa8yckpNsLOyX8AIgETMPX617yfIQm0DgHppACgirIJLSd
Kv3S1FCfD4W9VpSFQAeLd5C+sr+t/KkrgKFx1cZtaSqthEaRXPpmK84Hosx4DC22
loo8xIJSw/q9ly9V8ZTiR3YfqOM0MoiGz9/kj5cqy2qPPYk2bzJxKZp7MDdILA88
yI32m31M3nZ3mQJaO495iz/nUOSH5+9mrSJgmZi9ilICZMWrveUJ7gLWHyjDfeRD
LYl4jt3L/FeY6RJ0g5bJn9dBNzmDah4EGwxKttvGPbdL1BW+BnJ91DVyf82ezdha
5pYAfabeZSF579bfNITiWZfZ/TnaeH/28zSSEEGeMrcXhsMGenBeBLGCgWL9xCU0
syNZg5p5U93kWUSCoWr+3BfntO0dn8Vwh/KLSU8rAIYhywu0PJtnpJ6XcODmzEVb
XlvvCWkBLTM/n9OVk4FPMnfcFMy8kSUSeV8KPhMTm2sFzN4vfiBUu0j67s8XTzzJ
lohwJzwakCI6UeA0WB72rIgWAePxhkhgCu5N0As2c2hgL2yO3kc36OlloES+ZAdi
R16GYqkAw1sqxgIlWcn5Ma7xvw0SNr/gOC2zlui5UmFPJ2snfCIQsRfrn+CcffGV
XI27yzScxvKkCGpq0bQr5KrVm5Tx1tyGRkAFO+ERAfUCd7dOIi323tQ6+jpPuTFx
EqYtViGirV/n4+I95K3519sxFboqGC7lnYxK/4VgNaFfqJAoZqyI8nz2QmtJplWb
ruvTb4yjq3RulB6Qp3s39VJPv1QNSfFVD5BmE8OdCNSI0+H/c9tYTte/fgRqp+H1
+DK3j+y6A0S6oUoplBmCzmIeQ75Kvsmuz1LVI/r38AR+Rc6mUdfYrFvS0efud3XT
fbOTQ7OnPXYAF+h9obCdlXxOjkbqk+2DVYB4jaIruz03wSuJuaD8mwE1cMOrJIWa
kvOjto+w+sAtbbaCDxvu0IkLjYM+McBWaWzJSbxurLrbmcurQRHu51X4ImFqxZfQ
sgPE7G+vRWOs9Pqq0ZARvyPJZPQNC/9bUp5tJVoJ7hqxtC2HyKQmgzEuuaC+QURS
W53vTPwVLEik68kP0BLm3pTCwtQMawEsJ2XuwxvIBxAExNTgE6VfdZknvEX04r2U
DaBfOg5i+KMQCDjQisWY/liBxOnQaKKpKQ7evDDsHjgagRH+HtKLJ8LzNOPBzYLj
xNK5AUQgxy0AFWEAmdvJQE5MtOHKbgRTad4tjIW+cpNmSSY64Mn8TLkEtFWF8kAG
lyFQ3p6SIv8LRiJOwiROPYUR3hf6oGoPIHHlawD5f3zKO7P1adarkeigfUTfhlMP
FC1EaGeb2cJXl0CE+QWcMF1nb3+J6RwwuC+XDtX8P2FCE+4ksVtyh3o5P7fhAtdZ
e+cITzz9gIGbxbBrRWX8k76J0zUyJSdLVuFqqXj17UUNspz5FTpyV7gbTj90pKhy
02Iyff1ETE/IvoSkobLJcp/ciPKdFs9561bGIteMNcJ11S+Q6p90znTpZ2fC2G4g
v3YNB5xhPJoVnns93EwLtoP/CSXdsdIqsqkiLUYH+FgB/VPuwfUEGQNz+7n/bBzW
jyllepv5Sl/48tg/nys4ZNHW36XQ8O6IL2z5Z4vJy6qjEg3clWSSh4zElTmgsO6l
ZwKXmQmQuD9//dqTd/fno3VbF0Xe9A2UPc8dP54dtYvtGbj4Tu8WbsQ3NcY2pytD
zXt/HDOHNF0yA9cQrEZM5E2vSLXyaIveBb1Kb/ZS/f95SeqXB9J1J93hNjhI767g
o6MX3RJO855eNgFUNqG+bhQop62VRk0sxFdiQkknTRIWVay/KerqNmGgwrIt5O3q
gks+lLUuE7aZ4oWUFA1Nv4a3WxqT5/kxfJtsgEelghSlMyiH7suQPzJKzRgwtnpe
qxmdVqzaghy6ej3L9G3IE2O+dq+aS3ljrHCGzaB7Xc40PUzaod4YTkSTMsKuD5yW
EpgY9L3qMSBi4r90jVUHfWvyWgIWEYLqOkTF7RTWHCrcSYbSsw+moC7iuHJauEl5
SnzkcLVDbc/ga9zDXB+A4ZX4BYciAfgPG2KE/qSBKLdstjmu7BmAvMo4hjzGUdxm
xDgoWlpitNuQjnlodxPTLmigeq1h7O9UNBBgkYt5sZBX37wyskJ21CWDD90yseNN
P3ocwXjVhxGr0btWT3h7zTtUoYnxAqkZqIBwEndK11HY5Ig9+RLyDrmZ9TCDtA/3
fZMyhj3OEFW7GsgtFpVL8OewRhDThfVriy1ZiyldVNE5AdvORr6xhBvq2oFv/Q3S
WXe6K1ShhTkplLOh5wF5BQhLlzitteYkOVZYUdOJO8b1kjmIcTkXMjl6L471lou3
N0W/5z3sOPRLFYO+CnNg/SnXBN+PUq0BziYz/VLSMriGxN8+ojzHVjQD7cPs9lgL
mbKxMOJ/FnYNlfYAgyPpn2TlQ7MMU0hIDIFlWkgG4UsU5/kYijlJAgMFQyDjhCEJ
fZ7U+N8pXdedeIJW8sCyZ1aHDzwHfF7Rxj8poy1XzRxUW0udvrtu6fIv/QQVfPcj
TehxLejUaJfP1B6AR7hrqxCJBxlzxEWWS2TX7hC9ydImHyNVN/9UeDYp6USZQvaJ
mgFs2h8ADVlNZNXU3YP0YlJck415sQHboCu82OXFm8eI/pAImX5FvgMP/tIKZ4Tp
4fLUxDgY/U6KI7AvdUClHn0xcHYjrxJK50VrZDphO/aSsIA9+HSpUJI/coiYZe0M
7VaKhV8g58nHxLNwTZltoBjsK4DJmzOVKWZjFDbDEIpkjZdoLcLqlPYPRZn4o73U
69xo1iSnlZpNE8m6+cJoiNPMMAY8eFhZEF2+Z6ISH2dNzjNZ9B2aRKgBF3HCuM4A
Fg7uHzV2aY4MVGEhc60XrWMYNWrEAXOvct+fxeRRdHzXEAJNYLtC2ITT+rOhrkuL
fPLNnHFq0xgEQhyettTdDTt9wSTa+aJ8ZITQD/8cM4AQSwpd1F5XYrt2wxp6cirF
G/Yz9zjA9tbL3SYXmG2IPxcBzY03BCv+6uhgOVfpn05el+lg/RADYki3yJmNArvr
ugUjm1eiAOaMrwqQd6RQHQtbF/m9Mm8e5B6U6YaRdRn+sElLzbd65erTbtrSs/BT
WEDiscgcN99+DXBhOuhYpOhCupiQTtc8+Pvyq+Tsj/oipU4NOS76DcVvBoGn22B6
zxEm1QgolLxpf4u4vHuRfn3ORq2nn7hg4OrRUB8y/rygFRlDtepSB5Dk1SXUXGbL
IRrkf1nYzk7Pnt1xkFLwuE+ra7fsOwgOPMlqiZGAA1gAArBdVSHM1Lph4LKqXzi/
RnS4m+93WKeRS1FyxypMkkn8a6w/96Uc4h1wz9Y/F0lvKBSOF5d2CN+qryIVWVQv
LAA9WLzkqtTdhOzJn6DSP6uA9uFhvbD1eri1hnoE3OximFg0C/lp4ph4FnsfrlhV
qjJsKjzKvmieErtnRx3RvqalIyNGAtfercurV22NTPPwpxwkOjzkITVrxtocZA+U
Rbfg90X5Xx7BuAjYGnKe5Xrf8PJKgI2j5KUEoWDJOqsvXA7m65+ntoxBHsJMPYV/
kHG9mUuD1cB8dQ6ZW3n1vO/QhvD0mF3R6t2v4jfpP2kJA4nAmu8ZmZ4nKW5VK5Ge
sqirfIfEwGQ6kMDSr/frImKEOTXmNUX9U21VsV5rqISx3l2QbZJHMkqriH/C0crR
TPQ6b4aPaeSIY5Cax4r4j5dyfFW1/PSOoZ8yN5LA5ol/ZQdmQQR3ou40sHZeSAaV
bqPZJb7V4TVr1yYoOZ1JtBoJmzOyG9j50tGd6N+stJY2EM5/7Bo0J857cxTyKtu1
Lxd4QBjCF75nXhbWjIs2aapiicR9x0AChMzA/8AtSbT4dkVFNwS67tMsTU/N3l4x
LSRGyODRQkxjB6YYvx/LfCfiINwVgK7r7GpWP/srwqN7rmA7FcFUdeQvx+MNjfnw
RpnbgmCuqfjb8HLipEHmyAVi+1W5wDI4vDWOefr7bRgYpNrlZnLI7ffvrfPJ4oVD
afzPyuHon54Z3L1er+rCOe4KnZT9P2ZeJMRFAKrHl6h2Q5chiSQzKRl0e9NpbZDg
8wxctDeNz/pBt/GkVUekOiUqAOqDioSQIVBA5W+pM60aCCIQ58OPJytDsN5NRQSS
SrdSPwwWFiznm5GQkHnT3ah1ymgNtMUJEob69ISfJNbfLBSYRA0j5rk7wJdqDPqG
rmo54E1RS/Q4AeUG1ghRzkumiWQ377osz7dIqPlrnuwpVNJDj6AHaVwHWQu6+i3j
Ghqu2pMRhx3cqq/k+CsLvV6V745xMFP9xf1YJ6oJJefXkyo60Z03fRzR4voBbQJR
bP8WX3CW/Ec9oA8+XMbilWnqtP/Z9xsPb0ax2YUixPzrTvn2AHvr9MdZMlnM2t7U
B3QoY4c43XSeEOyEP+qwKYiKfnZeG6OHCnQFknSTHybRP+vDJ1mKCIDQmGwpxZ5o
RSvVTPgVD1jj3Y93GNr341kG5qEOcD0Wn0sUo2uhrvhNohuppBn7S0QCNaZyCvLb
F9Vog3RmSgyqiONbrZF+HUclaVpJe67TkNwr4fJFchOWl5ADuh9jcVrOdjEJOSJN
VWsfq4hxhZcT5uTQrEt2wWE+KcBDNfPpTzRCWHTMYLzl2VJohsTFpql2i5dfilWC
iQrq8yyvw2S0Tk8COkZXq2tTfl+EJevvJU3mqRhTEFg49EK9go9X+XzQ2PN7Xonw
9e9+IufuP2aAzhSmTTmAD3eLTTtkbKL8muqBYzx/ATG3Y/l01nD6csJmVvoyMv55
W66geKTGgEM+ah0FCX8tj4GgjQVojRPERLgNYZh7M7kFsACFTTaVV+zoRcODiK2t
grSgoSX4bQI0XW6lGpm8lnIpLsGg83MmlNWknv9vcg6QHX+xEaKsUrKjlljJxy+z
V9oWIiMzJq29NcE/AwwBHJfNG30/2pXeAQtkyBgS90fo3TraOrx1LaMCcz+3OhCS
mLX5tO56Tw7F08JB2GMOuvCsJ7agqcc0pX11ddwnX0B60seJURLpbw6uBlDu5jX/
fWz9HoewAhKncF0R8su26Ll7Y/1R8GPhykcNkferxMb2qoURRdOCuYcK+i/oMW3J
9EdCKhfEbZwUmULiZYb4Xp3QvFJgwMCmDLZr5hbky4GQ3s0aC29eDsBoKZaAUb1a
sZwDdhz1FMvWGj5ZNLj0CxO3EpILMgQ5U/7H6dnk9d7y9gf2ypee8ZiNcBJev65n
B6M4/C4QuQ2pZV9Hpk29/hq6ZYiGoiqJQIezvpTIe9yyhL39BOU6CNSvoUEzum8K
8XdJnWPwNxezjvLCNtZ6OL5EPj8AbKw3+G4EcpIAHai1BC10Oc/1uFcYpVkC3xpe
vP8Ewx93h7LX3yIiRZQkPytNseHXvMNk2hCQsJbe68kEMP7EdlMFy4U8KgPt8yat
lbAQ7A1jDOfVGVdR6F2ly4lEXeQEa8rLWmGuRq+8lweMOTAulo95oIBPPOLCGuw+
0qt8FSwET3lLF4kmPXF74/yYk0LT1040vqf7YUkcM8OUggT7pCMTqWlK7IOTb4iL
5RHMaRzGyLtd25VQNT9ok3jo2nmshL2wM6oLWsQMgRU2x29+9/OGHGi6lxUKG0Nj
hEkov9+bQ+X8ki/LLHRhLHbvnASTtA8cl+dnqYeYIBBwkLJSg3V3ghUunlP4VByy
enbWzgY1B/YUaxr/rzBHG4KuJj/ZRcNiyOrVgcqJ44jhknZuz4l+h4pOfmWKn5AN
EDVvYfnHjDpt7SppyH9U/fdCvhLbuzLQXinYgEmTmnpn7j35gtXijZCSycCC09BN
BqLQ2HJOPtQJDuFnE6RGxYLYyTewZfJnWQgMO0qLjhu9YiqOl2B2H4glgMSJAW8E
I33AdwqE+OhMNN83dq+y8Wmp6yF3NnSeZdDbjVO7kFcHk65dOftGZir4csSbLk5H
+KVkKwbT3bJbxyVFgbpbHA0Het3pVfPZ0Vj3CK1WJ8SmsmsOhEsVgW+osbghEnnV
99XhFkwd5+vXizJSOKDCysN9GYN6YnHmNYwpFgaCdALHCCmOh2UqUXO2T/DBilq0
pjKz43YPEPli9EWAEAhiJaYdyTLXZcyXLGnVzjr/JNI7dfALmAw3EkTZDvfdpsiz
RfRVp+cfH209EuNw0vojUjFoW0cyjzuQptVum2ta9CVHS69a84kSqwuzXO0uKTWs
zo52D7igRtlkjvNkHAXXtZVa/GyLiXOwTgeia36+3C6akm8Q0qeO4qm8tZtp6Hay
1Q4Hg4tOKmK3PfkR4DfZ01RECKzSVKRDDnSGYnmOjoRnDsoSou0xbo/+X3B8DC7K
EMzbC08a8gjCruywpFt4eUunMeaX+tdjMg0w97ITkjWb88nszR9Uug3sMHkgfdVz
YFTlUeah2a0lU4WgQyc3jFMkU0Y+f7uxfJXYI2AMtp/TOhTf0y2Qs2De7T9D6Rai
14z4JR67EI98wg/u/J57hFKVkjmEqG80THqiwgzqLJezQAe2JlLL1jk0OshAxXyU
rbPunJy5DajRjHnolyFiOVUHre+nay5lH6PQJtkvbxIXdXrPhv3zewg5NoUhg5GD
RVuOd8jQkVl0WKISjGsHhMAlqkkZ5s5/XBW14kC2ANDGVufY/AiAh9av7V5kGE1M
OIE9yOCShgmLzQEWzAUNFWDgXeT+VUJuhs0vnomhrdaO+GHp8NDhBxcHMNSq/rO+
+lxIzK9lgIdXzzFS5lhvF/qppOkeWwE4OcQ8OpYWN1FgdKatOOk1UzMjB/RxQlEC
NkrJaBxMMyO2Y2J5akQ/CCw+LuWn/aL+mV+KjNDlaWraAMEPbn5adf8YHH+Za7f+
aiNZei8iQW+sLPaeW1XWPjwYNeTFQM9e/ewKGeH5WwgzNlsnmEJi9P2CHZgOwomQ
+iq2fKBgu6K8GE9lSHbG2ifTjYelQHqMwqGXlK4bAnQGX4oD2bB1GUkJWcqaGDdO
9o8g+GocwBN/OEtHNHRI6k6SsrXohua9RjckXTzLhJPip7fnF2XPG+Xr6jm2TVx8
Mx1fii9hx7hn4tfKO35Snl0Vnk8NcsVB1DTDtBih5sO/FQntuVjE/585gwaxz1+j
AwEAZ+JGxJDQ/uMEB4wadklizpv9WNICeYEpkwCYJgour/VYUeZ6/FkfqF6wCD8f
KQYMkehdUt40sFKdKY0JbPXjaCVPe3jGRDrLecJpMneOwygRiNNq88Ooy36gwiAx
FwUzf/0xo7kloNiVwf5++HAy+FG/yqlpO1rXsXd7shVKFbZKnZACUWplYFnYv5Nt
q2+UlPwqENYK7IZazNh9iEjkNdLHJmDjj3slEgB8iB+JIXnH3NHm/m5YL6G9F8j7
rD1CU1Ic3FWRtW3dUIitKCtOF7Ry/zwLjayWJO0OaSEezFiViRYYyhNKziCYh1Up
DsEDRfXNhDdjBt6WImmFCzdds+8aYZN23jsdOoF6Sy0IVzGaWgHI6/5QPzdz5Oxf
7wUqs5l27T5I//Yn3ltOsDIhRw2nsOmuXeMnOyY2ykse96hpl/h3/y09WmiK9/xM
OPz3N5O9mKvfb5/mVHw1Tuahf/wVHVZKq6fg2ijZifqeMd0u/MmWAL8XYRm6p3vn
dyAgJJZOSWh6ejkzMJfnqioea/LB7R/AtA/vr4nBHldReHbhEMFDnKpjcDKfKNWG
P85GIV2NzfiefzZoEJOAgrz+18H0BzAqY/N75TRSqLoeu6D60CHq3+miiuNASDht
rse2kY48R8dHrf++ekYFTycBaoH+RmDlk5MgnRHkCl/Pf1hjjoLV3rv0j/kfLxma
BQEktif/sCoxrsj1jmakIjuK1TMd7EFtO+Q9q3AwftUpu1U3r7w/RdufeX6ODMBA
lnGzkRSIKuSIe+mG4ST6BujOMvYBO+B7dODCNXjfYU5aF+xhQONen0ie+kngTgqg
if/nUrPzr1+7GVjO74281lbsIBmVbNzcTCZfD51Y8tFnIeCxwp3VnsjFr9ocJpMj
hULtP3NF4hdAOwzEFfS8rfKROmc8662MdnPI0ctzVCDXnZZvE/huCXS9/XJjZwqq
3JLMRsx/Seph9G7oyyaNBEFELZDRhQUdPuuKt3lXHwiFfridSmvoOOVbwQFh6AdN
rlGv/fImp6I79a7UEgnMlI8TqfBPK3F1D5wFpQtQ5RLLp0agj44bb5X7HhV0v3lg
GCW4vNC4WeUJFKSQS0TQ08pBqegP8TmpYTyTg4FyMQFugGC8UnIky2sgud/sYgTX
+3Ec/9GypRlUlhQXyo8xRHRxHVJHGopUQQJHQpzy8LcLkMmaHZEqGvur3YrCkaLg
cRfx9mag3wsyn+67ntCwMnwJjSgPLmXfKJVvjNbxMHBGP83yBRJky7QURqwiyrXs
zTfe4z+IG3cIozA3DTttDbyP26UAUjnHfXI5QnwBnEoeRgvy25uk5EMMAfE4s3Jp
0GyqFZ9NppV3eUD+FB440CzwjDj4+ZCXvFwyynATdXH8wwOzrrp6ROo65/AuCOcm
M79VCoaBoPF2L4mN86lv9kmjIdr3lrmnOEmMt+6N94bgN6+uOPBhFlqGqWSVk3Fp
jGa7VX2tiHoVpIthOpcJCd/UemUosbK1mW3seAumSVIm0z+kdQ0g7KSUmVBkeYI1
2IahSQJovp3r2w0Lrg4woeSqVX2ueZaP6zKe7sCYyRZqw9OCq0qCrYYGKfgTfa+p
QLSa7/BkRLZ2H92HYRhmWrjkEG4Su1P1n6F8/G/yBEgpdAo7wiaLSmpkU87hKciK
ECJjabGHzcXWoKtsQDV1QaoMYGlwg7dbycQV+tvkXUl1J1EPBzG9ad2cKiuK3W5X
sj830/NLPVy9HI1Lf6ynEjfIlkglTWS1XLLIdAivWOTfLzcI2MLQMGVAx7IsKOh8
zgjHuRvO/XVOJ20cX0DW0Pgyqx8wpXtimUGHHrM7/T4SWJEJR+yinccFHLLfJt/h
5buyh6+a742rB2ypDEz/wNcXX/dRsBam/OPjbjU/jWuu5ifTw486ty9Epko1VN1v
xEgi/CvAve+dcPH3viJMtej84lwo1sYQ5rSH+0JuCyxw4Omc96olDvsxGrwKpugB
ERZTjJq93ft9v2iWpLdsJhs7iPnRX4M4L7Ozvnh7MslZSiq8kBVHxFppoQqolX/8
wS4tbZFW6NoSmU/FYabTvJpSGHGw7oIqO3/0bKqP4au1+cAHlIlrGxd5IzLwSG8F
65v8BCtfnUR/LpdQgsvhWfxW1c61WViLjt/lhW/Uu/2eZsPNbxP3d01SLF2aLMAm
hlje7L7WY2+VON3Rv9hRVcWkFb2UU5YroqMP7ZIbWup9xXzKc6a2bDsqnCxE8a24
kUpMQSo2fTqU/W2ZINInvyKgTAP2yHE5i47gF6Difko9kHfgnBW/FeZDm2eW9gtl
vCXMAFFOLMp9WBwfEfhaTbHsGDRz/MDtQJriMyDChQqGIKF507DqPZykbGc31BlW
gXZXPv2HeelDTF05DBPaDGHEpePQw9TDQiefmMvCoRNWD9Qhg6VHdSmyjFKm2b33
fgYvW4osrx4xaXRPh8KArXg4lCF5zQ11nMfcgMxJFxrYYFEn/lOZGoCc4/EWOQHP
HJQDMEfrorDedR+eTJTMlqDkeq19CRFMtVdqMHkDzkJ7Qcu3yqnKScXDZauPs2ra
0JeOxVrKecLyLzgM7qOEWNoCrHlpa7iXmWZ+R6xX2BcfyZPR4QQopMN7e0xxAYhw
2L5jAv3c/E11ex+YyRxYxCGVMOPKhMyewG8xPikNsUiXl5uf19XQVgtZvVUD2oRE
iWsU6l7JNVI11GKsRYBFV3bPZL+E9xPHKjxKV18yqUAdhH1wsZY1hNI9LGtzmMcE
Iw6e1HZ8eV1qBtoCl06ZNwMi8BPc1NXnse2ejf975C/fC/FK2cvQAYFwhEEQnwQn
DFfsSvJiTTs4Bn/+cJ+Ca4NE5fKTjK3FfqPQGVmsYaTNhQVA6oNYXqVMMdX3SvHk
6BXVdTgqqOz1z781l3H8n77Pc8T8PLS9vptHrI3aQ9wqtBEdVhTzkTB8MkJAQtru
8btIq3EZGupsIEsMU0KVMN3KfJpVg8GZNsDw1ZovwEz5f2eH9nHd0J0V+yAkn31E
S3Qg3rTyyYYXzsV8vc8cBmuVdUP7FJhajnv70d8BiSpluIxu2DPIOXWA3hJ6XNIz
D0f3cgjE8AJ6TGUUT6lH2pHWZGGZMX9qmdNthQyGNoad1phX/3ZhcAFsX1v7OVHU
BsYwdTr33/5g1faIHx053H61YD3a3JK0L4MdcpsSJHp/DyPCz/HrVz7Lj4BuizBY
Shxq3WfW5VIwqOsHAlE0kEkp8q9AmVeJMp5bIKYJBkXtylt+Anq/sxZbtxwtwbf5
uF8pc3ECm1v7MChRKTiMfMKdCVVuu5BDGcdPEQSbu2usNekgLMH3NKMZMvA4HoKr
pDBH8fznNt1tv0Fks/k8xItH0fsP7jlxl3x8hxLVI/sX82EPagA0Nw69iQLkZtoA
+8sXpYX0/ckOngNZ0y8gsdRYUkFfIA4IZ7NQpNqMHw3ai8Ut0eTFUafXzVbstepG
Jx/2Ms4UNE6o+H96FlGmIbfsaZ54kLet9TG3odgyX3rqirE+4y+ryXTQ3+aAQOtP
vIPUJO/sv9UTNWQDZV2efLVXkb4Rd+baQkNSnl75sGys+3AgbXk8ZZrLDrz7BQbs
uOqJrsGjBTZnpGHSjmdpVEoIs0Ippn1UsArxpDFaeQGgWzVo9gZ7PU+ydUr49aHr
aqfRX2X+ABdmJMh0+/SlRK+EvRtQr9rT/zJKUV8VUITxPigcXYeEcJZMKbJwwtZr
l1CTxC3dKVBz8xpyv/UUqT6bW6xPE3tczE1PmiIkn3IfJ4AxZ5HEyNql5hG+MWgd
pfzwPiMtYrmqKt/GaOCA/nWN+kCbGAwor8LAdvG/SjFO8AM/ez6M8uOF+EvcwTA9
iPyuGKfWDNz6MW1u0ygxOjPDQIkoksUEHSHt7tsuYe464ex28LeEkk1lvaLSb+Er
q0wzRPNXIODIhBqxSeB5tNGiVSa3pKzcSJNdVlLgiuLMF08M8V+tV0iyMog+cVt6
MPttwipSVOKtx7Ax6vqqwxy91HP3IsUUVFy37N96RN4mXHy4rCrB2e88qkV5zDsJ
cfD/VhMcuXtMNvKCTJhNyve4WY58YVCVTqfNmui3cUU=
`pragma protect end_protected
