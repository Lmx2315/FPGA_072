// (C) 2001-2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
xllfNoEjMTpGqbjb4l8azp2PMzmALJETaj46DDPQM968nFO26CNrrK5Kje7Haw+J1YQCBtxFcgtl
o7ERjhbY0jDINIYYWU1qLOzNxaAWIVZw/v9O7IuET4PxlNjs5N1nl2zN+NVO7+zZY2et+vn2zyh+
wvljNRwYuJ+zhEBT5+TRjXV96Y33Bw4dYhinRRELpIB46DZHyAqAkYfkzok5khmhng8dFWHOwO4q
+dcfh6ZJg7o519m6Fi3wjcEkncVzjQXY6caAJjxe0vodmIeyueBSgxsPLLEtMfEdyb96KkcscQWF
+4SuCggVB29QZw77lWA2lIdxG8SuIn/TtRH9og==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 1984)
UEIDP/WCZX/RNZ1OwAeFFRpDPfunC8hYwvJC5nHHXqgM93bJ8XEhXVUKJ7R/gfjN6IsRoCRhegS8
ujuEN85L17o4jmuCaLPevlqx5DS4/5vY++gUFHjVMlNNZceDtWmjw8HgqzT35OBO37snXnlE2ak/
QT6v98LqP5PjIZFSFsfke+ifDwhs7Bg8CxH3kSS3k+hORwL6/cy9jCH2axTBEEqgXVx5AipoVNUK
paFitlIEzoiHTonl3UVTb1MEr6s23fY0RzPcTZHMrmdK22sZmfmS1T3LvnSW4lh5ls5gWokHZC5z
XzE5QLN6zrpFQFh+t8zAz09sklikDR5KOyHvLsskRExqMM6tkoScL+cs4FthKnWX9AsCcH/PV+UE
0eeJBDgnRD/77sJnTeRLunQaBYJN2tb9MAtxmtBURO42uNvicL9lRoHNBxYQtY2UkqdTy280JeJw
WmkysSBMXWCWai0YeQ3ogK8J5H6AHakxr9yIo6y40VL0rVJy1Iog6gc3Sha/Ps+2KsQ7HVi5Upu0
IOhNYgOXVZDoRCLKlhAC8X2Cx7uUpdZyffzkvOYLBr4BLvL/rInCDBNfjBdeofLPQzHkvF3ok1Hn
9TPhYBdcw0VDjyAVGAWaqyGxUs114JSPIdC2FzmoWklnBZUdKBvvHMi0QjqPDKkf1Uw7QgRAAOVa
z4zewAQOGdO6Iv+UWTMPlFPppAPnIuYxGu3IZuSu1jqxb5ttEgZQt2xJ+vZuyhw9TTAO/JNFB5Ac
p+UVHyO13uPiRb8JMQKO2+7vF3/AvZ0NJxt5Xr+gdSu+g/mIVUHKFlh5HkvKa/aUhzLv+JXos6RR
/YMSyE4kCvz1kSh15wHPlT16iOmRIkt7CrkWsYq4cnnybPUGsM36XgXfNfUYkuByBxcsFNYln61u
82jngiMSXd+F5KzaQxjEjlXe2UqYo/Ct9+JAj4K4U7jHWvpyh0miIUkaLxKcBzzgp3GqCtUtZ921
OgNAKEAPht8/4a9+h8WGOatPC846LiwqAYWQSGeUUo/gV3U8dzI/iozVwGoOY1FWKTEVX/9O8Tj6
AkfGnNpy7CW65cpbThJo9mDCaS/u9Q50JcfQAI6XDWcsMOlGKhW2FspNCWe3VYuykjuxC6io6sVo
aHRpEIAnJXszvznk58TvQNaUkMzH3/WehQL2zuaUTXmSAuHpYunw6TEa6PpianUnaGv+UFSNcEnJ
WOIkaHzZO2/dvBxpkFLXm1NDjHLab41Aql4vlOl3GcGtMJf18lbxoYeOuuWWlqvohmDRW+602D/Y
pSEbJWBQ9UZsdyTC3lyaWWA4UIGEzUuAQs8cxi8SyZETzpafHoUv8weXQVEb2gby+iA+YpO/w2Af
AHREVw7wM6mXXg69IunG7PwZt7ATiN6r4k11KFiCsWZvDjlFohs7Ppz9Hvv7QSbMdqhIN/kDrqc5
pB7jfGYm4V29xxe0vmdy1vb1Kus7mbnLaaB9CFlgnyKQ0Sjuoe/q/epSZ6sn5Kdpw9D+GXJPaMFp
dYLCd8MdSEsH9ixPa2THiNKRSQ3P/Tt207VSt0Bi/QRcAymUs6VErCzLS64biJqryXY4KzaFTdPl
udEjU6z/GP9GlztphUcOwUCBL2CzxgM5V1haDU+kBOA7TOhbtMmHzaa5uUCYfb4tSpnbAkHrJCpq
qXLqSPd3ADw4OKspO9CiIj1H3p8dA4joAT2MtmwDQYbTsZDMvOAJXm/b6UVM3VdKeFyLk4bw+lBK
jFUv5U0up7QTmRVrjPS7/qBqAnMPtbcTy5jg4W1nWbivCtbejydJP26oaq+X+9AXtLO8qyvdPRHc
9T+/v+xz/qtyQC7w+iGGyGxshp20zwn5kPzE0qi/jEvidcWUl8bjZKR1WAEts3/svGB9ZZHVnVSY
ufCnV5Qq+Xbhp9cAqzrqRceswURR9hBblDj2nwGIgnHGKsNn1IeHlT9rZBAEEG9vABaogPyaPeqW
EcHwtWogNbxwq7E/Djl/umImn2fhnvcc1H8pntiASp6zWobVzn200xdC+NJn5CpALTlnZI8Js8o2
q7gskJerJdkI2hr7JJiieRscArQUVMAF3PdXepIoCOr/tCKxK6aXwDwwSyRAhYlSOU1LsIOpfUTw
eLdV6V4Yhz7fZzxajHtYMznUdIaucjqtd8hLWrMghdOeQ9o54uEyFScY2hfrbVqPnlQzehEGvabY
XPqjiJNzywAEC8TtHkulgwl5xgpEvSNuIJrloEvV6d/ODWDAk5jmQzpEll09m1PSm0g3jb03Rb9E
paU5P9cAQlvDQgI5t+3ACIWNPIwE8wbsYl27QQzddw2aVwjpWUVWzI8M5ERHhJB/fJqq9xkNJf7A
rtQlPnoVkac18SbxYm9flCTxQl0CKky7MC0CUWcS0RZzDQ7uueGKySu3Piv/k7u7h5O2Tjo6WbwO
vQy3YnqvA/hBfIqlYCbDCSv4AFpfsR3iBHesT4ukRU6lKMuL1WfysWEqgMxsAUdauShszj03g6Uz
cJu8ZAjhe9L/tPxBLLLAWkvIogAsIiH14vCaKC1bSK1T/zU86UQzaGcwn+FSxr65ejC3p/CdKHmM
pcjSV6Zs438w2dau7Nzm/DTE52NNAEHoeSr9dFrghuGV76/u8IESGZHBDXzqFA==
`pragma protect end_protected
