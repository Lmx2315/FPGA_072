// (C) 2001-2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
0cRLK477mBC1J/PX8lLhGXjgQpwdTh+UQp+vQ0k3xF6nGGhZoI+Y9bJHvmvLwk76yZ5bbzfcQgHH
RcP5CtZ5lzWEhk/HLSLO3M20au0pbkMgzFALjeZA1w/7xKZCyOLkCZ0TKa3OIXk7+ARCJLHip9Mt
tgBGQzA8DQ7+i64VoSuzUfH6Bm6KbIYM7REA6UQN0iFdY+wdyn2htCY/rMNaPAh2hX3SoCEOTrAr
2TV5xi97c3p5k9IKq6PAX/nJhqKRcvE5uDN4Zf9+yQIir6obm8RFC7aS31981id78ViZGTq+z97w
EIHNsqO+pBj5DmYgkAmFfFexkzSYVHOIZ/SW7g==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 17280)
wN92l1p0FQ5CU5UOLHtSGmsl/JSubMu6rOyVd8Q1o5MY/F9F/mye8YkY/h0CaM7IJt58exSN3lmd
Xph6snLdYQGwntzx82XXkS2vTNdVMPv+D6B+zqZLEC7XbUkBfxNlVPI3lboef7B8JfLldZ6UUFKu
7GdGFebVntjoAeNKYYAO20C+L2i9dnidrYBw/BSd3+fq1qC3fTAixDPv/UF5wB6SUyiiV6c/vULP
ecKI6VbeH772o1n5UM9EgqqpQ4y9iV4MWRe9zgb3FI6XqreTvd7Exu2v5Jdp5ostno2xSDHmk30n
5+N+26lK1Cru12a5Opd8KU9rX/saah2CQ8lNFvxJ7imX3c6ej18sU+K5dBQroX9lXJc035x58jkw
sHhhNsauHIzju59MbWbRSeJQarT/ru461nqdMFJctUWJjwcTV6lJh7foPecKVFwohop/RW3XsSwa
PIkkFlrn09R78BHBNCPZUrkiww3zQvU5DqxydMADw1J/F6+IVwydL7qZhG/YAjTZSjGogwDL8DWv
EaWEkmjtrmKe+fMS/CQg7/XTcaE4WhhtiLo8mEBnAr4Xhbys9r5FOXKPnKVD7xQbQrfnbtcZRcbI
MSHVSNd5HiAvku+gxoVNyUnZHgw+8TKZT1Olb/hy/VUv7kcvWZGWEvwiqnd6OR+OIdlSitAkwtRN
ZioVz7k+MVOIN3/+n1TJX1bmdQkZI0l3w3xr4ez90EnrtvPvw4qaHaAGb7YKrzrY9mHDE+hyDZxs
WuNZDkQ76hwBtpGnNAjmtXgoOSIAQInwVvemmyGe8AVPorkW2CniVbPyBvLo8m7pwaxXUJiE0ZlG
zQJ78Vje3QaNmQqE0FnAMIMmhZz3MJIvjX2TPphchcRDH+RFPcr56WkhF/nQUsvcee/f9GfN9SAi
OECujjCcxnbWQyOk14rwfV/sG6Q6zB145cuOfix4AGqxNHKDENT7TH/9yPVvh8hYOeJNHILT0+F9
VPk/pzFO8GtElq9t1JJI3CjGTYYuclZR6hQCL0D/koIjcW+kZ75bt4VV1zIi6GUsaU9PDvGnW3Nf
fQsNTGfhYuWNMaZ2WG+6t/7qBMwCm9iIdFHLw2VENpPBg4P+4bw8+KZowESQEQj44/exn7gyeaI4
I3DvohsgNcpk41S7hPA2dWp3jFKAMD1Yrje6FaRoAmB5LPYrsW93MijY38q4f85WYNH18znnG5Z1
6x5RWEx0o0bxEnFDSP5C1RBRSkr6I37VAM7KqwPoN5ox7VD0tzBJbN3yS2Xfnk33FKvV11WbbqcX
Fp6CRpPlKBZsGjGmDr8xCIOzQsxD8RYhiFrLRIoD09xsq5fPWxFdVEFZucSo+LbmrILN8++igAZs
LipO7dW0OXMDRooxI+b7c+PmxwgGTPfPVr7EJh3xN6P4Og5qEmZHBMTBCxW2tJ79k1SVpI0fFlL4
r61GryeYyXpNXWwrTg3ZQL2isfarpT2KssuxMY3W6KLVwuRX0LwfvZ//6qYwn4Xf5sT/RAMsfGIx
2lxh+n1eKHfJz4uw+6dhmZHG4f8lOaViaYDSSJphfI/qOhv048m+johkBhwUxfDoWA/HJ/Jc8cV0
Bt3wetlU0DC0wCpMK9NLcI1E/5+4E1Epc9FmSw8R6D+FMgZ6V/H5y3dzRGnDLf9xY3Xyq+rye0vu
cWYng9eR38qTs1yCnUZwGfoWpNvDGY7ddrAJPVHz+iIzFNp2Wo/5Piioml55qwAeOAFmNd+5fsBc
fTZbujim4bgoHMjlvq8vGutfoTQJNkSODOvR5fnMzboB2CLORqYd7SS1wyiXot6Obmdmx2suM9MA
QiRzq1gu/o4JxSzJzlOF7wzOCzmDrrEBTVdhUbQnq4H1OMTEPESvTxBSjyDzkydmh0PXyXYx2zpz
qMkFgAMoZV8m8FVX3NWFURvHo9PYLbaPAGn/1cLAjzEsUSVLdG5sL0hxvlCsLhaIN6ZzVV+MwDEV
iMJjC7d09Z5T1AiOUAI8HFm9arZAEQE0wMRDRSVIryrGqr5V14TGiGRvWsXE1UDC3MUSrxEF+7B/
RWCrsAo6yV0/iiKtU4eYEC4OF2bTIhcAUvO4vt6U9u5N8DvRJGVkW2UZ0N+c/PzO0KKUT3TlnETK
4Nfvf4V47XAFX7xUHIBeA9Hu+ll4or82P/pQkKvxdLDCwTmuUtyx/zBwzMKoVZtkKwH50F1fg5WE
nQUWdng2mXVk8hJkjq7BM35uHxlYUuatkc4DBTEePtNMXaYzRZMY6ZRfwsLOFkD2j+qRSTG8nXOG
Q40IWS1qV2Us2oPav7O3tYPYD2ZXSgt746Nzv+pmhNvC0yeDUQr/tL/hDhhMJFJkj+vi10SO2GNU
tnarznTeGbEJ8FQdIOnyC6qPo0y5TANv1vgR9ww90uGeJMBxn+dGFbH1xRM921BVHoH2bFmOgTUk
GpW2lVfPh1GWULdBwxNWPGNFlDr7fzcmd7BBYdHtlbVgTTngmvB42eiBaPyf0XDg1Xg6GUVpRur8
bwWlX4ONLavqWW+xXmcQVM+A5fKy/grc6tOyhYjr/ksh73OcClYm46PBldmEn0IAyijYsV4y9h2x
6694cPXbRxXYktgF0skWRZk398XyRh5g2ucWF+O6XKAZH13CI6qNnVx64uqVxOwS6xAVC+owHFx+
X/TuPcOcWMVid0eRZa250xCvdBl/vb2NWLrNHdSsFPOkdm395BGXicRzGGc3HkO3Oe1fQNVr2oaE
BqOxZlPSJqDrojuRfgAK0KRhO/98t4pTVts+ZG3DwAhO0G6WktiOR8SBfYP5oMYeI41tjZS8Hj6U
tXzKYKPAMdnJ1aILC59Uqn7idJJPjYLlt5EF5YYlYiCHtfsVTAxsW84H3Kt3+mSfpcsn5gmbCIB+
n713NYV4k2k/rkTJhqJQVRnH65+XwjzOP4eX2avC4GiyX4cuLGghizmIwMkmkk1UoTab5AvDnfTO
6RDSx2f0hiuELrwptPQehYaW0GkNtTns4uXvjQSqzewLDX+3ONn/ZgbhgzfbhCgeKYu+ezT1JaXm
tDXvMRqfQCSYLkzf5+iN4Wc0Ax6QfS/2tCZnBUpvweM2nlzeuphW2dRYfySQI/L4GcScq5CJdi1E
8vtsyLPEgPNYK7pTU+5dC0QzkoBJZ2QkGjXVcZE2EjBpHS3z+xFRuuIgpXSbC7WIDbn08KTTImZQ
LBdSS0ownOdaDrZ63akvXptWb/cDt6SVwiRGJLokq5Wfw86uDyW3rUAwPG+3AYQi52UcVRCY/gtJ
KmUN1c1SABA3UkeEp1hCgBDOfY+WcTvD+4VRNyB9RsVWH2ick2OoWqeA/RoYdmll76S+xHfkVyhs
TIDznvifQjFuCwa2FPTLvOO07N+g0GpJvW6xF/nv3cSvRnoMUpewg6r9Lez5vF1jJ1GQmWgpsAn1
tYaBRrUfjhcCn3kG3q2+kSiW4kzDQ0LftE3FyvKgYnAriqYvzvwk7ZrVCC74pgmvFYSyd9VRZ3uN
vEA/Xt9QP6T1LZ01fQNinHXatV96GU+6SbWnCdRG2fTC9sf5GdKH25q04v1ZUA/G6oOACbq9vv1m
1qXTcCsmw7GRmjgUnv5g52Dj+9ajKCcYbNJDrBvN9+0vSTorhp1gBYJxoGCXveXUCXFlOxoGVAcr
cZTCvNEMwjPGyOxnM7JO/p7yM18gzL7O5gq8gMR+Re3amTYX9LsAQtf35XJCGhIYxJ9qEgcy033i
wc9/Cz93/p98KR8psShEQ55kxEMU0Q76fFJz87d9AP877Aex+w5SSNZgVv3C0D2XFmkDAxAKq6i9
PXduKl52NgSFzKioorleCJWdonxC8inV2rpsfPHx7r3wb0qFXFYrFvmoLabu8ty/MkDxxmKf4jJr
g1kUzcD5vxOrtijWkkC3jLaGN9qqEyEKDoOcA4KqCmAtFw9+epT8vo7iY5AbfSJ9dzlznfSkrCjJ
95lVI+kVttNuGnQNpVUfBBnGu9+fY+cPtl9tnUORx0dg2a4zW773PGrvniQ7c+JbBN49lfxKHVE2
2dGvTOjcJy4/vrZ9KGdlZef+zRS90HeZ3AyU+aQTg2ZP2y0JtU5jAEe5P200D8W8sxmvkl1f3OIf
/+RgI/6t9h4vAQzwY28rLb2zns74MtHdwGk7orMr5KDJRDm6UyTGJM+bsrzGhR8B7+FlchE9fDtk
yD7DcRK3iFp43MyHGtLbXLhFMoFdIx7T/21sXVNf2fWsRhu3kCOYCliLv1bM0vbkMLQm8Wo+OZrX
qBMa/28cZoDBBzv+vUSl09yt3DgLfQL5N1931eC3xPDlvHihfZ5DMGgpYis/ix3T49XLf9/7X4jj
DCQslNhlv74OojlLACoqDO6AdzTHGlYIljpkiJd7q3av5wDMsSUtOZA66O2G1s0OUCpJkbmJdD6H
g3ootzNzSiEgDUnKlUyDh5LiJIK7obArXuF/aaYMSXM8/wLbGvini5xrmWYGKI0IT/aYzmTKcdCL
ra/QPrMFTur4AgWWLitE/JKf5MRkY6GdMTKGiC7PApBuWbzC4qQxZ6e7iXRNmHN95BsymjNLaL6c
czJWu4AJC+IDgJwZLB2lBMzCMxeUUPoQhTW44v2sMksTTjZFb28ZBqJPs5om2ihzXPKwMGE9iiwM
lwtNFmIjkSTQ3w7r2TBX+C8OeB04zLDTuJccIkemFX8LT1Fa/CFGV0dmsQPeUWH52OOAKBQrV59g
z5VS6xbJWReVzmAbQc0I9IUGWNZ++8Wwy7ZhsyG5IK7K60IiT0F1bFo8b+tfDvVebsAjeh2MEQ9Q
X8aDp90sf9X7FA3p7gShlzgMGI+zpMVFW7OZUe3nwr+Fwsbc7VJzqrCJFyOAMW899kl3P+HsY2o4
g8MIq+LF9L2Wo6d3jej4D7+AboK2nxBGj9TXwQe50iJeA/QsqkGFl/YZUIMK6PAnh+NyzEEH5l1p
4netnl4LI6OORPsJDxh3uje55uZ9VXiwotJoUlixWzYTrfKukdWo5sCRZb2eIe7tT8UvhNxUIZQr
Pfj14PfKOZnAicOQsI4rj2d16n4U6WIj687aLwtGMrxbSxUZEDKshYxwvDxeCWJUwK1tyncuclS5
YY7G/ZNdfwi7AfFYe8OnWJagsSL2kSdum2DzP6vXFFnzLrx5kLFnp7ozPUx2x7IzasJrm5mDhWVy
tbAgmbF7AFrOwqGcqs5r4x4/ccYA0ydpHAG1R1kJJ5ZZiyD8ctTcFFo0EElloDDQC6RsMWUwVe9W
U9pcu2WhQ5DweQEhSkLOQO/mJXx9cQL3WJKlIMtuss1pZaaq1qYwGRB2xMcki/rbTS8L4QQ1JxoO
JXkExNlzYeumgYOfDhUY8x7jgKkkV1s7nE1AXPjCZCSPdem6VWtyBrmScc3CmV/SiReykz0jsWTg
3F2P4j9ME9b73Xc4toXWp2mPmhtqnqjFVMMTFuIGLs1AJHdmG0E3w1DSaQKbHB7yhr7t86kQEIQT
Y7Mjjeb2uJ+GSBw2oOpjQX/wqniY/N3CIZghQoSJab3pKa3Jxba4QkXaVfjX29cpROi/J0ZSFgKZ
bqukCp9wRY7JKik/vxEUqHEctkxSqDEjISgkBzX6NcdPfZAMNBNXx+HyNwMhzFR1TIiHoZw0sP22
aV/oWnPJPRJri5MEYWzh2JhytffkEVMtcb9w0Gsu4CZAp/duWKofNml2AySDyvl+Wk5kR6XJNGIl
IpEWsS29f1QNZ+Dt89Jthp7Yrd9oi4jyvZiIo5NBytQHGFeJYPqSZNIF2e0TmKA8OFrwZ7g7sf/8
hwztO8LlKYET85PXkUPxCOoEi3Gudhvb8O/t1gSvvxLmar7xHtYDeI/jgZ6Yjgte43iFUDInLVHs
x+qjQvlDraETo6TK50SwgbwK+uLzyQLbXOg+mBhxm/Czf7kTVF8tMYD3cMuer9l6AwYCs1Z3f8wT
09loDy1WkGhn20Xof2/JVdPe36k5qxYiGlD2GeZ6Dhuzo8lmW2i7MqUhmXU6EoRRNx2U08WBJ0LH
f3JXdvcrncdbWgVLU9QbgUMQeyRsGvk0dkgAOfEfR9+uI2TZuBcPvhRidffptldb9KxFagf4bw0y
i0+6xckCPQVnffuEla7nVS6fot64ntOtSU4Ek+/IQe099odf8GOwsc/iux7CfAi8RSuto26++PqU
nuBFfRBwYNVPFyqTCI3DZ2a/Pt4GGXImgolWbI6eINlNanluc1SbWSmYl5844TiXYs9yZswXr5eP
vkVdTjRgmp1ORbj+Nc69C9/RooY0EuRppt7dUv2BgRjRxG2lYWc6YoIyZsyicBX1cEhncPYnEhCu
eRqbVW2u04I6tMiAQlt9hMJuBFO/gy2nArXFx3xZajUSbXPZCv2MbrKm8HUnjKXxcue5ZKqU7w2y
FgR0gAlfgrT3ihDQGooC+FqWPtjSc995m0PwWloyFHb/No2J9EFGb5mLCdV7JK1VPQn4Xc/7PKgl
JmcPF1qRy3gxgkHDT0weNRbwLMbZndJ3P0o6yWlo65GMnbeqTaQM/JXewEIVQLvhQn7jyUsIwB9I
tZXD6rU5mdOyG43RUEkkkXDNIF8VLGc0igl5swlBncWrkqorcKtY2H0mMcniiHAdfeUbzltSXxeZ
OIFiSOL688HJY+ITgE2S2NElFk8u1UBU1UmsOdqqdM7BNbqWkSMXUmhyl2PlX0kLLBXzLRW4wpPn
AOiWLb8fvlFUqj2xYCkzGZm4wfAI+kUIrmwrKx2u+9nrENNGe71RykgGXCzWchABMPnHOo2/YO2t
WoyU1RqyN69E3Fge1vAADBPD2RWEMJavfv1eQ4t/2U7zzvlf/uwZAp8nPAflupRyDWXbLgI2ZIEP
OphKe0JsPlq2uq4Xip6NSCk9fE3+lj0QjclceYv0uLaGpL6GU3scQxgOyZg2quTQN5MAlmbM3T9O
fzoKRisXGtvoowjK2OU8hH4L23IcDix3Wy+cWD0+ggTgjsWYms65GFUvUh35RYGq+I66RQRwaY6I
OYyfZY+aCPG2EjWzGOjNQxTO8EiJ38w+sw3w/i2GfDTcQ1mkAnVWwkFoyyoqN95fE2PeVUeQeiYj
IORa3w8+rryy8DDqkUd2r8qQLxWASUFFSbMBXtZwz7lUatv87TJO0Khu6xKmEheTy3zidHrb9hlv
993N/h9tAmVQKAsl6WWsnp0yiUujUGSCC7qz4x7ASUpEN04bA1oXygJS8MB2jlQMzMSFCluu1S2s
fkSw/mrVWY80fAU6zfBUtfFPdSu08FYoKGe98N3ZhpRs5bgMoq/B8O7o3lpB7wdJsfwo6UPy0Q25
n4A7EGgdlDbGld72ypYlOHcufFIhgJ6dbxPmneytuSGq64Z3fgOXWb3numKbt7d9rdnbWUThUNu+
CRqs1IPonPxGqtqTs29Famh9PCKP3+4fQAsXYuvnTFv2A0q9MCIHup+RjoW4+XJbiK3Twxs3o7sk
WflffiYM2OaieRLkwiArjyhCGf4H4T/WNi7cuE7nQ1Zs9XegaG9U7i1w0rYT8CVaSrl2ghuFlSdk
kuADgpnNw7DmsqB7Qu9/9+nKsiwAe2IQ8MOGxZIE8XdrsFuMj3FMUNOuawRjdmgLnfP3caEZaLcQ
2r/4bI6/SkzN0mOz4ndutO6fcUz1J+0VjGGaRgJAFOT0jsLUeIqEsLDJCZSNavSYbb3/XVMg4vtC
XHRGDn81w8IteYh1TvT89PB0uIWBWh+StG7qei/27uI68duQ8S3yx/tktTmfCAQH+UwWWNg0zM1g
b1m9VcmDkwzio+U/S6l8jSYbbKRTNHTNLFSUV8hngcjKYKH4Jk+Dwmu2I128XQw1a3QGwmQIHdQ0
HnuioObeZ+hhQkb3+1wcu0X8XWsVGIUlCKi+nfTSz5zKAfQLSdTSo5He4QzFcvbH7j68AO5MMftL
1tJKFb7Ewyp2j9ZKL3TxXeFI/+hPtSkbsyxW5A1c2oU3jlzEopFeR88kXoTaGlWVh3w8+Y+kUt+3
gIF0s3ddJEY+aBMsXFS3IGaDIHSzUaTtbt5xPQNoWJt4oT5PTnCu89cWfzhBHuVoxfaNwK2RKErs
6pdVv5f0MdTgA0nHfQJ46AOcasfrEXqoyjXOvYFC4yAhMVw9EsFvmfn3oEKRKRDMuf6CXdpkOS4W
+FSCN7L1zFBhbb6QaW2jB8AmJMb8BvbCJ205/0erfdy7Bbqj2iLQsAd9bCgf6cKjk5DWPhjPCzp5
7IpZZ7OUw2ZIjSWZnD0FefKs0zY1rsr8HcXobZi75Y7vTuV+AqnbjyeeuyVeurmKx8ruDOAMfqcg
4R7X8mrjJ3O2GKJluMC9MjGFzk1JT9GA8Sd9bmQ6pb/jjPBm5ttGQPMIEcdbRBGTyQCVM1Z1NVra
8NLXZHY9pS8EKa9dtTDa5uJhtgj7xMb3u2VFJkXMn0xK14e9Ysg374cq8XBQtoHsel1t/afxR+M9
1/i+Z0xli6OMezarASIxlMBFB7O4gKPZ/tECgXNx2/6/B0qnfEt+vsd53fpOuF2hEV/S/RpmT5hY
dhNCgMGVd1z0yUwvjpKcHHrMjaIzQTK8YoN5zU5e/X5wvEUM712b7L+ElcVDGJvuxogynfAdp13W
we3xQA61XICpq8o0NyeSBm48eHaYmrxZIvzfj0pXewsAcH8UQwSP2d4QvUy9Ve8bjoHk/dnpZ0i2
N968nhM6PQv5cEAwNtOv8AIz4SbS/ZnucrTbg/FwPhaJnnFqLbbLLFb7eicQnJwKDcER664X5WhW
UKcGPp9QLBI9anoKpxPWZNx9Q4m+7cwmV3F+935xdVllXjilJvfP4vDhJ98XTDcoAiw6X76mehxz
kB9PI5TcMuJ3FGj9LGxPRxBSe9AfymOmzADwUoXfdnzWJPAw0V8wp+Ud52zRJjiB821HYK2wl4BT
y+bwbGZ9gtcT618hAPlxwhfgGq0nGXUmj87MwA3Tya7nXBCq+nAuwjhi/goWjPSRVqFBgNEYpCHY
6AxnM7JPZiA+i9xW4Ig+deLb9sugxgAbwmQLRrdj8OU1DFZHOKQ6U7tZT9/ThE9EXw0Hc8av8F8a
cFt9t5bGjZDTbfmPRhLjvohBTO98895OhcwRzRZDKJ3dhaFLbPTJjHF8eiB25KnBfig8N2RgTt4y
ZvACEimLIjV79daa2oIFaktmsn1B8Vi+MP0RdLRzRAM8DPC0J89vt2kV9fP9MBd6aBCH1DOsjqfK
0ILs/rC1Ckv4+QPhHUXot3A9ZlfmTn8YQsV5U076FuBUGJosZe+9iqIJxPiU1XBXzlWUnFsbn2WJ
1B+IlWXjWeyhXEIYBNZK3way/vTWcHlUU/YURlvM3I40Ue9ieccIs3wGISsfrkZ7N2aQXTaeALRs
1i3KdLXUNIBZozfjXVnTvJ6P55FenqFiyR54iQgWFl0KUmCAg5uxVwmIuuAaPp4oY9VNbI0W6z0S
kqZyxS1KtQfdhyQrQ/z6zxPGK1aPZSwZjLL1xsyvup7nwYIxrRRfgK56c92hqFy/OfVDO9NJ0QHW
5ljBylloOrYGjiVcm1wp/dhLY+DOBUFMpwz+M0r74KhVtSNK5yhRV+QHUTb/YUKrVRQratPZb43P
DB5YJ7K1mhKM02kldye09oO3KOMmePk4O3IVOyJlygY72ge8ENB9OwMTo2r5R6U6XGGgLgIYf+yt
3HGyGCaYebNi+YLxYx6/hrkcW6w38dHj+gi9ipKEzDUEDTBOzEUWES5K24t1gLSO/esmlz2iwLmP
KZO6IQuzyt1MJYcZGaUUJ7UlL9hPm7Tl/5ahm9kfgNwu7s1euKDoxw8isouyr+AdvvaTOk2eMp9o
lzjO0FX0rKk0FhvuwfyHNKIWoBZRB84TwDF83I6Rw+ptdb/wgjZBFHStZFAj5j782GdPrQhfOmc3
yvubEK8WlknlBdvx2ddWeoRN073yGQOtvT+tO3CXHIz/8MAcbobg6OFHHKMC28KGsA1ifGhr6ExY
7T9It6wwIZX6xvm7UjagtPD+1HMcSyRDnt8T8kwk2/f7XGlTFXTluKw41G8D/R3CCkTs2tBdLv8J
MZQKTDnYBSz2tjdCbjGcczYaMtyVj8rcdDPEAfkm27HUWT7GjrX1g18ii85A8aq5eFR7Q+nfPQFA
t2LxRYMrUNq9ydsmaJEDi70TW3rfY7HNripXZIOEygsov+xtspQ0TLOckt9ieUV4jlJltrIerkRW
p1KUID9inK4oC8R7Yp9HMmTrsSu4o6WYsp5qGhTLbm7BRV1fOs+H0LdR024jGpO/U+VC6nHSDTGT
kUB8sQ2e6+us35VzutTHuzP9IIfOd+g8UvsEGIoC3A7LBO8VJboi1IzgZGtJ6Rid3GYbiW5y1c7H
s/SiXxK5BJ0FwzHuaBoi5fy+kjRhkTlv87A+ObYNawwq+UXU1rbEgriBXi7bR5o4NHOGfIVEo5o3
zeI+Hn2mB6XcUbCtwgctf8Oqnx234i8IVoD+1o9tzAraSz/l7bu4DV5QvOeNRRCap71RIGawmtei
GXj9LufafQXWHhbl235ZCmeomm8fReDgYdROsYcYcvD3eTSb+/V5RPePfkiiQWIdQHc+VdBDqbZg
M5GanBm8JoVjlPku+xOHtQW4VqlmdC7t7rXmrSHE0qrFjneXfZ2dNUBeJygFu0L2LZ205ykHpYsg
nFWyDMF7UwsV84Ptx7L/RoZyKwtE/6qwH8Eb4K2a3n2M2fLu+jV4miPB5YwPHsMnVLj6XCpEHe2K
Cvi+jy1a3AoHrXuGsoCgD375lm7CgI7vF7D4Ok9BL8oaXySyazeiZ0Pxz62Q4LMGV17gsJwUa3V5
rkpGUmI8Fs3LwCrqaMCzNeAIxyt1Za+lF7H9C2Z90U/PStF0H9/zbq7Qzz0wZQjiDrdHwpnurLaE
HIPBJLzlt+9HHfptLsijFk+2JQiTayYseanBZr196mLjb96v+rZfFv1qLaVxoB4+v6eS0t+0ozmP
Q+Xy15DULQf1pwyu+/9ZFDDaVw9NY7G5SDq10Ngi7tKQOSH9A8nKNNWnNfbrtfiFDAkPCqnQuV9T
yrdIUGhgxW907N96ZAH+njev/KQK1HymztHzom8BQPt480wtWIiIHSzrNak530CXuu8m5g1LxQX/
MfoAttXGsw0lIBxGNPxZw9c8nbJ58eI7NzKkjAGWviHFL2PYfTBZqWPHqjZPqlF035mdZJcd5ZCZ
UYQjfEo/cPy5LkmkAZJv3BZTW4lCYEm00tW6v1sSKkbt7j3TCgZ5robzQ2LRA9rnjh6K5POvBnvy
pF5HQir5P4dNyCIZ3XXnrJh5VlvjFb0jkVF93+PegKFs7tgtZabqHIz1g+Icq3cNYizjmrHJAta5
QV3KrDMwhww15tjsWZrZS7ynNwqz8ze+tsQCFPTYF0c/SXG38GZ3fqAgV8rbcW/DM71xxkomn40S
KWwBbm5ZhuZllvknc/3nLBbo+PE2kDRhH3AmDk2JCVfsV1iJK5OLsRxjDlQsvZRdlMv1nXsyPAJ5
pqKl3sbH0vfGQHWCChMPsuYqsFxWctezumdzXB/R/SaUsz+jcouHDRN8h6Z6s6Vgdw68MOkjhA6P
bBXYhlwIOuq94vCyWDj20m9N3EKuKUpd2XZzmpjXJQvkPWgh8DkIWQQbnSHPiTuqjXdoDNvnmBtM
zCYhr1p5M1W8yKHkF0x1Hewi9naVl9USo+3t8SNSWk3B5exNBk7QVfFejDSTrwCFIzZ/pz6H5Uqd
M6+fvgInsNPMLRYq29bbJdtfJLS2IL47SmXYlFttkxOXrl1r1rFFOQMGAzYIkzMJNCU3WlbeTyvD
ab6yu2ucs0+Lpf59b5jgE3IU/ZARl2gsAw9mCSjlxF+f5uZVDT6a4AHH0s21IfNhR3sVbzZSkXgW
gWuUM/OQUM+4qIanFUJD7usZxt3RE/pCEWcT+kh7Gsu2IPLqsW7zxplDsdggiflGxu2x5CYyjPau
BZIFN+1dT7QfugsjeT6beOFEugH3XzD1+ydUwHUWtYZm/0SkUlkOx4jfdN+CXjLfhjhQ8ZiFctV2
EjONjSHjJQTaUJ0CYmY6TgI3ka3xxrGdJYhidelv2kWMI6PtAtEhKgaKTCWfXhaH1KqYc5Nrqm9K
eg3dBPEfjjziqx538JGv2XOUbHHYoXSh9o8MFuX3mVLXI3qqqIFvA7JKKKY/Jxmx8p0+1RVK2E5o
GYG9m2uSE2R6+k5DziJu5AJwgU1GZZbNOoR6Y1tkEfYt3RAJ93UWofce3BnxOh1ibDrBcJ/3lch/
wdzvOxsK36EIji0NCWS7n5StZxnx88OLILtmujM89UrtvjgX99J12nn3ir4XuFyL/IaO346ek1qH
aCgExXhnzHFsysJb7lfhW0w/VTmCQtBrxM6uqp4xS9uRWvXbhWps9dt5YzsuIdbBEnC/1w/8F/rF
P04nDlRqyESq5Aj7fs1dO8F5RkqS1FIkgRLobz/lmYeoy/p7b4iHy5bcj3Z/NQi/Y5mmSRsFhns5
u7ui9MgVw+tlPlqkVsRek4Vn4B7YlU3yM1F1/YDTJPxWOFvj61PbtjSYAO4NEYII490r91zT2pj3
xEfoNrhq7VGFzhDVYQvZ33Ob8VmnrZ9NmnEHy9PU4ZMwl/xLqB7/XBOqrpuIkhfLkfQEv2F4aIhJ
ZUNB9k7L9qLBI9c59r1fghrRFOqdF+xQt/B+HSB658z3bEj3WR5Ib7z4ejay6Qum56DOHCCajMai
ABZ1r+o+X+H23OzhHwdzqEyKZzw5kjJKVuwMWIetB+xCiPmwjxLxpduQ+PmEi77WhCsRozCe4U1/
krhdyAD/2KdvppyG4oWNcfrK3XXu8dRuR4Wm951CcYd5RXtMhOlniJg1lEtFA72k4Y55qaDKExCE
oKnnMPccs8/bf92z7Gd08NCNPz6GaJ0BUO9B7gcLjbiamEehLMz4s045wc2FFjdi1lFsT1/p4ei1
c90AGjxMCd0dbeEr5/F+NXRbFLMUR9hrg4rsz6u9JVGP0YXi1xIwaj+f06IC5EKoDNlhbr+2h845
5FAmVotL0s4qyQRVkJyYN8dcFgLhqmodmXSKNtW1mOC1JNWD/LFSvX2XbwVe++u9CdBik/sqzOvt
TXVHw62/GI509gufzY8XbRm2zuO7oHxhLlGVdxp3IccDZvgcwVh1BU3FKyAx9Ey6OGH0vOEroXh+
VJW14Dq1HaopWzgP1eyXvFiFIUMFfEPKFyLMNRYkVVOD/cxkz7gd+ljkziwxsqDfiQcQqdrKcCII
imvJMi2OiQ3otKMSHKjSCxBikYLHR5alr3ES6Do0F13ixF0XQfLCq0POI20StWX74RzfNCt3QdHt
oQedFsXu+XuLPJDH3vnj1/bTuK41y/0JEAaWFOUtrY8THTplucc6ypSrO+LNJzyln2y9p8w2Fhb+
y+4Nk6KJUIQ235IjZTWZ4y4wc+C/bY4FvlaSY+fq4NuPVnpdl01I0RRBhImMU/jwHjJs0SX7DDST
LO+fp84NVXpfTCggd1eBoCctnasb3EMsxxCKrSFePhsN/Racl4ZuVEiN4ABXrfcJCj6RRoUXLGm8
sAtzjdqgjxSxTXkKD0vaKG3rPnu5ucHl9skqbVeGHxAT1agI6YtWCt7pN1m0Wdw5f5+MriKmmB9s
7XTfB9I16Gs0TzoxGJ9T6I4nVHn9/v9CiecCVizqQX4b9gtJNNhDv8WZhhZS2syLQIbwPERDbs6l
n+R2uF6rxAaXliL2/vSRMIiTVpUKsfKG+tscNqehybpT544jMkoawH0G45h5kAKgjY1QZ0syKAvT
a9CyrhL8K+d8Wl6oJvySVx/+uQFchsIF98MxK7Ip+yJ9qJ2BiYQU8Ui+M/gu+ZUS+fnrMatKpImA
OCyIyRVtjgTQT/zAxjh2BOxA/G6W2pRZbmrEyOXSXVOjDsY4cFNt6s0oKCIVPlWFb3Go2uA71gX6
S6mPszMzdQSloP3Qp/9KfZmcVdN44sGmUsrLIFedtNYHpUyO0O0AavjnX829t+wdVJI/fKbOJTCm
v/NEDHXiQyPThH/P4vKGipg4WsQM39X4W0ES08z5IRCTK0qIpg8zRrqmivhFfQQcnoJBG39zptWy
MgTU8J/DbeuhJFMe1KKQmB32RKMfVjILH6TnBpPOftsEx+0rbKTnYmSArFJw30d3DJ9/1aPnqcYq
XGRSbI6ITzZP61FXVRVRv6Bx4yDC0tnM9E+3PM/5gXCMt+zu31pbGDAUcB2v5+6WCHkO0MKsumds
7oHTX7bjULr9cEUvJUz0lAXrWr9VyKWM1NNoAY5dmwDBAhj9jtEawBwpRHLNPGsnt84LUK9sykfs
QiY2a7GZBkadCrwk4CNzBJq633bP98K06XwyPRcbyYAD+KJIr/YSJO96B/8PHY5SEXUtTGF1DfwQ
/Mer7a7M5olRE/y3ad91rhKVvnggu1hmICkGs9pzOEbSAlY1ctsiK/iOjwFLHwGITBfvWOa4Jfbr
/HQ7D5QYGre+qWIVpzwENcsXIJ66kQI+s34vCPx9LLIwWZJt0vKwD5XRH1B4rxwAEIfThKwo2K2W
nvz9ZFqFZbaqRS0KjOxTpFN51LewZDwNLcLFWIM1m9SV4/e/oUq3iZl/7lrDdBhZSv/UBp2hdbXv
wqQ46dD9bse8b4v/cReLj5sK1T4L8f2CcTjXfnZzYdBKzbed9eZbq2gC9LoJWRanHqAYM0n6EEo7
/ePyifRPvqtL/cSSD5vHeXbPPvNRjIdi9GWSrc/Fs9QGAeXXbBatQFVrkoTfyTlKKwvOueiPEiIQ
qPsUmK/s21ZGJ6HJeEVC+yYiRf/Xr8ApM8JFQLW6K1jQrm7JamGyJRxYVz+ObU8frYy+BzaosmfX
jDO+2HsiW2sWBNBIrbcfk9dT0CMZA9rO5gqnY8jKMp2MceXiEik40YK5IzLysqNFh3Ie4F1eA3dO
84fT0MS85e13ZHRVAbUKGRzRBr25D0dSFf1Qu+0Z/zF8xN2bAtiTFhDzGQmlQ+/MYkbEsEL9RrPf
QHAJCb2UTpKOBlnOs8A37q6iqK5eJ6ovTrOr/ydj56CJ5RXleeGcH0clAWpjcGZMdSuxnAkrqWry
49Z61S7JWZZc+sLnlLZi/CGDHeZk9XIdFXoow59FQnLjR4ZDe9iWXeMQEmkw52p1lU1ZpX9x966B
9z+WjlJjfbMnIm10/w8AQICIOCjP+5zb11ZYRf4aWUx6R5HHxcXhUnntYwqVqyISlWKCRCgOCqp5
JGNkm+jXBpf5uGPKZp5jAO7bVAwqEYvsHEaf+wjrWsDJVflpT3a8ujWloTFxNfgHYwjlOz3PgXSE
k5FeAlsKe4TN57i53tqrA4yZ+IelsR0c6acuEVXWPxm0a5xcn9EM6FMPCvz3iTHKAua+QcvDd7cI
SBQ1/KU7Xy721nDfcOcJUkArioFpEej1XQ4hKp+G4cd4yyVmiixychyU24g3Y3SeZhE4xBrf74Wb
sOHtUQuz8jpbQDA0jP4kaDN4sMDOntFwSq1BgaSXSC5MZC2SG7zpWu1V5FHJxrtt/Qx8c/54VYXO
WgBMRtF5iBHZHNJPQ7LZMjNcbKmIvQAblgVJad10Hutm+EkokrAwVsUElpmTYfPrNiY/Uh6EthYz
n4jg7yxN9ZyqQAGlxuyCzB/jy57hOtmGep6tLTEMqv33Pv+nrgerQGqojx2CJvm+0pfUpzjFdZ1y
uoG3G2CvtfMai95cC+waTGvtVtpLVkpAkGy4a/qSPtWaMgeafXqbZkCEN84BM/Da5CigIWsp+Bfn
EPlaOkXpSO+ezb9fEBw/Cmba+yrrXWel/OlcyNY7X4xpO3TTShQWbdV7P4X3gyg23htSljuKHwyx
lYIDcbnfv6QzrpDc8QwsqhZH6JqA0gXwCJCystrEl6hUUHGWOefSfKduI9Cu3H2iDzFlbpMh7CXd
10KAx3LCUSMWZ4Y/WmxQVwbisytIn31bqibKv/Td59PD37d9ttPXXDkgrpK4T+lXg/az9VXSOAef
z8NdQPRcprgdh8HYU/R9XchJMfkrbniFhe0wJa7Cd0GoWxe+2jFMfeiCVoHjCczZAVzB/lu9TZty
YHBPrmz60nxewPF6MdN+QOmNxk13BRjvw1onTkod1/YkPMcFgYTteE+MaAs9oSTncZPr3WZ1zGCf
+HnShAi5NMwSjq0gIjLDjLKgeNtarxwSnxwMUtViZzeMTAB7KvGn606dqucd4wMk8whFrNP2+bRq
GQlQvSPq+GY6of7Gsjy20QE4JBQXQOzhdwCm68ijIns7ew/SI/Zh7JvvG7tcc3ocPrs5zge4OybG
EeHbMIyZ33FVUzr2SQNCxAr3IRkHYxnBMfzgBjecF47wZ/F/+Bcu5bWqyCcxVUOUWpzwZWbd4otW
0z20i2fNHJzeFjil6FbZQPmPDTKXpfP17mQHAo8UrQ5Ztp2SwT/obX3oHZjTgUF2kQwD90eN6usi
aWvanY0uxLeIo5wd+8T89GlIx41Hqc6g533KbID5C2KwQOW/oppvs/T6bsGuxgxv2dLPfV+G4uZ6
nrub9fnZ99pZ7kaI1J8O/cDrYFBOV2OQjie7rjio3coHyCaCV+0cnzSqmuBs62gZvsOmGjmFyCoD
R/8wb2uI0yzkky8DrkLhJhjKX/JuKd+jKv0wAXYJlzihdFmvbvdxYA7jhl6aJV7yV46EO38ZO/z1
no0E3sXcuy0p+Lpbr9KoXQzjX1NLrZsouVH5h34zjJ2YAuBdBsfnf7VzTc2aUS2AEoQ37I761guQ
2YCX6rFp5dhCzodFnmC1c1V9iAZNp3wG0T2AwPVecrt30BP38wDNqbimqIsP7Ggq7asuzdrzEcHx
9utQMS+h7RI+4XMO+gWWTLptbmec0NuvyPGP6z6AswoyrlrHqyfQp73oOXoufpL3gtsdYEzA6GJj
RiuS0S4+UKV76JUqAPRG8JKIRrrvEEMOFDYcN8PuqVqzVBoN+P1m7KtMI7jTz+YtC2kWjr0w20SM
OgDUe6RPKG+qqXmvpQXucB5FoRH6MexUdpzcm/aF27Fd/e28bQEZfEZ0FhhWej5clooelmMpOJHe
NnzfsgLKclofL9Hm9XY9Y9miE21xgKiyJAtCoCfnIV1P+5sq9qY9EVboBUgn75ugHOuuHqEEOUyI
aI9wfNVBrsPiw1qK1xwvaiWREmmiDJNyMLiw/7Krar4YtV6e36eXKz6qZH5/0cmPznOdmRVbd+X+
qaLM0U+/A+MYf6ZAbzxI/JYMC6830Xo0OBiRDVDP5MVI1EhhAlmNcSJZJU05spOr9/z496x2vTOU
NNbCILwkYo2zFqYg4TjRROZVCbS7OMuztuNEC22pgG0mgJD1h7Mh9ao8PwpE+rqSH8jTenjlRQqU
rpRp7cVkZcNXqEic5o8fQmz92jPSebBq2lvRcDuV4zlAomnuadgDwC75Jfms3fYirWluY1X7WEwM
OtdXuUFn1IEc0ipXS8L0sL1o70iqEB5o+CVaRV20NlvYLVgfNusOWXorStBDkGw6LlYgsC3SEw8t
s7GMoUCV/a9bJoGcOCUm6wHiBoOZa9GsnLPDxX9jfLRHtZ2nZc0F8tyYM/HS3PpTnyoIrGC2Bwrx
9i90YQdOBkCFH6ImGe2YRhq+JHGT61lf3ArteNj7WPVM82eSl/eTVBQeWbJjacAiCLHoP2PZNMHS
bTaKwOD/7mVb7jRSkASZ1HKJjM/TtaQs/cocuhExxd1d1o9YB+9FU26Y9d8GdkevxFghNpxAdJdq
Qq91TbbUJ1UrfF9AXSJX1HIDpDDs8INTES+ojHYNrfUFB1psZeBn/pWI9ppUkEmivLPH3V8wUwyq
XZ65uMQT/HcJlxK6E4jrddbK2bB+BQ/l0l4+fFlSp9MUD2xUNabGJ2mFA5fDtq+MZhTwJCGqyVtQ
uNT3sTPe+Uqcce5rXBZZ8mcR5WHYxXlhDu09CXuZOJ+0R2axSMrWDlXU+c5HjuMYensTsy2UnX4l
y/fV4Dn75SWCRYYp28I7VwMFKv8a/4YWPXJoE/RS3bjZR+ihPgx/hDN9STIqyKIzgfc/Xr72kfEd
ONyz02fA+JzM+KsG8TnMUgwCElxWbJ962UlGC+Dbin6x+pNKC2rc5Om3kMXmtCXx4eUov143RVc1
bSofllk+1AIv2dCy0wKxyHcmv7uidMTt3MeByoSr879lvsE4Dzr0n72gLwwwu347BFL6JHlzQTay
jcNvtGmrfln1f226lJUjhk/o+zgq2ngUpJANJHtuXV++pVWLRmUjGScr14ELv/NfQrRm1FHvzZo4
bddu7skuTNJAkIfOgpPuhULusR3wl1BmB3p0Ktu3ELIk3NZwcvJgS2WZp7S87XCoWIXM60s1nmox
V8e39T4QR+Lw8rZ4VouQlZSacqCCknKE/YWW5wl8hyhNqYfaNjHBzrWl9cOL6N80XtOHckD9cuTI
Y1y3VDR1E+6jTSL7q5xLVHK+EWen5dj/s7sCtqwlKyOPnHjy3eB7Ezw/zyZqtffOP72LhVwLjjTL
rC9/5Jzmz1yKAfi7/sOV5dVXJ//reuqF/2wrhtiIfVuts8T01FsGl5/YOIR9wCZjVsX+ci2QLAMU
ipyWalX/aTG3fgUlfsW5MQk7AdCrWpnHdvdD9SKmH4ddpbo4sy1owyaRw2wfW104vB/DY7uVk8G7
6wvSfub5m4if9Eoswzkr/OFm3jmILGWftINM2g7+Eq/6sjr5PKxxkNzR8p1bXeUtt5BmDSeFL5PM
HXVYNtgDIX7aZP39eSEACpJxgaWmT5FxwGTxq1VcTRuUeO8mqQbsEhFrpbgmaXDMLCUig4vzzLZ1
ImDX57Sz0ys2tv7xFFhUl9hml8MKzek6A9VFuw2C5UmgKbGeEndPeABphBOW36G5/cx/8sbLIiNj
bvrStTYB1pDM0x12DqYxBWFSXy/rvy+1c0dCdSxa34NAK5M4I3FVU2OTnStbkDg4yxm3aBGHN77x
n1/6gy9aQUi/yT/RPlI9hSa9aOAhQs30GQ1MAnsJg2jXLaOO7gpnwoF16Vg9Yl+RGUbrNS9z6Xvu
EtOQ+xjOZttAVX1Lu1/M3c4d0Glvre9RfAzOLHpG3gGYWfKMTpq2XU1pBJB6dUwkfVPgGkecGuXz
6Fa+ctsfws/M0gOtlQYdQhEwIoestzNzUR7dFLO4FtNwbReOcNNlg2jviwulbWSL0+5H13Ujzapn
VWWNdvEdVTnU0bGZMNe8wO95GYLlN4PwLrX8PJhHzIIIeDospD40nTWCQzBypDxCrVk0yK25a+t3
stbJuGkr0gr0mi+OpYjtIPVBri8RqJyg8HSJiQgiunhUZ6UDs3xKvle5nyT5/bbSokUZeL6hbJKT
8onAjNE+0IpRGgZl5LyixKpeJuNbhqUupFdwgmpIWmIFPu74E91kMSuiuEsbcjoumyzIXo2T/lW5
Wom/on3RTrY7mkln9eGy2GRm6tH57qkSo6qNeS4j86snD6vT9/MpRoJMirHC9Hy9tbhOJS0YmGG8
0f8c4qachs4PCD4BdP3WCN3E2Ox+RzwkCmP1opcPhcpxkaeL6TZcmDYrFol6zZ080fECQjvCnErb
7cYSB7hnK3rOSwARQKieFoNzwRVuU/Sop0nD2BuswRq4ZdM2m9ztpgKwWxcfMUD4lIBfDYwpFdnc
nNrRg1by04CcKW1Pm6RUZOARX9xjE4pYyMR5FMTErBysyTiSatXEph7wXBbQIy23GMblAShDl2MV
OfyO6L/qf8KsT6WkI8NPcKinFGH4boo7jUra8UPIMzWYtcyfV0hyegajLlBrlJ4mJbYr/+FTMN0y
xpZexUCcxctbDTj7TRBHUSt3W9+VDfOwxj/mDzq1+N8w49YddbwJnv+TUhM/8ngv5A1eRZdWLZ67
94UvSiAVlo/JgMZHW/HYhyuvCb0fuDufyZTmcTDRR7zMA1fXvCr9GDc1LcoPv1qUNs/IdJkyDAjg
AdoxI1lBdU2Rroc9+BndJgA5Vo0/DGJ4iQbQcsjVKJgr8K/o3OL/rZy1++CTs2s1GpExeDC0vT69
o+352W/Yk2HHIzSIKLHPk0I3VmECi+jW2RM18FLDHBlpsGu68dRXyGM8X+F3LtaDNqnA2my8Hkop
oP5zQ1Gmd/D/UCVyclpt50f0Kot5eKgvjh2kl4cdr+Se6CJa3Q/oh6mOikBD9fD8YAbXxCgJN1c1
wTsGRuXyXAtpTvyQ0lO5pWUlduRC/8yB+7hc5bncm0dXpf5xz4PGBnbPgCdy29Junbk/54aB/iu2
7XQQ+G9rYgBZAkZ5ntQGQlGlYJ4y4g4llyGDZRL+Ei0suiD4eiRDJnmhDbRAtWuA5bFxDdZVPJAB
ydBto4X8o4OEVdI50rNC/la6LAa+/+jL8W5IhQlLoqmfxbdbZM7PpowWABXMuogjOG8kttZW316H
4zW0IQakGj8iBQB/G7eCPAhc+PZROa6enia8Pgfnm0Dt9guFXEW8hiax5dYxXI0Za73dWXUmlSVP
+/gszR7D/CHcod5CPWRpsvumCbbqc0YPa9WXfdjLgZxca4hVabAsU+rbqAO9E15aPFCTh4zbZAZ/
ksCNowwf8zoua5ixjoWBj2YBaQ0XLR2J+Ort1LMEQHr7d47Fp5Isovh8H6z1u/Y28GHGxTVHT95H
t9GYn1O7JKI4ti3LfHXYyWUbTUmdb2Hy5WogdqzjP4T/tg0WKsXNDe5WeajrjaDi5+NgDiCAspk6
a/+ZxaWiUMoJ3QomeTlvYTuQ9kaPF/r3Oi5TzgqMbZG7Dn0Hn5CAkMoZCckupKKXbCUXQkYrXXJz
xol6ujGyb334qQ3/PGmORBUp2Ir0j4zPXiCFvdvXaDiDDbYhS2Oh7uHw3u0OgxPdBIUtbei7dMFJ
XSfnrtkuWAlIQPdpJRvUxEloyRWRi3wTmbo3F+f2/8CsQAG0ubp/5V9Lyon5xI3CN/5lhm+F8Pv0
nhnrkKJba1b7m0q3TNojplw4v+RXVEVAd6YTmKSoNHKUCfdNE2Q4Has2wLFj2EH5FexvHM6h+NWY
XDghJaNB/1uPuNvvLY7YjRr7Vxy1CRGnIE1PMt4NSQhrEn5j9NX+VAk3c0Eqj3bYlC2UJ5xTF9mu
H/VFxLPft/Lg28Wv9dkEqVJZX9is47lARP832aPJSkF0c/jLivUFx/RGNwsDO59TNkdjUbdJ1XUB
hmjWNo4+bw6iIFFu7tCCSfvHLGo5AE2O8mc/OQXMnTuHc7kltQ+7YwJBLxZhk1pkEsQWUY5rRRzE
fAguk0YbTFY0qiPyKnVsJadFYnmQM6OTIhykCOa2t4RTOLqdV8VU851YeUg5Bs1rsmV5BQLxiYF3
+VXvHRF+G0spt/NvyiSGav5F07QVoEWNjD8DHlba/tHRbEgO7RiU55PwRjsdJv/42VSOI+cF9i+a
jOesZnlI3XVD1aA+CLyOdB2izSCMgQ2tc8fg77Pw952dU/uCjoJpdOjS1DuD5Rn8Wboi4TrnffYC
NM2XJa4KUOnEWJLJhxRSD6UKJVW4dSt1uvtztRCqKfgUJyvhZWG46GVcVJdVXRcrsRMScWPo3E/2
bgMLWbGiL9uU/I7tCHi7WnCKT0jUw/GlSdLieSr45YS3clsCI3RfZbr7YiFeCNzG6zuJmdt5QsV3
3GR6CvIf0MrQsDHrxzTldBabXAwdZ4S06/3f31RqyzbxrLDg0y7Pj15yr5pLyCvAwpSB49fP6e+i
FBDBkYPD5kAsoF8wY1d879HXLsSYFL6JHq4BgzDutixG4tftydhYfu7Xk/684RUkJL4a9wDaG1EH
8gjDHxOxG/chOKIrcKnuLplWSu3zf04/EOPZRtpP1ry7qYfCg3MuiqNh25x0oWoE9fFZXuHODTR3
sQx2T+WHX+v9jbU4Dzh8RNqn7cwX7OJv9GNRZBF+YOX6+sLP4B1pevTE9tOJuHzURNzcky5TT4s2
4EvZDw5lXZqn88gzVcDr3XvuK36925MIQVodSmKAeRwM2VIkBEyXy89WNMFk/NhE0e/I+0rnoGrH
uoEoLAxinHdLYpIazqs9GXpzgv6iwYj+3WWGc9p64/k1mnAaWXNoM3LXxSsGwWIo4KgwAAubAWRa
0K3+9UtBS0EHh1BSPEjKo6uNXXUXsjhxgGApXLJWQl0kUaMbmFsa8Z1DaEDxLzEiw6uxCX+w1olp
FIdAEGO+048cp2PCmw9qKYez208+v9JZfAx6r+uZnhziPhXtqTjeZJ+K4PTcuEwBQ0LXtDOQvtnG
/WR6cLEkOm4Lv3xpk3qYLmOlgW84AnfV+jfjsvHp/411KajHlzO9PS3MGxX6KmKGluxLHCZhANCs
DETy8wdGSDmtQu7r/+sxM99pnkuYQps0xNWPtvfxnS2tRdJDZTqiqL3wRsu+008vryFAZfChdQPJ
3yo4svxbuwJ9k3Lkd/L0rkEOjmxsnCO5J0x+Aqumx/FbGBvN4UB7Q++YJHWkpZBvFAe+bAx9eXwS
ilmz/cco/CkCrYO/YZT3zHNG2kP6Q5PNp9WPDAlGh6SHUr3COXdRM0WNvKY6D2EQEZQ5ygT7qmo8
DtAD0xsZ7SSMoXxZ467B6TCVnlHykK48pfIOPrlw2p5rxdrcyf/+7sGNFR0OfhiK7puNRLUE0rv0
lEDBQEs+mAdgxjq2SpNN68ytJKOvaWnEwvMsy3WVQGB/dQnjt6eHXfie8DQZKifImIotdNaXcN43
iEDtQEDSAddsNBTm/4p2zwUsXGKccHXOf2bFhx+9dmIHSkXsLuBz41OI0XUmf43ZS9PYvKz69A/k
r+Ob+0/g8h89i2M3X/0eMZOD77P5fRDuS49fsStgmFybszTsuwL5/ZxrPMxSrPkV4A432X1hZkou
mxxS+xg/692nOlLw4YPvzl0hKmZ2GGMEc9F/PnJQItuVUgSfXV1hGxTiljjFfBidl86tTMbaVjup
Ip8UjfY31TK/Dr/VB5lM2gd6UNDJSwEdbv4UDv9/h5Qb6Rx0KJbr57iUmlIr+OfEwwUKDr1/PdVm
7LvtibXJrLQbL4QR+jgclTNjqgv2PrG2io9QqZQRXnHcp5m4mXWSAHjKzjOcr22jLOR2D4u+NDDi
8KqnqmrNfUNb
`pragma protect end_protected
