// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:36:46 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
db8YfMSzUIFofhjwHncMH0k52BLkCjuPJ37LfqXONTf5eRudvnTp4NlGl3uNqnPV
F9RfGbcrX+DWxr2EaDUIdRKU0sQ5u1kfZMxMuWEcyNjpRy/WxmSYP2kOEPTTHVtj
4UNhN4slTDw11tp7UCUKA7645pX0adBL4wPJ3oi0rBg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 46192)
nu87pFa4fKdBx9jG86chWxnWDf1DV9DZg6VDXlgccVWjvM932fP+he1542t08M5r
4g8Rrojm0Nb30BG4WD3pM02AfJ7YPHILLdvSU+m7DlVuWlWbVYicb4KV+FZnXnp0
uynaPWNVEYu9tnHpdqrlFJ1qJANeQTylWKg80mi6QjrlagKlHNxZWDXJmBi+UbEO
5MiaAHpyI3TIS50yfAaXY/rpiS4f1oy5zKkpKIdic3tN0NzyyT/6MoLOxOjvr1Hb
oTqAH9xmZTWfs9KaRjnckugPvszEEBE/+muSF+G9t8/dbw1T7j8CIvFatjYdoUme
fjL5YTFWDhxThf12qMnsbnGS0AfhM5INxoYjkrWBbg7H71cCqNEJJBHJ8CBp6LYo
sXxu9cuXSJ/NtCDyMZVOmyTjBMEJrFqALkU7+oSkAtmwP7dUhQ52TwZsiVgNmDYa
zskZUwl0gtd2Qb/ABtqkZy0Im5LOZ8Pe1jrP6ekTHbg3zzAZg6fHsyvNonCjnxa3
HMNYffQTnhQA9CrfLAUUrtofPsfP/VTC6poZ8P+NopZQYf0jGHoY4pZgiGId8rLz
TSdy4TKTEfa3iSn30cMTRWoHB7ieylwusGFDiqziJJa6U9m7+F9efDPqSVxA4Wix
AVumVK7s1KvpEGnwsxHIyLYirDGYRNyOaqYor0U+GLBiM2tpSdOwZb9L/1LCdq3y
GyFHp0/Kl59dYxc5bBNflSjZUf3tBtcUhJc+F5VP1DiVnE9NVkV2x5sD6OzprFD0
Ysm6EFzXfL34SllmZ9w32d26ilHfDXqg+KAvGHH/5+brga+0xNchMmcTAV6ZONFW
5jYh38KFvHpjBDq1yoQoIvm/UTTLMus/G1UDGjFGsAhn+gr97iFyD8zf9+8JBX1K
DugavyZbZ9CFb528Wmxr0aIU0LUmRPuhJJPTuO0UKuvxljWxpRQxmPs751wuf74/
WpmGC3WnUHuYHzkTSFCRmq7S4hk/Z3uM/qFRmitUn3+4Baslklgd16sWZUTUDDPu
Gsm/zK9iV032ox8b8xMJEuyR7lnQmfMT5T7XeGdggRB1zVveuf4kw2tfGFgXogna
lnfx65Q9gJUjrDPs94pGIdpok1u9ThmvvXSQOCCirjL5gxSELu8jzHPZfN4fKF1f
s4qAOY26+2o6fi9UL6DiP3/UmZizAz+MHJ6zuRmyphdi25cMvMDWd+f/v+zJlnrN
fHLV5uA0x253lIrOOcXPwT7+EWbB2mbxAU67gd4X2rtYobH4gv50MBdSo1J66uP4
CVJUyrlD+f90F9oRFz5ZWwSKw86pbf/HAmgzoAVvXyoqyb0tNhvVc/n1Jn6hesxk
gwwH9EZeCPe6BF2gpEi0uD6xst1qyPpEGQh3CrzD/qNP3awVSdnuktUX+6i4GRil
0PqR/CAvKlaBMeECCcBRYNlsiX+BESptAMyGtQII413wZ1U7Lka28P7/Ssg7A+5i
z8FwoRE1oLS5Qzv6NLQk4GFJ8cWs4h/w1/b08L20r3cXXGWdYqU0OH3q6iNSInxS
OXjk7tjfC1u+BV4nmzOni2CSOfIx1C5swoPVeLUGxxmMYRrbLnP1hmnGIhtl5twg
moBdrM8o0ofxVfnImL/JGPk05Xjyg77vSUWQH24ZxMx0jGZ+xCqfbV2+s55Uj4qa
hs7+65oquKQVqORLUFayw7tmyY6Lpb99gZ3llbKuBJM1170eEPPOJyl5Fk08OQQe
f5d5rTRRCoBJjdYPsybk4QrHpWbN70T1b75AXNOpDjIfZL+Izo0fdmOmMugaIQbD
gN9RNCWnx4R47+TmqAXLf9PtS0JNVpKODSCBdeG940WBESAEY+pOKbb7B/3o0AMk
sU+PrCJoO/NzCL1RaqeLVcjfVam00D1ZxnuEumoFG5o3mxvI3NvwVtCPJrtlVqUd
8IzmblN9GU6mhXmXNVDXY2LWRmCeJ9U4eqv1NwTT1s200gMPRZltL+gr622+gDlj
IVPSW5bQWu8lq48KT8dpq9//Q0p3NWvVUZMDCR75gf9qU8VQOAx0pTKeSouja99K
9w4odR6rZFJaZLB5OlgovLWP85Y5KIR45xNQ9b/oO35VeUDh9LXVdn40hcCZOJ0v
K6869/KxrR0m8e6hHHbIlBttmwt+IBuAJdtT0H8aM0JIvo3yUsHi+qbuM7O11l+1
1FNNYtlHAh5TwOcpu42kdewVckuHnP385Qk18GmPZFmrN7Tv+yh7PGZNGorD37wh
hVhLuJ1C/yxqLEDLkGqgutH/oI7Rqh+I4imntNuany7UUB5Y70PocpYC6pD3ta4I
1zWqqlRNNelC7+Tv1aDRW4DM8OSvHxncz+UNkKpv8GBxAKX0d6V4RRgM2Z8dgwEP
EW2JnZeHTvPjr7EMaWbnEDl2H/wKxcIMb8cm8T5Si01U40nwla5zz82oeE30jT+G
vnU4G6TNdZ84v39zSAn0WpPHN6D5QsUUQA6nfQsNVPoFbw/VaUU9qkmsYu6f6lJ2
x6PtyXhZHgAA6Ozzbd5XuTgeurey69d4gKyQGw+g6TCDDlBA3nc3BsnSFMa0mYae
/E8Jhpy3RdtwIxwSO3YYfMA4l/CGMD3jPKS/KniiP38LwLvwtuW0KWCrxYwDQ2ta
5WQgj7a7RH+XVnQbhsIvtK0E194bKlY7zn1jOZvO+RKKxe28ihpYX86/Prw3ZgNM
9Z4gNGFKMZlrITNFTMJuB8uBGyYgdQthA40q/tK5bV1aUiMFGh6MMK3fxlovKi4Z
TWeVyx55pT9jx6AyIQfndbj8+/Udan8ndTqFYzX3jhdDi5xKFzNUhBjkfP63lqHx
qZS/tpoquqssOTPna3rKuSJ3n21bOMGg//+wrYwaaKbZqe7bVYKZbyFM+VNnyGAK
FdhPkio+QhhUW26akCz/EWFMJNdVK2A/axi+39zgoKYvjUjQS2rWi1XnVRsmK59N
CEfC0LwSiU7Gb3C8KDurVYpoomD0HZjjiwwJdqw+TUVOlU+kkhgHs4BgPXDZZ1FM
Ev8IIoV1rht16wLse0ML6KG1MGhs5fn/FMlLWPMKh1zB/Q2HRsQIv2Mprt7t+uTc
YqLj+rKVqj0aNTbje2X3Iza58DcwfIl7GUNXSA+8/JRmJuAdjNn3SXJnJgcMEDYj
REi1X3gp4v3aEG/Um13h8K4xGcdkWA9THV1Bq6lsmvkix+ZvItd19fv3M0zlQira
4479iDtmG9qrNdjsjHsLVCsfal6jz7umioq79wNcPaFauJN3z8n5+jyJ+oA6DPtG
OyU2cZiVXDPke6yUzV57oNaI06P+G25WK0l/6ukkKy9KUyVsDUWcy6FoQzNDmPSL
y7N9NLsGDgBtXg7QclWr+nVtE3fv+ddre46NpSTErNbqt9NQ8Yl9bh10sXmQdlnG
dy6GG3I4qpjafw+f9GF3wXOTdv/suKXk4iGdP7DDeuni+DztI+n0s/ocisnozYCR
gmbFjgvurAo04/hhj5mY+/YGTiGo9jlLoFDf/xQIuz7isEv3GAriKJwwnTTKhA5A
R6Y6d1jlF5Y6oLHiun9rQ8tAoJ4oPSsPH2rpI/nE6JsNfOmK2Jk1EyieHRfcVCK1
lWpW2zpuHCoMKa9AaLd4NVYsF9tY+Smy1g6Ok3hrQ0k4rl/qT91Q+Dv6iWdadqnd
5TJrbz/7DmlRp1T5KuHxVO4bWlDeYayz1rnct5DcvG1ognRFk5xXNSMrOIjXYRH3
We6OpO1Lgfph6Kh8aikL1da0KDkV3wsG0qrxqIJbxtGe5z+BQlXi5P7/cavlLuql
k+1QaJXdEnH9r79iylgC3DscH7ydUpkIXw15SllcIL+Npk/Vngn21KRhjIN/peZB
LiYwQuvj8D8y7yY9nojXck6xLiAyABdpES8GQU5YdavEbzQQHk6xFIy18faH81S+
3/HVbe2SntNDoghyTJlDS+N6SybC+ko6qoV5CPQH1u5e/P/J0KTw6MnGtJQvfgdO
X0xzqzZjGUi3yW+Tekv7MEKORHtLdGaxuaufQCoZZe22V+Kt0VG2Er5fMXYN6G1r
8foYmNFytWEWddUYEg0skBG5FWonnsHcJ7uDo3TTE5E2o/XC3S2WAZqYptImmzZC
JlVcs7v9svB3m0NRUkUujMYdq5+n7ro00iVjTNNhqosrXV7yT5j+XH0akzTJW+HS
Xpqq/QQQ2viNLX0+c8/UrF3QTtlWI3YxCl81qJ5kqihGbuJjvF/dyIrYTdHzoLjX
LaN0NJFANiLto14813mvBnwOOLusckOsn9bHd2ei6uEQK86kjeSr5JRG/rvQho+j
8W2qO4Vshf7dxh9eUk0fzaVozL3yDNqdjL6QYdUiB3D3NiUrMmwYO1ophPLpvmpA
dTRLrDpam+1pcqBSgeUuXzy17xxSTq3hPyRjbwl5lRrbQBp0ClkPRMAFZHNmSSkb
iRVwrhIyWtZHrlPTS2glZLbdqjrwY1v9eiNKRdRUm5ZuyF29vwXLTllzp/inDyY/
+PHWVZkMO7H1Axf2SSUl5XAIVVcQxkof8lK+Lg1Rul2DydLhTEfOQ/I10UTDp0dE
e/TfVCyssL369xHWv7eDZfDsYhA1rjDJdgD+x2Q1nX/XqGI+igWgIeXLc6ZsXHmX
jdomAdrZLONHL8sTpdxH4pFUdd1ihCzGVdCrtR1uzTJ4SkMZQY8CSx8XdKqYpyON
AtTPdMxIBWBCC4Z+V6jRzSjy+GBOXuaZBuFmOnJWZwF+ZnCakNWIfaexbeRKcbOb
iVOjCi09q+QBkGuHH5OxK0EG3z4PakT8oLh8q2jgtaWqh1ZqFeSjUIA6FM7jNL7j
qHgVUz/EXoY6maf6PuXp7Yg2eCQHWZj3rtW0O1QTpZ48HfGrQn1Dp50v/gXOQwso
m2cyT5xn6p2U6Diz3LjyfyG7CJlekfXh+qGBJJiidEbPP7Kju7AfIHoMHC6uP2Xc
NBdBDIgxzpBpxufG1fH7C7kUBwdgmiC/p+QsqJPf2Ep3LQd7BkW3VnVM5dqSr6VK
QnnGnuZBkaiIlqcX05LsX/mrgNBlGVJJWJ+X2Hu52j9qpZK07JgpivWJpRxN0gqg
qg3QAvM7IpJlm01UPyy/h3I5tjSEAaU4s8eMDC4nLkIqNECrrxPGEMQCE5EXsVn9
9L1LO0XLUtfF/4jr/Wy3acQy7j9v6o/75q3oI0k9CYHd2FHq9GgZbpcY7Z0ZTtix
yzHimLNRBQGgzjH/OlmT0WDJcMXVsLIfq70FLz2ZwmsdJYHAGnPXsfazjtjJOmJ0
/PKVKVyfEGmzEecj/BA5HuczQr9OfNGTh2RFZ+YZYEKZz8dqcReEib/aZb4JzU96
r433IDrMu7agDujAnZXEocKPZRhvg9kwetvdaxEoETjh7NIm64EQfpEXdLE+/hj+
nMKlgjTWwMoUBX+cbhBjbsuYdymY3BZPivJJsT7Q9Ehm4VRU4TaP6Pnr5m+MDqjq
itcp83tySRTatHwnRLW6997CzGsfjGsaTiJaaGDq8tf7Y5qMp+KV8jEzYvf1BhnG
20r/vcFe6T5ykZblzEr5pJ2mwRi5xfQutGtb58D3CGGybheaQjDEJWwHpbsGl9Pu
+LYqHjT9J6DaoAbMFuJHpn9OT/yCq2G13FP1ul6GUS5kvyNn0ZueMSJrsX+RsoNg
vwnsSITiMWjS9rGLW8IE0E/ljugv4rIhPyg405pa2QJXMXDVH+MdH5wh9HY8h0+B
Jb4Zz0Bfs54rjCiOR51w8nA4XwiLEe59hF09jsYBRhdcEYK3DNHm36UnzJSvariz
VDJAMQK/nt4jgP5BiVtUhLgn/w10y8JMQecKy5KVoqk2XIXe4X90MTT2Lw3E7afe
rdJHzpnZ91ax008Uii4sJ1kdsph2nNt/lZvA+6oEK/TZ3pIk8JVuSbPVnbasm5ph
fEo39snjHiioEax2ad5v+FLMvZMzLDjInrUMpmHk+xPZvyNA73anHwe1oZ/7PXdh
RlUgkBnmrFdyElIHCV0Gw8ZAzi6WRvcrjTkzmBOv+03kl0l6H/b4XHXqAlzkEfUJ
cFOyZOUCT5LD0ZOG1/hiXeVJHlhvK2wWQ7S10Nl9nVEjfcimyFKtYJTgzhSZflrD
dUCz2tsv+1k3rvs52MXJoWVnTxEECkdNA1VsxdlupdUMI/2KtNL1yCFaPd3OzMZu
KBVlEarr0cesNmBi3nZE4H0X/4clAN1R2srmH2hteT72eEFL3vfTjwvhgHMgBRQK
lPzM/NrZBsZf+g+I58W2k7gcNYG6o2DD9NoBizBNNiCmrtRiSDVq3vjrXL+Pi2RD
tYyhES19x9TlR0zcrQCFDyTVjZO+c+s8K4Mg8XObbgTU9azJXQEeP7LR6LkkSwnO
C9f6NK8f3pa5ntZbgsN7DdabtnCBHlxzlzLTCsdSHXfrWWI9BaQM/eTxYhHG74Ij
jj4L/P8JJcjhv6pfgkURRq+s0r/LO0YdICY4H++8uYre3L5jPWOhjPS0P1/herDZ
oSqjIGWPtMYnL68B15OVfIULxTaVaCKj04/aP3EnPzsrpNZp9+55NU67URk+loH5
pKJ5E4rIk0wcqWvmg1F+BsVWMijwZ/E/obLAvufaMO4huoCS35zntkijHuDpqcgq
603RPThuDtSF1M5RDYVmhGUhMC/M6SHoe80oIBeYkFbTXUcDh1EsihlJmCKLmuI4
Ke9+nqmd0QCqzbGte78FTLoRv7NW3JW+zHY/1szUcDwsLiSbGSsTQyuH2OmcsXS2
qGg2awp8NwGIqvW5VDKsqG9hqS7DlNL5oO/+SS/z93jwMgnKuEBIRLY+TMl5c5Jg
V7rpXF7J+SMB4uJeBawQqKgt/tcS/DZYv/+oh5K++oWstsQpEQtdgmokr7WiEINl
YhbMN0YasE2GaBsvUfSWmfb9qCLHAwaAjdu/DkLeBoto6thFrodlGd1XgDMuTn+B
XICPimZN1A2aXA+Yrz8l1EzOUSTmU8WemLg2CSo/j5vkqRNj0Ojk5s4Ak3d+e/wp
NYhv4rmSAig1kEO6YpCSGJQ96oMv3SxWOUaL6HqTrXDgxkjV8jej4VsgVn8p6eix
CEmwMjeW47hrsLKdXWqlK0lfIxLWIWqgidS/YQGQPRZKqi548tzrh422XvUhh+ad
lml8BcDeE5CnvOe1cBnJ92L0C/MmSFFPrm6j3goEpDmGhV+k7NVQjYkyFDgRS1GF
2+LmzS4RAoo3afm8bFbYc2i426UY7x+V++o32GuY7r1rDr1i3GWb91nt/VfoSKDY
aOdV/mel5uRnUmMPIkFY83S3SgILDv+b2Psy5AxvYJy8E3/IkmLxw1/qrarafgdj
SBrBEmV9YwLUD2RVUW18XWScLaCjvf1/zL2CBxdiC9teEOI3QRiAjLGM867a3G0T
uB842fp2qDba7HpXZEXPVLFl+tdj6lKxRvB88BbZUsTfDP5OwVwSd9D9bAQZhbfF
hs1oMAD/BVGPWDZNZsgSPZEHJ7vfy/Db30R2CHEOGUaK0fI9d73zA8xy/3aBdrvz
Ay2SKtJlYAFcewwWlXddCjtr+85jMst8EnwB5q8FmOC3lQA3PezKpDQg/5w8LYzh
gJkpVKB4pcE8TOGKUxdl/PdZ8mEkfU6d+XH5ioA0XyxOSirxC7HiwSNI2GXTo/xC
myFeZ5DH2zEx/9ZMwGMvSbxaQ9YWAEueHZABwZnoPHKtI+sIDPrfbMGg0sCgts2Y
PeMmCTnJSnKE9XbQT8rJMmrvhFRDRGlnzTMAWJm7bV0Ig0OdLtB/6FWlrYj4XHGa
PXVwTc8wCdmaR8EMmY30F85Djg1ZW6ZPeE4xhciWvZHyKrBKhzWDcF1YY93sMKYy
dneMJFKO4fSHy2ETrcdkz84lGTnl607cZeyQQ+aGapoTBPSe51LIu3wVRcILH5qF
tkRYqa3IUvLneLlwpjZR5Zv4DRsFXu/l2tk1F5rs9KadF3pphBX+1PFlsjYxDwpu
ge2/7Pl0LIACjj7m5dT31ddjcMl6w0D1qDHab+79mt5xrjUOoyQ5kQhdtkU+yMxf
kC8VPET6wOOy1EIfflfGh0H9DVjbcmhBeGEuzWdiWP/dH1xPmXUuGmC6hUTzffHs
FFaDHr7ehTKwzIvCQu7MUJB0hmwyrfP96ABwGOfH2+9ZAsN8+zyTsCayPUIczUA4
zUDzVrrsT517BifxoQ/FLYrS+vrFtHkf8AfCvHQaaAva/quXBmgQyP7c8NlLbw92
oZEgfljh6nJ5XqF6NugH96GV3bjNA2/ebOy7ErgBOBbebkQ+juP4lbF93dR0nYKo
UJFQoCVmxz7JONmBugILIfmRLtT2wuio4xoFio4OWNivCSKdLKnsV3BoJySzuUae
Cn9MF+Jg1KaTGr0IkXBS8cHqpTMxb5KSOpx/vi7WMlLZd3YBMEBE6S/DLrRMDwdi
pVGBqVE2I6oZX6ivnXGogxRXPtf9+AkH3ylBlnopo5VrFG0EjJ2llxvAj+fc50mh
/8azJY9hZIUHPZXFdjsh86Wb367NyLB0Xv8WRgvN/JTjgCGKVcr37GfeUssdD9Aa
6gfesJzAg/yHgZ4Ow0cvQPfTjQtotJcDODyrbKMLxbkml+N0+9rBaCuLE+Gb5zL5
8OIdg5FrDBuCMBH2BDsvb52bbdpifRwFCR5xb0ArFTykSBRn3qeywngFYfj+/To6
lONiKfdHsbbwz4DtByHQxM9KwzkUE1rD1u9Dy0id35XU5In1Of272g3q2yYXz0pb
azbNhRz1LGA/IqHnDEoohMaVWJuIHoDaSEwhVNLrsKHtc9X68xTnoHJSpGjyzlF3
kKkRuAFQCsNZTjeGG0mKYmbtRCd5JC2iP9sZGHLdRIE0iXx4yXwe71tYLq/h0fz6
xwli+5u7vxJGzTZIA2nzrEzqWBK5wWsI1nRAJBr7oU8Ue5kwocLpXIEF0qyap+ij
7QucahdZMjyq8i2knYyF5swMrhoRwmzTIzSl54jbV5aeIy/1ow/9ihNBPdtUcqAn
/M2UHHF3wiKAvkdeLlgoAu2ATYCgDeuQjbmUAuiA/q8nXqAAWV0aOUttXqSVivfj
Ujr3LOFouTkK6bqkTCE2uKsKwd+mE9n8rNHKymr8+21hOkE9GhZaDT0B1CBvjVGi
n9mcWZknF4Vl9F1D2y8TQ3Bd8xG7VavERNtRyoPGS1BXfpm7qj6QkusdDnprwjIc
YGaE3m6sAdMdvAptmfGfJLnSjuTlEm33Y0SwTcJLS3xugQJ3g8MVyEiTrK4sG+24
TVGS/YaJoPWEoapKGFlg2tX1D9in3sqC+QRsoRwjF2/cwMx7WbIkio1k6itK6dfk
R7RcrWJ8dkyw+3PTPhnxD585aRzroa0XjReWmyXwnUdy8nGaTpajeuT5gh9yUzcE
hCX2aK7reHzmsyW8mbvEQhCpMMR8/4xQcAtkP663M45I1z/b5HzMwWGAOnaMaEAk
m6ht0xr9R0MHOU3f56QSrKE9YIU7w0jFk9BarSNbMIpOF7hByAZ2KQalK1EacvzR
R/iRQBlWoavQdx6a3wwXnPyLiynqw9o7StRm5naGFrvpDZ8cpFZLwy/21xS8P6fC
mVYPjoB8gdiYR1znRzMwp8A54deK+uOPzzKHxrTPEsladtajKgYoGoOXw8UdXc9S
9AiI0jSkIUi3m8oiiNwnF/E86DEk3LWTJwWyEOgM34B9GOYc+YhHeGrhEEQNM8Sw
mXw/UUJU68DN7YeruRrgxyXsgw36/x8vwLGdoJfKimIidPXh8vRaFEa0m6itsalA
uceJ+4SUTVB5K2bKkeKNo7pgqk8hhaeoXObJYNhFBHpoiJ9mCLCUxC1w7IPKLFJo
UMgFEK6UIeAaJTUqQh8HRl338C6/W6AuiJ6IqvblP6oOa2epOiJl0QYsyiL65L7h
jkwCR7d50U7N01g34weZs6+KaviMGc86M5Dlzj5hLVsbYHNIJXiQVVoJrNdYEkoE
vHCjTVI32RcC+uDXYtGHqbC+7KHpZVXlz2P5V3LRZOt+S+bwqyRhsBtPrc8q71Li
lmbl/Mb6l9kPiiTCPITpStN1PCMuqWFpY5YVVFhTV8AEY/oMBPJPsdIFxcRLTmQH
EIiFkIPRsm47SMbCxenW/KR7f5nnly8qcyHpCuvLC3oDQ4lhOxUH7cwMEUoelCRS
oravWUyppmVEDNbUSaKj4fmn9bOXclau98kZMmFwOMYa3nUmbJdM1lmZzlHRtxL/
IA9G01QICU0s9nvQUFKBg84/rh6RN81jYV7OwHMpS7wq4q7dEZAmvKdywYxMEz5E
NFh3CYAL3lc4KEtJID9Rt8MXIJ1JhkDmNYlMweSbsGJdLl5f8iwUn/yJVI0aZB+S
W4A8fV5RIKjvpwMc0iSIgLd63FnwPZ2Og+PZNzG1ufw0hs6OB6FJ/hhDECnJqEAt
JVK3pj2XHa/1qF7tOCEhKKKHfdejlpicMXeFf6eX0Qe+TJJ7r1eJQc3i/y7f+/28
Qv/5lPGgzHYWlywXRf9PckuYHBx0qSjL3NeHDt8Vnm5WuI2vCGcYWNqxyfHOkVD0
zsWvsXhTHNT1V1euYB3zYQYW7x6tVmEu2I3diPLL5Pv4RwArm1jXAZCLkl8TJA2M
0A9hmxpiUIkms0gOKM3456nl+4DRHnrpJN6zP9uDzo7MQgmrxIU6Wia1V31xBIGq
HgsVjryE1KTSUJ+OoeE41EnKeMvoh9FCv2bVqMRnwBaxDtR/4QS5tGxHMZQ5od6N
hJa59R+73Y1jf4jQD2OCbehXDD9MsR24BSJM4SVxDrY8JBU3sw7jyrZnCxuuVc6W
0YEbY6dIyG5eKUd+4VxrZb0vHcg2GWkx1769FJXfKufoS3gUeOqT3HF/lPhJw0ni
Lptz2eyy8OkLzi68bnQ6R6sHEdNH3CaM/6Rw2q4A94aDIUP2w0Q7HSJEdgL88ii3
d4WsWzBQcp+UnDHUJZyC0fccyEe/bvoPq+ABtluX2AyZ3emT2YxqZ8DNcTWuWWmD
B9aL67bW76km3ZC4SQn49kusHEA63rNmIDgMBZoCGO+6FlZJcEV0+cV05kJydKar
Rjbwn4HOC++cDkjfUOBwlQXcVUQneQcbIDhjH2HO9HLdE6pZcNEV+UntTzadGmHd
hC/4BTsgAzhpMdUPahoQTPaIb7MsbJPF6rcsO8x6JdJPQLw7A1tFjJPiJxw9KNPh
1iTKX2f/wbMcD3EUyUYW30NpTDzA1QG+EhjAAqry9WJ9Cs3aOcp0kW0RwRzq+k6o
190BESPomsgCQ1nvI4G1OSCDD7dynHK9VAZVWeVmAf8+eOELViXiYC5NgsrXp5Zv
WtwTM8G2BGBXyIicvbI5lE5wrC9Zsg0vv/PJOiJMmEQaEOxqR3FvUbJgxnMhSAwr
huVc3nl2fJPJM01x5/vovYhe68ln4WH+Dq0vGUQIAMQrTE2R8LkVolHTS9CP+XBh
a7HuhEAVm99zVoC+lVcQj2kjAwPisPmqqidGb8Kg27R1T+ACJ4qCkbcdW7SIq504
2XrgHtIB06qE2YIf+6wTlPGK1Br4cg6AwvpnPAansF7Xayk1k6HjfUEMsmaId9PH
qDr+Ach0vlzjPT9+ZRfmpDmMaUZtJLj/vtenZQc5nLMX4HGFXNxYlD4eeF5QLEZ2
favLMn+gypG2ScC+/SvUkDMR9+K+MG4k2nU4lbC1NRDaP97FmqIpMFUz68Crafme
99WaeYD/DGn4LFQhd/SVIsWeehfLD7uUDHkEZJV+J5l3wL721hPiMscfDx9rxT0z
2A0JtGvHtKLcSR2L97OxL2qhBBy0zeIaNj4vvNuJQpls+TAQLzGBAYY/m+chtLbu
daUvMvgGnFk3ozw/kuUTFXuRvpRYbTmfs5yPzoX6kerLCVf0INsy3npwId6NHrqo
oTSLnX5OQoFxkzn6twQC8evWFJpLGYssaxCtl6AUVGUiNKelLKope8A2iRvOwN3q
1De6a6sccuswyW3RGo289RDS0a5Z7UPlBZjpllWVLoahosBcQXn9B2qtPAmNpEfA
GnnhbgNIQmxujg/qrXJqfDexA8wJwdXxSXiBIOiC5EHkSfhHBjSQj9CiqEvkxK7L
qvY0XwJDe3lgEIHPMMl728DK9FQ4QWdyW/TdzPgEkmx3SEaxjiqyohsbT/mUnrHK
jXnotLbaLvrsZyAoH1Ue4agrtoOUk2WLVNZYp9tu4HTt/9i9UsIOt9Mhhv1FwoZY
/Fh+PcOc0E3NxKZJhA4+qohNqUOZfQzt1RIbtZwhjbAxprAcFRoNDI8sE0HCU8uV
BMiGZdExEgtIvBNwDarGIsrvMRyVHtg/53n/9CUbciL19fKaw18+lgFNX2e7AZ4N
JH8E9d7LklbCOmhwOjTgRCL/iCK2sx2NVnayc7wMiGnoi2MNGHVVUisHsxo9KC6H
Ihhi5c/fDjHq6ZlHn1UJ0EPK5OLYylP0L8CqpaHlZmtmWZTvrA/vg9KPnXSyLNmW
NqHQ3fs1eBw/whniQ6+sPVVpZXovwJaZD4pmIzHLNZpWqWWyHDWLFVdpQiNB0/33
R+GkpC1Jy+arUBv/4+K3tsklIx0L8uWBRZI45ujhkeLv/dBF7C+7cnq24TLTeExi
TtWqde5PacYimp73BVtV0G/YCDSd6/kij2Gw77i8N0bLxXQypbOZCIJ5du16ouee
YfES0yuODhbGG95dPiQ+QMfapySCNaOSZI345Zt7uNI/uV1Df34BdddXYPsIApYJ
nDfkrnZlWmVEKV7mKQNjGsfsuFC1mqUrMNEttjVpXoO1hQepG4FDTzRM0vUza6JA
UpUjWf863cLibac82SpIWGB5ma+n4jI38uflfA9AnI8eyi74lA6kHyg9qCWtsfLz
Ieseis90YVFIWt1unHCWnSjZPZEOd3gmx/byaFdLHUAJqAcYd7c/AA8gpPo2evPD
m9v/xRQ7jKYyk/yzjTSxUkmWiF7aY28hiZTpUKsa07TDxAOw1UkgpTZz03/5sukA
EVV/R8L5AQHI6oyfn5FT/rOemuPOqynBwp9daHNKxclit/2iF9zz8Vx2Bno3W6mn
1sRuxfshGhB9xQNcXZ2A9sU91rYBchXFI+WvWvXQmvFKvaIjH4is6WGjlApANPvm
t2oZeyJKNzIYqvYmMiEFcxSHTLgnD2yqbP9L6yBjNq2E9MQUBj1ssBii0qLg+2P1
ItyzZia0QdmUVUfN3n9MDs4InbmAypYWp84eAlSm7ERex2r/76SCxoIxCuQIVBcz
fr3pYaHWW2E0lxxq/7ZHYxN81t/kUXOpnIlU8RgCKtrrrgVHfuGDZNSHE9KSsB4E
qYmXZmHSBwSWV5Tha4PjLhEkAt88rap6vZjKu3GUW9opXZB6rvucQcCtwiFIQ2Xa
86GB/CvneiNtPHWMDmH493RRr3eo5qxNfy8Mgfqie07ZeTmWEHhOGzgtgjWddGQk
PB0sPzwV+vT6BY1hU1KV2wtPLhHhPvNszn+1lK6ea6BwELC1BB/4z6sjc31ACfi0
zrJBc7UsqNWOVBqPv+kTxGSvuD2jBbxNGZNIBsxiKJK0OvzaFfaTP8TXrEZy1srq
r6pzrn6yYrpQ3QuzaqmL4JMu4T1ZDfrHXzk5HEwewFIJaMszq07EdxKPutoJP2LQ
2tJOL+/+xkCr9TYuK+dA5iwEQix42BJ1TNEb7w8HyHkcE4//gmuge8eN+pw+Fs0o
ntuW1/pYq85/jWlEdQ+z3dW8fFUrlxl44yvpLo8A8jA3LQgUJWSVaxnoD2Nwfkvg
wKDd1Z5WcD6rwves1QD/fWnjt7B8aLm5J4XaH4gnnbfXuSzQ63X6DFPHlkdBQ22I
WHevWf+fQ/bA6ULwP+CZZRfN1+LvvzCfpy7XipypuKUxslNsT5Y/t5c4idqJe/Ue
I4XK0VRKbFLsx9PxVg4JchnbEkCUOQ5o+syawfZ1F1k8pUMi8yEjlznr2eOUvOR2
EXah4ZMiXIXCTN3vrI/AGBJZXhFYztJJGwH/eJzgwhSkvbZBnc8inmqG/i/8S3nT
cpO7jyJriFFDPLFUFkFS1H/6I3S5D5xXBFS2RIiDgjc9cKZqqABqI1PEkY1949ig
FhzH0KxUlVow6JR5wNRR5nMqzvxckuGn2HL0TvCE8XP8pvSy7j/mxfMo99orhUpU
ZHQD9JpUADwUVUjDg3IuYkBBkyOIELPWSDsIgqSdZjQGas+XP6bP36jIY5yTL9Cb
9qFQBAVQAI8Mh9KiyJsQlfXcu1zGCdzKslbJdn2Rqkiwt4/YNRc9TuZxnPhsbk/s
Yv4KCXRrZZURMjonyAA6XtNlRkJYrDbCtzX56ZuBCJbp6YwjiG6AMcnmzX21SuQF
WQ5TUikUWK3y3MNyN4JxQ6yS9ecExneYsLbjrCGnofz4vMrGn5v5OkfSIaFRNQZm
4l9y44tCl1L21YkmakUFBUMUBvmW3mH0wY1go119KijPB/DJVvN7aQXjzNSIBXCx
FMh2hBEyYzJ+EGeep9HA+10KF6jjkUN2mSnIh/aTgN+szW68O3szrd/dHiD4pwqo
LRXZzAmUz3pgQriaqO/ljgaT7nxD20F7ScUBxoJ8MQgkL6/C8AnoPP7MDUrS+nkR
E26EwMPMq/OTGxDAx+sImC1Ox5he2Xos6TjFVlMQ5M1PTlH8+aSZj5IFTpIqo3A5
pa5W5ymSBv5YT/WmogIO1OKzQ/dD3FhUsDvIfjSJeKjFV1fYShsjVYHB7fhIWkub
2mm+ElLWf/t54LGZ7df/wOx+kFMF+rLLp1QonpBaPr7CyePtW6PV0RowJ1PYFASG
NvRTmna4wFNUzIT7ruG5WHhsY0RKhhHXE+Lk8ouVszL6AvijrjOZ5Z9NjJ2GHo1a
EGz0ZmueyhE6EiINTEEnYkUDw0QQDjjWyyJXzTq+Bgua0GEA5GQLBGD9HJTzhQcL
y2ufeVL8oZdLmItAGilxdV+e3lulq4RZGrX5FOtxWdi+liP0lEgTH/aCgJXjjfo8
8VRtjZCUyUglZaKCPUyszbMPt9Whqfn4EP2SLcWK6HpMmjjv+88sB9dciaInX31l
0lmqROlTqyKAqd6wT7Ur4wH7Fh570fv7VYkHUP15a+1/5I7YjS+bT/r0HPuGUZmJ
icK6SpHMRGzAL7t9ge+znGDBW0J0xgv3P759j4pqq8+wV6gltBB/3KnJx3pUovJn
B4XYu51MdrELDqZh16SOGmiP9iTtUBsErSL3ePpehmNEvLNFqlwx1YwrlzE9WsAU
TX6pmZp7gSfDEskagY13yIMIL4c8PpIw6JiP1D9HGTsQJFDGa35FORJtnksj5OEP
14cpFxIQc+AThZurGbB+akPuHgJAoj6s4t6VJ2WbgAqtyz/bubvSfuAf4aAmKfxM
WRozpu2/DYnP2IOwbf+CEIEawOpVpJtoh1Onki5yPSaDAlrhpOaeJzoidW492JES
8Cj0ancnp/smSoopxfhzeDSjztD7ypG3Vrn7EiM8iKYFB2OPmkFXZb/XQ/j6KJGI
JHUq6bzxSPVtDhKxwo81ByH0rYW1vKIs+0CJPDw9DCEvExkmwY0HvZYq5qsNbES3
BluHKqVZdGjPwuNRnKOrXy1UXKzEckjHQHqbPHFUmfXSsskb1j5HuP+hPYYMi/Z3
YtaKIfcc016bXelJuU7ZLOOiDTsOBGX9qo6ScvrTDTf6ILm0CJ6MCIr75neElmJu
VPRWwe8Oi0rMIvKccPWNvJgu9+KnyoXqiU6JTOsTDFCUNG25dePeTYOmTwGwZ0Gx
wwRkgeT/6CUP3VOt3JvNN9af6HkNGEuzbd6JLo9JlG3Hb+DopdAy8r66UozZpsHH
DnE89RJ9QOd5wTf6psjzOTgEkzhGtSmGskzvvEbVqqCAf2EdjpjjxWobGJvHhQUb
BYpfj0sb6iImkc/uM6X3Ce++qItTFmnxLhbYUjAnmOS3rIIz9IfysFimAlnTR2Xp
aMe7DLyLhCZoEwJc8uFyj1ziFvcdUHW0dqyHGoVtSnkv0VLWKX8iV14rhBBCa+WF
XqZWYefxkikqltkN31QG+kfMeqvoQZXSZ8RK3WeXUN1Kfynq2hVbWOqLup+KgWIk
wbwHwI98q9iT2wutnLP1FMWkiLiIlr0MQvvQW1XkSP3ujBOUKZ3PINHoXbINvfxU
cYoinQ1//PwfNU69D2yyW0s6JixmCX4k/ABZJOjgU740jMieomrFTubaGKvUchzA
OVrE6Yn8NJx6+N1xPZsqtXBRncdLiWO2qHilwUQzvnhYvqZjnECmuQbnKAxhaY5R
crjrtVRFiNsIEKHJ1Ve45zI1CFakTu8ORPvFofXUw+ACw68jJpdSNsHeEgXUKUOA
6nujqF7t2MUk4WlopjZoOMSL1/BTvpW0TZgdf+4CirUoFTkkt+Qtki44YKtqAjNt
MFyrTF9U/rMB7YF0Ny3xd1x06g2kXYsE5YTgNm8+GSU7bLeWTggAH6I21Qa1fCri
t5SCAuFXvLzkVC+T531XP0l4lTWWkK8+W5R1XxuFNtX8M90zOB0v7BVF36fZsI8e
ywoO2IzRGWas1xqgEoX95juCenmS2lhz28t5UbEbVGdaLcZR/SOkCgTcT18jvzK+
ioYFBehuTOZw9kJCv0tRz++QY8T2L36AlYgYxLLI/5bMm532o+NCL5aIBYBcgyGg
F9dVQpS4/7AyiHz8rXDIgC7NhjRxfU4MTeFBKSzqNN2tVUHjEc84sHr+GLtVzR1v
GSfS3ANK7dFhj2YA9FtpIqrpvm+MTJosvSu4hLVLEEnweQnqaB0KUV+fYcJU0Acq
Ir8Yeg0zgnCjbp/7KcdTBdFpguQHExKzUDMso2JzMhoF7bJ3vqmZBAqX3yBK1A/Z
+M96JbHEWOFOISBgpWwCpG3lKDnYnSgvC0+V3dICYyYZf0bX+RKHx9VkpXRufMh3
RCXo/MHZinEhUMnfGQK2QwjB0tqHiBPfJR+ZIysRO5oRJehy0U+chJV5C9QLBYm8
AMw3U2r2NtENii6qzuW9GQFNUpO5QwTonPilSfwstVc3n9ZK/6zX1C4goQpfu1oV
pBqVSqhJ5e0zImpuIZDHBKnmMybDnmTHiU1DqufUxMVcFZXGQk3dzVTPNnjeQbl6
l0VueW3y8A9jH67vMebx4HiekGo4IZKdICfkr1PeTnoeipInb2UzV2d+vFdyrPUC
FKfrMYm4UbCKuIpaIDaWX3/WvUwk9CVv8vUeCi0jm7nS5ghCpgkfb4tR5Qpk9A/r
3TQfNXD2D1TekSlTpMLtG3gIHNkW1t9OQb5LV1tQi9HqCWmxYpoFTTUJQt11JYVg
cOJgKsFcMztY5uVl+gtnsOX0+lpq1ZI8N6veE0qyUM/fDkbqqB1ArDzbcBtgyEWf
LYA4F3jj60QkUyWE+U7V0JADNFWxyq4Q3J27VBM1HbuENeMwGgSHsdGDNBw6WuZT
Qx6jZq4NxfVnv+K3LSUXkCBfOUE26los8SAdYK2GVWF89RIHHB6z7Dt6C65C/uSG
UZXQatoc6lACIeJEpxPGtJNEZnGB0ttMlPKHHQLl4TqIKoYWE515HR4fQOfXKWCM
zcii2Ihy92v1KvuXMfDhwvHeFiTvAfwGpdn2BeNpqkcPtfCGKS8gPpup0wcspmh7
cjqo64vhZTO81RCuULnNcM+SJ6AzbEzUQWef4X8njh4MEtZcRTUwd8YAIc19qqHD
vw3Bd49XaJrhc7Gj1I7Tr41Q4m8iDBJo6sSoELKy6mQJekn1TsSOiyclaTi2VNun
kzNCFXvou4WuAkT9+XAqJUIWed+eWKcwhpMBAwoHffk7S1o1tH0GJLMAKJF9rEqy
31s8anmq1OVo9+39IhWUhhANvltQ4tpX65cDQpGIQ4bXBqxYPhY+dgHVAPZhAefU
PxwmOFHL60tFznJt0MhQastkcH03T68VomxFe3EM5MsLoCgJjUYwy4vtg3IYEGRm
TPehlQ5LkrEZvlrmD2HFPjWsX/oQeK89hb7jtkbEXsQU8Ne0qWWFzWO2mPxBB7zR
zf12sXx2OU3g9czWf4HHbq9N78fEJJ7QTG7XKJ5zxKeslJ4NXEzk9b+ZFvRGZSna
XdVP6jNYoJVuhnTsX2FP/AG/W95f13ZnxtX7S8K5FeXi2+5Q76GCKwJBBGuSfY4C
Cntm32dHiK1aJF480COV2aVMtrHAP1iSwEdja5s2AufmaJ9hyMaEV56DPUEIEnXv
8NivSWsmd30hk++nGZd22iYMVZ9PRn/1ZJsM2DUVQWLQximPMi9FT63CC/OjJ65O
pSEwVdnq0OkFHd566EwJmP2qim6keH1bv0GdyQKDKF5oWGrhg6hof79L4PhISFk5
noTitXa3IrYPfH7+21jwuSGvwbHCFN0LJa6lFLe4F4SWN81b3SeqEZf8We6ahnfi
yKOMTZUilENY/9xMygW/R5KYInQ34aGkOcjN3S9vgXQOkM7CPT406f41NWnEVFRT
CA2R3JvScECMD9EyzlYZ1XjAlaOlZZymYUYok3XJceWXBnYmTpHytUAjx4T1ycGA
Vk4pTQ7k2xJgiJTppCr9MFdfELDvro52d6aV8cmh4M07CzAKMSt9TX+lFR5cKZE9
HdiNiKI3m6dwXfJ77ehsRGicWOQYaOEotjlR7ReQUt8MOxhw6rQ+IoZIGqX31K0a
kXhfgLzGoxfqMrxUyP9xMVofeZL4MDDS1zVkizGf/aTvaVYU36KfsXbgosXm6ma7
GZ/UCBVz00s4YeIwOZZg4FyQlxgQ0NnVp/dEnfkbmYdA+dtmWTLPAlOyqy8Eoqq2
24NzgyMsEhZDw4iZRcyVmE+B5MdpJtcA12wKkeYFVe5rhq7nGp3u//tAPukcWm0p
LbR2akFMm1/VrBYYF0Y9TL55B08QlGoeIywEIwgYsU/LDwFDTfUpuAgl6hyiPUXT
v1RGMIBF1MTUS7ZYMsbo80I/4mx8kBaOwTqCPydaI7n43D9lHjpQPJIriPkRr+Mq
PQ7lX7YjJ3YU5iIpgcNIzR+ysDqoMyo+2d78Lb+P0iqB8nphjU6u+Wm/T8j1t1ul
iIUyJ9APb7KzDsFe/T+iqzYDvOZSXpBWkTQOf+f944rCXW3JzDFRhv4PJiqOya9K
GkQg9/ukuZCrjNUgwklh25iqUkeKHZlmVaCMm0RsvWmQpwhUJ/8R1MZuitukhAxE
rpCiNjL7+oqoCll+npnsKhQj45wXdvmO4F3jRxnptGE4JeFcoxwER1N9TfF2+cKG
4oy5mwLVAo0pXOL+ZsN+QOLxS0zGd/YrXkGI0X7r3w4GBk1KaKBKT6H7nVGm9ksu
d0t4R76GXoLzll3n1WyMjpJZp0PN6clQRACteHhUUfqlos2wSol4E2Kncb8VJ/Pf
MVDy0QM60aAQBUOmvQfVAEWAtl87vHWPfoaGWfnvHsQ846B80k3SFekrCalM6J5b
2J5+gpG1I6goZPNX2hB1yIrNzVBOoQ3ToI5OwkkhxAI0cWW/dUIcGLVIy2xJmEEh
pLZI2fjh6K1+I1n9wxKBOzBhawqKvOoEhEEhjoF7/U56KiZhKAGJk43nBDgkf7Ew
FSid9AiUKxe2FzKGKDRyk0P1Zt3i2O0rH8v2/X8GLJnIAJzrNn5flXbBSUnKOiV4
Z45gWX/QWUjZW1b7N4OYIWijyuTNiGzZG4WJUKcdXAMCl3sefJMb0QxEXEeoEEQ0
m6t48ckkc2kFP8XciSY3aRgtAxyh40q6zw4wPG0ghv0uNolgWVbDeAtW24bhNE8W
gegUFCRB6WkbuxrPBssl1q7h6jbmliw5zOU6Gu2uFOFAoND8Em3fWisBfUW0gdLh
MN0QHwdA3dfUq/gI/9p853xlap+ySUUVH2SUsXFFavTzferBmksaALQORshY7Jaq
Lkv8NEA8DYtEMKSr50hOO3IjUrxDH8wrZt0asIe+CjMMEkUE2rFVi5yGdeFao4Go
GlqaRcs6edL0cirk25MbIhcfjoncsatuZYxBMg5IGEg6JyD/iSynm0oV4Al/XrdU
5BN4mRN0ypyghEz0xdTxR+WED907arkpY/xVgFJoHEYX57xf2/amrpH2K6/urYh7
Jh/wNOI+Pge/9BzANZ2CouDvloDNowjxuR0qq7zerjgwpNQI3dcuThRKgsMmoCo4
DRYgTf6uWvO3LoUWC5aF1HH3RJs8nmT1osvn85LKkv+mkeD9m/azcz976Oa1zqJO
gDbysW7dBtJ2VUENeGFSF0p2eNlmw2wq7epL9rAMWv2jEnh6CYkbInuCWxjVWwm7
3BTwqHkFGqlhbgccRQuSBnRADnuCDtovOqTwiPg+hzT15UNP3DX2X213ikvKia81
VGaoVnFLaGHD1C3PbnsiSLqWb/gDgdx7RERzT5q1rgOefFFWVV+lm6WejQxb4Gvp
/rZI2XvYvGj0RTCCHhV4ee/mFlF0lOy4zAI2NpOA+6t5CPouTq155y76yCOldWDu
LTWnSWHLE0lRKG8uvHKiKUAED3/e6pe9nnJi4tuOLD/gRmmHKinDEiLe2YMgaUZ/
PJki+DkiIYWimEAlsCORBX539Okaz6YcYqI9PHJ+W5WKi8BCfkDT8XuE+yDp8eCc
QAWOa3RCvR37M2Wz0R7A4Q346JdmW9v5SRgD1TP+1X9QDdx0nIz+1EMX7hLCrBXw
lvJUoIAfsxjqWPW87cbSqG2aFyBT6Ab81EWF4UpxAXpY5xa6Yzkk5KrQ35QuFmKc
oNMsGgJpAkvmBe0Y9p9wJPQdGIvrO178ubNGbyaYgTD8eqNMBMZtfHlqVdozq6or
gLNS8a4G6FtaTQflVR9CKxjFXEJd/NRzzjqP5oiDx8JC4y1qfrcTr3lZyL09GNJ0
/Ma8YdqW9KBCoydiK9F4J+qCB9iLguoXZZeLEPIdNS89n/ZM/Q0oZA9qIEqya/9w
eAoUCO6KcE7CAQ8rZMOMNHksYzkGmd2OXwK8786odZV/2AoQpoG2jaaaZsPujw80
U0LdPzei1U5E74zRB4V6QMvpp5jBT42oo/+wBssJKnL2LpEavzVsl8RC+w0E/9In
q3UnveuYzrXcoYK+prrZ/heoGPhLxnygL2vM3JzunMpU69fbp/Thyumqt3yp4xu8
SV5PQyAJKzGyw5+6CbN5pLjCdALIpuP0IL3hhKMMC2EiQlJeCTBV30TP+7S7Atr9
R1jc3qkxgbe2q//Qt1n2cPqiq7KJqs8O2Kr4E4Ja4XknTp+P1yF4+plrWzFB176l
K8tLEeO46w+xyFs5neeNfL9ZGrIuJgMIQH1/h+lUJAntSW1zqZczJW8Hev2Vksy0
/cv1QUN5Y/JavWvZ5r7O8Ip9GqK8qsa2iBvQ0JolsDj8Dtupae29jUM8xoRBaBeZ
ad7UB+vxD3P7q1v8fA702RvzlTB6jnJJcVSRRmo62cBrgJLJ9O+6N0mvZox3bK9/
AulJa19fjMX0GErRLQeDlWqq8izCYlQiEwl4bzGTpz7aqxXUGwOvPBcF1LrrrTFz
+UyNmQbCpsG1ucasog8492cdzU5O73Ca8HCNYGZuB3/q0WZogVK1uCH9K1uvVgCM
j3zV9cXTEBjEEKmRVCQmdytxyd4DCAkm16mjiGmyVdQtMIx7HyqJs1iR+4irLXSF
eKdl4KiXHrhGagg2h4HYRHfJeEwptabpRmbX0TGST+mOzS7PUz1ww17gtn6aKSxE
EvYy5WGOSOmzhLPdMFckCdS8PJsj5JIGjlYfWxZyTr3A0bPyrOIoWeyDGENZpDWV
ZObW/zCbxfALxDnIBq3dwcu3O47S+hG7pq5VcDo4NmVNVRvXz/a78qke5/zm0kdO
Evi10iMnOU2BZfK3oIxxLw+TKeTMMpVJXCpYyt3FxgIGU6aAY3pofbt1c+N81W6H
KqZ6yLuAm/Imxj/h/YWjiZy3Oy4i1QQsvysHmXOQ6JleHvSmIYU5kYKbhf6anz0j
5f+l07sV4dmXqf0e6S0+URR/UTmVUApxLE1xWuG7E1Bg3HAw6uf/EGUZ5hSi66ub
knbVYEjd6OeGasOixqsuR81dLQ/G443vIGgyY0q5VHhk2SOPpBQAVmILRrGExj5K
dAFCFDgIUW3hT04OGDZiFKzqa8RMfawfvuhUoPShlwyuqRZk6pGNv+TPeuEMGxCE
kS/kEsfSXzbtjXF5lbuRIBJRimTtDYMozM7Wuw/4OOUG2EYPXjmA/c1V/aJkrG3y
oSyoMJZnEfNdQKtV3ND2pMeZMQdNQLzfJj2v3uP+0sqsolky6Cuj7jOyn90TtFB0
sRKD116AYkmkO8H+m4Uj5Z+Qnyiph1kiZDTQA3ZEhl3do1Gxlz/sIM7JrxbwGNFm
HeKyzKM7b8dkRxKXCGUjLZrQBiAQOa8f+nM6hMLSeK7JoZp7NPjifX5lprY/PmOx
kVjExKT6u3UY9HWoa8lxlywynvfYlXWIEQQmikVlzkzdi+o5sXKBGJP0jB6H02AY
hfYwMrtMO86NoZMWdEYewvWScXReW+WGBdoOvr5WEPDFEGwXHD4tDzMVoBQdEABl
mkm+wGSJw0vRwdTYM8hPBe/6ya2AoalkSiS/x7F+tyFD1JuTAx6kn9HIqrPmJVYt
BKjjPqUQzEm9tnqZhf52OAP5TpW40HB3O+5cXdgiexDpFgdgcG18hdMVPK3lfWRi
jlDNm02yqTFgIre+H+tVCrBl28d4U8Tw6V6yZbQCfJ76HpAX4AYxgj59xMXaSdoN
iIspVSmcJTXMzoHh4E4StRQFkInJHXTmPAiwK81prwpvVxbdS9puFH8mEANrw+39
Yr1XQmGjQUNLj5ei2fF4O2/sAkhc0RBQxUe+E4gKyMyoUCOQ5ZU/fF04wruLpoWv
LmzsMm5InYsMR+iCd1ZQu/HjpDZdrKb2W2JfYcuNHt9pANWm20zd7T8cmcH45m4o
saheJr/KHHvOC5a+frdiDSOqG2oxzGr5CZfp5ckvBeugKKj1g+5kij68WLIqypaW
pgKI2knp+zyr5wFqIi7EVSw2XWuCwC6g3nrdgA81z3tCAwD8f7bak5AkDh0/+Q35
m9dXUEZe/m7fM8xTQ9cXlBpLS/iGo54LYCXglRUHRNqvjStnPZpc+dHTla7QwV7f
dumKil1OU0y9WkLY1C8onncAAp/Or++ikusBGtz+rCfpvHTOAr4dGMLbyrP7dIrZ
6l0HjVt1KNXBU9XhKlMc77uywnw1c0sBPxica1I4Y48BYF5ZCipXcxK4CIJW3VlC
g/VLrqSWMuZdWWAzqA6bO7/FzYrZBZlwl5du8Etkt6fTMjPq5twiR67Yihd/trHd
LdaUcBVQsG/Nhj07KIFDwHC3VsPh2tGscdXxU0r+MGPsFucL8q9KXfvqK/UXQ6Tx
fgJPyNeMcVQXP9k0QTU8AKNP6flJ0pLrbONxrxmWdiAkIdXmVrWIljff/OwBsXzV
QqEP8ZWyfZCBMGX8AvIgQaIVOLXkOI2Tt16b6TSF7A9t0CnR6hCZYHdUCxK9hA3R
bS8VXp4cAeFNUom8Sa1lTEfqqqCH9HQd3r9EANPP5BJO+2/lOAAEfJWBDKP1wLkg
zKgghxXGLeVDWK2sLx0UU4MtFHBt2oP6gtNx0Vb/y1uWqL44ieUcH9IhnqvQqtdJ
HjRm7KEwgoYAnwW/LJvGAyhSfM4y7wsnx16fZYpjnu5DbWloTOu7ZjuTvl//zaot
COkHS4BKDougyVl8uzvkA2la+EXFE1xMK2d7CpoXClqM8i13BaRZ9VEmBP9qV4Oo
lML0mJsN6+D3lJggc55GkbFHJwAqYwsCvj/7B9M9aX9XU4B4zS64cRAu5BTOqU/5
TBIEfp3yNVeFro2QPGuxLaywQgmcoKjpvodPFgPUx3WX71skcDdHqycfvJs6lnVC
iKO8phBMCQkqXPL3bm9ekSFH8QctwtcJSDKMFm0vgdmWx0yRrVDYpYJYur4e4ycN
hGX8CGlH0wRwu0MZPE/vdMhcQo3OzFc1pp3Dml8V+CdkWtcf75/57XHOmu5xdn90
A+Rg7Rx+2QyoPfeVQKvsizoRmUECYAzjzIhUfPR9dQyRuuxfqW0/JKd4TV43KL91
2om+ZnwKIRXlpm7Evv6pkcdlsK6l1y+8Bzyl3zgtht7gNXLZVEMbTqJx++A/S+9C
UEokZKPhCSyX7R0B5WmD1w6e56K7UYc9WlR5JxPfCc3vj+kB5F7iLcbi9nHsXL+5
Q5R711aQUcnGCfRbVxLiVfhs9qKMpnN1GV8L4iYyK+EwbjXW3I7X0S/z0vBL8mrC
4ZOWGGThnL5YqxnJtFW9+jM0nM8npqa78l8RYX7f1AQ1ePPgfXXf7x1uZZOHvpp4
1yDigJyUH7wEIula0rZl3OxjIU47EPzVuZFINaYptyFoHe5ejhLkaMEzaWqrZxjL
KPQSv1jlwnVLBi5wJkzS1thBb/xtTJkRxwb59XbB42GMqje7+ujr/ZSo+7QAmnLg
YlUvTHJYV0nxxRG1wiIpvnkq/aQPARtJTZalvvWzRlRgfvomLHho++T9waSslkER
ObRqf4YfYFKJoTYGxLWcn3cXlhRQrQ+Alf3odveOmy/gd6evnpW9kT+Pe5Jmuf7W
ZTBKN1b2w1yda6cqnREf0oBM8sEnW3LEDzihmjBjj8P35UpHhzVVjWxondZLfpHr
8JwhqfUXVTBi07quadTzDdoB+rebxZja9fuN0r9ADSM8boJ6Q+mimNbAnqh59SZW
zICvhuvONMZqevVqacJRe/D8Pr/c5jQe2IXfnd3fabwbYLH8i6ili0oji9NnZinr
jEXM+RX60p1oIpyvFVvNivdTuW5Ifa/NGtlNpGWV8XMOVkxwK/lJfWRNMPnHZdLO
j+BEU8NgqMnMJTFt8DGvhN5rxVlpPPuC56rfJUTW8VeJ2TRPAlPBIedcduOCvCVz
FMAiNErOrIRAGwU9pZ226wLy4nNsej832ugt4vH2nOoni5L0Tq/25/cQ+DqaF9x1
48ANR97UBwUA5E5StElReojYrvmQKHWKSvAFQsjqQNEjU5pcX7idT19AvTeZCQWv
7+0KEYpPi4aSUY7QqTe7z8xSFPamOoiS9IGJNyu4kM8Vv040prVpAgzxbdfgnHTQ
JTQvVn9Jum7wIH8F5Xi0BAb+MpO5yDVJuan8FaUcDqlU3I8H9K2BqwLOBAjp/rtp
IebzgF9GNBFc1jkKQkdEni610wmtuxrZwilC/f0CkgzisTMm2fpm15ZvW41tZN6K
jZQSUA8tWhgI24hh25j9mE2KKtwQpXMohSz+3rr6cRustit0b9rEwIdkXCRQqi9Q
27z0iTg04adGe3Ss79x2yQ+uTPwJWd2MwLp5D5yVtpfXQ8t+KE3RT7yGFn1TnY/q
gnRmYgeEQ81aP66N3lpw4gv7UuUMINBO5ccAwBqcATnccLKNFaXAoYH75bRiWudl
7vSxiimwbSNVCFZB8adbdPstlCXSdFj+fljMitebNvWe2hp67LqLTQRbhiOUWBww
sAgeB5356ZFciczZUPPHdUptOCd0+Q3KI0WDqA1UqFwRuE22D+I9Ro9v57Ptau99
ZfvmArrPJvZ5W8j57pOS+9tdMVmQbNXouVK0hzLt4CBq4NsMDcIr5cFqkjxt5uYO
7UKIwJViyoPTBtphRdY8TpeczpTouHXcKH7V9k6lVs1LQV+kQjYyhwn8vN4XeQ3J
m7j0cTE3njgHAz7JpwtrXkiveSZMdp0omkB11ifWm1+UQwYCUtKxWha5uj7AyPhm
17qRuqnskJv86abzQoPXbTfXak+VdgMfRaT7hLxhAJfQ5HyVkUmAHwwBoYwmV+N9
IHqBzrCnIckaaE2jwfzZz77qkWd7X6UtauAQLnuN7/RwLD0KPjWw3qExqtf5o+cz
N1Te0tTEioYHJ7WuGbrOCO/kSWXFj/o73aDP9F3E0FVQZ8pfIB/38lI1g+M+tKqd
r0iar2CemqmyH3SVGWc6IKJpNvehq//92yEBTfnFLmu7xy3w91sLrR1NuGXpJFQ4
yYc/m2jKR/2/sssCeGfCafW9Uw1whDknRuGpKNvXLBvGplG6NyEGWIWVtB1RgM1J
k5iXr+LQiv/OOZb4jd5nbcTfOcniY4FMvjM0LtOX/7kEQLrXxnA1wxOe84N5YE4O
uiiEdcIizORnghIoY2EFZA30Th4eedaQzN+NhEJ01ki7ID1wJbUnjIF8a/AfnAfo
EGBWKR01CJb0PB+ok0ipcFwqZUBm7QavCR0Df90xIiD3JUu1VEjkQ+yQbA2B7qsC
gTQKrsM8X22pWAKW8is6Tp1qnJV4x2aXQVeY2hWpD7PDSafQxin1llSjtJxVLHA0
nwjPJtFJXWL6Q+kbsI7gdumkwCx+EY6g/eNtrBA57BdRobX17pa8k+FHUyyW4Iws
Mjn3i5hmaNz/Hwz9TGh1dB0HebzFYTaTF+fYSQB61R0e4UQEtMbjtnuF2rV/zGbd
W2YqEM4h92OoNi9fJY2WoG7ScGPtOdnuOVH8z7jyDk+er0aavPu+vjmI67hROg4M
K0W83QJ6qRgLTsZmApyCdbLMLoz2rRp3jdnVnvoyaoAHVK9NVwe9gf8XbM1gdx89
ykJr3LRJbJGWPjphcAX93ToHUU/cocIdoRWb9AZpWWbpY7iXPa0u/hzM3XRdyke6
q5oDy74brTdr4JfC8ggq0IFQ/VptDh5D/FRR43TRs0R8grsoY/SqzekzrVwy0t8c
Zl3Z50O1fVzvStB3TkazZJunEzXvq6S1g5RdmTC2kJurqzPTFjcijmh9dQwzhuDJ
Uaoxu0A1FY5/B9Mi4v6dsMM1Q2eoCVaL/blWfubgRYeersro51QztvbMKaNqAX9i
M2t+drKIVnqBDae0K66TNIj/dKelNs/RvgKaOxOjfkXOQvkS+hXNmNqAutIInrOY
WWXhxXjcgw1W5nTGUNwOLK8fuZdc+mI6RHDveprPMJhEQqpEy8QfcziACf8akT/J
O1yvP9J/WKcBIlMlxNfBW2cV9zJ5eMt7EhdeMG3EDSyBXxcPxH9E5LiOlYaXkSbx
7W3KnA0xS3/7JYA8W0pxHf+xGZv/hoDjM+9NNj9Ag2TyjJ0vo5/jeKP0Rf7VN35d
MONnIBpfp+5HCmUYPKjlYxf6h9pQLYyX0bI+zLhB4VNKJKPrrleJ9Qh0ymYZv6IP
46ulcBFkaUSX055dh0rSoYr9RIQNrBhVw0hjOfOhI8ggl8UEzl90ZPBXCBlyu2lC
4xQBYhjAlNd2SEmC/P0Qa9IXH5ds0QmxNHq1WsVcS3gKhgfPH3bRi6giJv8PepCI
YB9eNWz6SRKOQXBzBEiXxi+ExmnMaLnlzsqkvKS7lLO5352Lfc4Nad5qVJd8aqZM
uEQg6VKA5FouUtgk5Ybpmz9O9Ln6cx5VFOQ4KDvFS+v/R8cSwZe5uab6O0flyLNl
uB9gG6yDbmfOEEVzXtXhYgf1NTxHp8OyZJ8irsMTvlqaXVYbLBGYCFCVil1QoVwl
ULbZtjIRFp/f7Fx2HG8twnvwEIy7VQ3gANG7P9tuVMl6ALB8vfVLhAcbjQShXHL9
/LxBp1ObVslfZyUei3egL17hHYuE6MGcRqKCeqUwl/yRrjogxFS1UaP8HK6HOMBd
PJhfkkP1KrUWHia0ywwx/+Cclqbhh5GefkDMbHjnyFjZSlnc2xmkipgb0cyhyHMs
jzTSPhyzs/I6uwZ0ansK0upVWjt4lHIqjRRFQ6R3cpzaiYALV+PyXQZdeatxguTz
+uBsUj+/BPxkde0xP17xg3M6VyOuIDI+5NSFeaB/sH78gJ5aFggCpPUWCrarq8Gu
QPzXfpg7RCGVO1LAKaz428crZMYq0r8WrEctc8Gj7jDcgrFY3/GgNqTWyanxSCI7
Zd7b5DJx2Y1kKRIwFkaJTYRr+onrohAcSjfwg72FAv1UHq6kvNHluxE18s6LhDTx
k2VD+AKvEMDxfqnZ+EZ33kVEWCsxWRBwC0YJzxglFQhKRuJYpcMVwsW7k2m01l/r
q7mx5n299RGGBbL5FqcPMf2c//Lu0GGEmrQZQxlbVyqQYAeb9e77k1iGbg8UGICs
xA7O7dwemUj4LdRJgeeiYqL+B6BaNekZ+xJozAbaJrEog08QStvtc6R3x9TbgU6k
EVdSGWO1hD2oNYIumSHBDRLuNIexMUXhnXPkV7eDjbc8OEdQ1+bz013T9GjZdXSh
Ukh9y70cEru6QkZxBK3SLK7/yW8s/9Ty45lBbXqbbDLPVRN8G39MpGAr3CuIR2Ic
OKixD+mh+WoihobIu1xypRBeIwsSR4L7gUp00e5EYzKVfgWlXG3pKp8125C2lVex
Kx0tX3GMhzuz1LC7HVvHEeTp4QY01XPEeA4Td5ieUWs3yzQRyu8q5IpmkOVEvL4p
MS9HD7GVv4s9QJgzz4x3Lwro4OpmEN5xmfyMrx2HluthQoKJLOM5iSPx9s/bTzD4
2C92654eEyhC6Rkr8HKzTqFqHQvtNndV18sHylwGbjZxVWWfUU5/odTFTpIDCVlK
OhhCdCEEbmhmzmwW8AgHEiK+HYexfWT2QbMCyXEM4etXksijVPhsgS9CXs+BTMIo
7RJheOWpVHde8Cv8EsnH8IB9/bO9FkaGMTJO5mNGtVkr0pC6ML+nQoqLR4rJddeB
IvA5/bRT2SWfgUHeM9kbCKua5uLK3v03a9X+j75sCywVavaL00NihyFkXMZRCunT
+gKpZcdJXh0TblZCCr9R5ov36mBUfvDB45lelEovtpEhX7sEhUdnM/BKYbS3su+5
O3qg3vh6RAyvfQX1MB95JI4jmXjSU1+B2MXS8tWm202IVJmUN25Bj8EcfKjHPkGK
sb8kP/nnQfBs2hF4UP8LjeFpoCVRaz0x/Nyua1tNO6qkHav0mv03nOvlKdjREcFT
lkyazYeHsZYI1Upj2Wy+8Cd1P/8NzIockmujPcby6fs3nGksou18My38t486OwXE
gcbz0GvmQUgui3A/aL2kZXymoKYw/23ScYHQAla0szRe8xQD5a3xmqHlh6xr9Sl4
iOsqPk37N6NpohTfwOiE6rbLTGxCjQ3so8iVCBbWmRomX11J8iL3KLbCcjHFvZ49
wXpUWlTkVfEB8txaMhC5mabpJgZFDDB4BKHdurG/cLV4it3HZWxzM7xvz6aBj7m9
sqkkbvGhUXroPCjvoDQcGdDhd5xu0Wp/dglc99jwbYnTtVYTAknp2gy17M3Qouc2
SmXvXzOELdNvcRWoIE+gYZrEq9KFkYgOtZ/FqqodYF2ms2+ZimjyXXYd8SRmgRKu
VJ7gwRwJyPd10BNuEAtuMHbgmFcqZbdMicpFMaBmhtbEs9FUUW/oG0Snru10O3g9
fHfM9dI/bGzmmLU5IFUJysDX0kcCqXy8SNy5CDEWo6y3eRZ4bjxOAsAmxZpiGF76
kua/cHkqvRTmb3upxiU0MqXCPZWFA8AakFTqLridiPVkl79J2I23bJtBkf0JqWbf
x6wtxBpl4Fy5hltlvJQ5tnEIWOCI9u69GxZmBiJYamdYgp+yemyxITMQNTpODoaO
rAzFaAgWeyHy4nj0fegvyZko54b5p3Iwd9DD+lwU7NE+lHqZ8MThXWRiY1gP3Kbz
XHR2TXKyPa8oq0w1Wr6FQYGMUixqs85lHl+AeC64V8gxv7SscFO/RUxWiBySSdoV
c2YiC5gFswmO/wlIig7EPXd3KKnQTg/WCH9YfjsxTpPLia+zQbtciO4iQmxwylRI
zSxdQfQwHr8pt/o5GwtwO4W1Fc3CU7UO/t5fXlka7dbTMrY07YgIzbQozWCW633L
IIFI9dpiH8m/Puzt+1EMtkSUvPtHj+delWFtihOrELddKflWr3vvyzT1RnQk5FcM
MJEW0ydHqMBGhOWjS/xB9GdLXliuMSz651QS/D+CU5T/wILU/NBhli1WhFgt0pfF
e/bocutu+VDESkeRix5tCyoQzNQifxADy4vzLZb2nEbYD9Tsrno0ucAwE+cGxKZm
YuXOvelNzSqhdCclSguR4J+pGeZBN01DbFzerwa3087XlNxwQKoF+MR79W0zyHIU
tEHflCu+zlHXIOlS6lyZSONNQCryQSLat750yaezYhOhEZslt1eKoAr5jcmfSsnz
ae5BkUmCtpqYyYJw8P+4nWx6QcWcMURGtw3zBqS+lwS9Zc6lYqTraoCvwULWC/3b
jnS8iHI+JLyxGAcXp1m+JwB5lm/mF+0z9YElA2E4M0sZ/3KqyJOeB8VIKpXMMvFO
EDdBbcXVmGlxKRRRWynVEKOlFhNIsWYY3u9nEtyen1m1MYf6GZ5Mw3jLJ7kfHBh7
ZsHcW9MomDkmRkmRPptNUiGjMV0EaZvemTAs8vDsi5FRItpvYJ03AVKaPEuZNq7a
/wroXMpzl7A2Y6XlS40mmRXrg3QkaxKbfNBJDQWq+Xn/174xeVij8sCwAyIYpJU2
5pjn6bzhEk84vjj5Z/T38wY6mjt0xiaz1PgQQyalgbRe+WOsCz4/1qngko6YKBN4
EGFlvHZBytsXoyaKRnm5HkRb1D5jS4e/f/8muMUseF8XD2Sz9/nOzopOFcStO0rP
5FmwK21ckpY/uQO2+CjjGvpYt2xVrj1zJX0QPr47/Np81d5PB7iX7hxE4aZ0gZry
kN+o1cD2xdhbvO2hTAiZUfpn/vNthtxDz6LDFCF6mGD36DmgOrhsYPFzgow5S9Yo
7patPKNeWGfaCEkUCp31tDRWCGBDLaD6nEWW/dZ3RUDCeR8dpfRb5rHJvka3NCT1
Cw/EE5p1RN5ytUKKZPPXDXxbJrP20nf+7Zb6KmDwDe7BFQu+YsUCu8tx1c1YlbtY
l2aoL/aZ8KUQdbKiV4tJcoRthrKcnacwtysuIvYWgg/YKeOVKlP1JZnpaAO2bydN
kFYXOUDdQthbaQovKfzZaAAo/wlBIzyDDtD9RJiS9kqCdMOjNEI4y/5NGngsVOLY
csRKWjax/OjxTBljc3HM02Cut3IUuM+G5WN7dFfwdUeaD3OTMiiCXKViuC/u+OBY
dsAMcTsZy4DSESFp0d00tV6VKNbciqr3JR4EczBmbcRTWdXWZsbo2QarKAckj7bY
CU6zvN7CF6L38G6YFAKR8nQ2TPBrDZr++7D7HEu/woHT1nlwdo3g8Id/9/JNn21C
2AXN7LUlRsyQLUsssDfq3+37RX+ucKfJfbLWGQmZ8IY1wGWIGa/Qm/l/xJdheeNh
kYs43l6FtLOejt+OjuhWMPPxnD6JUn5FOcesr7RV9Vk1w0IxwaIq47Fztp6JKET0
bOmvzwgwVnXJt60/i0vd6rNaJyGkhZhevUGPHbSi/N/LGCDkExtDRymjJ/YOxCvi
+T4HzjzFq2jz93qX1y2hJjaT6UCWohUEIFkM30+6RiBTp+8+rDSJvwwAuwoullRx
ep7J72mXw0Ent1bVpaoQqDFY8pcPxahz6krLT14+MsXFEdwNiikwWVQOZxOuXXI1
PuxWcg9gjuJlIWxdnJfvTAbdj0UYangSI02mGgnakv3yvPi5FibxrbAIuqquLcX9
vF0N3uaCEM0Sj3VylJxW8S3Bs+E6xrGhikSn08QwYkOg2By1DLjCS7gpB5p42IsY
CRRIdgbQ4n7vGBa+1Nb4XDeto8UuqRDGieZBi9/dE3i71sxalezn6FWE3D0p2lPD
hsBI1/VoHWDxuFvB7WBp1nOOzS8KuPxKt6WK6da9cg9R67DR/l8l4kBE8tQvQk2c
L7YJO95M1Cymwrjjy4EUgba0P0WOY/jsjq57grUyy4f/jq2XLkZHaJSZ1e1OgUVj
8OnvEu1LSyavS4vkttPZXELnAImZWc8sphM+UsIUhg+gr4U5SDJaU6Xfezml6cTM
dFeltjiJK5PpZn+DBXJ3BzReM9hI32RMyxW4GzFh4fUZfsB15Kx3+fEb50ALc5A+
RdgHLNmkj1XpSwEKNlOsXX1BGSZvq6xGVA64d539WU0lE2acHg0ssKsoqKQ2YuL7
4dsP821rLT1senMqzv3c0xYue9yNUbt2lmxPIAklliW0Xn5pIa0zTkX1pMfY9K60
8h11iBBs8xEAmHsy+oH6QO2n5oKDEWHNuwRaKewsSBqs02D/hH/SXNnt5ps464k9
N27KCSolLABwtS9CLs99k4FBbJ/uHTT7J4H+3Pdzp+Gk7iTTeRfono7SRSO7SgLv
gtAi9M6Vb3F+07LkC8Z0KgCcZOyZT8/0XHPSxudXQt9G4MidwLGWvmt9oEW2O47l
qWsKThtJRzEQ8tAeA88N4uH/rT88HZ0idSb1a0Vjc4wAr4xJQqlfGLcb9WxHIBnj
i3g6UZ40b6ADuYOpCAHEIGLGnnOfw4pqyzhr4wK+YiA3W3MvMonqoRF52UD0dva2
j/yCdbTT5j/VuX2iEtpQLlpJlDrS/Y5Hs5C6WjnMUgyLqPkW3yJl3dHSsElX+e2v
g7BbJnwI0tpAACeqow6q0sTtsMDG3Tlds/5t5n9lpRBqCDl3Tc4ksApvPTTNiByh
guB2mSysV8w4sIgdtOZdzDlGaJp5L1CeZ76AQaHef4RjYxDWuyNetDwb73L4rLEN
b6OBH4uX963EmOBK92CCcjfQP6s0LwlyyHqqPTPVhf7MwDriNAoHhZOXektCi77r
YzWSo0PnL7zg6opK2WPNYcW18OXFcsfCnuwiSHbzfXT4sBxZh5R++73vhDMGHZD2
ZlivWvk0k8ejKoxZmLjTLBH5IFEf4Qn22nevKDCbyroNmwkMNbSRfMRPQV0t5iOV
zEH17LbIVmjlmrlGO+s/uRePoDcSBrOqBmYbeSh+F5+/Phy2CmDpGCRAWgRfZ4uN
VVyBWZTWxdKGoRj0GxDmS/C6765nqDteiH2MozaelsH/IWNa03AvNh0Ov10FwaIG
RfRvnlGgssEsmggFbfp2i6mS483DSxfCLqCkJswPDpxBNvFOwdOHRWHfcjpQfpoE
JfQJgqbDJmkjX+uivJFUMXGFMcCqAo+2KZDfjtWtHboNMTqCmrNOhjqX0h8JU16v
5wN/mymwNU+GKmQS+yT6Z1Hlk3f3JsmnvHWAOB9FM79hTW/Dg3kJQ+0nGn8hw08W
fDTDqpfQEwzYMy9X7/wU8p5dPlPtlVlVb8hjQFmPjizwmEyj6O1MNuroJtWqY1kl
yzWtuJ633u1ZSTtHDb94e+cHhAjpX0xMpTvlkATl05FznzDay/KYTULA8J4EOUlH
0aiSeZTEwfeRKCq5R3ZBTg7CZHWfcwA1vqm1mtR/ZqSeTzU/esK9/SvcPxeQGUyE
Q8KO5mJL+tQAsgIOI8bUsrUh8NmCGZ7te6uGR4sHt1qjcbAuyeMC78Ip0uA11Hrp
T7++GAULUbf7wB3b4utopmvCs8Y/zgdmPiReHJshCnXnu+uBmtgAesRyx7+ruoSi
k15iPWeVI7FKn2xD0jq4ZUOI+1MoqOzrzfL4Hm+ftoMWJ6ISR9JMcrVPgqI8+tE6
0ntyT4n7UNRdJuXgTs38TaL1dOL22MyJEmMmMFCre3FfwTHG19bsREntZMUHmHSJ
/MZAyy3vAgNqrTNYqcTBn9H8iA36z7p1dgyvOyTNN/6hbw8tyz+AaCTNLPaS6wo0
jTX62AaxVQnt6K2yDguCcB/0fc7Uz8HWYS4EnlIZbEK684gj57kEUAUe3YKt6ebe
HO2oxgCgW1OxS9JlH6ZrKNxFDJih5/1bqThde/Xcb3T0BKV/aMfoJcX3i73G/p5b
IipNQ6th5nfz3lB31vzuO+QuX6TkrIPZME0VLGEdg/TRZ2N5UN/W3VtVGOGCFrjB
hJivfg6fo8AC/2iGIo79R7qF7/WVF2uPgFoqVQM0/IpKiO5O3cDNEZnEGST5hW4Y
K/QvdRnBYH8e2NPPtvmyKp80fYY+Ki5AIYfkBg1BMGF8VKehsPA/W4hnAw/3uAot
wfstymgtU3YjDfaXlNv+WgaimEQpLEyrzu9bfDp5QsnDQbkmNUf6PiQO8axc/9bU
SYWn59YBl8uRXjuoxwquDc6OUN7b5zHgUyD9NUAlmAEDXCcHB0r7wPIj3XXW/cv+
fIKYF/kcCdOm9Efa95FqFOn2iTDCst+dg1tWC8TukgVDNyAK2iS3PyRfGnfaUah3
8yvRa3DVC6C2bG3/Ml7mIZZd2ikAcDJdATGY2N/O6tTe8LMPyiyJxzzcxK6cLKDz
qZLWVYjh1T/tloENLVn0zOiixq8frhCjlQlWfeDyVa31D7QFQy7WD7ZFrxoFZFKu
G9FSO4PC7wLf+9jljUjTOPeZqh1QPGmVws/GSYxqahyI+GiRyorXiiBm1UgZOrxI
1u1j+R6LLM9BkFup2J+olRXrff2ileN9bOK7GoLkYZc3LJr4m9+uE7Z4TVTkS/S9
8Nh5Az1j3iBXw/hxJ852TE2PHoYIfm9WZRbtKzPq2LlWcTUTFdobYwd3dN8v+b3p
ssJkFQWJUqv6Q0HcDB9EJHF3dbP7E92s56E776xsA3sfgb+KS78w+FCIHSlsAQmh
MS+Sx7wRbq6qMG1twMuAv/6rmZJWxE7E3C+NtTGaqet9XC/4rnr2ImTLZ6vrae4J
jhQhFvOEHAkwfZ52C/dBd5hPWSpwDfiOMFMO/6jHLMb2gEOO1VdrIJzSy5zAgGNF
k46e7V1PpN1TeEEcidFpiE42xdli5AjGBBHsbF5yL65zm30eL3AV6W8BDuGKqL9F
abVt2s0m76/zNzwr3l4MMI1RaOwSRSwWcCs9JKR5+6nlO9z84RzOzlPurxnl6Cni
lng9vEntKdV3rJx+tMEbldbX02Afx+bEWdHN0QgE3lEl80EkLP4PvE0gC6d/J63T
DtgGpMIpCT+54+YgKEw2fKMAplOrcmzwC7JK1+gbnDCHD3Hx+ZIFPE63oodA0ZWb
ntMRO+IKaNAp4kpsr7CwgpHRSZGDvYwKJuB7IXBFwlJSytVFvH2F5gt2oLc8sLxG
zmR1gv03nMFPU+vSP9sJB83qFMzE/hhRG/giR1H2MH+qfHf11yVh37poq2XS8UDE
qSePMNoOFi3ZQZa4ndHsNtYuRI0VN34ir0fBLrbXD5oXIMqRw85EZvlURs2U2aMa
7IhX3Wnjb5oActkPw92kK+iOUryGZKupDDxJq1mAAhxFHrISSn6fHtl5krD4Z/tn
bGIFh4x+8pJxg6mIjaDHwXVdNaTX/lSiPH8TCKvBd3cHhNvNtJHqPeV8SFUV1aTR
FQfFgptmJkQaxFP7yNRh4mIPj7oOjSdSXGav3LOdUwCraSx1dHTv6rkrkoxcJTG1
/3OHL6Z42PYTAkEERu7o+CQre+Ouvp8gc2+hAoxxHpHR+d1QvDtOQKxRW+XmUWJn
Rk0ae1wPpizj2ONjEYqeH399+es+cVkU6ClXGffif5UGLqsEUKRDxOhsL1WsMDXA
5PSVd5EWQWQ5blamqyGZSw+fNhXE8aKKHVmqFiUd/Tho5SoEgn4nfuDNhvzA4p4c
UCvZjMf4/I7f8/wfETLXa2x1anmqLmcip7qxBrTa3Zlo7iBjNu8X3pm4SHO3H9uN
LrJYo8WVge8ZO/vaU+hQB6XYWjeIdTb/eC+NqzdHxAkfJrrQNH5oelxhDClWULWC
usLAHtuX/ynwiLrI8O9ciO79Bd1YKMhul9YtKfi6VQole6DAb6+7fNf2V+aX5MMP
nzELpTkjet5OztNzpdEgtokn8o80MYT0LaVcMs/u9LfS/jDqGgKz861PV5XrnNum
I7Q5LJjUkMISCeo3LcO9LrOT4HnN/rak/0UmvMJvgruHC/xsPaw2Ez2Fml1OlYWC
2A6/Ta6x2ok1lV1ymlkXJ9CcNOfUiUflv7FIN2fg6DGd5GGymWFQeTKSFrUo4vlI
ST4T7JeWEn/vjclgL5r7CYGSZa4uk3FsJdSp3iKRlR8IOgfINlX7hWpxVV3bmDY5
/96Rt70gCp9lXq+MFLvbWY4fCZJuSvDaVpcIqAH+P/dxa6cqLVNkbdlox2TqqAmE
2bNsx/P0RHwRjg632csMY2EZWmBpPxlE92o/d8ZkjURrs5CbbyX+dBmm5njbyjOc
f0de0QFku4ivXn41hn/WUy5SuOclJpUm+RkXerQ8f3zx9E1ZJHsBSjFzgOImxnBY
jvKqBd4OJofXaijvB6q9kBOLJHJeqfqtlGSC5XG+nF6EbvEcM1R5VuwvZL9/SbXr
fHJOPsskHq2EXM1NMNTuGoJJvB3lybrFY5QeqqFUSKTg18lTAO+hg6dzeuu4pwBz
F4QWmvokMGW08NRzwggx0RNpdZYFOER1uxb4HyhZpYiTTX+v6odjFxyljRMmJsT7
QuTvkUdeXG/bwiGXvIcSiZFHF9X0AeYN30jLXsmP35+DAjwZgk4sNKChs1G1LB1t
F3UNUjc1viMOg229vunX93cuw+hpVH3OIi+z246DZ8h7XGtzYmNuTHq4JSvIJH7u
xdlgRbCYOAzhmlM1S/VQRXYc7bqfbhBBRMS7VT3R++PSyVqWnFYLzBIXSQOs/cHS
6GRJLzx57DoGr95mDf5l6VaKPO2ExlEfM8ekgf80iuS5oky22WOtrta6sHAfzagC
p1mXx+6QQne6cTZJqshVylIurgPovjx6ak/Eok5bCsuDjIEWkI0RShXw0Ky1lHfU
I+vWb/ldLN6K8L8zmyonbIZgHEuCpUmeLnTDhdFMaH2tuLQ61fZ7jbEa4vZD1DgP
I6AvQcIYMNSOBVWQY4eCiJHbUWTEcYEwmvchBWXmvaDyF9jS7qbc1WxDUkGl5i1x
O40o8z6N6WPqi365UHJ/yEoRlUHTThXguohpmMDvVuerfMZd5szhWLyOAYqfWWiP
SXSZ5pvRpdIEN0A/Oscv30DrtKnmW9/9PdKMZLL4hRB9GCTXYntchi7FtlU7fwM5
IFB0Te6eF4VHPfyyrthtxbcP1V+wLJaL6x1eIvK3MC4UFDgLzhjqVVTQib0TQ9Ny
m+/V8G5H2U5ptCD0zU9Q+zzLmxejeXtkkeCS4X624RwM/w2Pqr3oxWjgKazETKma
Gup3DVz/9Ly9VP/W6pSFtHVQaGKtc3kseb/tq2YKaKGkqWtGTVxsQUTkvJqUyDdA
oioOvz0Qcq/asR1CAZwC9veNEkmytgXYLRDVQsEdnSi0nDeIkBRX7tlBrikviwp6
l5fJf2NpJyyrP58LeO2jaSeGBhIt+nwhZ7WItZd6n8pP852r8BFaM892SkC+I2fG
fZYshF9O4SZdhNdkqOJeES9o1fiePByiJ1N9qvn2X1OKZ5RKkdCk6MCU2OAm+3XT
RlijAUMU6KJeS6F6z31LbN+BN0taao6OthcNLxQp7wUPm4FitXRrW0vE+4SpT9F/
Y4I92ovb08c5rKKt/mIRAhyxefpzpuRErkW1fEhfPfcXlA4efbeaJRNpK8SDreDF
gdyH4GmKVj2RHshgEg3BBloWPQnNsqc5xiNcGp4w7bgCqhUQFA1tQLNUUFBElsGk
ByHena1eiiioL3p+9lTKOCU/4KRYcQHvHSB7H/TCXe1ISkaMuEohxVFp1fOFs4sO
qPV2HVZzjvY0/0qbEMTP2Nqc7ikVFe54JLnZob7l4UEnqXUmMh28wGBKFRmeRdtX
E6VxtIjzqjQbVNiiDGa4LpXyfRixAlnoWvP/jqi7xv7Wmk5jTRMEt11ff46QgDY1
sc9Ws+9C0JerDEv5J3UsLv18ZoEw439SB3LM4MlbNJmcjN5KaJABUqFz/pklyP1/
BFbMSBxpt4AllBkGWY53dkye9YcDt7D1Cc7PQ9siy1rpxKraGOWBIlkxcltb7u2G
oalAzZGls7ABPzw+k5d+MLoqc0zKWQrSxhlqOnPfo1gTVbueeuoVvpngiBIH3f7A
Lw0qnY15LT5SCC3TCrJLbMg7AgySL0Bcwtiu8UHMBp0tGBy+bCAwLkYqjRG9jTjp
OvS5Sak5ZoeYXgqEsOgW2gZflXQSTpJbNmzkx96Ikfn1Fl2jiEs7IVw6DNg0stO1
URPFFZWkRcQnHY8DoKBgaxy7fLMeVa8Ec/xTTz0/K2zXLXKog/UP5hVHLuIpNu3f
PnE6sXerW0/wQbcjkAojoUBGHkzrp23TQQuJ19CX3ib4u27o7muc82vN4vPu2EFu
/s3QDLDiTNlLdwBqTOrEU+xO/byxdTUGJHJIfadmpUgrHIgXuNIHrmDrhEpwH2rG
wC4Th6AWxfv1XN0mGbumipL5zkwSlXsAbmsLMJvtPzpPujs/tEDJ7HJLVA88jPlk
5aKu/0iqqdlYN+a/7BsNY44kOT88iab6rv2bnrqJAFRHj6VteSPIbVQvmnrw27lU
n52x6Xzmc+GfDSezbAv5TozIR2k4OqKqzTzhGd9664sPGgu2WEWk3FwOJYzG5ElO
RdHaAO2fUCNxku9g9/soL7fgs8exS3pPn4rqPlQfWhTxg+CdKvm5vLFQrl03WUhO
kl1fjQR3kZURdD9/rQBiijrjlvdgxhXxBy5lnq7bilY9cM9YX41qc4gUZIMql1oy
Dghd29btsbFP4bcdF2tfK1Z4fJLtRPXW13qDF/Sp0Y0qzB65EPG1YY+3egxR5xQ9
BLtTbZ8smqHR4uYVesz5WBWuxAWK0sQhKdWOR325mqG5MH/wDKkCQlr5/FvAN0Ez
+Ak2v7xqIBzixWS/DZxi4kdv5Wm0kbFB4n2tmIW4bnPTk7xMUGznzhjOZvb40tGC
4oB8YwY7EatSv/TuHMMZLknA281VMRyFzARffSVLAMXnH9s1n1UpEE7VV/jVqXNO
pEr6CCFUTVQH03wvVxtILswmCqvtJHtOoOfX2m0D4Nh6M5hslhgxtMEUQlkaXcXo
/hYH07bcrPgcGNje6z2i28VDoqD4RR38uxCSJa1Zw/i3IPCDShFBMmNtAObx5l4E
WsjAZtwlNZTRW+dYXe3nJDBILzIzp63OBGeCk66Du8dsSP7PArPd6Z18JqhbyBWf
Yz5m06tpLD8UTIZkZdbBRdAQ4HUhVPOn/aT4QqVJ8fVOetK5ieF6lzo8pc3m0W66
sDUBZTLRc3QxwVz0C7VfX3HFFyMFUySk/vHwegKmv5Zp5X7bJ/iof8lE4CFi4qag
kJNv2SQmWOTRgv4W3bYjO+IVKXgMuh7eXG+i2eLFsDBgdY+d4awnePeWErBm4/9F
ZbZTcv+GHipbOxvoDD3K9uMz/vcnAUyaGrGhEynw6PByWwZLHf2df/bLC1g+8mNW
NGpOtBbJdSYmNA+yLA5pi0YHRJMcg4npgDa8tqjnLQyvSr24aPESK0B63rFElQfC
TtNgJay0ByDhJ7SvMSvBChPh5F5S1FzCz8Vfh4cBDga4aIFFRIX8nNbWHJ2l4EqY
9pU2oickR+OW9IED9m6Yehjn5dexZcKowWjJGzrcxaRPXuaLq/w+Xu8a21+kPAsl
FlkIgtqJBkFsMzqcpcn7ClwOOsB777GkmTqglPx7cYT7zBAbYB3Yjc095PtEcTfM
2kUIYeH2LCnROIRdj5fiFSFn45z/C5xMHyBCicSxIJGAovjbsKP+ZJ9Fwkq7mw6a
QizFWZP9iOaSmUkkhT7bczOIOZbmFgUYbECbt0MRTeSUgj8/2krYddX19cCB94YP
2YqnHotzRjDytwhCTm5efH46vQqd8KqPyJ5iueERW/oJz+dWxkwsOYWnxg/r8vTK
0UZJ/N5olSBMNtlh7NYXlZ57G7X02fnan83Xmu5s3Dh1Z2tMWH7dLZkSltj75F7E
Om+aBM+zb+wdccyxvIh0bSgtU6YhL6Zao7dEGc/Kjl9MP2XRAdRRAOvRY0x5QC3u
XzoFiT4clDpfEoQZYjgNOJMF0zqX+gttD9MDO11lMrIl9hStHBo9YDelI0ANsU3X
ijUKm0qqYpaJ72JrWUND0WPzmtShfkfn9ao8eCR7W+ckVpEkws16N7jHccxTI3s8
u620XCQvnAhPMO9jy4RhasqCYKI98htF3rRWryK7cXgXVsV+XEDZpekAa4X+yY8o
sF/Kr8O2rXUdqke4L8DHEakTguHaqqtNzC21xzSsY2/Jh3FBiG/FOgb9p4q4fa96
SJqH7V6wL0jZeH002FkPcaptAbevo10qJVBz1Dil0DCvnWU4imje77X/taM8GIXx
h2loixIdN6OCbdV1L5vi9PJWbgxwwJCmAAvcmHyL3Aa/4d2i2dUG28IHOvpY8c6O
d2earggtBF+JBxSvUlF9CgmoGdK9IRHqsYVtn5bPYF1Y89xdxLy9qnJg2OvAxat0
VyFPUUlyGFPCEiPAsy61AHU+FXMwNSHxFHQs7UOVstQwC7ljlZQzBpJTFn5bQKxO
UlTEoY0/wRtvkSY6O0smz5lE328ahySOUFESG1u2bXffKs2xjGPhzC/zjrX8tpRZ
/n4S3P++Zaj2SovCqLfz3zG5ZuW0EqS/L6v3bHtZV1m/oVMVzkJcxwkP0ot42zh0
DfePHS8tGiV5BQBEtJYyIwW69pStE8hCvzumC0V1uiIEGLQrRLV7cYosxuSjSKMr
DoSRV2WCaLCGMKyug6pm0zWHPFx6w4GBHGWyt+BOFJFyG3TfbmQsOj8v5wGrO46/
Hd9jMOsxvtMvSc5Of2gnDQQ71QzoXezu8gPtxR+Jmx0RTKIEvoD9Tl7gm9A3gJMi
3dvdIINZJ2mrmbbPtLo6hB2W8Dwy4naIV1lAcXTmzC2UDlXfIN/rPORCivByUBvu
4hIzZRV+BOX4NkNJOgdtYJ0rJi2pdOB9Jw+SHeYY20A1HaeU6pomh1bpr6exN7ZF
DnVxcDAFxY4kftw+NmPRXNZ/dEAxle5Fwu4x2K5zlRRSa/brkiYnjUGZaQ4/E/uY
oq2WIptQ4GAXn8cgMfXeRNmC8hAH6kW9pPem4GPc2EKf/31cCy9fEHOuqybPwCuO
97zwu7JDVDeccQRGpE6TEyQbVvr9MJE4YUb+SoCy+uW8xAomNHJUla32thqGgdMT
ETn3m7dZ9lMNKSVvdYE1PO22cT5KM4w23ppEWHDbOR4IdQoq4Ne159WGvtZWmjHE
CQVh17OqNdHV7YnuSGHJ2iiThzyTBiychh9ULplx8WrtfxktbDXhQ1qHR+W8/1eg
zN7D/oXza0M5lCsgvorSCSu59UqULdTAtGgoDlhangjYgbrIyo0R0E5/sNKFzl/w
jht6pbBESCSKy/mJHb3i7naYWscv7OMQDr4it2iOfMSeNNiDPlmLGnD6dWdTvh4H
BglJr4ZNo2PuD0NqnsONOGy2iPKxptQRZBPB8KZ0LDVpPgD/neX70JEuRTL+SbtE
rdHhQG003X7G0ePOaXNc/GnONRylNTCY6Op5MlWuw5QbAp1308fJcpiOI8tCRcb9
dwZo/AUvajIrMbxaoCQwDu/abWNc7kykbSNUcsLPKYMviR1SpCJg87oyCjHE4hzP
Wv4gEQ7QaKOx5IkeAKPmHHXXZ8RYqznvRewmslfbBiccAUEMoMJEdtzDXO3Z/ckl
pUxAAX1Xbkkc81ZOZ05nBea/xqjTRLeusC4v1ziClAX+BXaj2lhObfuP2hrS3xAX
8dWLijoNMG9Xn9F+ExGBqvDL8Piqv6GfIYXLTB4ageBlHq7dHlGjOvCzrJ0zaOG1
M8LicRZTU5geTHjBzzn0i36nkWF6pXWEZ0mrv4qVAytvrCdDbs0AAnhXRMy9DbGB
4XKj3tCY9XdyWUlZAUJq+kELvssN/tmeDZKsVctKM+SVlI5rF64/YazFYB3rWnwB
50DQOFyc/Pup5x0q2JflzKoTFmTZfUCeGbswE4HvrUEcY7iYrsFMgPtLo08v4bvi
bxMLV7HQCNGYStL60wQOX0g4jSYsAAE/n27mX9vdivsZSELlz88Rmyv+Dq+imsoD
vj0UOL9ibhSVlsFe2I5wKf5z4rr/fzxBd7LCl9JGbq6IDMCVbR9jNMLXcinW5HfQ
mHb6bPasBf47qQub1S++xeabIibQRBU3d56J1hOfOfF8NCvT3wAO9EMZ344oQgVp
GWjxmuRWB6bm+mIBu8wFw/2lFwcgMgBKb/H1xuts8hGZGK7u5uTkIaWn2oxHZ9HM
oLRHyWQVU5Qc6GWMRHWCnCMMXOFpweHtiiDRiReEbAikHe4j4nreNpHoq0HuqGrD
Bz5e+8YDxx/XvCHAQnOrHMqmtY+O/ZSnvJomtthavT7qo3n4pkI/JPPyYmdlMS7k
c2iFfMTIQO8jPDdvZOLm5v4E3AhVz67MIYaVmq5NQCVbdkTWCWoS3HElcop4wgDY
s+WAKFKk3SzRYI7uv0Nny4hvbNKCte+F34UG2o/u4tnOdw2z+A3qSQEtOPM8foxc
kSVrv6xswnyhWvsLwBpl8s0sCb8Hni8sJYtBod48fL5v+kctw//kKgW2Ad/Znois
MiHjp1EJHZ1A/Tc0y0rh5ylF8q0PlQr6OzrGYvDDa4ArhqF2q0JLI/lUna/gOXuk
NfJrZygyh7PMXMjnbmKFMwrEwtd2KP3l02XDPGzdBOQwKpjEj9cOdLm5wGnpEMxJ
HWrtAfuUgz+AsGckeRv56pdTzSzh3uMP0v0UgYdGIliJk581KVPYeTkjuV+Hrir9
brTEoS9i2YO6S5BOJv2JIuxrrfnXk/p4mMVqwsw9w5dsLBtOI6VfuE1A+kwFqrZ/
GeKySAfKezrww5GWYC9BjdjEsVVBPcdE1Wqkw8YEEdj7jRFGdsdOJfLjiN9Ygvy+
k+qCSoo1wLLYxt5ed+CF5Hov+vtzEIeE+LawcwSV9nzIeO82EdA5IsVN/w1+A3No
6iGruBfGhvZ4+ca2TgBjvsqip24I5bU/kAymwVcmW8l0HP7K9BGdD7dQfvNWxjHE
/JtLUw6bXmpHwTJITmJR7GvByadu/wyHgDI4Mu4DGlWeziIebsNpKRwn9P3zfYNc
Y5yKacxczbcZtiHqSXDc11zQ29gphntlqB/gUwuJdzM5u/OJoM6vgZYuow0X3DyJ
zrUJ3q3VyCCEROW+cj8ksA7RI3NBpf5BqN5Bv7OHmiphamM+x9E5DYX4oBG/S1yX
1Fg8L7WeR4aG9ArpzjlOUsuIpmrh6XLKZmC4v8a386N22TtQeT64o9Qo423MWLxT
36L4VKNJz2kdvUUzb2zmFQjr9giKUcu265/vU360040V5LTvZoZSFK56eEPJV06f
aV4iwP8UGxDK2e7u/k/dEgD4JYMJFDAJ64rPxi3IUEZ7T0U1ItdHUEb7tlpD7sFc
Uqcf5507gplNtbAmEmI9GP5F1E4bxc12sABk+5I5Lb2627ZDyp64rwhAhB2Xf5Mv
5Ozs12Fad8MXNQGGt75KzrCACYwxrZJNyeL7dkuZ5NgEIC3GQTtkV38g44ZmXmVj
2YFWtqhvXntl3798ozpfThzUpiUZQTet8O4ok3FR66L975HUZSLqoXCSswt8O4EO
ypv+P7t64qq+7y+DohpLip97ZHWGAtADRw5ovyeBZB3DAsNCJ2FlJNrnLJX3+f/b
nqRE5xq4WRL6f7VcwriCZSOHLNPHrinRJWFokBHiwI9iTp35yzhZ+ZQpsIvl0YBe
UtAttbXvjWqW6FwypG0RfP0nb/zVRhvkcI7MQ89s7qjqnNrDTW94Ec1iP3aBRYw/
NCr675h5LKYujClr55LRZ3DIhLty0QeH5jkI0YJhHtZJLa76pfQgG9VBS6TtbkWA
QIj+NyLWIKl8M8saK1Fi05J2xq27R9rpprDW9WiZMiCKExCEcUH8jj6ayBOVNUzg
MOqtbdZLJKlhNhzvNON5StLBzdmzxnVvT6wjg7W1UarTf6zJYBfVqguJg/Uj7pjt
u/CUCWt9EjyaSMr5jldLFqdDtvXumHUrN2S1AkkjRVgBR3R3oTHmwbjh5Uj/sqH6
Jxt3XBiBT0ig0ZpnEZSAkoMprEBKekOx88bqQhem15+zuAIQiHI+4fVf19b9pG+x
CZF3iK3uNfZ7vJtqQkorsCVsWVj3iS+ytwVygezEeNVXVmms1BgrfhOu3WkWoSBb
Qd+zGfZTHX4yeXn7uLcmvmaJKUDBksaZ2P+0F1nrsdPTMndB9zfXbi3AVjdO4Aqj
RXFDw2x8iDVtAmsvv7qllhU8hr6bF5dUEzAo6SnOPe6yyJH/w6PHycOj57dBYJQx
41sYDZQxKYSARiUsb6CeghBhD3J28xvotNKu0cxfaQMas4t1aH4tqIhFEoMr4RDf
CTyjF4oC5C2PDdaEXnrNbAN39BH60puk2D5GDr2XUB1pL/plMduTwmt4YGJKY6bE
/aLByEYevjjcRV2oPpnrunVNDuTL4m87EGalL4r66D/ZjL/WrgFsf/m7FwA+nif7
e4OXcdSm4Xt82efYQ4kmCJl3D0ot9ApRxi2NjDGtI8bcxN9gs4O7BJVbys82coJ+
nKazQcZF5N5OheVrLp9zYRkGS4q10h3V4IHHYw5d1/COBT+T5s6XEe7xOcjnddCy
T094W8jjyINZU60CKdXcNSUY7ExjwFTgQzC6sHhqCW201aAEU6UP2Y6AGpXHtJvV
hpYbuEd82LRoEdQ7zDIXJLr8fheHhY5vFgV00tYaD1ON6CmBwCYhXHRY7Vp/CKoL
Qpqx7uh115S8c59gm7d3Cfy/l1Sk+lv8TRTul0ACR+LpJzCPsiQMTXKSA/TZIlu/
tY2jKhdfBAnHwNI08eYJlJtfv9sGaqQ3vZMJdmnOGIwRM6HFnYJhNxA3zTawwqTn
ao2w0uwkgy9S5X8yxrNkhJVBCW3NS6HLp/g8kV7yizRkwvNHzunuX8qR4KhEWQFP
gKD7/0N6TKefUBcwLmUuejgcuSAyz8sDuM4CAPGL5/djICGXkhUxTYyc7uYYz4rG
H8nBI+5KwvwJVLjndWc1OpvoVhE428FlB/ZXw21l99tw+XwtHjYsXmZ1aTW3Vugt
uIX1a/NuNjugpk8skSQHJmbdXyZSWbfwMOOqlcyGWQsxvyGC9Zx7Rwm8M6yDBwwT
LQH8JoZxN29jPXp0UTO4wOFtj+kGEF9mESD5ChpfJOmZZox9jUh8D2kZpedxp1lI
+5g8sNjKSfrOE2v1TGHnXkZ6DiF52QVQwnWU5d+oN1aPCcKm0+bNPpCe5rpyxJ6/
nnlynhVgx4CT7SJ6d6sLLH+ZTUXM/EHibVHO692YrAS01HUYup9l1MRqvP2JaCLi
UxPtKYfyuUvf4rrJSZXZAUBtQ5DltmG4bjtJhGkCAQ1864eXcnxZiWLuT7fmytpR
Ojf4mHo5GF7kd/w/H/pRQt9DB/+4MUdo2xjd1iHOkU24+Y4sWZ/rDlvvo6ZFIxZQ
vxlm+fOznuMIKF0NMqOILSRiw5Yx05Cx92R268X+xKOtC3bA1gH08mNptjbQAh7x
MJNgkfUQXj+k+UQ825vSef3iwvSROnUITayNqnEVUjn+be9Dc1HfSObI/+k8OJqF
E68cndfYy5CDRCgjHVRIfVQSfqxsjkVNca5OXU37nhqzrHfMJlX4WWV3xv8dXZbt
Jxt0s4/iXT6aAYsIZncCjS7G8ai4fQHsU29aZjDvcT4pxjCdqKNbEjX8JIomR2EQ
c+FckxVqTlvi/SpRIiWwVIMKaF1uD8o6GUQtBubC2+Uxf8MDt18PW+AtHdPWLJeR
MElF9KLILJuvqBBVmKPfWvqcHDLLnqpmIuGkj4PEH43F/NAtSlx5OTJK7TVEiima
0IX7C2o/aZ9hKnhyisk2ZdycAk9RIYDrhtMw7E10uloqHTtMyW6xI3qAyrlgIxyv
vU2Qsa1pDWCVk29+jBwthRs7hePs1O4QSwfEtS809XPUZFPUaMscEwJ9ZGll/gV+
OPTAmfC8kU9e+4MFMG2PTadJWdgyJYQP0XqTUlBvycCdCh9Z6vJcM6A27pDMLLZM
4d5q7S8fCtof6Xxzds7YPvl3/CPBKKmFAp8X3AdCkKIhHMsqyFYqkwtx2KZqgOGe
a1n1RZUCuHKozViSnRCJw6+FrrlTk0qh+ZGCX/d7FvvnrgT3Yv0E2bM48aevYLiU
sShQ8NP3S/z4O72o7WA0mWV7LwQoidFdp0KnjeiS65+ifOA/v2SFiYmx2F4Uxxzt
vTBdijDh3TI5lPZQPUUWpMaG/5slM9SZGdOxykjki9DGpWoWEESJYlQlOQQWQFme
NW2qczigH0LFIkEtkM43KXDyhgFQuxItfGa4B0Wwd+MxVvqv3I2ZEuSJQCCknFwD
s+Aqsl/rxHAtn6Ng3ZPboMFCw88uJpt+jFnK4NvpdtiJrJhphKmOIZL9O1oXVAzc
trfSKCyfDTsdlt40S+iP7yJ/+T2Cf9HeaBDs99b4A5eg/I45jp4OEEM0PfzgQp/4
YvlRI/E1RCPx1ZxL+wD/1OcJICdotKgk8wxtDCZhE9YPPcuw062cH+K5sre0Aki4
n6b4u3BSjfENjUzRLNO4nqLrU9o3w+nSKX/eqPGMKlSSxPm5YkO8oyRLLQfUCHCh
EhZEiifu/4lSg8bO5B63hDz7Awn3XTb9RfllA6aQPP8Zh6nHTXbxde2Xf8GP4g5g
0AnBeWDKcUHxl0gqPybNc8qEfuvZZ86LNBcswsZIdJS2ANSDdzXPfkoJO+2e1xUS
m1nMy4tyF8eW+jy6uAQ4Y+VMlWdZ1kCa/WwYvQMj9r4CSi72XzMnulshsTopPKJt
Ixa+r5Meuf1yEmF6pZxR8u/UCfIxUUZkanPT+dFXRdAqdGvs18zlbQHjuupKbTMv
oHF8FmT8F4tDjpIdcFH0IV8Xzq30AppRnYkeunBT1QuuiHzppVZQr5eG4L9v2UFV
6olU6Zpjsv7B1fnpl5ZDC8tGp1ZL5zFHMCrsgdRSQazEKvB2w3lK4ks8uTghuCWa
R/pJzPzkOCvIxyOL5ahfmdtdaQLeDl/pMZgntIJmUeMctMmTWNWcUAeNKjgisVpb
NkZFrxIeP29NBhj0kxQY++Nol6lDGuwiLKtGA2BCGjPcGp2AHCAoEVePMmv5EupU
lq1KYaaK/MMCNuKkE79vVuCSwLpWI3ZNXaHAFxF5QGMw/1W/GGFe9FUevs0vwnUc
j6P/34VT1xp7Xgn4R+8P8q22qMp4qZbke0bQ9SjWaCNHMjORTZmQosb/mqPbwtw1
Y/16AwIZnE7YzW7UcBrWnH/GLpBDU8xYo70Gh1do8NGeGGGOOQVOWBSfpxtFkn6u
jPYTKmTVKGdqYzBwYBQnUPpv5RSjukSy1v7E+xuY/xmP3M9FAACU5y/uGOX5TK5K
vGOQu6unE5y4Q6C2Ni/x/bZV5fDqPRILM9qIPRzElTM8wFvfJqzCD/+fpd4kxIsa
z/NJpctAaW3r/rOSxbCBuKDp15dryjzPhw4X2f8NteiDSk47Ukizf/p3UuOkQmEd
36cPN2W28phIVDK3/Rikz2T6LF+Q21i54Kf7Uz/aLxhziDhcjqZ7mAP5rDVRYU2d
Md3q/Oro1sEN87DarhSJz7Y+bhqXtl4JrAZeMdrrQ/pf56CsSs3fDGsB0Jt130bD
gGcDMP8sx3r6TXb2T7Hdz7LdMYI1qEYs52JwYWbQ7LpEv6E0DgH+i7W1sJ7jHbMN
d5I7T2QMt15ZdgqMs1VrXkzifPp9NIqoYRvmkFpQt/4Ox+II2vpogP/1hA4Ztl9m
uWQGlcIm59uK1mpgo1W/mNMfIZ0xm+ASZNG3GjzIgv4gwDxCYIwynX0l59mITlJA
iZk7xmUIl4BV4dIvvkJs7x7XPLWIdbDZxDtK4l6pSlBKm6IgYjPWRsi2xGr9GyuT
FiNXzvN8OP/T8RL5Ckf0BiEqKD7FFEXZ9QSCSYU4G/K1BvynCiOnrybJKvUcpS67
7cEPjWJuM2Q4T/9FgkTWC5zOODkvbXAFfxWg6/6RSjvg213UxmBx9lxPVwH5SQUQ
7/QraCNd/4j/wdy86jJDmQ0AcG1F/J8aR1tIJVOLeYYsvDo5S/CQjK6GZvApGglk
56oa1f0E5XTyUhiwJONgXqtvU1AYJjTdLipYApqdUAx7GguR57MBIOP6QP7juKPg
Rm7jiLmer9QIhHrsnwCcZXn1vrd14BmIt9arM3QKXh4XahsAvnuh50mV8kv7R5d0
13V+xXqX5hXy/Evcy4N1hnTYeTGiILi1zkLJi6rwXaKK4bQZExT8X3vcr65OuVrj
khU4cwU2W8mrp9Ge2954RctPuFGoGN4LUN7WKS2fiBYP6RuZ1FfdaHVjwAROj+JY
bUUv/AjILt5P7AVdxAvBfyYXDS5+jX2jJ07qCCIw3P7J+zx7nZLADlXqY2BUtHe+
4Wi353kH+sbQC2zCkmx+x5TZu2leev5eScNLNQyOIvoNV4rQ9zPJhHvGwcHF8nU7
sX/9jFAOHWPKRoGIF3BrX4WlW3M1g8/XGDSGpGbD8fnXhtoom2X+FTMgqA7ozvXA
jWBk8CifZBW3UbtXLMzVQrjprbSpRrCf8tSCxm5o5Wno+UMXKrCdfPy3IETPcTfG
MPxhq/sHteJVImvkY0QdBVDKFyTZ+DW0orYIPRYkISLk/atsC0nsnqAJoi4ZrQB+
HXaLoKI6QRvepg9dNM3MFtrUGTXXbvSNcrqcqvp/4V4W4PGcl71v60PgsROA9jeR
ox/wMAGYvp/EkMZ3PSjLtIX6UggjkcipwYV6iGRksevmD7ehLE+Kb+zmrEqXvRYD
rVGwdNVOxGfex7SpCc8c+01F/ivomU73O/Vei+rd5pa5NfvJubsPcIn91arl9SX1
ZaoCzmGd/jUNcFAbFLFFUUaS4A13Nu9qJ15MQ2rpWbuAcZS0+uPCQ6ySvRTpmove
25lQU3e84ObhHfTJBavCZ0kSeUKg7nmUuQHfRLth/TVi93w35KHdxkI6RxSUITEa
RGIBoYL6Jo78uwtXLzEzIDB+/ZLBpPDawQ7tG/ct8KUDv2KAFihDWiFBAVp2IwrQ
thCNZ4oieih+c1k1qU9RGYvJvQzc1RCUTzo5862Fu5A3N8uYcyJeAio+6ArIthzi
MsYqtvsITEZC/P2fanC9iHIC1UxFDVO0hnO1QRSpdjCdaAlY4mcywdD5auY1m+uh
hM1hShimMBAP9X2YdiJpn70lZqybtRvWbE8T66dc2uaLGQ6RoporpwS7/lVB9CUi
v/1maOuaWggsaqTCmKcQxY8O35kGFMyetIFZOm80wQhkcKVJY6gGVglrJPhQG9o4
FKU98tplEu5TeviWCBR3zxSVDxRVe3VB/89dRscNLSq2cu6nf1GLbVL3u7ZPkkJg
WTnGyj0kTfSYK77tIm4k+nza2Bb2JYAMIefMJqdySuJj27Y3BrBpuSetFxY9tAcd
iB8uThq88c2w7Vr94VYdfuUDBe4W15DIp1b+wkAF0g2GrW9Zm2sKC62ggz/DXk3o
hzASonN1Vv0ko4nTi/fg4ofom/YbMeiT9haXgb/bTkAlfReKp60Lm+wCEIURZf+f
zxXmIEy5vS5qI4RATPOk/yZU+arLE0QJ0VShwVcyffjsZFogOztPc/dwPS48Joyb
ls8KHE9DwVyXLCIIM00jw26C26V0Ftb+3xCoiTikrhja3eMF83xSqIHj5+dVEFeD
iTDlcPiDaS2LSNIFvVfy9Xk+IyQeX0jAeqMzWtvcX4uO846f6fRvCtWmi0yN0Noc
QpQPKdKj+Pn0wrHiEInamtbstu1DOLNB35046xBCcVhPrBXi8xe5+oE4MDEuwMjn
PE9U7gx7szJKgnu2AI+9K42fDVhCtCT9rKmKmpIhtXguy1czMsX9apzcOsBJEiVz
us4NilvEfgcLMROTcE4bzO4H8/8JZh54xD7DANMyC75nNXIMt8FMmPtG1afEeNPt
NuP3UskbrSwe+cUbu0aJTy/Yr9krJH3bNiXlOGOVhlVYgV965r+PoVq4W7JkoV5R
Adzxj9D7nHk0Yt1Ayd7uBz08TEMe1q4zm8J1WqxqdxwujsP7/70VA24mXUFaWV3+
VO2IzY/LEL96NKuBFGzOSFBnzR48O7MwVVAKW0ottz/xlgG8lIQS/pS5axXGINKO
BgtwhGxmB9Z+3G4WDj8RAB+4/v1zL2NEKStxVODrfJ8Zd7KF5TWcf5h1tqTZl0G4
5Oaisj7nMpxr7GE0kOhizQ9cWNXD7rMw9P/+GnUwHMuBtcKe5qGqfBpYqOxp5gVz
+gsxjuFoLga+F3bRACS0TqKlBdMXGakW9Gitwa3NiBdlBYxOrl5mPQahmvxIMaSb
Gk29ajtXcMXmLNMnZ0j2nfnWEja/05jaJAZSODD4Ajz/x2kfHtNqU9VZuQuFVx90
dhvlI9UazNByvvpsNr96nKU9oVP2utw7d+cdICtk/kw/TWvz+00uDQbckXPZGaPs
vB9FLGROp3i1ib8mO7Is1pgnTABVlsWN75RWQOq8YAs00sFpaIjXZWLP3d0K//pK
yJ3+nIkA/mQc6sgk0nrf05RoLhDya5wUCJbkkOksn9+y1O3sQCxoOvZncLplfpvW
u87SVzP+MZB5mAbC85pDgC8FufR6A1bCsbvB759G2MNDU5RUjdw7XDLS5KH0aMIi
iiYzQ3P/klOkATqcWXQNtq4AhI5jnI+PR8xNVaxPtHytKiBkcdkDdfBziCXNeTLj
qJQ+uMxB2ivapo9PwLMGT4xTBD5P3p8fpI4IwgIz2loMj9U4ilO46hzX0s0DT34a
WumEghzzivRZUF1K0hkhtF7J9UuqLQhnwawU20ZxQOqEv4cgX/y7jHxGz43IdwUU
IfG2AErd6QDqlXxx5ZmVL81kCeeGBiUA7YGE5lABxON/nrHgGLlpqdFKvYhhwLWV
NSXVmquu9m4U6DGX3bSBQvTG33bYoS/hKWvsvM2pwV8JddXyuY9xQxJ8mwAEYmG2
bKT5QqO5ax0ROei/axXZDyUd9xtz+X/YTQ/EA/nK0GQ7S7WsTF3hZbQCqHCQk1eJ
XPhf7oL81jSg4gRLPrATYn3uIHmYwDYhTfzjDY3/AyvYnBSL9schOMPPMEI2oMeh
BGHdnBKVgscPQNf+wN8XE2PulZ2Ra8zD/AjyHhLkfy+uhs05ym8J9fGoWPo8j/b8
onPLcxvKoH5rWfqEIRNVVRcReqtJVeQMYiY98TFFGtKmG7MsIysoqrtBimaFduUx
mGd1l9uwqqH4+/rjH6CmEb0POl8Ro0AoOlQGTkDnv+c83NA2f+Jj/y3h0wkMMvmR
wgFVSFnyiDNmMCugdQJPe1iEhkcVKVu8UBnBV3bec49cTKZJLwPrReonffqeXnys
R41lTVVaGRIWTlsIWFCH9AVQaGU7qx9BousYF3BQK9LbJigSzDXdApHVeJU5P+xy
rDmbDzuWz8mmBWmAzrUR2VVyp7Tb1sW2HjumRW/TkNtczQQfdLNkrG+u1O1nhu6a
zcd3Xc8JFPdkolsWiTLNKApEV7enyHiVZGDbrMu+wAyTLzsVCwk0nQWkGbjhQevs
MNoi/879llrPHDChC3noC3TQU3gocFwcrJAJNjiZ7Qqrv8d7XHYOVrKRgsfXYh6h
LXkTYsrEFv6KZqvDw7gJi7syq3DYaHpOuuNTjKsAW16cmrQO6dgSnfCaJTE7szW6
mjMX/7JZ5ak6BUr52P8hB7M5UKMLGa5YM8nyKCAXsS/PPNo4ZJhlTqF5hngMbl8L
VbbEI6OJBhvHccsFOtHzlJyKhaKmHciDsgbf5rMjOK+vLUhkXQcheuh1EwCe9/+T
InO8n9/dvjsxN8EVQxQ8xW+vD1YFHdrdI9VdKXE+Gi5TRF2mUj9tJqca0eFgGqSS
/drSZ8QMTrpl0lNEWgy2hSmSEgYjT04ebuGpK3R+cR/LQFfxfisSSgqcsL2vX7gm
pkFBpM5WT/ILT75dP3ab+6oWFyxLyaV7w5azj7mBqzgDky6EoWiJ1rEtz+b//hin
RPfR1zM0MYILXY80AoI6bWHrkXAMsAQ5Xctp3RAI7J9/XucvZVMPonqwi9r213pX
QzPF65iJ7Iq5mTKY25LaAT7a4F/RDiDx6hJyPEk2pADkM65x70v9rIyU/oEKDds7
FmdCXDJjc2sYI6NpxTRGQH7BoRbvHR/Y0Mqlh77kyRdnAkd7OD/Q4QCgT1ZC1sYV
jCjueSME1w4v9PUZmJ0B6KYccuIDHzm9aZdckgvXjjSUQO1bjzZT4b+I9w4m3UdG
dCo3WU+s9F8TL42z/2lWD97aIGyuswXNP7fcpQM1k0eHeyuswz2u7bi3AKGNVac9
fbR/BvWYbqRGbU3hAPUM5OyPce7EIR2Z6tmLQ4A9bO6En6SchLgw3aLEe79LTuV6
xQ4pxYSpBJb8M/ab7aAlzyDaVNpKzzI3ktSSL1klQJWvNPjWzV/ry5vyGSTQd4Vg
xa+MUx1paH4fPTw0knyJojmT278WUrDd3JaWktSNZzsp6u/O1afg6el2QL6Rtm4k
9zV5J/dki4uSKreDxXHqRC+AxraEfrcj+/Ak0Mf3nqlO5xrgPA3kU3WsVCO7sWwa
h85TEcxkMdBQMW/jURJ8nsM5G2q1nXeL2NVbOvyQNIBzikWeJP8T744DqaLgtH6I
1res0B5g9gzz95+ZeARp26VQE15jZhNAr1FCZqGN9yPeehqUHX060p1gvQKSkC6Z
/6SxYEjF9Mvqxv5Alw9VgcE1qXn73k/9wzONGWevJQ/kV7MXEmU0Fz/XiFD2poO9
ZhNIMrNhVRLEheW+idjNSnfnqNg9CcOBjE1xVN81in9bA427GZKi6E5JOlWPGL0s
F3mBEwYEorfWpyaZHhfleaEuSygPTWT7FNAdsIOvRoZXAQvhgCiIgKZqUxvT3M+A
KCdtPkrMjVzosqRMo0evZGjrJEfoV5AlVUrMhmSkp3LKOijRrntEQI0Bs8i+/Kpi
bt0cXTCM5UX+IcBESvo4kaTOA5k0VsPRBpcGmZPCoALhPjgRM8xl2GwmMr8Snf36
U211ay1iAsj5dxiVBgEHhBO8oHOCUDq0Kaqph6t3V6AY3IT+kiguA/5/0r+C9jBK
IsvDn1BU82dC6bfjhUNNfSiIp5wtyzKV5XbRG5PBeOS9OxdlHIuviNXVGEGd79HD
CrT1opDnFP/YpJQT0AkrYS9zxNgglY2Zygl4I71yDyE3nepZhl1k78GbQMITuTP9
3hPU0IANMGS8pkEeKNh+h1J+qVQYEnNY0c+6OkhzyLVtf2+ZTEXetmolZmJzVZmE
4uSp3OZdNUVjPeTx4zQec7varOF3768bbNQ1zto5QsCIcjL2+vlgtRChw2RLdaeB
hm+AWrQPio0qqdhxDbUHHMNiVtjYKDShgh+WkBJcGnrOgSkotjObgg2mK/E2Lrmp
B/5FiKxo8y4zd0hEEF2BoycpQLTpZolFqbO4+FjYIMS5PXZQAqtAK1mJEkgmZ4+D
IxSYtJACCdKqm+zxLAJ4ahMkgYvpHMKgNIEf+Ah57mdLdtKh/gIYEDLH9F1AgjMK
p5R9vbZXr/Jdg0uIuhu13IxYt+ipq0bbsQJaotCFnslltJmTrrOHsUenawcbcXOa
Wucl2fGAa0/RNBDjaM10K4yUGNvv1cZNap9oZ6FSSVN/4eFo3UR8bGR+x32DZ41s
VxCMaZSb+hGpoylyII3mrlkYHIwMJSTKZnlLHXZqYA5gLCmvp0TgQ21o1uitjqzY
B0H6pDfIFAzOcFaBAbX2ipg1tFsPQfhfcv7zv7PpZWWDL8bqNCLPIE1RmKs7BIrK
h/jMPJssMihU1B1WnAokaC1cRlkhja3iVIrWLYTzfxD5Kt2/vkhj4lkten8eX1tM
n/dAVlCSYGwGOe1CMHXAHOSUVqo+1hikEF2CvmZwK9qlYZIu4vmiqb5toxFR0UWT
o5f7BCCfRvuT9xSm1KK4R0nW2kVy2niNUchB62CRljNi9nm8TGv9zZP22pj6coIt
f+Qq4pNQwfhMYPj+m+xbl9q8gYg9T7PeAIp3v/XUSfITeNUIVBNW3kfUxvOp5LXc
U1p0XrGsd5DJXrg5i+fCYsE6l26ggSSto9NXa5geXD5Yz6aHEg+GVAuCHvpJrdn7
rP3nt2bDXxdAXLr4X4Zflc5eHWurnx7ntZDyHm9BwRo2NkFhX46i6f1nndH7wU65
pmt7JcztG8TDjFz7VyAouPg0DhEWefqGDlc13hzbqaIlKTzlgNfBvExDCPae6kzs
XIaWGWvuSvjaTZ4bNtsT3o2osjfdeMTE7wqoywIbRTzbqCo3lUAR1xZiUJoYMSGi
DTrtgpT3OtS38bPRfoOQ2CL8ciooyhzhOU5rsgh0Yc15B+E98RykPM8WxA4vp0/t
Cd4LqOJqCPq1bZQo2ejsox8NjprPkbVxrMa3mkjtGHhPM+A74bQxI7X4v35gF+3q
ZLpH2NNi1Hmicw1nZnp9DKT8hMhsG+z82JWQsm1c/okdoIYy5Pwms7GWU0w/N0xr
8z+/ykBbx0O932Nu+07ISCU263lv7KBgKxIUxaaJD6SgmvV3ZmfsBw1V2qLD2E/5
TF0vGTE+BF/AdTxkVeHKu4BNoaOtiAsebzcINcKyZNqoB70FYrjhkENsFczZ98WM
ErkDlfWgNWzVGcugX62OoRR4ivwQD0Clvb64MRz+ahBRpQOalFfxDhUO5qatuIGg
b5dbmaS6ZXgk8SydMUqtQimtjR5sVo1JG1YrQF5gPvRFdGja9vhMsmmI9mc07QKS
Z6SfuTeSGMayAyMq6nbPztj27dwu70pwEEhD6OpbKCcqfLDbpwAN5BAg9jRDd4Zg
NW0yBsO81F+6te8wz31Zb5VtWu6yu6Ks5Zx6X5K4KkCRGIBJoZT34wQvtkB+gGOq
C1H6QNDo0FTHNBnx5OMzk4UpoRTeQ6JiqOFIoSzb7MIi/PETVTT9G0nZxMm/oI4o
bc/BPJS5+WWB2I4/Rwx1cQzdG48IG0JJeSysS1VTA4t9POaMd8rvKhHudOAquvjo
DXRRK722+SYjXEgvpUth1Rgf6UHuXhTTHsf0K10MyHbBEtL7SYc3Y+QVkbes0f5A
gPNwcuuSgVGJKFkT4WpmlysahlkyDgjf+doK1f0ohXJ8UZDzCh6GVpzI4/C1vepF
hrSM6DZ/ONxsCkqvCV1bEzIqBhGL1DeLbXCugURpckJ1+2Q3HrFxTV9oxIJ/15OO
H4U6wBI8NUkepomXlLVHWAMaHcDFZZSWH+rn1UHDeX+X1c1AgGN/ZS4mi3aycEFR
VfDbdJUJBPRwQsvNt3/eIJc7Lq/jOm/q0sP8/Rdwv8i9T9bBwjm0EBdKC9IvLqi8
U0kquWsHxS8iSogrnU83bn3aTQFjEWR19HFWn4FPSTyOYtjsuPkpULl8qejcV7R4
jKFeNAd/DIJpgW5tNJhtfrPS17j3JGSyAg+GRd9AB0Hy4iV1mZMTrONEJwZMjEHq
yxG0J8Hx7CrRjMRTvR6PM9P8k3KDE2skZTxLvS1q3JzLw4FLdX8FhZQ5TS2j+nU+
gCNmQ8yFMev179lIfwAcRP5vbhxXdRIc08YsUjkL9ZtcgXOqfeZ6yRhyEzPM+Osy
PcMmZF0Al1Ln34EBpRBbjHawl/ZlpDWgJThuNNa7nVCe0PBPhZSERZQo2WK2He/8
lAwliTDA1gkuWfk2HlDro7sMx0bFSbqKxgLT+K0o2rNYGX7MJ0NmnUH7NGsN2Wx9
CUxmbQLPiytFfpuQ1jVGf9OH0tAS1T0mzP69Dpua7miDOCEP0YcRTu099wMwVNIO
1zZbpdxUllrkunUfp4aaNUNtyXgdLfqTEw/C+qqUEObf6HWiEdEALriHfYHFC+Bz
xFs/uW+XORU5La7UEOAPe8gQCU9pgUy2p9HOuCFuBgBzVnIvWc4VjrIMPL0MTqGm
/5SuQrjgiSe3wqGUIlY+YQYDQk/YukX6O86SaiQ4LzJwP50YHSM0QSNeQEk4oKFK
Emn9moMwNLJTaGdlBYqNFK7ZdEqPZg9jaosa3q22KiUXgS94epP8D8e24yT46QZr
bZvVFFF6e96akgdBMrpo+7nT+JdkzPftR/cGAB5QwMfz7F7txz/tV4Sfzu8sXxbO
Ln6oX6U9wjR1DaTJuupLKx8xsphSv9s7nFIAH9OqrCVyhPBw3HqeshPV6cKlYeW8
3MPgOhfI2fX6I3VbZ0C4O7SBv4NI5V/SLjKkJKdE+xVJvFbydYNzLdW1q0UN8lDx
zc6F7jQTzMWrDIeszM1SWL+x92SuJyO6xrfOfJVDGOQppEYq4Mlbv7xvwBuw59JV
3Tsp7p7GpYZ8MQz5bOZhei3ToEkRlOhbGeys3X/FNt6l/1JutAkVPsbNukMbWoc/
njiWYqPztGSYUAwm4uGVVL88tUbEupOK1W4YQZP5fhGfI9xoMjglPpN2bqARk1WU
wHjuYJdJnlyWpAAfAl1PJo8JcxIKW2CSu1bzjLQAUoTa2kqgfx/S8HNUISgKZmfV
KCBvGS0A83j1ptGgv36PcPt2Y8c690oDpygq+1EFoJPtWq7ChyYpXwtSCC2C/onM
Cwe0dYhmvscHPfY9H3Xji4he6TPBhw6SVyvoJWS3oaqSVeWKvzXnHy7qaQYZIw6I
9ps7WC/S/5xUu69yveyFVdCsmzcX5hRDblKB73lLGAYMXxIvJwcEPJu51fcDnayv
5WbtPqwMAHDYFdMQXUVPiH0fyIm9FfsBa9P1NA2xFiaC4SQqmnWEqwTfNcK+etwk
q3Dj0kJKsRCo0sgAzgOvKHmhv3fxM2ZkdIiZgGWLkIsxfJnUnhYC9tMqOgr6gpXV
1sxVfO+OfbK8/tDDl6t4NDQ8tqOz/9SaK6lWYopmJfgXHHgdL6u/roXeBFusrvV/
WCWQTEgZ4TTKs8u43C99zoBj2pCxzGZi63izQogzp1TF3McLksWDi/KF9D/4hng+
Vk3KtnXLGoYIbPNL5W0/od9DBT4TajovyUWZ7O5M50POWuq+0oNYWGj8WNtMon1G
C49RT5/1uveQrLEb2wu68AuXgkDl+dbo/zmMVLSSxlKiXxlzp+3x7vfik2g3skM9
uoH4A7d8d2Ay1Ar1TkEakJ+Hf7Y7K5teAWZQQexU94ilZdbXThwOgzZz5WW5/lxq
BYHGMwxmWcXpY1XOlVX/hCf6REgV4cJWyXkgWGf7+0Qub5voKU/IPSiTQdZos0Ay
4u4u35AsR2KZ8E3cjjcH0lc58lViohA2s/Oer43IVxWec2fbQYzPgQypbNDCVDQ6
+x1JGNWpzO1VNDHKwTndp9eiPswXTNjsvXGWmpA2h6e9nDazzlNohpN4OJFyEabO
vB3NbxKm1zts4bo1523vNOhK4hyd/x98iAG9QToH1TFA5q3C6yM7DUZttxs02QPg
Nq0g0nPRdX7JT6tujHVCkcBRQYWhrYp9PVEcs3KUDGinzqrgrmzhrt3+Kke1Q+nN
j/Ye1eNXgeyb47QUyhzxHAa5qTeN08XzjBcnZBYHFW8Zdjpbz5BU/113TuEoDwIl
gVCJf43WpC8sCjzP1WmuWpA6lF0E2egYSO5q5NO4Od6F4Qrc5d2+0BSLIoT2yXF6
fm29Q6N9hTEJ8DzKDby/wpyjhcrBqd3fQasM7wmY+1OmJv2z916x/AY3AbPjIPL5
khBS4gbcEKYPaGgw5Y7FgwUJmkzYadLiqePJh7YvKnAdlQ3xlCwPQ0sF93av/sj0
KSXadSOuHKxJv5bpLkBbp899cD5Byj3YM16dc+jJJenyO6dtAgvimu23MDP74PeD
+o1ac1F8ZZyJdHbbwTNcfC1YhDviH/rHKf9rrkUiNm9y3rjre5JGwNW1l/7JdSvH
k9UCyCBQZ1Q6L4qvHblCF+55zkSnnduhd6uG1CbecBpgR+3hQLEkgi2NqLXc8equ
Y2dtkqF7Q0LYGdUUhD79tKUTkupQazN802f25f4Yxi3C/KAYPB+N5FbUAgCmvouN
0vZ6KOn9W2gNs3gQLNtMMe0YN1igQ8spZ1X67OvJXPQlXRvzAB8RXogRW0YdQxtj
OIJrCiUjVNcawb44gjnk4f8ulVaEPMP+0+WaboEG9bWQVjSYbmAqHRc7XkAB2JgI
4R4Eza1BYRsMPK7ZSmUX/HPFyKfEvHVbLigEAmZtqy3JjUyj/vfrib7qKNCcNwPz
OrtYn/8ARCPf54P0xUOu6uswQvAXdU54yx/YGt8LnFK56ClsBPIIPbSg6ZBpsCop
6Wz+W//5Qdn/jyD/VYvs5WQU727gIP1RgMy4j/4r5OXxHT0gTYlqcS9V7p/2Stmh
d4f4KZ3yq92Tw+4FyVk8t4PpfAKr5BiqL/OrRsEUasjVD154e+QwyYgiDXV2ySIT
0NuV6/P/JegfOWIBojqrlPW4knId0GW5GmbgV71Lz7i5PdMZ15qaiX5L0oOAVypB
vtfS6vsQcXJgTvCF74qAJVd6+UI6UDLww1YVRZJmNsqBKtH2eMfWJXrASk0vHgGH
r5s/QjukTUyLYDD/2gdGdIVqEs9QbmG8yyQ87F0X2oDobwiEYAXQHnkOqJg+ZXtr
YjKUXTj1rRnB3eekhCxsejs0OogImiq8GDiGUKxOEeKINgGTRxTESb5XyVfadHkc
0JW0j3QVsd2GZIdMN9L4zWGyiNMB4U4Ts2JnCWYaQmOOJmV/UOF2b1+xcyhvrivp
LZycBybsikXR2cXDkCAncQGWwBjZG1w39hlMXqE+9Xr3lhc/sw7J1pcIpfoBYktb
CHnRSPDp//F/59PZJExfV5LCHtpJ3Rq3ybcr1qHgnpghKDtOmu8HA6L2nfl9TOND
FX8sNVhqvAIkqMDyfWn6Fm/kBU1zSTgvElmlztIv8MFOnnbkCnIW8V6LWbbVNLJN
hgPldbpDafDxzx8Fp5mLZRKVI0ZKlj56RpEI52BB60OVi3S9qhOM64TXcMceYFEF
Usk6j3Fd6UWF7804lIVVXx8TGQtirn54r7wYp0wD/a9szHtDN+66s2AH8yRPyLqC
Lr80GD1dq3l3DMJwNumhXkHTR4u/8IeNPe7rTDUvqKqX0LpJCCSC+nEBMnBevpC7
A1pWYXe4y8LU1RBZtGGhxUesRTMOviU6jeFTnd2/3yvbQW7bi3nMI/tprJ2tVYp3
dxIxriYICqCvFzq98ZYQZNXmZs3nZGa8otTBcz/+Y1jGdL/FxZqueu4cHiqcGSSC
wAqtDIKmIxeMIftrWX3rXA0JAulHaH7am0iMCESu0Lml36kIYhMh30EC9sJ0cAKs
5F3WtfJwTcWSjFmfp+nTv57M8ZPjHXV2IkKEAxPdyvwm8Es1vyBlD8+cstrtw12X
RhoPVgC0MT2Eb+x9YgynXRy+9zqTmj9K7nhNMKPVxDB+xPrynQDAf+Qsjvgpwux9
ugbwPwpCFvoijRyrJcMilOsDG4b8XE7b0zKsL0oXQHxNMSzJeVxb/vF/RBnDTQRR
8ZWJkLHk1bzGipeIzJeljwLPDLz8dX36SGlwvGt/5Otaf9S4e7lzSb0Q5Lx8o8tZ
swSD+Z05v6kV8kALxXR+WGj6SvwLBew/YeXEXy67E6KhEsQIBifX4f/HJyMSpavZ
PYVyMCEZ5E3DCKq3AeMklZ0DbzXLU/vEsvAMwJ4fOvYMs3Wj+YMs44Psa9cYiOtu
SBUdUknzk+4BkaDCTmETa/dRxi8XkvEKpo1hZyWdgCrR8Yp56QATHE9R8arAeTTJ
1l5B+PrZiINT2GZ9PmY2kIP3oPo5tfIkAOuLG5NpIKzdEFPT/er5KnDwJhU3G1KJ
vP4i+kapPm3Dsag+vKQD36w23KRpIZU/lqADpttGDnqafibW7T08kDviNic6/Eiz
eTWLDLOk3FSUqwm0yAdwAaOBEV9EbVEkjuzHcfuEFXTw9cD9TeK2flfFoth6uhD2
6O4xTYEUAPQzL7/6PB9i4K4NW/Z3YZAlaRLGvNAm7F76N9T93ANKS+QKVcnug/7l
TSosKiMUI7o9mXodr/TElYshQbKw+8T5L0RlJQOaITiE2ME89aFoZd+kwwpwLbBt
ez5XcMdJTK4ATcW+k0Hi9Z/l7sQR8U+WIAHjDTJusHJTaxk/m8oGNmiRH/6iuuY6
OJ+tF8/EEfLz2CBZua4XzhQQemQb9cXfiVePg6JzwFXsTT/Udoq2O+YxTkVz+Jxd
+erQSwDfaJBjkWStdxBR2pGuE4oh9nm+Bi6jlmHn+T2AaHdKeW+f2HCJG1o1DHHi
5Fi6jm9miDs/rafLU2YlDGRzsQX0MB0qYb/EiYn5HlVH0ZvY7+j3En5jM4hUTSCT
AhVnqYfyZ+LlfDq0e2AWqXCH/X5cPlPv/lBjUsgj4BYFqMmL8/x4bmTcJszYVN6a
k9J3knANigRf/98gR4GNzfLBOn7x+XosXC7QF8nHLvaQXDrK3yXVfcbiRL29rcNi
DPMMMGAwpkEaqgj5b6vR7gbUz2mB57hDQxfjY2UP5VTBZSd3iW0VWbyHe7d3JlYo
FleUt4TtJKlgDfKS432Jsk8/XkkqW31HXy+fjqSdnqhTEtEwxaH7vtwt9YYIAjka
7VW8vQ3W+ZJ4jeAaIAnkItI+Xj28RGaPtqsKgHlnAxNeeiozk1xKueyl6k7Zb9oq
ems1Q1JkdkpS0T6YXT6H9IKqib/Z/Rgp4fOV0D+OQI0UYCqmnVceS0pPptnZZQla
KBrnbuXQGEGNA8LMDkcioqMVBUOxOYjFxWg2kM6MZaYcGe9WeR7fztZ9DUrGHmr5
BE2wxuD2AnCDD8ResKlH7TvaxR9ZnRkIRNOR9QqDvLpGroAjnTAQOxRiMy0C9/Jl
dbxAKwtZ42Ktepv3POchz706Z1H4X4rpNnSAIDQimrGSYjjNz+ce5+14lMmhdV+7
JmLowipY3iK+WQghG32W/WVC2lF+B85CducK65pwUPaLsbGGQUEKKBv6/WzweDuH
7sJbZCSO0eTvUfwxcDyjTRp2tQfWxBWp2aX0KsVi6Khf1AYLUhpWu2zgU7R7LqG4
f/TMpwOht3y2GbJ4Gp8d8m5yac+4vK1fPsRFxLVWeTgIHogmwX1ATjNvanoJN/hJ
q0vbhuzEdnoBvPoIouWvvd6raZzBx1ku9DB2pAXEAXkOKbfeG/iUMG3E6hMFGmc6
XzdBbDVu7tEO7u8HDYr7sR7URUz5pAPA9U+lNEV9UFQ59PXqke3kNvJLoOSbFPYk
cAVvoda+6TPYY0sBhsWpyLUqJAvm0w1mgDjNF6ruOCTqvdHxldOdNbaT1zws4amE
uQ19FFwTFiN9wXK4wgKM9r0oU6YMUyyPAkfTTvlKBKZ8EQ9Q2rOg1mLoAFePhX0G
j5txhhylxmwjc+CITPFfwC0sKM32BZ9hGQspkuCSh9oxxvssrSjeiMzZH8HTQYlU
AUwjTeq4bmB9B02IU2lBZJ/Ra4CmR9bC45YwTiisWBLeWnXSOGhdw8wepXdxoZ7X
zwCoieDgKyeNhzNjM14kahMWZxKx3Mn2yJWt7jy1kNPBq80dgIKztx6VXoeWo+hY
DHICEwNiHjKF3drL4q31urdH5qUoG2ofufSJ34c5OXhgDwn5ngI45p3HArypbtsg
IKR5cKG7XTa+c1Jg6kNKNRx5SkOYey0zUAqfgCaZcoYIzvNc+KX54q9GEAVzyAe6
G/039HJ2Np8bdmKMGlB3tf26aRyqYD+j7yVUblnmqTI0+LH7xeS9Uth+YdyaTc7n
6ai11nUNmfJoHOK2UtFTJllCV/qBbUrowu9RZl4/CIzGnKIAHvRjZaFVlO9y18+K
JvFa2jUnrlpyOBUTr0dq2v8f6R+Hp95z1jBI+F4+ymjg/20sFIXfQDSiAGhdWLT3
Q8lkLKan0wfxO/cPAV8qUlEDj4Yzh+VKogJGtuYvRdOHoBxf8q09L1ZDbOCIRWo/
+Xz4ZKSs663DCkimHHvoZ4wxBhGA28TXEp1WJ57x/eC8pZjh40vKg5rvqk82wweX
Avt4Db0r6vfivfcoKXP24kpa91PkXJt41BAvO3Ru+dR7v7Oij60zdU9t5DvJQB7a
F3HnuOwNmC1zz5rLq34eVsIsWscmmJV3xso681eBAqiFamvC2Zlw0xzEjg/x0Ux/
3CI6VYcU9JwmA+B8Mo4Xcg==
`pragma protect end_protected
