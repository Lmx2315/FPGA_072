// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.0std
// ALTERA_TIMESTAMP:Wed Apr 26 13:33:40 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
gOAk8P49XqTM0MnQ9QIRvzoT7sEdvMWuz0q5jK5d01Xu+m+0pFr/BYQFvOtmkQcs
pzUNcXBav63umIqovLbBnDOniaOsgTihfAH+/U1ECCyMTR3nSAIFL/2gdSrUf0rK
Ro+eZ8+MjTC9OuEi5G+9lpvaQbuPZKCjhRcU2I1AYaU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3296)
1eiwWncsRQWLLDsrprpvztn+FVF2wSu2NosXsNsm+mk2Kjp1WrXeTmuESeeTcPd1
XWoutpwyLZ3lqhAZWE2oAPIHvbadtc1wV3Z6ui9DWFJv3rZXpBT8ZT7oEFPAVWLI
9lYrSIdoi0Taj8ik2KPTPh9dS/lqMezR3DyNYR4ikRQ/qYq8DBWH+w4PwduXngcR
AWsaI0OgxTn/0tTvvfd6SVemSWrb2iJlC5L0FXXLRX+gEKpaS9SJ+1yKVat+CDTd
ouk1hn/M8IiAa42/xkSJwV9DL1UHKqbaPba0nrBuFHAlF0Sj6TLqkeZiejUTsNe2
XS1GyCD/JZHEp4+ntiZTYFYO2fRB2pEteZSekp+N2GiokgKFHudw7BHCvcJ3Hg6U
D6TJM9bp7hZiOG7vsDI5UjzTUKUqEjcksOTKZAtRz+h4YWqrzFc+oOO0wtNkp0BV
D+wweqh5p56uZ/kI7hhOk1Vd9+uip0wYIygIw6U9EyDj3LgGO69HtEbpNkkIEPfx
OD0fxeAJtCCdhNI4QSFyTD78alkbfwTQgAvI3L8s2bLlNMfAcxa+UqZgyxtYiS7z
rSsD++l4W1jZa+K/HQQUe+LzSxdr7trnb9MljYus6Jr7XzzZR3QIXsCmn+kADXZG
3E59cqKwgUsBGwpU+XOFNh6saPA66EQ8sNxWMih7CAhh/PetH72vpWkJXkg8WYWY
Bbn3wkHRh+KzYL623pDyv0CSUErDgst31EjwCaVcD2Qf07vSvmudzxGCzsLa5qFz
KsXvxnG7/w1bOiI4Ztym2+fxDig1jk5EIeMPrypje68XDFKifXv+AeP48E2ZE3U+
ZSWo8Cl/w0yPiksulDHVa6Vp/KK/fbPOCQgq2VpBq1MuIlnhEMu+WbeffVZIWtKm
ocler4fwbTkiPMdSGn7NnNneJTlxn/xMcMtLT0lwMVDThPjenMsvjPDRzo4jOZNk
DPe7M2UYA4AE+Nrt2pvbuNyQlOVnEaM5ps9ZgaDvnQgk7AwQZ0FAEhng3r8tMXKP
G3tvkJNAMj4BxrFCxUGxgFM5P2sEG0ngBQMT6DSVrxV+dAyWsYj3Zkk7sDAlGQ55
hrwZphLr2K+bJmG8Dwa1f8DisHpYreb+phYPCW4TTeLmoosBlRN0p+CxSEsXCWlo
UZd5LVC3xk63NTRjn5qk/k2F66rK3hXekgbmOavLhhHuB8l07zf6riHRqYf93bEC
JnA+4h16Xi/X1GWKgo5qoCnlt/TIVJhSOz09kT2x6aKsYBdPESd631fSS2nNtovp
t3Zhj5e6RMogsrFXRXcEB7egJ2I9qpPjYLVmFs1THWm4BvyegWx35de5xWAH5jTx
z6Oi4Yyv4Y6ZtbH/vodhtkfZv6VYEOxyl9w4D/wwBma6JlrCbmKUQFlwQRdlJcmT
/l4h1/Y0ffBVrxBHaMSO6qRKq9OrQIpW4iHsH4AcW0ybheyMRoRYS5LXZ6SgE6aF
P/t8+5MzUUVOCrF/4orNfQW/hxJg4JNjT2kagCkzf6+tiTU7j1ixLXpC9WGyyw/w
g72tFOz+uDAwwKZhLf2YsssweMZg8j7r4TT9QDK64JqO9LPSZi2QKO5JbLD0TW3F
GQc5hjr5WEdi6aFSz4m2B8xpkZmu7jAexn3Wsb88o3zuFWt1DY3ur6HuU7xqQp4/
H2ZQTlf7fzWbMxKL2P3tbWpG2pLS9vR96pkq68wguwx5EjhOpTFQqF60mLl+L3E/
+2U5J6gF1cROOKlV4aM0AVWWXailZXHpG7wyG51/pIbhbE3INnYbaRq2iBSc4INg
8Fg3eZHY6JgHhVQGMSHSUbhc9UsixrFNSVUWI+ASz6u/ez80aPVH29NLIVnDy/xU
Tnp126mgcV8E53g3ATEYvQ2Pqz3qLvlEaec0uEDfJzXEFIuyH2khXKu4FPnCYkA3
q8rvV/Pnilr8o4gFCAvL439MN5Sfy5csC2boxc3Wi5r2upGIhUOxK2QD6Rj1z7BO
mpKJ7E7NP5Rq2YQKL3TkZLCa/k5EONaimO6SAYTsTeOPVKIuy9dPJnS3UmOHufIB
h+axZImpNQldHMWxqeM02tqj0Srct482/2UMgt50ora+UvKi2E/FHXbCXySbiXj/
yDuHjVvOLN+aoRTNmQf4bj8UmenFY7m0W+Oui2ZkIPHNpP/C1iVIIHiPdFNtssE4
pTCtOZfnesCqYXSAE3Ce1aZXYZj+hgYgKCXTa0xGzSUNmnVhiAa66uBRSzlCUQf/
ZZok3B3Kd4HxEC1nOAQ/FEZ/QNvyZ/hb2jQO7DxOVaGmo6qX79+dlJgEZQLT1F4U
RGhEWwew+LFKhgm849QjrRvSp+OcHgd/SoZ3Z6wB4WXTFhFz+E/XgNcJ6N21JogS
YbeeJMj8dGHntchWU0E+nwI47IDNwFMJPoik6D81Mve63cpYXPAK189raOqRONOD
0gMbYPLZfCM3VobodBi5Le2xznQ6XO1KZRHde7f4iGDdVwJPLA/Cc23vpCfjQOfE
oPeCrw+5L7u+FHkrnCPsdhLiNO1g/674fRBLEvhsCswZ39iw2+Iog1EtYKqUP+mQ
kuSr1qWibGxV+RBJjV9vY3LVTeqBVFRP8bedd+R6zSQ8cyy425DWbEaxgHnGDSfF
OxHYZ1ukQ74pMbL3wDp8L/4Vb6V3uL5WDc76x/mDJLhOG8r8WmpBvT0DxmUT/wVx
mHMSFPenU7ir7yTiiNP8SUKzBOZzvMKJU0Y9uAhlNC9f9IhfliocAyHczpehWGtA
C1KtWAWRrCVsPXb8R6hVBO/mopQ1WQuxzTs4kWfzvs0KdEoHbU3lqsW8Xij0+VNr
oqhzvj3Kyleu7DNn15iRvEY7mhWcKk0dz5zKJDVdLkdrHKesXDM1mmlw3Kgw4VXH
XsR/5p3DQlqJZlclB+4Q0/v9J7zdRggcFxbvXH8aSatALqeqQEGunCYVvZf66Izn
6QpyR45/r2I2zyzpr757ttp145CD3HMGH1fLpZ4DRCyq368jNKHYJNSOnIGjICLq
gi/+o+4CpMykK7agiVRwWzwzOYkhCjBdy/saBclc9aKq8i/DM0dmxVjBaGNUE7nS
+/9XUnt00OGB+De0mtm90z5TLVU1bvtf9JdQz2V9KXE4F+LaB3QZNaDVVfQ0aKVs
gtQG5WBkjkJdvHhvIepwRgYI3bKe4UL78EF/UhNHmQ+5BnVDISp3RQEDff50DUuG
a7iIQkKotsCltx8F/IRcQVUt/mZ5hWCKcBV+e5NvO3hkQ5EADChYQR0FF08UBioo
ShRQ7+4fsHsbfpHy+ixVBiuM5Af/KOMAUww+UMDen7226itChVgd2DJ87NiGeSPc
alChKakSsBRudefD0tqjD785/bMU5KuVdNVeF9dR+XfuBMrsxQ+fP/PI2nsKVas5
waH/wRNNC1KTKiNUAIjizCjbD7pDCMHP8UhRUxhGH+q5FjTSiYTnSI4hXXJC5tjC
2TrEkHnaGhf8mfjOYHlygzHJ98TtOumkVEe7HjTjP9AjtqlvWjKIfeG+be+uFRYm
rGnOtjXV7UyaFpGeLUDpsEGWZ+rIWsVUNTtW2CkuiEYWLWOc+5SaA3tUZj7iKnrP
YGyS54lgLb1O0uhHNBcIvVyKKc3tHr74yjLnHUA5YCDdqWKIgLiab0DkCsVbW3dt
tdcZCZHIP2WeKXudPKGRzYlqLYsbigEp6naGUKAqmnO+hMOttFgjnTmrVTS1HIOl
2bTiySCgkLX0Zcl/IlNKTacxWLch9hYZZjZVfIu8cUowBpEY8NAVPMRqX6yeFPiZ
W7CJFgOTh0SQyQHU/NCEd9BeiK8vUZJ1GNRhF+GuOkeiv5wXiQOp5+Z+XNySUk91
RPBwyHYTBOutcC3KjFFdcKHoF/zGendbWHdVgwIyweUX9d3YJFVPhBwW0V7nOuku
FI56KEdQ/z5HgQkBUk3/YtrItTpO84zyskPQEdf+Ijj5TkbIxjAcAfFRdpF/ADNp
yTv6rlfN6coFUwyCX2oOxAcnie83koWX093sNHXryaakwkln1bIZCcEfHcyugEnr
aHKHoy6zDeWU3gEjF4i0VR/RT6CTW2ArMN3jT3jjsDIZda2wNMYPC0wL1U6Kjzpl
rEFDo80MYMpPFSag385lEhP6HAG15AWgr5//dvyqISNH8W5v7mDzW7NfT/oYsKfv
eV5UDFAhuv25gFgZHXMluSFjgXgzzZCZ5MUo9cncO67bv3VtJNEZmYs1D6J/drLF
CQ9lGp9I68S9cG4vECqy+aqn3NlbiNxkUWsVvvc1ab2rkL7kXYkka3tg9VucphFx
/FBt3YnR/pmpIZHSK9VvtgFdfc/GURnhmFUEW8dw2kWw9WNLNm2mpUiUHs8wkAfB
NVF8V5jGqHjEdZ3RPtHhq45iNId/VOOAe+7cqiKSdJA=
`pragma protect end_protected
