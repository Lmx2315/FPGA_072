// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:32:41 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
m1nagb2+09aHVx03CPgEIeEYWkWwTI9KMz/RRMuC2hyVNvS7POOiUDYxVOY6uvRs
XLDpsl5EdFet4uo05T16BgYQ3zkI6Mj0gWdjEWmST2ZZPTzN3X00wdLtkQH0wDaY
vhZLJc67oV+lMWQd5n2fe7EvfxBl0WoIrn/7XUczUXM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 4192)
qDtLlhzMotgofLkrbQkIPrQkUnEx7PXtdgyOC0RHWZ+5XxogKymS/NQrOBJ+GqMV
inbxHGvc2keFeM1OBSjm7a1Uz0N1yVyqj+KO4bPB983IcoHExY7+/nXlh97HdUlU
3EFh4QgcUQJGCJHHzRzZbTu64ddlFUMlzYtvgelnBMPPCkhr86cLKTG+SmdgvVlk
ZSpTTppXnkQJJ6d73BGjOFKR34L5QdaxisU8Nim/DEX5stxngwnHCWpcQULf9Uox
+7G065qKcRmtB3Z1V/2tzsXcyR8TEVs2KhepKA7J6/1Jvft57IKCjAjINZ+nKiAU
LwGdDy213L5Hknw4VZQMycJrOEXJ1pDoEpBPhzQqcXA3WX9LMGVgaVQ8TE60vBfO
tVAyoZLNY7GgcGaWy8Tu76QvswFpX4I1mFj3jL7CEsRbGyumqI4WDss8ML+d+7Ro
3M/A4BfUVAjKotE9sctM/v38UysKNiDfSZymogGgSSJbXNFEz5+QdGN2yLACK67x
UzF4ohWRdfN8WGQpX6NoVq7lMLR4Pjub4vzqFeeI8CX5BKva8C9u5Zje6h5ISa8f
wF162/EnoByIfZuFpaAnCB9/kDQG5BaDNQNE7O1oYKCFOjLmKYr+RsAdognvJJUF
ilCR0TKNSoSM9jus35TRrOecX6ba6qD1dLB/E688oxOykrPZp/+0gIkR1E5450nD
gQpYfgaQts39LayjdI6AYqZeNiA2ll1vNUouTsX0XNJu8LEbDQkgUxRqZ1xQ021A
CFbRTGmBgXaoplgcsj5s408rrTlxEFtTl9BJfrzdxqD30R7XCg+6v5a8U1Gi5lkN
1JkiM2+errh07990KSWPDFcCmBCFbniZMVw8iUGx19BUy98sMkugzMG/ccckKYQ0
T1dzyqit4Dn3eZ20BDpGM4osgLSC0XHv/UmL2S3f6dVh9GvKL5MUoqXMv70AlXHG
xg1vTq2GVUKPAdYlZK3U4hU8bQw/128p/Am4MsVgcikZY14St9lyjPYGBTmeWc7b
4pDnpIz544KdKi6wLiTmQhmQH/Vd0F/QElzdVDYIlihECyt5P/KIHKd24jcgRtDn
WnMhYA9nu4sxuuSD7sooLdMKP0EMWhdfDibKQvomsm2h9qQPFkFUSsdXe/XIpyiy
wlaQJvd5vqKo4cGeWbYp7+n4AN91p82xNxmA+tMJ9T4hH1YoS0tAGdm/r3MilCVk
PKwNq3Diii76u5KkR747FjMG2YidHQmF2WqfrxH7vtzcFqxoRuBjRpLsNPKGALmw
Pnhj+NrKbHtS1CHaU7XV+U/h91gy6jq/5Rnd+vYAgVSKqtYJEfk0TWWdv8md+SKd
kQI9Hrle1/flvIG4a3HclzVMdZ/Hgyb1NFAqxWyyIZq0WGxTJCzbvDzWxjRnNHu5
1eTT77TZFtGwmr/DdiQIP0o/kRv+bSPH43lq6OY/cOhyWlbBongF8yFJCrs/GdR2
Ob7y+q060YN7CYZ0B3svxZHbyex1xctjBHQgll4M/NcY+I4IJ0j0wfA71VxbYyhw
hvsyFVUHhtxzO3b3gBmVhb6nGd4ndkvbm1G6UrvEUqjxFMow+SCmZ3pYgy1c6APm
8XUasRshQNn5pZmLap0QZC2/0KWhid9bhr6Z8jDiqUOITHms9kGSDS6vkHvWi8v9
MUN3/h5WV2xqZin6ujgz+mg5le8b9iWTc8sD2gP7aNH23xbeBbNQdArr78ogeogb
bhoRiV2E1O27/BtzBDyYnZe1KcleWAqpQwK6m+g9EfyfNqGB5OzaJ/z1RlX8l2G8
JaxLboxgCGhE01xPPuCiIksoH+xFzi3nWPDqrxpGFJKUuqnxtyC0Ugb2W+5qfDCv
7oPKzY4160dvySfRor9e6fD0S5b0DODcZ274u9/6zn37IGU5uaDv2nQJrxt7T7Ng
6iDiKUe6UxLsf8getjv4I4D5S0chS0M3gqFvEyFx/bdfFXzY4IP1QamApJVg6oXT
TE2JzFrHYED7o79I2DmHqKVB76t94Cu2YxqwfqKdthfUlEjdQZhiYStUeK2CnlBc
qT3Vbtt1Z2omzx90UMVKZSTj13U4NJ+pCfdm/2EwIwsQii+oMBbuNSLmvWMzL7Sr
k52aeUX+v6WgdIJYGtxhkWcDHcfJ7hZjFw80Vg8njWkLAWPiLV2dgnZdziJ997ZP
blw6dQmwBeJZBblFLmgCHZDd8O3XnNgzLDN99A28263UkeaVstEii5l12T7Gjbre
TUH5r9Mn6yr89FrAnKW12Oqp03yP+HoiQPyOzOBVyJf+hJnH9e58O8i7t0ntps8W
370hntEbBlW129nJgJbeTzhGBupMMIPu4uQLf3bosRMd1QJkcy9hkNMMVwbAP7a6
AKuNcWvRw0pfBt7wb7MkQRuaTqQiCmwZO34U98Sx6mcOtfHQ+xHXUceXIc+D9gL7
wnythBn2ucF59/Fh4/TqrD67p9CsA3h40aeZ0BBKDrvv90f3RypjiBBCgeCmXZJU
TCz8PwqPowWQmzWX69eAcXz0kT6xu45iuRapEp173eCeC5oIxrWmHiZaZT/aXuOm
NiOaVjNPsnYudSy6z9mr7VlFpjiK34qiW0G7fYfhMzd1yQ+GNrnMNHiOBQXpW5zk
1L0mqLb3kcAoGByNgvo+hGfS54nOjd7bzPBwO4R035raiUq9K95B5eJnczD0ZjwW
v67+5ZIE2Cmpcp20rgA8B47vTXPPm2KR02sz/w/RclSNtryBYB8z6AGvHAdlQi0Z
qtDuVYvum95E4qnwuncKBSsBBIiUUvAZBH0sy51WOkKpG1+mRHrW0aVizWoxnS9S
BIYlQlMR+Mdx7bXTI/aAHvsjqiGgWUpqnDA544Qs0FePWtYPXuecLqxHNu7lNefe
Av56RO73VB+XHa9juYYzWGExpKqZSiVZRhTqxROjIGfNdh4214A8LMn3XxMWUamT
ZhzKlMXpI5o5G1m4pRltfLoyoQ6zb+cuHPfjZqzyovlCjGi+LNRufLmmWU/QtrKq
HujowjD+gOzhP6y9TPz5RoPGGNier2AREEaEqbCrh8LRUF2qyRKYfIc6FcEmrKGm
KycRrC1SsA8nq+Wv/ABt3V5/nuaOOpflafKZbxO77TYf3szq2Vpm6MUmapO4EE7H
Lemu7DyVl+w2/Czi51A6EVh/pdyi82lC9Ei0Gs/cYYOaW2ihlHQIOGx0fBnkXdjD
D3+jWbn0jbAwu9zTMbXFGatZwpE+JhnhXn6HYzo7wM8/cIrGriBbfndGEuvydzBX
EnZ0IzPvOCi3uvoSI6qeAhpb8368mHfTXQF+R1eaqkgVtwvhz9YRGQ0k/MfV6KJC
D64C0KQq51eb/jSjO0RHBnliBl/wxWLK6qNEEGQPebvAtyCaJqS2Oe9l8P61J7XI
+6aknUY5XA7Fd0uSyNvV9qXwUpOBoeBDiZkl0WjjrcJSxxzYbjuprgVi4Fec2dhr
leQkDGm6uOSl+kcCLAmXso5zo6HgCwzNQpos33usOTE0SQb7um84rrtqghE9C0yl
U/S5Ghwx9/d4JYr77px9nHV5ndNFuyTuubG/lenn0hclOlbAgV2oCNQ+CoK++mvi
DmLnWDxBbsAdDwIQkgSq8wL0j3JtbnFoqqHMVmZ0eoB5yxNLKW3+5ZO29ArIPpTb
7HYbJKnaWYxrfIed3Auz+DrmljPE+JCKVxInXqCwyXuIcP7DA5acDpU4G8OAS6dV
YIRFH9cKR0cosYpiLEfmU7n0vkYCPrXrUmLXpRpPpvRDYiXZY3VPXuM5fLa3iZ24
prOTZulKlbwM9vQu0ueJpm+km+wclymWAjqU0T/O9da+LkwYZAl9CgX55B0m8PET
mjvuDSq0PeNDzHoOuSfJx0Lq46OD/VXjIv83PZdqoy3it928LZu4Kbrgn7ypS4lw
PZ/pyv+1z92i/+LXDXulh2TBOELryVdNsnrRPU/uisL77DB0RupxYklNV0S55+Bw
v8xefKqRQkVeuI7RgSSTLcPdsmi1ttKX6qiMYiHX/1ttoaNPGTylfSy/UPOBlFBF
TQhhMkGH+p+xgvLRPu3M2GDh5lXUWK+EIundEY6pSHnn5DqSQdV50vRKfnrrCQuR
3a/qa9OR3H2XGIrywTU8yHCFvIXurTJ2zCRh9/948rdCL2QZh02x4+O1a38lNbJn
Cjl8hmUIwixgmN+jz5yUpc2RcPz+lsEZrRCjRZCO3viIwNBIq0NEg3o8Q/bHIQan
C9wRYMgmj16IBXPRq8/q/QuvKHp78Dnu3b92VeFYc0uJEL50ZWxVecYE8B0UKEl+
Af9NsFNMUuWZKFg/nR1MOqHCTr6D9TcqhNlPS2SGJtdK+rb2b85gQ6rInKYs/2zC
SqJd4D7fbJZjoyuQKgct+bYsjQacII8EltPMQW0Fjy8PUY6V36qA2yVGWsBNnD5v
2h4ojx5ONlyE52F9K3rn6o3ccr/cLMzXb/z7Kj2jHzIL2HNt6uCWvMTZ7UGRI6BC
7EuzQVJO/Lr2noj5VqHc3ZuXBt92WuhVg+3k76tr25HDs2oASHno8lmEV0xpW7hC
F4OO8uyn1v+qnHn4aYxtBAY4G7wsFtQ5ecBntSzQx9WxPauLzumh17BT6PrjVrhO
sIOjQZFlR5jIU0VoddnbGT/bL6sakBlagqMIRk75rvSrYrbjDIcKoVyUv2BFaVlR
LPZdKNwTSpRg8dt8JY0VqbxHJOMJ6O7+8Od7XdmBMdamQ/CyQlLIWaCWx4r7Gbcx
HFkmNOiuJYfFtOnCVhWJDWAQ6CoXj2Rt6F3Q6XYxvd4Kr4fTwszTbGQP6BsnjLyC
47yoyXbk99pp221a9bRZiCLJr7FwH1629LXpLwPpjmxYwCY+1iKD2/ZQRlGSxEya
Kq6muwbT90Be3tjiefqbkSBgVn8LMqZTZQfUgiEwHdHzwpaHTSyTJ8/ysEDn7erF
vUyFF7uG6pwYf+Mng4Zp4UI+N9MpsfnFxKUmMprk1w+51ucou+Tjyx/fiVQDzDR9
2dKwAu0pbxsdRUzqqhq6DN47mvhp9uqE7VjBvPChUrpajmthDbI5bljWTDBDSdr+
jyxMl2NO/TgicYdsMVAVuIOdpHAVXjNtZ6e3IhUgglBcMCBhaSLSFQd3HchrDVDj
C4vcJ2Z2g9jx/ondMb0tgV+3Giuoh8CQ4+xONi1RdCNoEYdAcwbqoBxUxMDgQHSO
/rNdYATdC+Nvc0HpP3dalMNMHBrTlE5TSuC5OchQ8WLoIfbDLCGcMyj9KO/7FWF7
JnHKUxx2DwXwUeezieVki1K8Z2zW8+AWJJZdaUf0LWrxp7rMkkBsrM0h2NLeuziK
nwqis6Rv5JXzWRmSshUJght46h3G021g+YDNXuoBpQyQZ+q5AoZNSmsVORaz6Upd
oWCQtY4O5BtoPY4OAtENXqthQ1+M2dKtSLMYPgY+l22ugjys/o/tyi8oIAnPPUiZ
SklvN0fpiCQ0yuTnf2SJ/KVx26rrrEkGVxQ+zNqi5hscgGp7wAU9exKj2pcZZQaC
BszczAfae7+w0M9xa/ne7cJQ1mt+7NLvvFTTtvUWTobKQKfnWPaJxVpHpmqDgPaB
HPS9aNvvjmPONiLzQ5BC9Q==
`pragma protect end_protected
