// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:36:51 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
LLKGuWYqWDFPmwUy8KnDGPO/RA/F2GquTPgCe5g6YNjk93wa99i8hKaCq0PvVec+
y0rXP5OvD0eglBVhjhcfFTNKQ9XSX7nyPWocFrlK6QTPS/lkTWGQmbuN2DwfTcFB
HM45CGxM3hzDHF3hIAhGcdc71XNcKxfVAcLUBjrN4zU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11312)
v8zBdgRD/+0e+gu7Nz9djKUnR2xzVkRsI7oZppRBmnuVmRo6Lgn5nAEx6VPwCo7D
upuESk19k3sUOr+t2NYvzmruzYC2WA9T37wHLEN5SouVgGcfwHSX92RnGPrM35HJ
EKIedYK9+KJaYHw7yCgFn9Ayn1ajZZl2H16rVpqTmVy91UFUlPDdd2XbXFUMMmC1
LmXG28EC5oxQsOdzCtimLvIsRJTBE5q0IE4UKfGAwsgjbQL/D0x9RjBivNSWveRF
RN7QomrvooXQLPZrl6fHC8rqFlglpZv7PJuqBPlvtuuC7wl39HPuC3JvtqN4Io8W
kR4TaTMYVGWDJpbokFGhRngZXKmhZ8+t1WkO+Xh86jA1GFL0/sSwT/1hTtP3Pjkw
ppMj2ir8CHG4W8v4cydJ3t1fHA4GcsbB6BmbfxmpwZdPrXdkm8+Iz86gg3c7ZPF6
5DeAUQL3DrGnFttSdaV33OT1A1RD6/q15q9NyDYSgydmw9cLjcx8EhhYtNVj359r
mW/SUgAV9yhkApNLl98oS0Unh2MqPn3ldk6fAoJSiz2bzTZ0tL3BZUnaN3UVtfnk
g8iDAtoe8MR8arS1jXeTUj7w05TtM/0B1d5fvFiu17Bn3Loq2YR5wfK0oSaK5D/P
C2yQY+CY3UPjnB5JYzuIlolC3SBXrP3onqDGHzhzOEEB/9XQN8/x+y+RHFQtdVin
XDoYQjLIHqUkWaedR9oM/kKOYAF4NsKUwOWhmqIdYPgH4Q+lnpNdhtZO7hFjBMYh
RXBTAQ0E/CRFX5HqAOCMrm4DRFkLv+LSuyzNvgIWd9iZYCve0E6KzKxtHjOXPTDu
/QUDuR6Jj5OygxWk3JnezOqDvHJPDECrfAguj54qiSSuW8uaqH0Ky8075nj0XGRg
tO2D+q8kmoecogIL/2fOEm4Nua0Yd/mvQDHdQXuri3+/yey12Pk8GnZKvVSRsiIW
tykZhq/ed2uORq9feV0fmmV6OVyvAK7X5Vl6HMr+72DYSxjkROVjmDYKYPqc+CDy
wk6Z6Z9IriMoksaYEuU5H5gGfZw9lo2tBAqOQQ6nC3AOg7uGBWebUVKLtJLgkGNZ
hv3nHhPHzrtbUlPPHmWNHD5xeEwQYTn0k5hhO0PnH1JW1BzFFt9yf7fS5lN8GHnA
HWYu7r/nKu87+xOtBEQri4ryHMGEutxvBUDaFo5v3cBJ62mzqI3ZpksomXWEciQX
qMYgpMy8EwcUpfvrjzNAUYuJeo9NGEAY5hxxLMT38CCN04QVnXhbal/Vc1OQlBtZ
HGJXLPHvdqhVQnXaBATnNgmqh3l274HoXHsHY/vLD80hi1RceGZOjYk4zPlYItd9
kGlq/AtdrwQSmgOHh76J8aRGsw263znxlpFe/DXxq9/W3Zcdt17lDWcNurpq/eSX
b0r7BhkJmqbe/0H+wZ/B0j6Z9bD6Vqcrs5RvkfspMOrF9nAfGbs4uz4nmC2Hz+Zg
cZbL0Cm550WNh2R43OOsIZpWn8fkJXip3Olb+rAgTSO6Bo1eUk6VGOnubBrYpqeR
1gdjKkz1ju2GIkkkxnWfx+1cWkXYZf1gwtQvuq2HJVP8BIy0mPf61OWdxDIgWa+a
vJS2a1voSTtN2hexNCx9mz1882NilOm27ZXwyLupJCH7jAQV3WR9dX1WBkgUm3ht
P+g/BgfOB6sW4GK9AN6XuyMe17t9FWH2amE/58gMPL7GIMziZ9fArqj2xJZd+462
t9f4p2AUBSJoun7g5IPP3kI1dM97zEjUF5zEKo/G7AynEgWotnF8T9e7Xh+lxbrV
UVJ339gR3y9UrKUI2/kgA1BRx60l9EjtV69qCzDr8tbJAyUDm5ZEZRJvrWAHPngV
ibStErjJKtYGk+k50L/lCeqSYZ1QjA70jCzoyfzkfDKaWltbiZ/4hEYKHzCRTfo/
RywEJlb+l8DngYCx8pUIyB0CC0Gr7APFHwWCXoBPxhyGlZBTEoksUfW5IsHtr7tP
MCPEmQQI/mNwA+lCmctzaqhk5Ja7HSee7dFfx6O+xHXu4opDCQOeOUrAK9k+BZJI
3X25Ed4IvfczKWLCQyzLpjKvfBhwEbAikPdwppol2ubSKAnndYl+SpEtHRniZY72
a95L2di7mNM8A6wravY1eIo5F8OfLe8Vg6VdNTV+dv6IUO9z67UrS+vDqdVcMbT+
rdWDcwl8W7FYvLsIgznujBtVzfxAWicv61XdUqh6/vGuoPzIBOLCb/a4qelM0V46
2AQhXXRekKFwrmXP50P0+jcu/DOpiZ9CzBonFDEOzI2ORJSZBFfkEZqdzrnK08kt
NVwMA1ZnpLpd4qj52GiyEYf58nj3TH4ONSsnG9BMEFs4weyhXRgeFPeWB/dFW+ke
/cT3gNEWJmcX8rCiUYCBuaJLmZXSM+tyx6CRf9BuQ8N+tLwvsO+oOdTvfqh9QfnD
RMLbJmyNyw37W+4khlTJT0t+nwSkQWYZCbQg8cdKfMAmnlYkks28iPqk1tRdO4Fr
pEkLawa0LDXre0J1DmWyBibB5J0BrjLMJd9idMkhU71uZhT1f9rQsxlD7yuBAW+e
FC1KU9/ifk1yhbsFS6T2UARFZb/ZORpepXZZCpkkcxtO4M1cOP2PSw1FYL1/paCj
DAjietc3CFQNmGcw2MohYfvcft9bKVR3gpZpdK2wwhc7JoA/Ya1xxx+AyDiMTSHu
v5FGsLNEDLtxZg6S/2dmnGIP4CQzs6dkCoOhGQ7nW95aUpAgp8bFt/7G/VKDpSXv
rDSd98Cf1UTbd42eoMRyf3Ws0+Vq+ESqm7KF0ELl9VRfwmOm962FMJrkiOXTyGTI
VLITXHZ8lfTE7VkNhBan1fZLEeluajoE4Q+jDKgfwqld5u/4k9IBP7JTx5At1Nb7
lFwq7zSn2myxXBWSQfXmYlzNWqnAmEZj7S6IfQEhKNAT75Z1tKyV5TbTVc7aGTQP
JqoaUwFMwf/SdgU9rr8XBAFjSxGI3jb0sPQJ7ROoDW70gUfVmpiQ58L+MzutJdUn
7nIqgIxyGJcoHjHPuxuPpsmTWpA/kxSJJjppNLjdd0wBB5d1Iz8rUhaVXO/mQjs4
igilNt+Z8nZmqYC3bAiri6yZkXAnzcud9LiWzLduqp0WAQpsEEs/E80hmT8Pcf0O
lA/eLcACFS79TT2+0lbZIjsKb/TIBN0DsgT8H238cMeqMwI+MNjTNYNwYW00B366
Nt4dZRQ2KVmhWrCo3T5TYlqtBcjg5bwqm+/LJgI+sVcYwq4yjz2A0rBtwpBq6Ufu
R6soG0QYYeViGcgJunLXzplKs9musPJjTSLVlN7Zg+C4QBUT2OWVKy+wbook2Yh0
nSbC42FE/3e0IAI/dHJOSVHxGJ64fWguGMl9HlfjP6IfYky8WO7TtuecKQja5THq
ywGFT9KUtMOUBK4xxfAfaiPJ3r1HHUGD6MNk2x/v917V3/lj0og9viXzPsoz2xRJ
Rc2LqHumPrWORMQO9131DwNxnte4TzsCK0e10ebWPjQlguqTajvXvFH1ayHHvKiG
85+IasIAi1lRWOM39IuzPVnPX36TeOmsAz75XblWn13NEl0QcktoZ/pRlXcLY0aT
0WPb9QwJQUFWsyTeawzV3acYGbjfWZfyxiw10MJDptRTyMHo2Z4r7sT9CWPmQ4xz
qksybuupLvWVKalXucnsUOHNHvk7WeZ+3bRodxoj4xJhrv3z/wTjwuQpewX7T1kL
i3aWivXb+RKQN2h9rszlv04cTLpNoohvNmu3jDIC4BkiBpSGs+HUILAePBzqrEfn
GmdyeDLQJRtiHWJ4GXLu+FPs7C3yVvCAvV8Em4EV7W9syL9BtFsOPjbbV9B8dRks
dJFCTM6mysfo+laa3GXLVNghRv2nni1xOZtD+XNWlVbbL9nx+n2LIZb78tzSKj+Z
bmIdUPnMtvCsoFiwkwUx9aCh6F9B8fHHjrFFrRNonA7R9CeLa0quBOrThortaya6
Zey7aboaAqG6+T5a3XTh1hjnf/veAnpb7fhE93+S1P+CP7ZNOKEMot68sDxer0Kf
JNzK8gJ1Pv2YjecO3uP+B35PPhYrgr5yrNmn34j7b9wqZvLj4yL08KSU0++qmjD8
DnfCTyAXEQjtJHn+2lXgXlZkRxDlv4fy8A1V1Rjf+J9FoaFizNMs9QE1SbaDHS1w
9fdZ7bq10rJKFUCgnaXRbxbMBJifHGvWwiOTouHx4vHfl+iQXP0agGTVAhSMuchr
jDlFg6cLfwmrU1LWLOIeTG4Ct2KmP8285Rn55CEIgdL6PXRwZE+L/ZyubDqXpJDW
2Cg3ot9MlRTpqostEHINnT6qT4Oee5s+y5RrBtWLBPXaBp3XvoxYAgzVIIIe+WY1
OShnu1a4aQ1sVkGMyaPAEUFGhACWofI9BblTeBJY++8BXXOw71i32xVTwQN7JlIP
5k2N+nVmx7zb1dl32m0x3MI/qUHEZ6FtPACFvYtPfa0kTsuU4KiDoLQ0C/46KX3V
A0WX5HzFXFwoaKPqiQLGEFDpHjGosS3iOhSCqhnD2dOwx34NG+HjpRVzI19b9G2h
VL4U6TfZ/9PtPcouVdmH9Wwc53/fEjfl9E/4wU3ZU+zeryVHrKoC3CjdkdlhHqge
/6gmuJeEFH6y2E5GTs8QZ/A3bbsU/aukeqTyo4TjLGfRhjJc0ms2NI32lyqiSFow
FLUbGBxUqfF5a7tXrjwxVXT9U//ksWZCO4CLn8Ej9KSoaFxC/DCWgbw4lDjzP2FG
gGbdhy5Tl8sG1UF3jbZvw2QiNrfvXOGQntXuP5hMdUIapc2E+kVQ/4c5IuEd+mGa
OCasiYogIviGq3HzFKfEzh93uu08J3YWVLSQZE9NkHlYxHbvfhVZcj4EOILtxFA/
KfHY/rpIpf9RXQZ2TvOXYKinX6M26OPlgmWYfGow5nTE1aRwrD6jqq/O9OlgsBDm
+yc0p5z5L8XWznHHeB2djtJiyUV7coFew72l0Zy+QMrB4swcqTzAUgt+ZHNQy+Gw
UzXm9eKRMecftARPwVvf2aIDQpEE4Cq6sIpx/Wp3KQAeA4Z413Nl//gIUz+XSJcw
1bn7+Wz6Pmr0qBJXag+s9Kn1Gpj4DpBd8PY9/64pz7xXY9a1XMRTLZEQewN96mGC
bexnRaP/EbaC+vRDwXVDV1wel/bsENVikTXdWVTrlOH0AxBgyT7HfWWS+R+FLm3k
QvacVPGx7jBZ3GWRtyeXr/Tdw4wweMB51Aqavzt0Ikle26m1Vw/kS/OYQ9+Ubo1R
U1sYtz6eTuAviBrZVCpv4YpLF+51tUB4RDRP40ZcxFDVrpMU5OBqd6P2vnhtmIky
FfQdbm9eYf2UPkYkn4ya1V4AW+eaMw517lAtD57Rs9hhiiE4cwt/kzhCshklu/Kd
OaTeMT5fGcYGf31DZyKRz6K0uuZWEGrccDP7f3UMTzaGpqUm08R2GWoSgww1xcPR
lm0Cmay360hMkRq3KZR9Jr+/11ytSYbJq2yAHF3efMajTAOHXdbrnUyJtN9jwOpk
nBisQ5sF+HG/WwH0cRERRLhIzjGGiD5bvh9IfMGFkWk5OMI5TA12RU/ajjzeqA4p
3i0EsB+lmlp30sc+pXWSRAJb1KONC8FqtzZbZg34zms1oQXWWl3srGpx5VTWF2I+
jQKJn7Ty8FHWXN5wkqoESvylsmwTiOOtvnuF+9h1b0dDYeirZFfwf6uWGHfICq/h
Dfz3m8nPeiC5e6rI1nPv7+ScwRqj+Z0QZAGsSUxWN89hJeKcc35I8elpM9tUlVw7
dH6NGkL5F0ALKAMMxpVt8cKah4+5mg5275ObQbkfM3FNMM2Fy3G0bMYNxtCWpAAs
vvSkhoU0R7RW2kVrX8BpO05/BnnIGiqy9JoHGExfcJOJoIaxH/xI10dQdMzdAZ0+
9GkQ1EFqYA0UWhrYxP6jUssRjxt+Q4f3m0NTjO6DdSoAAMhqVCBi5vFTNC+WiTHB
miWug2pmSmNV/Ic+irnZrxW+Nv96POT1rJAYySa8oFEBpR36Ke0QGQ4LdnmQHhTc
7yviKf5mrGWrPhpP9XyZ694LgNNvio9oCLU/9egLCuvxtertQz49vMIpvDSVJEAI
tjJRbk5UXHhXvRQ668EnJsbtDuK5msJKdCY9dK9xtiA0+oVOF5xFWIAP68sW5y4O
ZGlKP7VFK0HjYnr9355pj7YpfIGiRRgsXPIYmPxGRdNY5zyzousjdxUmpqpPoIqP
Xo+IQxsvYFaOHrBxHFN4Nx0SaoDuX2G+GN+VC9I3l+md4lqBi5K1oSqnQgEN6Tom
K8+gfR7ADrMmYnPr0pikctBHmDzzMuH7MUSZBiMuDtQzLWau/N7zmj6X/TPOoA2l
/K1vnmdl3GqLsgZ+hMlUH3qwaO2rvF/T+Y7SHb8hZOlmtQJCnieX862+NHc/PVHa
zep5dt0UA8iD8Sla/Zr5Mh2caujdNlT0geMwrU4idl9Il0aSEorS/f1iZ4hA6Zm8
bQRbZ75scjPL1q1gipSkATTz2aZ/B4eCIVIZQMRbFKTw+e3VCwcPJ0DsAuG0E/4d
mEkJ/5X9uMsEfHeVrBRXRIXrD99gwY/F+hhlUGxJH1HNQ4s+b63S2esBvwWV18Mq
KDf197smIe2xnJHMHjFshAGhKwKmaF1awYXeX77fS5jXmYram2MPWpzCw2qxFLsh
HmWGVx9tklscLCpoT2Uli4N0OD1pTnREsR7DcO9Mklfuu6Hl6SgsU8qXL37Ms5Se
a6oYgYoF9XoUMJHXLObSc9QFjt++ngVFpuHXosTU09mk9Bx/BIzRXQJ0tfzqyIt+
7uQmP8zDn+ZzgJMpA+UlQPi1wdEYZ/N5Heq5IZcRa4YEmrNsTA1W8n1dyfgaJJS5
6+OMOmZYOSpPK+Go0x61eD8EnUrw0R+jFCgOWhGSd9KA058jo96tbHK2KnZgaI1c
odHUJP2zmt6XqDgwG0IFY58DzJF6sl1ERflQIklE7GMWoKcSxF2vFdZit4BNMG+y
xI4up9tLfL602FqeGXEmLFgVB5an6mcuSlr4Tn5a+KJbBM/Q47x2wX057W1n5y4O
JJPF//mP9YM+PTLJ6toNdn/MWqSz+/tr62zRTYBxv8JQtf8J8QJ6HnAUllDDXeAy
nXwi2o7BFeeZsIfET92heUV3yDvotYUnq5avvJ1CLRbYi+7kZEwhgF6Hwz8r5grs
sC+AawUJEsn8J/f4HgMyzzIMUPIzbFhjghZtSuJACNpnHBlZn5Sd6l4Nbhq1yL3W
RqLuO242E1XKvVRZG0y0ue5MsLrMWB+plU13bp4SlJ8L+hqmVuADq+OXgrcf3wlp
kgWvwEbkev2Kh5CriNzEc6GoRYcwUBQArhfxiwNlXEXdH+Jgsm2jKdUDxum6eypu
PybzJQl/5wDqmgBhnD935GeYGdcq/KK7tbQ1XQ2q4CaOVrwCp4s0or5y2qTV0rbw
ptFe86FKhlBPmledSnUNxiqWPIzrFT4W86+WcUCTmlEOOCe1pkqPhcnCpu4KKHSg
WuA+9g1M12toKgk2Jtt06SnDSMVW7EDsrHz9n2l+tg9IYJAXenJc7BmcR3SBPPhb
75kFki1C3WvBuWzp/0pMthtMSAi8j24e6Gczs8c4TyzsCzJ0OgfgFGl52htSxYpr
8dyl2A30Hc4iJKwle53QvDtNJ+alPPdpnHxwpYeMPZPecwSa/xor9dt5nGrt5XTS
hJ0ACRDhX3S+/8E9MtmJNx7pjwlNYYATi1HUzqOi7lsxwG/BHIPEn9jNDrvkRTjw
L17WOLb9q4Z8LvCEhdA9J99hHIXY3hTmiBe7GGCOZDkkTtFk8vGK/dFQz0T6vfn4
ESmCMNzgdIEPBtYfGxkho8lan81CjSe1ardowJWBqVU0ygAKyICwnD/oJVW46+VG
sJ9193ur8BAjj1+ti46PjQlk/KUWI+M0X9Xvj+ZgB90pEPVNAAaVvBtQdFqBjjES
WCqKtS3iP606gC2ZVooyxFUZrkTJiG6FYsfHRoe8Wgtexp+QC5UbtP4ZOHxJLzEP
7fqxkJD81COOu5vDPfPrNziRRi0yuFrMgC2CUUbIE4gFTVWG/JsnqtskkOy/LZ/E
mFrdVQ5fJ4x2ST6LrbUEN8gvZDnkQjNIs4HJP4XQNgGxOdsGo5WK6GPhkSE5JAgz
Y3cylkFZ9whAG59/OqddrHPHmCVvkyRO3tQ9zwZyA0FbYXxGWMYO8WA62HaQrmr6
3iMJVMXPY/z+kjGTeMHh5ipQh5lz7meaSua7rEXNFPmiAwV4cfVTnbxboG7XUM07
y9fL35ECgpXOtKesQInWqQVvc/yw4/AWg6gQGJD3WRMapdjql8dgUDTocwxwV+97
3mwsEgLOysORYkV2KURJP8303pxhIkh8Pq31ZfUyfHvoDZbm/Ia7hNauHgf08rBT
t9KEAbYdLynynkvXET+NUQRXKKZbnrZTC/4lWLl+E+xVrO0Jy7zwHDFnF5mVzX7H
rqfdmx/RLaNLR381lQKQV4iGFpotfqVDZoR1NovEML1/OzC/m6vJBUtMLL9zFfTO
yTZ4itQf0tGZEyXgDyQHCD0X2ZWlnJajr2CvyO4+aLS+PvdJwRN0IeE9NBQzxKAM
q6uJ4vTRQ7NBtwSVLtncgoqZdaxBIujObhCkKjUAX0I2wbkQwnGDaddd94vnsgmZ
/EfWC2xSybcqFQ/ECEfzRs8WLi4ccT4ye33xnRbX2q1YjmB+d16XUaKr+6csewnU
6Ong5x67FYza4Qwf3FhYU7OlyQx5qegn//4B4DuZ2tpdGEd4A6axIiNMwqoacrqv
YImGZ2hL3mZwqIf3SvtbEcaD3ujXdiN7qiUhveSKqgD1uDfjN3Wa7nEbWcp6cPd3
J3hRG60TafdqayLpHFqCjT+T+U2QW/P1Vr0k39xqzvRI17BMTZAnl7wtbdBlygdt
2TqUXfBclRdbgTaVom3arHQe7u95NhJ5WKcM4TOjtuljorY3BZsCi1flQf8hQ3Q9
CxvObVnPbiv3gS5FT0aXyIyDtnDW9KA9/WFAz3mWfunCb2uIsPgnyriXfjVYpCGp
UHWOPTucqlTMHHv01bSDquwOcsFVoQ7nUXhi5dz9bP2DE+VHDlv4COaFcOGKNrZi
kJ20ACEq+xec7/5SbvQpSzjdRRydrMqLmsQEvEnt+eyFPCtA8bKyIVrNS/tiLVHK
ommAmGnSbKZl3CO2CAiRjdhjjm2o2HOQKQiAECH9eVSUBr2UZJMBa6Scu7CK5VNv
YDRXWvNtoBqHmEqdeECxHocSSVHm+Kce69Kw9XvM/Bgq6J00TPJojXJHSo9JVNht
Cq8V4prFZxGywgIL3EEA7O9urzy1GKbipkgoOzZW4QPhjcsXcH0Okk8aFFquV/oo
lDlVA1sL+t0w54qrfOMvSvRxJ7qH7Dty6zzNAcyKr9XH4g2si1Ykejt6SjTwM47M
vGO6PSf4NxpCkFSKjRF3cSchqF46NOA8VY+cwAP8AVW89AEGNgCbsnaH65Rd/7J+
PCkDFW5wgaC0WPN5l7gfIEnCRuVU36ea4D4YoB+yfTrNFFRB/wVOcJXHmxncZeqU
u2R3jbDJ/Wy3pcnZQ4UMQ00fcT+DVEDYooM+2kYawDt9SwZ/fVH00jYTKYveRsQb
L3JkhJYKqnGM4Pxg0/FDRwlMaEBKDRAMvXzR10dC7TiPbbijmtm7it/qY0hqekeW
NXgcY01m+nnkFkDCUUDLvPScG8rEv540HfXW8AUOppjxFjcDyYj07dRCCB5COTOz
OhPW0DbLlRWtOJpYtWl0CsZp7InSq06oqAek0Bw2mN/iPVfO9yXAH6Zxv/FUi1Ku
zGLlXkKk63eH3lLkgNMYHVtuP4x5Q7BQSGKAv4Vmc/S7KYULldGERM63EGyqw6Vk
+LvrmdLJcf5UXWfiSgSPv0bZfhJPx98ka2vBLBFCy2OR+uLxCVOOj0v4epmmfgMX
TMQKlu7v+DwE3DabFsUyMyA4WDyp2qGBxwzR1kJhroV2ht6a6Lpe6+FsS9Jftawy
irAk+oto41bMpKR9pLGzz+LF83M5qh4vDv5DSvVxMJshUIoOhXW3OW2SHnwCFbfD
yUwvuQxRQDt5YSoCJE1kzfGkQuBu8EdXU9FZjJQ35kaWcYr+i9DhE1NW+rAogELJ
ANi2wgeMuzUnxoDIA1pEZuv+7fLz0J0VXpzPcUFkma5k/LyLiLyvpCt2784IN4NA
IA36LLJ2tzvcYa+aIFD2d3kI6hPnuNyW27svFQxeumD7t6tLP8v9j+lsvrXujm7l
qepLfVCic1UmGgOFGbZkEA+UxxsmIZUGRGPWgFTFx9ZFJ9n+NOIqFmS9IdlWmja/
Dna7sJac8a6A/XXiHGvA7K98mnMMcc3zRZLGuI0B3ROtqwqxENWZYBD34qmDwCgC
Y9tx4aBOxHfi63fxX/jgipM89Zp5hNQt80DxGwq8bBxI1Zj/5P058GVTTAurymM0
ZJXLcVlMAkeldE8mPGkXJCc0Evx/14jAf2w8SpZoSm0EUZQaNTZMu2uUb8hV+uwa
PCsXAHa1Z3eoHnSyHnu8WM1yoZcT8QiqVYvIqPJ3QZ69nunDU+4ioD08djN/vU1k
zw1g/KYp8AjPZCKHRxNaaVMAeEvsZA4lXsO4IIF19+aJlMngbYSVE+ADCJo1IdT9
JBNwqFBwJYsnSNMJfYC3pWHRPE4YDNg+qckahoBbBIuqmQMaJYtz9We+DdQtPA0s
ATkUJQoLDpVqzWhBLm/kNRdY9nEh2vXLHKzi0kFtn/nROCyEbdtLfYkQn3R6iWXz
A0EZnWAp4iiROkr+0rOlRfKXNMDEU+IGQX0JSU8s6kiNK9PZ+JvnqAc42Hty+nD5
58U3/8XQzZ7NedP0RRqgT031x0FmkUrEr3JMVOEU0rZq1R/YHBqPFM1cOB1JDFtq
PsAKyLTFOIcFfKgw4I5MAyErfn7OfXmhVAhBY1jOvOKSuhR5b3IzljfZi4HmJlMN
y+WXKGrX7he6GtUNBugzTjlh+6Ehk+WbcPI6iw8KwCS0rk48pdfwmoiao07KFr+F
o+X+/JcLy3xB/8SaqEVLn70kT7I6BP+NlLHaNTEcigUYqElyh7FVNmXi8Vx5M0RW
yQii/bs9eiuEYoV6II7U7iV3tSoNMzcc0cRCVcYHev4xdpS9Ms/oVZkfZXkB5dGO
cTlQ/fEhpc4Pb/JlyxvEMSOYPtYeAvrxfCh5ZDcfYUWNmj2WjaA/MPNJHa3/ydkt
t8nD1790rploXaEK1eAvHPBX0wkMkCWqtRUy53ufpS8HSlILL6Hii68r6AFn1NAv
+2Ws4XiTw+o8tCh2GCebwgAREv0Dzc+NUixpmv+GZoSMIkae0g7StyyqBZ9xrrUh
Y4cjjXAE2LkNNZ+qUHTooaVTA3kTtpK2i+T47FGWflgXArdANUVYCB1hip3NyU/e
taJmVKxwhxMKsPp2C7yWzWJkyU1sIFY6x6ssPjsgCUWedFTuJpsHHDq60s5oAW8Q
AVzkZV6wMX2oUZm2GPaK8i8t6wQFfRB4GWYHnJJl/fhcCvQu/UE5I1Il7Xsdc4g0
PzBivYenzR5l2OIRqSs3/GdlynqAzHsdiNNs5v5e63ncT0Ub2orJ+Wjeqhz+ooRO
mIAbaFFwwRkRxeyb3c3GL6nJKDltirnA6OCidssOnvQ6DdUtVenxLPHDQKUPQap0
nxdNtNJKo3DS0YLm1bnd6kND4/BoiwHk76J4mNq0Zs2im8/YOHQSySw11lpUJT92
/DJl+pd4bs9l/YfhyyLuGDFZmj+YWnjPY+3/QfduNT42OLFzcbg6vscDj9ZNOt4g
kERTC/+a63unZtvo5ilQblJOYNslhAMPAhvk/dMdAEcW8RBZKeANngUSydgv+uYF
cM01MD4FhLm87WCAVrTS9/itj7PRdmEbmz4nfDtxlvodE3gabWvaw3ct5Cgz68wQ
n0hsogZ60Ms0Iq2yzVtJV6Zo/26d7RDTvZ+/NuEZgHKTgQxC5hspkYgm+M1r6T/+
5I1Ne2+72Up4yt3bbpxQPRMV6L2ndoSDBXPK42yXuuy1Ppi25l4Qltvf8DrqqFix
frl00hEe1dqUfqY+3nfqL0k1EEo13jn3u4cJnJunwElBN69xPCZmnZ8WH5DQLl4e
iiAOQLc1CGUgbYBvOLXtgAVcjBlqBUezQzx9loFzh5FlMbdXCG3YwLdAiN+71L1U
8hwYxQCxLxJSnLuBVjXi44ID9foPT4UcevjmxXapFhIhCRFkB1WHRV05t1KNjXw1
9hY5n2C0D3LVBh/3oHe7WTmZoLYEkn3Zah6YUHXG3A8q7M2A/KG3EwhtE5UiMuQO
KD4C0MV1sHUa/8wAwbXl823yF5qBWrKMtgbuDPikrHs8Yd/q+pnqUgNzhqm45pvd
AN40Hw+GWFPQnCq07E0mbhxb9OJkyEACTLulO3j6L+CfEqG6pcf/3+ukFtrAxSnv
y3L65eYIcbcKTCYIndFQKcegirLRMt+j/Voemb88Rjs5D4m8qXZoGKD2we4FDPGH
efaADhmf/FeoSqgfX1WjfJhNnCUoB807vNmYXekDZZu9+J2JO+Po8phPYXMaWmxz
oGsndrhtnDmD/E0ls+3yccXzW0Hy3W+qIAcIdEnWgKeLNM6tD7hRdfWf5EDVln6p
4mU4M1XD0ksciihwqiK72k8qBwSy6CKdgrqMKjvg3N2kwwA1mk2TF728PcEdoPso
Bl4gabWJjeh2ZOdY4OGR+ylSD7bc1SpEDgyjP1O2Nk4FIY6EqP/w6SIZdkrz5q+E
ing6UUttqt30mkBy1q9ndx/NpELjwZhuYtrf7n7dFlo1Lflsa7FiVlytPQk4+B5q
Quc++vszogavZPza3cBTS+gNypkaXtQymMACc/qM96t1xKk5UM0sEXEY8W3EzM1D
89x3IWDHFKB3in9BQ8Rlxo42FUxtdx9leDILouZq+UsMkIPODY7DXT3YGmNok8UQ
TtHoOnT6frRNeHWTivIDFyqSgHQPSB+EY2Bupzdfw0vEkostBIoxVcVxLkNg6sS9
UNdBcAYivqRsvElVHg0nK80U5Dbq+a109FPTO+HG482BlQqBpm48AYrjMUCd54re
ilxomdbCC13TaiX96C0AHGxRQ+X4e4fbvPQBPipp3i1+uaJlWaJ7rVB9XgxFgl7A
owBYlg58NMrub7+QI6+XTuNAGr4yHkxwOb3b6g14EatdG+F8kDS6gIyVk0WBVqOk
Xz+WvMbBEMhKvWs5TVyG/TWoHnfTyw/njjvp+Jv+zPGKuseqrwo4XJ/xz6uqDQWV
ABEQaQNhSOh9rlZ5QvTphCIemWD5I7TeCLEwpEhxled5w0ihuJJnxnjrxMunml+g
V+XKWFRmEbmiQ7Vk4x23VbkU7e5cdJRuG5fuYJS6gQ/R9JtdeUD5iiAe17BPNKSr
OQcm2evmgn6Bbh3mw9aMENil74kw584dU+UWXKbx7+5WHbyVW/B7oXdOfQHMKkgn
pBBE4kFX/EVZiLvNCKyZX9kEOD6F7eQ5jrqfvJs4GhwtzbPQsuvkBYSxVoFKXbKQ
zsAaVSS4+K/RfhdhxbDiaSbSfMEcAeAeZproztCiERzQ+NTNGk3TWQneA8kSi5aI
Y/IZv6yo1BCLLE3NIPHjWX+GSfulfV82lTWg4F7ZI5V2//qp3rXE4NzUFZb6rJEm
8FvZdURwk8qzBCHapQ6/qjTBnzmepFKaQrRQsaZSfMZ3QWklyyGsr8DQi99eUAGp
bj88C0NxuavpuGk4YdT7MruduX+A0LN5RwCsmvoVhivmZq9ytZpNTb709rlxhr4y
LwSND0SBuaQ2tvodanJdwQqhmv47oHP7etmnq1jK7G2627YhTADsQU5YuRfvI1k6
MKErFf/ccK2zG+MEhQCQ2Pc9ufNP1FzQMJF6eA9b0lEhgRw+KhnIOejBQzAXTaJB
8yS0GAV9ODFot5/D6tGTlybD7ZX8fdUx0JOBhdJmWaFWgYsQUexgfFnU6xRjlSxv
T9dHqBMM1fg1jFQu865OPTpk16Xy7zmrlVTevaURgvypxge8q4jP5g3c0d8E6bBj
EOXUILM9qtPpMj01irHXqz/YjPPfj96gv2I8F+CpOxIJoctbcpaUYV1etRQ8Pjim
qomRI2s0/8K712kZH9QXGRL5PcusrQlE6n5V5WBbRpsS4rnUyweCYtfnBtlisApO
Mo53dGpdtCDhXIH2ZZQbJhdgIH81pKBRKC4eiuJ78ejnI2ehxTLPcm5TvfzHGbpL
XY+a1/YZmCZZiCZlnjRnHE4nAomJjUY/B9e/5In92rkIBtPeL4hcb9R8jHWUWsiK
P74GvRgJes73J162Hc81YH2BPqD3z8lsjMGCdWnL0lAHvk4VEyBQWi1FwQvYscTz
bfpHN8/WrVlLpy983u2mpenhsKNer74qBcCFaZfCmwUE2Km0WZV6LaSYFgbXtdk/
QN5weYnIGBhknUDH+zSxM+RcvAJjLJDujZZvLFJLDeA3h/V4hFmTxxx3Kr2aOVQH
ywn3kLQJJrk0bAYV7FjWEdWhTDKaD581Ve5VbwEdYrbUzBVABgtPPHgyV7yvdvGe
6kdvNU2welQz+hg9IqA6ZhWdkP96hBhuFXc1aZF4a48idGXbrSKN/qgmy07JNKL2
rImkBG0flUWIqr64pAU2u+PhY2EtcuhSnRlho7+zskxKNVdPXrpu/jy1YT0ky0lz
j62V4henQGHfyAnlEcyMqArXhX6+ZVpLk2KpDpcHR/Ckt+qsN48PIXsW2I7Ybc0b
8FBp3IOaJPausZ87X664aLGU4iElfrhY4zq2DO80HMFTFW2F1PAIOCALxMxeaj2A
i3O6THd29XKDyMDzxD0AzdGL4uPznoQ+4o3R5O9ixQ06RiTsrkk5xov51iYCTyTr
Ut6c8vWLMJ1L6HPuRxfepscQq2SaM/G9tO+IVrefxfi6boCT7VVqmuy3nvK9/U0H
7090lmHJ1cHiY6BEGmwVH0/Xf+vk0tXlliuvAWfbv8sW2YWGVRG9ZYN1/JTXaliy
o86mgNYrHbD8w2KToe7lmk7GRRTh5XZGar8AfzDvM7UQxkNf8nSeGOrv8ymdwzpP
ivrJYch0ftn3LNRXm4NX7PkmI4bfilkp1EexAInZjXQ=
`pragma protect end_protected
