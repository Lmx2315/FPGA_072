// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:32:45 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
X4h2d5ljsKXnQwlvoBeq6BjDQ2vRcpRuqSCm7EZ2XbnATOmNWGng1EEDnArHxt3I
pWOe18E/qgkOK/DeZ3mwWRWyZJ/sVGJrktmFG1bBePrUAR8LW8d0lvGFGK/B2fa3
P6wre/Hs5mhFsWKjk6Gd91vAjGHpVCCm+ckwnPmsF8M=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5280)
e/H0hWTG2ZEUv7v25XHP/Yv4S910WvEsYZGbku4+GHChFT0cn9NaKviebtC5Je2M
zUqVEBZbYqRkNDkICkmLQtQB/yux44dYfw65CGYpBh8B4NUNaw8lNaEZaGb+m4M/
+iOoCdTCI1uAuymypdEOJcH6XuHu2yeX56heYEOPKBhypKPrLjyCjQg920ClcNv2
gFQISGxgSIrVjQqQM+oXDzC8HyuOrR4RdHx2afTV6das5z5gGdXX4GcdBbRHOIqh
b74bSbWZhfdG9cRAk3vyEJEnPXPo+Z1Re3R0NKXPdmroK8zMCSWR2PL7jVhE0vOt
q4GmLlvV2sl1rayGNHK+SUnAKYN8D+6C/fjebNBF+eUCpfNOSS3N7yk7ssgL9rHE
5wBXxQrIejT54oyyzb4LvDo5hXKP7OlKYHIweDkhV9eh155PdcR3MZO0XS2sxF1u
iFJXppRwZ4nTZCQLCeYajdAc022lXyEsnwOiPk4BNxIQon9TnhwtBoQ88P/Bp2VB
W3GSRIUn7aWD+UTBZ1uraee3afNURZ6PdfWZ89yp2pIaE7tC21k7w0IEiu5upksT
xgoF7QHx7OZmOs537p8OescC5o19rNdMvVs6AaTPMqzew01B4DdZSYwbCqUFzZwV
6sUpWFYI5smrCRMzzjxeRbeO01+5zdjB33gDkqjxT6AfyM9o9jL3svef7fJ3ekmh
o7uIrXpjmeqT5I36sD4BxIgimEOssk7qfv140KDRgtveBliVr4sY825dw5rJXy3b
nWYYFXIN8cDLB3oss0gFGNI1hDyVQhGxnWzUFFsa9KT5SWbg9HNLqyZhmNoAEM5M
HYIQy3v7/vtR5tslu2dR4dH+uIo3QIPdLVI6gm+SbCo8L8TaPxdIgvmB27QireXk
l1uvEvBqDz3nm8leCOjNHO22kaNLOdmhX66iC1wNs4gcHsyOLQau9iPVvneVw6gO
HP1Iz1+vuctkTVwRXW1GV+edntBzTvqHA8nwug4mDi6cs02xzXe+IBUfNxlCYZQ0
ErSnbPG3giZbrFR2FyAsD5WROUF5DhziCyKs8FQRneXP6DZGKfXGDngxhinkovQT
uxClSna0F9igUvfD+54c7/Y5scNXsm7QGba+cIvrBbmOs5q3VshS6tfDyaOdLrDu
lrWG1WfYRoAf7LbcvrF3smmantYcqhDXehc6tvV362huSDr350uWIlvWsmXhQw0n
/T0G15rtiAIe2pVPwqy0dzvqHDFRQJWXhLpep3BnhvqT6mqwDMIZVJDWf5NElsWm
eyNEUCc/DgyEDVpwtv2Cvza3doY8zri7o7FJDLWjN33TCrznd/tbyht2lMbtt3wJ
4zkp0pn5zbr38MR4Xuj6iF18Zu/pprQKiSbddzFGkn9DhrtVeo50hx0dJRCztKcQ
WsynpPXL9MOMg4J70IHA+EFN8BdqUMABFUpfjZW7XSyOE3zLH3OTjrpDCeEjgKn8
NNSO8VDQ/hddu9spBr36sFkibJeXgH9jSf6bkMLZqxhqQYOPRVxXAgBBHR4rIz8K
mvCv29BjY8M2nV5h/R1mLNLhsZVOg/VtB5CO8Cd1IBy419d9XM8K8K8B+jYkTnSu
HXy+izEPIut6RYdmqTqBqsLnhvQeTvc6+kyy/lUEI8J0pvrM6ClKvmY23uJCHH9M
xPmH3n98WMkR+vWgA1TbHYhi96iwrc3+GVBq/xFq3ohqRQjWx24Fl1BUubzBJxJP
WSuPBBIUpDJvmOFkon+NVx1sF+q903yk7Dhu1yXndT7bkZCOuy0fCBKCnph1LHbT
3SR/5jrX7BWPZAon3D1OzIMDRpbezGZFqN0afFryiY8FbaUhUNbM61cj+Y+SOU5e
L+EqQPTTKUO93ovyjCBgLhfBUqOvXzw8n+hFjzrbrilW7S7njYPUQvxjiqlX0ivf
ZYdAwLxneMeUo/xQNdeTojMnGfU9gyW+q0f0uQtEEsHLDqPYdd7zezxgGHszct2e
HU3Y+juCFRLNbzbyoFvEkBU34TROuttbiLeOmqrnl2wGVKTe4TLNILcztJcHM01I
1tj5a13kvNt1MumVJx0yed4aGUXH2IOdqrW0vKK1adYTidbFtYJzi+qgtw02etyn
h6IcwvLETGQ0pe+dBppu2KB8l9Ty+C/FB/0G2Xbw60iQs9ybo/qjki5k2yOKKCdJ
QJ/miEA1bn7fU4DSY8GHwNDAYMb9o1YyoBZL9Anota0I0QVDkWtc3pyk/2IuYmE/
DTvuvcWSva8uUO5XyLH/x2yLhglCg8kkBpCODw2gEczSqAJ2JUNilPPQ0Bmb6BnN
Nnbx3jXoP1PTgn3ZDtiFh/3MaAeX5tlbseJLf22ECrqhJFr1dJjOCeNzr2CcMDFg
NSkjX5HnC6PbCCcJS65X+Wpe0g0JYHoNLx63Ca8AkW8+06LIobboUNuVUWsD1DSi
hWMc7fbwv/9F2BcQV7Dw4srACaf1wkHwdtYM4Kb4ur6bonBK2/azuKmq4AfMBP7j
ntZV8G/rfOpzYODxA4yK/5rW72sxPXf3ci9as/OPcRklds+7zqq5CEyXxWme9cIH
uqW3pbfetUNU9wUpm6rg4Hun9s3TF0jNpjSMXhfndgpHyGxFKY+vymOpyyS42X+N
VaJ6CFl+CNv2urs48he9ldA8S0BbzE/7hvUeEq/OV8HChC8564TtOmayRpODf+/g
Shuaq03baCgpR6dg8K9MPChcrmMQXCydbk5wnJR9YT30kvblYZA+9HacxyMmX/wR
RdW+BTEQlLGvDnOTfNL6XGqviANxS1ECHoMkFrYiXGUWB5YzYc5Fi30d+RVzAKft
m5UHY7gVj/l+f09EJF5iYMXcdm6kUEWIUbshCOa6jrRwS+b6P8b/h6NzojKZGlDn
zFzNEvVrmWR2Iq0SHXMHF+swnvrpvEoGzc7MJEUZBq6aTN2OVk6kxS/7XhZaBIS0
Vn240mff5//YoHVzc5rSES1vIYl3VqvB5IaChwFX9xavcwUCWTZbOesNxP8EshAH
etYnXx47PN3zQIRRBsrQK7rIf6bizOK84OhpNEG9E3juYYtpuv0+CYyZGyPwi+zs
0pPX3eUlvkBqJI5CRup1ruJeQ/2ieB13h7VWivFOu1z7YEex/BtWB+8pzDdxBCWR
E0KdEPHNDnxm/+j6d/+fAWGUZiAB9t5Ls9hr/KGz6FeJpdyxyIfNRONMfpfSqbze
FxbdHgg1wVTeSQ08RMTm99iXwaziV5ywMsvl9zNk3hXZzsne0auATbUOCslcSbhI
OZFZf/5gBUP0yuSBwE1LtDDl7fdCdxXJFOcEFCg1uZtJ93Jofu+WXEzEizVS0WUf
lkiGh3WN6Z3xXtL6Yx4vfZpfOAl2/KPJ4XIw9dJ6+2P1IVoVGimonuktT2z7z6EV
J7OqatUY4y6faO0+VNivWo5atIP3vtl4jGH6KxBl3NwaJ08dBVSJwXQGshOxe8rP
+q6BiRWDop9VeVmUbkX0Uhvp/QOEYViwA8BR9Wmjc3e3bkg0VVZ9hdOaPcnrDmXM
NkHQZ7nDJt43v2FIFW46VZJDpWnngFZV+Rqvp9pvnktfk7xZ9kQ7eexXd1rSIt4K
Cbw3ifojiUDNXwRIfw/S0o0KZVWW9UlebuQy3BG11LyROnFslf+usrdhmkb3mZSw
YLcB8C4NTRZ4v5o+EOEjVd5i07LldtRaHeFY/pS4x0+5s3xKbJZ8kEp4h2PjeaS/
cEQDu0iH7M1FtCYJEGB+biwxA3HlLParmlps7nOj7CncdCUiwSgykUrB8xa/16kO
zznSxM6a20bqJUUrDIj6xzNpEKg8rCThXkYFRxy7+DzzOI1mwwAZR49NLyP1IASw
LMAG0c6dyb6RO+vZivIb1q6ZIeEirB4cKTiu0zTD0foU45NI9poGX4PV+KXTsGeR
/xG/crd+iw6YV2aRfrlC/MRcKxn8h57mxD7FB9s+Qp8JznsfTMnqzVtUt4HpRWUu
Y9YFH6WVr5abDBgxyrIwQNmSxzSX2EcILAAL3SOk3b7K5uKTLb/ENSFfByEJEC8y
eJLf5Qe9reLwKs4RQg4mRJedlqTMKjrRyPO43TVMcurYp7ogbtSdxtnn8Ow/Qxc8
33+l5BSuIDz2KXfnEDUjw+cH/RwkmaFAhWwjEOW8p7kLaIcia/S1aHsSr4nRFX7R
TW8vBnxbqtpICwJZREOqA9Bf8afi7XWqqtF7BmuzVabhEjhrZ7EP925lLjm7juH0
8fIAqCOwPVuvQgAsdNSu5TWKGx87g1Obvj/P87E8Fh5nD2x9RKTir/X9l7Bh7QC1
v4tBoc++gr8sfMJfNOp4ochRRA0alrZHwT5IwKmKg9J3QQWzQJXFGYSw4YJl7VTa
43MKtIMEx6pOOgruJypYpTVdL+/hdcf8WR1pcX1nlpWNjRnW5n0r9uSX6eKtBZTF
ZUpp/hWy5NSXozkTsOGAtxwMc22/qVDrnZP73I5pE2XQlFnwbDLCrfIL0FWCPWSF
M8ErrOphs1M0sC7mWXSe78W6QEfoC+pASjMo0IbIALhqSep5oVZwYSrz//eEsY88
r79BBhog0FbYTo3dk9DPSZb5Zo29qEvXO91PpF6DtGa0U5yfIq8+Ss+0358H0nHp
Fe23531WItj/OwBQZ6RA2/+ivAhDlBzYVLUaVO7lpa/WvzbXMLkHG8t3u/2nO5IX
+LiCb7e1R6ijNEmrDh2sRpL1biB6K3cfRX33DIwBrMCJMOyRCwL7Kr4NT3HkTl7x
V6cWqM+lu3MZXwTLhk9gUcPXAV06n/hAT4mfRIJIdD7VGZeduES6HF09gzFePgaF
g0DRWmKbnw3SAUUQXvzHw6C4rVu2wBqjUd0fbt/LgqCB8UcXsDc+4Y8uZTGhmBCZ
mqlFsK244fsaWU/iyCCHyGU8hnfp4b64K/xzNurVtssj2E2sWV5ol5LAZd2GEXMl
cn+V+ghu4ioDw2ZImTBc9pmoD7ESG5vrKJy9OBVoJ6C2BTUTX3YR6na4+/rnu1ch
8GgNXt7RHQMgzYiXaLpOcPqfJLnhOOY0fddeHv8UEoJ+0ljFOQfeJsjWgIDKf70b
eTMH32y0kSqorQa0jI2IEntjLaszp6LQxAlBqNPiUxpdtwNUBI8k+y/s7p/7EysP
SEELaY3jWYvLxrsOSKkOEeo0ypOPwUoX1sXtPz9kMrvAejCCvi8unmJUzauj0BgX
z/auHXS0G0QBmSwjulkMKS8nUwteHtJkMPZeP6jfzSA2xQqOp+0XGT3t5Q/PX9Vj
h6jnI1OXQ2vJAgOQXioWYayWxc11kzSRkgAKeEZX0xQhESVWo+w+c9gLehONv15G
jjU2SvB35EJ4Po49UuxBCNGla5DydcSXNPjc5FfzxQSr1i6vBVasLfxStQnkI7GK
KitYN1zZ5+/Hef+zKVym7kpRLzFdos9s9Fa1sxsLzUnU9f7xxWoRoQSSOGffnCZA
1kZC0SVgFFGG+0D7hpbh5sHiDTDu+CKctd1olMwdYPZrLAQ7SVloIAV9cW8c/nM6
uKljWo7MRQdB710HanTgW5+FqaxmjF+pMuou7hLsWcY2ARc1C2lQPx8vNMXErPZD
M985PRuXYJgpprLZHSsb8u9OD8xyhN7V0OwvHXLRfBLTB00T+KYMSIPOJZWT1USz
K+koB2P/wcEbU0WSB9sAn4nTloB2GTxKmind74FF12wy5VSPbj8a3RdUPEh6ALcO
slyI7XdGuhG5YYkErRRKfOfMJAiel5+zvux4zLba0cah5qsPq9tnBvy5CIuagu8I
FFMI+ueg27wil/Y29b5taGc7AcykuPXA3lvpANwqjRCQVP58LIZqhEOlwErR6qMe
cfM6H+SpGakrUjHhUh3WZSV5BZiqgXpcji1zRR4PUjFyOqnFhoVG/TEbqqfuddu1
6YKLUBOGChTDRD3HnTzDz/sFM+vDgd0ziGjajvb6UmH2wdQjFdZQ6SplYJ59VmAK
IBBV+3cERkcuu3Wd2twUM5QYyZ4ikFjNxv2xR7Dn9S3s7IY0PM1GYxdSJN8Futyq
ZsWUzlgkgMw+roDuNhoD0Yr8XlA1+MFVHH9Xaoe0quAOAopxTae658ieS4AFHWz/
x0q4wWMVKs9CNDYgzX/kNXpFRfdAoIu80YyM/OEXQM95fERm4TRKHcdr2FKTX1/l
KvT6cJ4dUh6S/O36IbyFstxo7lyDO3ARUN1KfLHU52gDG3RDdgye3suUTdeSIYjN
xqHZPcpzVBTl8Fs86E6oPC8eP0EPutDDBGLGuMlyyuQHLj1hyHzu4xOzTuuHf8QD
jTyXo7vzsJWZ8CIrxzQr3vgiSTHSRkxSuqs1QhfgCFcz5ZQd3vAZlPHb/VLa3VeH
DBOi1ylxVy5J3wruqEPwevgh1fVXlLMQA+0rkXUJsZBRd7zi1vmb/Qm2I9vppBna
LiF6xNwS9E25PUTY7aVaVsc5QpXNQyhZ7SN0wWNEp8yZffbiedUHC2sCFybK9s5k
X6aZ1TX0R2kGRr8GCDdzKEB70kh943TaMXXOOXnP6cJwdmAgk1TAwjJxfcqgbDX1
mLvM5ShGIvaR21SbmP+detYqzIJOaX9bY9Vgp2xTYJnuZCFOTlfW2aqYbzv3aUnw
Vlco0xzpx7pQPNVFspoLxkiRswP0+ZQQlORaavUD9fLYXynaxbKkKbDOoFyxMV6C
o7AJmTpSm6UEKUr6bthnMNIlsLm0UBjEujpysqitU3NEGB4n+Ba8JjmFIh39SOZ1
z/vMVWdn9iCggSTVIS8/S0lpOJnGIpGSuQCPqC8FOJInh4dkds9RhpwC+rNvzppG
8PlzV3qJmqbIXGJYzJxU2wQs8E6BiBnxOwZLME+74KLsph+5ZJfaM/jM2n2mz+Uk
W/C1Q9BbB/BL9atigBKp6Hxa7XPoHb1Lsuudj5GoJjUosyZit7OSnui43Y6+sDAS
Wf2ptgAPJsgNLsBm39nmHchHu1ZcpCvZGKGzJhtB5uPCEr4JblNEwejaL6WB6jeZ
wYB/kAUY1yu4ZKh5LsqbzfyaUBse12+YDN+30xtZ1hnowz9jt1Obtm27tJRNexPj
`pragma protect end_protected
