// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:36:51 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
s79q88HTzKX6Jb6ZUCGvYZKDTEX1heZgb12tBdjjdmZRTIqn2XzOpq7l/Q5I7e+a
uY1+wdQhRELz0QH1mMYppAcSWY8n8lVy1TY5nALb3BJMgXlmjPDsYkDbXwJC/zNi
ROfR+auBK4wGo5HkfdLcKNi+eHfw2KoLq0C4JpZ/Vuc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7216)
zvRalmsdTs4SmwPdenbXEgzm+jdtszbCQwXiZzpNIwPmkREuTVTLqdgjOTnwi3JM
eiuwE/01zZqQbierp/EB5YpZsBzl7wlMlWrrGXfeJBa5Y0BqGBnvRJknv1bNMjtI
ErULWeJGOsQH0wjuCVHxfsCEJER0ClIyyTvaRbZo/vUezZpVoMiw54+svMZkYH9s
gIWjPr7EgFPBUO8UprFgH4qvj4/OW0L8bMe9kb1lwBs6XZW6QYROvkj95oJDWU6u
w255P77GqsmJC6t/v9h6T+8Ct9QRzQiLzIu21CX5BrVH/I0EP78sw+1DtNL/zRS7
mh7PXcrLL9wIAruzTtkSb1AShlr+cyuySDDcFr2nppnQ89ujI7I6aiWjig+hAs6X
2+wJQFJH64wKLG23mZ+VGF/zNMD0lGkStql5vcWFk14a0j1A2GIwdEFCdmlxPdKu
t+Q2DdsQrCkKC6mggXbRG07UEdoDmdLa9F1K3nNqWFJ2FuPBIqothdMFui372oYA
gfg672yYHgzFlbWBscGAt3F4zYIksBPeNYq6zJOxnrl3fpkYoy1Y2CGMk3HdiPuA
beKbYEome/aDB5LzEvYRXwrKGMoVbzF+Zs8k9ASvGUaNXSPHvxdWUMDzK2o+DWlO
tRpfvaYvZgnYsz81S2Q73lH2hi9VnvaHPYktFuwQd5UR7/R09aUMzhsOhgTRqNm3
D4ZwIgTPRplAk3E72qAqC1V86bO5LIiHF5WN/N1WUBcy8os2w3kJefmms33Tjs0m
pRQ+9B5V4RNF7baOesBWSBPNH+5YmKi68rfLF2yjYvyakMVuMyu2Ih3y4R0jEPpu
C4ZkvI4KRbjV1i/v6j2iqFI+sJ+bzsz0dqEhXCpUBOFe/L2T0GX3vswXQRH27pp7
oninY+OayOBamGifNtEkLubE6YfFFi/FFh98IxXMHmdN6ObCyJgK7ruQJpLxJmjH
VecEuw6Y1EIKs8NFDXzs7ptngAM91Zc9zJAjAwM4A3tt9IuNUBMPBlqxC39+rFZL
oaBTz+HKQnR5k1p3NLDcRxDxY7NbQ+wkqxHBSGD9he7UxM9O7rYLGt+PPLU1N2Uc
fG+EDfDjBD1lsmC2XCyoGyEeYGY8/o9/OLKNab5C312qAWcrg20Dhwf5YCnVXuK/
WAbvQwGeT6DlKfNmHLutdfES+dyjAJZ82ZdHy6RqNjGYHDegjbpPYqrXmOjcTWA1
YpchDOLQbb/tnnF+tCF+WiaJzgu21eK4ikVuPQKMKShbcEGlTcj6NLattAHEoFaj
dMID9ImfX6/I+u2ELHfkmLozGMgXi0uk4aCELsOW2O/Dzei4fcy8tNYgOrwJLng8
4DASnmkYCW2g1sVxa8CfXfsptuUezpnv/mhvJTtxiT1ar688MHQNAdrEJ7FLj9uq
6ZEyQGxJWStVTZxWGheySscSpYNNEWPA/sfRBiXtHc+ylJdneFmFrcC/KvA7cRP1
iC3qEodqxLG4KekNMNJGeDoP486RAJMVfbk7xF8CAFv9zWtQfzrGhl3dNJISzgIS
7sDkrW16ewrMcpXRzTA4KDRmx1z5vHmDawxVnkLjWw7wzyc7C89diWVGdPjYyrL0
I3dgcnd5i2blY0iHlwb6f0BmFW+CIzzYAimKyWuMU29JBK9MUjo3bc8TA/L7Ag7u
uW8c10GTMjsKt6wcuOfTKUQ5rABHRaRV7EMAopw5OSstYLsM0FBdL/oFPyQTnbDA
Vn3QSt3S5sLypbnEz1R7sXk5DzlS+A8Y5awZUlxP35hBwF3vShXyaKTwplDaV0EP
yUY6a60UY99LISfBc4gHH3qY7hHBHt2o1IN8YPSHO/pJgJwjosnXwPZ4GaLwFZ88
tOy9lom8TFZGIA1bDq5UX/4C/bh+UHJ7KCyaB8vWiUw0oykBn1gms4Sn48MTzhY+
8c5usx4dC0W0OJ1Z3be8yrA7nLI8zZG2RVeLF+SdJFdE26hD6V9LiuWX//Q7xVQn
4gypU1hbLEFYsG1h8wdkfSb7rEfBSN/2m4h8pvrEoSdH7Sxdwug3ZrRrCFtTC+Ny
hMZwfDUoReHldBPNovlwsUahn7LnK9NYesU0RZcwlahatsAWcyob9ps/btW+bd7y
zlgvVfVNStYmv05U5xLfHHF/6ApMDPmIAI9aWXMzfry5j4HfQG0uM1N1lbOvrXxX
cQOqIXR4jiSq8ZIAtUluHi+1UK0Zt5RTlTFdAYf+NCWUzuxITNqyijQdwOYAEOoO
/hHkZp782X9Zr1Lz7ssRS43wYYsIR/s80UUR2Fru+Lcmlt6ykTMyKKrX1WamloyS
qSTpSW2cl/sIrIlp2k7It5b7HTHUmsAGNByUqnnNChl70wbagbhb/T7E1HCP0U50
2LbiWMt+lIfcosIncssKphJbxns3+i1NZd57z/7j/D87E6LUPLxwXA5PpnWe62sh
W6jipYHtbYbD7ufIEmCPC0AQ5vtITuWxmtkpeIvq7LMVbbZl6f+ipq38XPsDrl8U
fmIeXDjySoIgiur0/vHPsaYsT3OvZMr74rix4/MBYrLKxrHpy9gYtOAPcrHwbgoe
a8dVohFHk4J55Ok7xABcwxOkcASOvnWoiGYl17bN3s0Imtw9P7a94xYrrEj+i8G2
w/q812XBFPU2XSkr47x2Gy5T+MVWfV8t6FGh+hfuA2IvOGGR2+GqKwDg9q85cd9o
tVhdrIMu7LSrYEE0e0iU2IEoUl3MSD3+chzzmiVZo865188Omc0l2+EH+eVSDw3r
kVyZfjVvdEGKKKDl9dJjyEH0Fqc/HmJI40RXeO8uGDwqF7O7dyeJr0SfQHa5Dy/4
vp8Lf80PFkMhcMwJsQXmcMjXan+rE0VfWArJ8EegcsmQ0LNoF+htw13/Vdsw7gpI
ZRaMJ2J4OGHi9YTxWnexh9VeMMEhXIgFYNXZzUuWamBhDT3+XZFNddHOn4up6IEL
CvyJaKWtL08TAQ/ZlAttYXADnQDVisq0e042ttZ/xqzhH2XAOJScsN2ZPj16jEv6
TSDMctxEd4kdCIhC13QwPNjHhXYxri0Z3emKYr3Ho1bPlxQjAuGU6buzrA6WQAID
u5vtn7QnFHrXJgVUFzaftuLqC5snS7cvEEp6+eba+kY+3h8Mw3i3HoVSPVXmh1jV
Qe1mRGcxISFJnaLIb3b+rMHABvrZt5e3VETBBUTIPGoeE8FFJjFsK3VhLP4avrkD
ppG6HD1r8RQKDIBXgI1i2KiumsBH4T2Pd05rkNqkLivV+u5Ty2O7mDkSMg/KtAtr
u4ovcweJgErsvhGICmfo5YMRvfCQPHwE5HmQKCH5cpn5md9RHtxmQf8gru8GJ5tz
vWQjfbh6TVAj/5HQFSSB7xKeYAXCxC3vCKeMOSiHEb4eG74w2Yt/B/eAxFIGVkYU
jQXcysB2K6q60il2qphgY9olevGk3zgiAW+TxaHQIHUza8OSanqcs3tafa6K8Iqy
C+HmjDB5NYIT6CxjkPw2MMSJMrp2UBgkfcEuoon/A0+O5Dr9MT/AHy/qFYU2mnEc
ZN0xeoXn9mXio9UUyqZkbz2WBIp7Jn1YWvr78kGikkEO8FT3gZeRpmu4UvQFTqBo
B3kdh5Xq4ATgfC/cFAqeasZ8pCfO9Zm311yBezTqF4aYWWODN0BbldHA/Lv00SZg
qs2ja0SWRWq5KCN79+zGn+RbykLIRg5nnTFM9fY4LThN6gTJEQy5L2WYaZDkyrGV
TUSCEDsDBgjExZgCx84NHOA/2+d96D65NTIaUIZDh0D/WZO/f4LZmV5CJRFcTwzK
VUGtehuLU6Ws84iHinW24PrFXt5dTvdetNavJlVQPmVFAgXF7W/wkbzTi8203OyO
EWoPOhpWmvDij5Q3ie+Npq85Iq9VLz+wRj+ME4RnwMUAhZnRAI3nRSg2SzX+x14p
ZW9vlLwXt518BrtrUDGNvdRbsQxsDylitP1Phwq//7U6e2neIpQEludxyfKvoMvR
ltV8jz7amUpUGFGwWI5VTRZEjrJUc/N22kKmakwhoDmcioYs16hs4j+hMRXYTJ5m
YDoeba46mi6j2wN4Iqu4TNuwTbVrZUXU0iGQsqKs8NuI6f0diBuQCwlXqgTjh6Tv
cjSajyXUZQSCokCME/Q7H1dQULsvFnJ8vQ9zjb8axQXJAhhR65HKYwlIw+IOarx5
LuAc9f0z4iuFzb6MKDrStA+omhlRFiabwaZ2Kj4MmSScUdQksznXFqxRpIUVU7yu
mYtT9xF54SwFrlF9vYQNSBVi/BIPssyQ4dweoumuqHVA0rUR6HpSB29BEQGdzaPO
2JU2Y4wKmM7HtbvmzjLEQHSsiZ1Q9wp8/YkWceVZ68ogPAL5k0JvHm0/tw8R45Md
TrUm9tKLATH1xPrgXXWym5dGJbxVR3760HsWFTHyIYYrDuJYaRoBt6dl9ArEEDkk
6DwRvWbDZiywb5zY/H8FDgLHFXxvTnvzMlJdnIuRSvwpAVPPYgvn2F9uPAT2JT3D
sXFhMm6xIe7t21PBQz+hSoPERYnjxTzJK+L022CogvHPsJo9embbDqiri+sXUR3/
TMYEimfP2sLIO6BDoZLBMPyrr9EzM/2Td5AJ3Z3VeOLYKcmjqXduIPzRDvgj425Z
0XG92OAbjBH31EgC6lrj19koWm4ltTi49/yPkuAx+V4ENs57xc8EQHvfTdEYzU1i
vAwHe24CJxRG4dZWGhJLq54v5kJEJCP0nidvpUIU9QbKXotx0zqU8ReEQye1v44q
ljyBV8Rkcc54IUr3eLdvyZ/FzV+gpAZEodXLz2eid5w9wbyl+RVGYoHHVr74Q7+2
X9ZCBJr64LdabKGx3tG3J3NTnhGWmqcOjKrjSEMfxCSeLkyyklNkpUe26Zhr4AcN
8LmW85IpOhmm05f8sXtD9JEaAszsyofk+AUOhGOMFCwW3cYCs1C1/5+GZVo8zLed
EgMjtpyHm2T5oD8sFc+8RZYmKD9b3IN+/O4Tc0wsR3Z2/7urFFvHhFO7GPyWTd85
KvKc+N+3vLoo3IKXM8SjpLZhK3O6D+v4ovaKaQOWPBntCkZxwhmougWJYboFdNLH
yapNpuedm3z8aPYzK+LU5ao2I11gGxbzXNGfnG0akZn9YSHZLMqe/qxkohEr4Afh
GImp0KqgvMPIlMvNMQd8SjIBwwQTLjpKcCZI2Ye5I72oop+W6m9SjaPcqlX1YHYb
fLLq/6eRohrIvZBcL55lnSqCzydVp9EzUvUbpGij2xkzzJtNuDjbKIe1wHMeoB3V
tmdkCKOSESd/Ou9h2z/O626D8Mk5wcRWw6GIPAwEQFsDusvMrKEGV2pLQR6RScxL
2H86UA9NtXogKbodhm0rEuHnzW+ZHvxRCBJhfc8eUPMLokxmaWAlpjacuVfkYb1I
fLVLHjJDQtaXyVxjNv1a97r7eEXCBLGo3tHrPKT7sT/RYLGyQTrH5gXUIl43Pelj
FxydP9VRgh39CgJ7LrnLeOoZOlmPp3vM14VToLYeDRpa/28frc8SyolOfgjCTsHL
Vzb8GJBqYTpiHYULz7ti0BTEhPA6Dl3PcZ76I4G4OsBlNfOycp99XOFJ2sKZHbU5
yvA9JFVht2NInI5o31Y6iDVWP6s8JSp9ymne3PzkEc5L+PObhoRt3Gjv52EYXKW8
+LyUhe6ZZdFfq+QATGqA6Rn16NqOZ11MakyIJQYQ6NYY1v7zHC3W993RpAZVbkVA
puRrl2J6w3C+TtCWCSuI/yZVioELkYDJv0K8MwrCDnvkojF3k3GOf95AEj4REnFe
nrxPMP5w/ej8PLBFNGidGutBhiJdiTSAYS9TYEjWcNqS1Umz4qLZcaBazr+0q3Lc
RFz4uX52YQmsTS3awxMlf0f0w/79z2k7CgPv2UfbnAwlkE/8muw4ZFxOUzYGalTf
sNk2/cRIdEoVCZZBRjGrlIj78JK4lfp7Y3Bx7cZA5k7i/uE6J7CCX6JteupZ6dV1
5kveYQpN1JThGJWtrlV9CqHaZKw1MyAVNJ+IdlLD8ECEXkxqyy983Zw9NUYeRCGV
ZbhzdJWMsp/k7PReNLPvI1W/QY+wdX98iujJgYbLuujxBt0iDwyIFdowrJ4r7w/U
lGqG+7kCOFVyr+aXZmmfctiFDF0Fi79QwbI3+SgdqOgfYUR7Z6Jc+35J1TipbBTJ
VbsSbaDmeNnRp3lE1zFBs8gIvnrSwryUn4XmSYzRb+pJ3r1Nx8I2+nttYgJvRG5z
ePeFQM3/GsZtrK1GXwA6RSVnQhFrjpLCVnMrW3H3TbG61u/qqJsCXqoyaWmDLMb4
q0I0vPnFshsXj/7CCZgrSPS3ciUwtC+7DQ205aaAxdeUR7xVJKps3y7zVlidfnZr
o+rPxNmbU+r2AWsAlb84QA4kqkOH3b+4xZMyX+p6AN9DRqA8EPy31ZA/UAKpswTN
PIT/BGDCLAod5XO9e9n4RoOz+j1zW0sTlsq1tGjNxgVtkxx3nxSyopyCGaWOfGGm
uLt7quKiWgmCoPdKyySjbSgwlZU0BHsqxsjpGtz5wcbkbI6tpeZs5lxuiLtZnqb1
qGFDR3D5tG4q7oSvU0ms/KGl1MTcSp6OmD1M5sInwTCqSZKSyqeTxKLFtrEk8fQh
YJNVBfj3yjEWrzQVyoKA/7bpOhWvwXU/uBc4kuZJbayM3BxzcBoZz5QvtPKFmmle
lcxYhpwZo2lxYXVZismms7AI2woxsvADxqu1zpz05qYxjsuOnyTMolzMZpU7PEXQ
pJD6O3EvbiKuQOsA2fhsZA86pDA0YY5ugDfWpPfHPGc/U640QGU7qJQ89W8+FBrk
8BScUvOhXpdJskZtDM1QYzL/9B58i2bxZbIbDRGsg0uZwXcaDyEgXlrfWYOMfZro
Y9aEJ3FZ2Ud7Nox61Imn1BTIWWwA2BzSMHCkDddq2OkhrzIGJ8Cq5iCPYACSga68
W1JxyOKEl3cLqRHO+7J4GJoC9b0hkiYaM5IupOzKfwEQvc1jCNCXeIlxwwCK3sIo
P/ro1HHUMl6ldHjQDtpM8VM1VQ5/Xim8Lw5SiJNOvzrZvd3lSGv26trnf7EIfWE5
dJ9guzpgfM4/M1UnrX01oQW4TmQ9buYkiuplROQOEyhs4N4e0+b6NCwDCCnyBKhM
3TMdEGw25D7fI8b3UqHXun7NWwcFDr8Lm+lXal/KCUnKcdHGNjpA9wEvbT5faWCe
ZtQQdulUkyHfB/G10LOalpV4DefqR638wEi4GTnA4Y6Sl+ygyhTi+0gLhWVLP1io
bcB216LuaeRpirgC7EOVEErrdsYqgbTfivgnIdt7JzznUBbHbB+W5r3KfJAfXtOk
ezUJn1l07u0XRpi6dkIU/iMt+LYsAOugAqp7W/j36mqa8mwt3HgRC0XMKw/eaASi
gfR2fP9rR+0e7U9kBzqPoiIOwQGLHiTszn6gUH8FdRvwcH+glQaFt+0T3ngrGgPi
MNoJpDLa32vInvwoaf+A9Cev4llDj7uJsxmKTNrUZoK3wZwhbOlnMcWwkAGeDsLf
ies60Ee37AD8x5f/CirZIjGHhf+KexJMjEGvNwR0sWvSpn1begJdP2vQZ527IMLc
LGIGiUXSHoxkYPy5ngnrTTJ2JGfsQ/s+Ww/dcak5U3ojRfICAA/RZRS6TRMN/fBI
91/QViZ7i4DBSNrX3olZS7Gmc8K7zFJssc5wcMl/1CI+IY9630gt95u9/XO+j2Cw
j/KQl3XgbR27zM9RUW1qzDbTrGwqrgqDJn0JkQkzU+amHukIqnRxK+Q+85K0cHQ3
5QxdZd73ulwO82wgmTAg1ZvUBCCvJ7FLF98ZExSr9om+Q3x6I10PXF5SpdassoAp
+ku7NMlHPaZ/C8ynf7CGhXq5lWFdU0cM4fyXYoIlhH8GcNgVlYM1LN0gHDHy4yiI
fhFmFyzmFjbI46cf++FwhpcjpyUMhjz0Uw1Q3u23bpy+/W75MELfbDpjZ3xTTw6q
KzGhGYb+EP0w5XKXZCt16shjFL1SqKtPL47NHy763/FVeWM/CKJ9nLc6hudhqUcT
Vpy/8OTOrF/gTpdPdypWvmGGqFK5rVKWwcUytdF8E9lfv1LjyuE6jlbCM/iCu4Pu
nmcg/SQMfDXJVvjaowt2LaLAYsuiRU6nNGNCt2/fcnP5JM2PPSweJTHipz40UdT7
hQ3p9Uae87NffAMRZ7HtnAfm4jiChPvqFf4NSeTn6/LBzz6I3KJvI5StrYWUzb1q
8mFTMl263urGWIXKC51+v8gGzcefUPAufHfaUvzJZd2oQCpTJVM2aMG0Vxug3owC
BAWFDZh4L3IYcMqxTtWtXbfvMZsuprIKnb42zQ3sJMGrWEd+/uGx87n2te3eD8KR
ANQLTQGbpedkq/FDQCeKGOWJ574VK+cBCQNBtIiFfUjkChDsg0J/OIMep2+avoei
kX+Bq5C/gkvC/jqwzALf5e2N69zdzOftS3xYvC0xfTL3vnl4hyfNUB7ZAbvV0XBZ
b+GvNZVBDIEeVlYObYEnRNtt0Uj/EuptIIm2nW8naqHHLvPFN0aAQzyUK1lpowzV
IkK9vMlJTMqdKtd6x0B6DhB8EQrk1ELu0KyVOQSqzBcrtoMtg8m0NfJYUgYMiLf2
Otv789VewA4NjvV5Isi4jedbJI4ihc1ibqrI7uyD+VNZimWyoS2Jxo51xfUPp1Aj
kF40S2KIpDOoaiBwfFI1k58EtNUP1ByNy/73Ur9ekXE6dX5KrREoyVAW2jB6KR3G
tX2vhGzTsPhoNuDugg9DzNhOQDhIwMwx7YRLBUJbGNiMNc9CqmLNm1VgjCYxQDIk
MBTEJ+b78pnAfbuEOJV8er6P7qMGqCJZz7HDou6urhG4Ecvu6ku+ee3SQZ8pAfor
cvN3cUTBwhEy96tgWvdMSnD0ksPm7LYlfRH11Xk/C+3xRJGfK7dcSK48hqjuWsmX
DWLOdVwIgjJD2VgxTjmkku2L9mlKdENftieH25d7nmvt+BusnAtB80YlSxKyGzPW
C95Ds3iKZRbXFfhP8Q3GCD5EnVxD1lQLl3S9LN3FK1vVk51hUQ5A7h9vdjgiWTXk
SpKQL6/mULqF/6A4sDXIBbpcVkFN/1RPids/zF4KaW+JcMJ+gRdUNBgpDppHmXop
s2HU3s9XeS9B7gPnyhWZ1aCgLPfCVwf/WhKGVsPT6WeFnSVoAInAPXxbsrqRD/Mq
utklw4xwev5koxuTpbD3ob19yCjlEzuPaI2cLLEyjTbTPsdaOafBXowEIHC/+vE2
L8K+dhpliJxl0fKVUoEsExDsjaoo/QymOO4lCJPiNeIvynPvdLB5sv/CnEeFvQJO
JbSQsHIaSaBQ9JPjuEKTEIz/qVZXcaKI5RKrb5SBJ09FNIrGKG7s1JI1lThLVpeP
oJaIs/BpQrakNPh4V3G6w3Yxa65rJ5Tj4QCDkoozch++qXpU1KPXBW3tc1cgyvDf
hN0HZ1OTVyRBmqmrkD1r9/jAzY0k8g6qu/BLj9x7yfcyw/z/2FhfgyC4zKCyyvQS
ZAmzSj6w4QeQ92cnePTzEgvcSkkoCwOijRH1NDE8/JQRfe9nBuRE+9XIKgKLKnfx
05dO1LyTeyWtWUPVcRgegRCHFut12ekgVsz18kLs99aMee/gnX/08n1gHuWvDBAL
NIakCb1VWSLVFD/2EBABWA==
`pragma protect end_protected
