// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.0std
// ALTERA_TIMESTAMP:Wed Apr 26 13:33:37 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
kmlcr86EFRkYQdg97m1CaclHIJmAypCCqgGxuV69BOTwiFkvbIachkqTqNvGyz7E
rqAQKtDz0nXz3XSBUmDO67btEQF2uF8bc4uJj87YCv04P71qFmOc2+l2Uhgk/BY2
bY7Mn/xrdkcBBUfnWDLVEX0kzsPdwkVpAQJWgdj3CQg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 22384)
oc59B5cZrCudS1Qx0xkxz3E3eL7CPjJZBdcz0ADzNISsUw1sf6busxHwKT49QP4w
CDBcxLHSzTAG/4xli7HpS4BMHNKK4M+/yKO7axrVMc/R0AAWLbHzov9VELcVBrf+
T3AnH76/L73BllCsYP4wHH7+ArJVBMniFaSKjnTYjuZ+KzOtAS9nXDMsaS7TAZKN
CLSbxZFGyvLFFiKXVvMLzmOfuWYQyt/29lFAL4BkY5czCJw8d78fjRUrDFJ2735d
tfbN+cTHPr7/I6saSB3mRXu8g6kIwozyWAeNPVftPqcCs3Hww0cdL2gzxidsvDf6
F3rY88H//DwAPZjW/pLoF5JPQjNn5UsDc5DoSvOjOzEr5DC+qH7+Q8wn2jwB5yAL
N+mLhg9l+V6Gc6WYfKvdY9ePx/g9OReI5cI+RrpPHvVMd1z8/GpNS79G6GbdIJQp
V8JfBneaUCRLvrRTyy2g/6WoWsK431CHTVhMlDLfJ5wzHGK4m9UvGViWvdBP2Lo4
GO8LVd2Vpw8OGfHCpnUu2cTiTc+Mmu2Bmfh+D7wxwgAgtcaAelNQ3/s3IfupPqZF
NgCmVYG0YtIzcLbCmXnjCgx/yPkHxHM8ld6NV5MCIg/EJG9266dIh5gYlmH4Gkq+
hhNs/xF/51KxzZdde5PgDuGC/ZaEyZ6I2rb+RH3UupdvH39kcgqteWTRd8lGDmf0
fgYWUiHWA9LNtQGr2Ik9v5PkQGcNxHCkgA93Xh7hpT8kO5HB7+tLXdmjIlK/i8kA
UbbN6NlQPMLD2CJ0pe8sfJ7iAw0uOBMcTgN3Ow/L3smWR8B+78S26+bO4wXxcM4Z
/fFsW0nafWRhongUZe9n7NFHgfdy9L4cTp9rlDItcvX5ycuqnBcK2w6QUCpF+8xx
/YhMmiotfYdcPSc849uoPgloclVK4ul1kcmHcX5MxE/uamrAgzvJoWKQNSBEVlBQ
wYVBG4P01QV4L5Um4XHpqNhUbk0x0VLQvBbVHSJ3vWuMevLYAXlMCLxj9x4KjRqe
pk96OJjrtBfxnLEaPLw1eD+HrYZ+Qakf+yFHB6WsfqaS+bMpeyWM7r4po/cmAtxg
LAUnS8NVkCJ1bjHsWG4BFoUvWyU1n/J1Uoi9th+MoBohaSkWMH9ulhbIHxRVFX+7
9yFEh5PmxdJVHehtDQ3M6TGJD7mw/tkS2BlsX6RfRYspthhAkWIr3j8i1DxZMptI
VQ7xHiJZ/rC19yN22hhgJXgrmXAnGzcsqRmWcQ3u0qu5L6gln3JfiKxzJZilmkGs
qWHT29lotL9hU762g9pKKj2t4sm/ILkK8AlMmMrAWm1yhyvTiTuJ+kjSr3VmZD4x
+BAU09IRCuSbxFQZ39yFrFvj116zpfDSIexOPkdnqxCKvWRfa4x7d30y7kRwGSnB
MVYwi+PSjfSZ6merFUXpjGpuD0XOhigISCU9aXid/PAImLWURZjMjeoXRhhmbMSm
pYN7aV/ywJLv+wbML6z84F0P89Ew9G29XrOxoZHIm7sLQJ1kfVz/lRTFyImFN5IQ
yaZSxaydC3H8HxBZak5HBN0O5oxK6E84C380dYlz9CJkUuLrpp7N//iVzDaG41yI
ecMidnjJYVcEiKAduR3bAOMv/lJieZKlmdWP0M5yvWCXdavsbWsdwFTHcRrkxF3F
or/JgjruRrUYAip43EK8nckM+Va98lmjnHWD2SPevl/b6XWMWyzhPyj7X0M8Ig/Z
54pmqQA2ecL3qVY6NqMR+PP90fXe+GgIZWL83QYHKYcQaLrwZIFfM8NEiNA6o/nJ
3PJerZp3o5d/TthIgzRL04xDFPWTh65unr4wcuPfKs1fL/DuDUCH+sZAGGwbZoMA
WqpifdzTSWkeJpyCMR5iVE8IX+nYlKBoWYr2AydUFLqguoywEgbx6KChCtKpyLpv
Nmk06aubAIhpGJDWL4CbEq/fyS0ke7Yd5mn1zJ3Gn1mGNCdCFAzQXpnRtkz1YLpj
pcMkxh0fkbg3UHPFyk98vz6305OvfWJdiO3S8tTuMfFRqw7RcBi+r8wDHnfQUjbB
DKtyM4UCWrkkjfAp1iGNFpT3mOqvmCYGpYmmJFCUHrVIMoFCINjvqoS1rB7Pp22E
XI6QZy4I3HAflJXtdCY/8aaIkwzbUbsLv5XpWjmoqAezyiR4Q/NTtioxi2/Bw+Fi
xTEvFbjQxrtbI6fcd6Z9t17pdReVsiK7XlyVvnFoNA6Vm52y1+clCntSWf46i1Mt
4bR3mfSUxoA4yPep2s0TKAYrGIJps42bIGjbZH9xze3FNPtijPLu7c1QpDp5THUs
aoE0ILS8ztp9wKJhIGzoWxsdnqOydW4pefvZcRFKL+gGcfb8pPKXWyJIXOqG4FZ4
igxdCcy3PbBpjqNpFlfcIl2cNqWHlI51Y8uiYdfBEBmqNeYcJF9NBAKoXSny/AUO
MPWvzcP9yNvD0CMo5buklmcHCCdqPdCey/MZ6qeYyRKgTropp5OnH7uky1QjVg5Y
Y+V8PRAzERKuQFUnYjeGsHdmXh8xmMj3AMyZX827gXljTSyvv3TpqnHtUn3TQ9Ls
Ig+IChp67ll0oYo9RKaBGaupp0qD1RSt6r6WMXYqgl2dnXXPkysX2Vh6vXzpc7H4
U2hZqBKY5TgCS2nMIU5rwqNbgsZ/rAtYsbIwlc28j7aILzLPXoP/lyE+kQmVbhxr
Np/N5wcRRni1re5rpi1fEG/HboHMkTczvrRjKSWk1OIe1T2o3+bTggEOSb2WfN/3
d6fZ5iYkJdnTN0ZcuiT8Um9wzruD+/aEFha/xemAfuH1y/x40QtDW7xFy8if5LZQ
Cm0oxlc+R6/yTvUj5temuwgOS6ZPvFmUOHNQY0Yr4KtrC+wTcZVaSlSed85eoonS
67mZgXEZ91/C19n78k2z+cUIfa1z20TFX3afYTpojRq79JUDNF1vuORcn4mp6mn3
//vBzAUhAHhPu5uRMbdxwPTGTwPNgyikxs/czM96nR9wMUA6Gf4rIrcAE6jMiJ15
naC/0LUzWfKtiaRyisOfoi3pjUUkkJi1NYoeddVsB3XwGkBiqcKJxdP3PxBymf72
oSD8wedHKIcuzJoWkHJHecgjz6pRADOv6VcMVzv50T899ROwy84OKjNKHIZL0oyt
EsAIf9+IR9tWaV0uSYh80jN6nBQOSzRqBCQz0f7BZB73oVPC5+zG625tT9SroumG
ajDotpzrSFXO9pRss1q/9glm/HcXKKluWOHND0fZeQ8vmXNNXnqF9kJmYWQHoICD
m122o6e7XN7zkX26/PYd5zUK6Svh5zOtLFDWbUpk9EKmkMB71K64BNTu0i7J+AGs
C3IketWWO+FgCzCK+T9KyXYRLxNLZy+O6aCn2x1NQ9p+lWnkcVpuWfur2tlcUxWL
cwxNxe92GyZzSwOZQzRLXDrvcrZf7WGy53I6urVT4w8Zrfv4ccPTxSrFiNb+44dJ
cc2AtVCGYY9ks5z0rv4ERNDp+plDRtcbWUMihS3W+zFwArqDOXI7psNxtJf1ZVJ7
F9BgDvNDtovW2xA9oGjV+fyRbrAdPI5zKeoie7drRn+yH2Eriy+NpV6XAI1o8AzN
GkNul3HtCvIKMUNIa5mtTQBCumhWcVwem68YA/lwx98Gm0P7QOIi6pWUk1JW9i4d
m+jwIMaea7mdRXzSq2hiyxY5lgcho2ArQ5MWrsP2Ui3kGxOaC4Aa6fuQ/Rnc/Ire
YYrnlyHe0aM5qxYbe7IZyIe3nrSkCLPKZPxc31PrEcbmOaueIUar/t41xNVLL1PQ
QdqKNHj/12mArQusi7alt9nD7+yiwE1YDeQqLSbHaSHD6v17kDG2r8OnjQzMwPgC
By2WN7JSCih99CDQv7HWM0bGGFTNNBmfDyNkPvHogJv78ZK/D6lUjJfMnkzva9D+
i/OuqVWp1xrpaoqgTF2rri9SJoPO6RD6f9tY93+6fhpeq84UA5yPGeOpO5Wk9OAH
kI6jgzRVBdfPASbr+D+QnxqO3acT1n6b6PhTeJVW+Zn1B6Y/UpNmIrkV63mBaurF
f3Iq+iyMx0x86BNePFdT2QtSi1v+8dbCri4oyuyZPgREjlEzMM3T2jTQ4Kxfjz+7
zBrujQCH7agki6DruofDSebU/ZG2K+lOkWwu0ay8ZrWXSCcHf/p1lmqL/6/V6fn0
BuDIED9x8y1EcNz1kt1UcM/sMIfpsgxqpTQrMRYUKjGuGV/HhRYeeVmGt2vkKDCH
+YsV1ajcm1Afnqm8uJNux18zvIg0uB4IouC0YZsoLLG7IUgtjmJPGggQfca7mXxJ
tGl37N3hzDty2dP/qer7HqKqPvzM72lj/v5iIOAlah6fD+a1HzA3zR6M93nlZCQn
KI7npmRCfPfPT2jzIlCFRD8ed7VR2PJ2eCPnAsEbSK4TRughJPYhHZVCZBtaibIH
xwkexJRh0/aC9+zGg9OEbpeRAk057ui3aZzYHV6ggIqed3ZIid1LwG90AmBQxdXh
0FnPNSarxzBDPmMaXy4wcwV8Dc4JCQJv3lskXJuxOzmp9E+5JFf2ldRRP8AxrOzl
t6FTqVClOxqhekuhQax+omftc0SVr+Wxw+s3Rg26OP5dLLD0NGkBpL+bBzdSkRgu
PMnYVaX/fgSy1spM0Rj0Gp+IsaIdm+Bbx4MjbK2vu+6dOtoe9K8Fg+ALdWEuR93/
nNBhy4AijaP4AMHQPGzu58HtIVBWocj4f78yMQH19bAqpFjJ3GF8QQW9AEMS3+D6
NhFI1Ia8l2tm7qZjUVp4kzMpvNybBlbYH/C2PnTmTKrEfSGYPFbq19f/JuOYBORQ
Tqs25BmJDkCdIYeaftGPKYA0VvvUGXyLUEYcsxVLnJFsByX7tmzlm5IlKgsfhZLE
akv0tjHyh3VlfoFfuDMze9NEr0t2IAnnMS9ZP6AlxXB9NOmqyCU6q2ZCzgWUSUa0
ELqXFVeaXbhFycrsymHQEcCAWmG4+c+YvJUw6hUTLMj2h3BXkRBIjkpBO3xCTkas
MAK5JGzgH3iAU8u9zyGrBGvoiIsuAXEsoJD9Eh7LsgIS9jKw/s5O21a1yzTVRoDa
KdIZeUuXE/sBYL28Llud2LiMHR97sy41AtgyjDrzTsIcEL7qt2zxmUKEsc1AeItc
VEJYmbSwEuI4tb+wjWLbfsdAKb5qqln5bmoxSf9DCEescBhPdJiPM0tp+vr2Yqct
PTCC+1veFFeYqe4866UxcCNX0P3VwSzgpNoqV49EskjXLrlZ4vDZZOB3PGuICLkT
photWfFYf6i0vmJUQvs3591ki5gjCXSbfs/qgkLwb/lL251mCgjiQB2bULKMA30b
EFDxKiy6auSR0yFP+TGv9ggpHEORQpyj+eFK5gswt40axiXtKtUFrX+GR6FMUL9z
a8NaUlIh+POIc3Lv2lXBfM88Vy2doTLhUy58owXjayBmtNeweLenLB4br0VP0Lki
fgYz277hM0dGhDn/Ssc05MmI3eAwVPWHrwSqFKUOAIJdTgTSJVqJIT3dqd853a88
nwSP4LoCMG6vDqhXN+vQgudhBdTdhUk9L6ogISZBPUF4Jiigwtjh+T8IwEr4lWDK
bsFH5oEXmsDaRzB4CnKa88CXNqDlhfFCZC+ExT7NZyjukWXn85lzw7U8EqaLqTOV
b34iKRH35y2/3vWn0UKS8Pdu/53rREmQYEw0ZrZisV6YcgRfg45E1n4XW2Xj7mAp
fdqXJkSohrV6YxV4+rVmPTifI9OZszJJDwaR0EA48gnAnhsq/OjRzIEAs7LbKw3T
ppcu7GEn8Xoo0TQ1m6tkwZAx8oTs9qWmSZKA3my1FtRWti1L9yFy0T2+C8aand7/
5eZf9Ixs2YfcqQX/cquh6+G3XBZvim7P2Pa/jA79RCLe6YK6GDSCeFRTkMwfdid7
n2loZPLX/F3JNMBbw2aqiunTRqtZ3QhNj8MjESovIzHzUQpOa7+jYtKACOUc1/tA
Uxir/XZMhy2WMVTbITaw29/WcWbNvB97r0pxOpaEUFk6tOq2SKol8I/FsEiQE2vF
0DGS3P/1sZuncLO2otPEqG5delGdywSepuEtDQzQya2p8xeLGGnhW/DF9ExQGXUd
cqV0s9+XENnca7J9QE2q6Ofia0RLCm7BlvFS3E3G5VpIhdO15XUJqy0hjawiikes
VZNMxXU7+Dpa8h75pvlAqIEWC0cUDbggAbAGzVHLE7RBWS9k0SQ9tQLcqNX41mz/
KgYvItfujobYHoA09jPGoEmPLgHLm1h8N5euDX6PRjTzzVZ1AXrgkH1a59eB9aDM
pcX9I1QBsfqlt6ct8LVMb7fqr+ShZgEA3Bv5KqhYHgsqSBUrhlGKckXeZ91dQteb
snuOtNsVOTd+XATZDS1j+ymiHpQZ3av+gOQrSImWfO+lGiY3kjowSpfl+B4bjLT3
2o6XfxTKBx6TOAva8XlOSSeKx63I55vKvbQyS4KqL/ciOpBHadHlH+yZ/iRhtw5E
oj90VizGrWDvWUeWe7UmzzrXjoQhrAx7C2DkAVvwUU0bBdWk0DCSeKluKNEBNzJx
bOMvjIHJiLVCPnWX0l1kOQS3v7hnbGnTBpyw/aNnY39NhenLPMX9pYym88xnR82L
aywXHc1+5t/EaAXJsg62FSIbadFah/Pyr+XDuq1PYlkOKQjiS1FptxUmstPM752G
Ugwqwh82xEi758Ctznc2Kh3n85Y/j83J/zVWKVQ8whm+S3D/8HHJd/e3pSBuqh/A
PvpvwburITP2xgQgwbmCj2wFDuA1LbKreiX5sVwhIXQ7O2Ej/+sHr6jVDQ8lhqG6
+mzelWWgHAlUeq6iCVat3ddRLsbvmNTejHxOReRUelwP9Vp2QSQPrBK+AHkC2Ucv
MWpYHS14/+trh339/Sm416CQDoyqx9wiEJ231vKj2HbA2CBFdEXkzTBGb/0tUMI1
tsqXURmt1M64gmTe+avQlyIPI3VCayVWVlMST1zoGmQMLwFl035HU+8iVq3+UWqq
N2Pu6AHzEQSuWmBrcpUs7K1z4i4CHdgektCIEx4sq2NbUGf9d/Afn2jJD4O07ApI
B9+m43Gd9PVp49MkTCJD2RpKTEOyzg/0Zg2Fks31jTWhHexe6BfAIp5J/OTs/AnU
Mx2fYfROsYXe9H1cqen+c93efJS9ZrcHP3DLFWd+zGXdUmv2Qpe8ZMCfcnuA4pL1
FHL3Uo7OQ3/Bt7ybw9b49ecx5GpNBk3hlol5uAkuVly6HawrW0q4jwvG1AsdrD6Z
JUhtPvJyCdUMQHkkVIBMnrJLq1srdawcEfV89hgC4J1PiHUfTtdg4wH0RDNeZc7X
1zuxvALklF/eNHNUKTskYzOsNlSQahLfdrNJz8CnOeu85TfXkD7/zTZmiphFNhaG
pXL9g5rurHPps8jL44eRRDBBP5ozFqVpufrtBEOwDib6KrWOQkahcGowJDWa4SIz
pTlaWSsYnlOY5t9rM6PzaUxG5v4gRYPHw2WyILMlcN7Ob/I6WZel7538QdZOHW3o
jdoSm6wtaBw/k74TjzTcT2Ln8lt2YNuv3sHHUNSMwkJYQOsOdXeAly7tdDX/eRSG
BaWRsm9unu5i6b8gkJgbYKssV9jcjVJuzodLIM4mEc5IGeLvAexXfhX5Auz+iTQp
jkzCVI3YDoM2GLMAC2ZrE/SpF9HIwUt8db2J/M47uNG44tEYDDtnPmzErLSiwD++
sYttleK/WGj7RPRYEDuJJ7sNIHlZBTO1wdR9qfiuK0pFijsJkvpK3ekvGE+Ha2d5
Ygin6bTJBh3dBXEzAmREY+q/Nu2NxkSy2L5D/aD7FyAaqZ0CW0tdKRKiKm7pRJP+
7lGezc4Fixm4yXhOwueMmkLBlivJoJUW9/63KgV+MOIdoPVyW+pC+lDgZnFydIVY
B4Zzs7j1wbfXRHzKh9yj0P7QAv4Yn+QiqTfxU+RkZ1vxWkAxZfy7EsWpajwnwkmD
HcChxE1KhdPW1mD/+tnIA4VyOlc14WmrQdnksUgRdiKIt/BYRCzfpnokLyDLDqs9
i81FxIsF+B/VrK8ZlMY4Q6rAFnxzomsHwkePlXPun2cFsXI2ICMJM7JluIQnJ2FX
/iznpg+uJG97sR0z5lcztibx/zWPjnJL0cuyrwbDi39isazvhtM9NUgeozyB47ry
w5JT2VbTJxS+2/gIAb3N0LGnfllIfW7rnEuDXp5fUWq1XsYV3LmDN8F8dbaWE5St
5+2YMLv/BfGgdtWO0eZV0J43vtekBznCekKwyC1xN9OuCmH5YCCUu7ceA0AAE17c
3bEB8gFpGph3khnG46/5dkz3VQkfXgLd5erdz0LyyMuDpE1Sj3/ws9NM6UhOqSSF
SIGDHrd167jcFraIGn9Um/l9KubfbOqy1mmXr+rzsNhQYCuWPUXQpKo7KWzZwsfe
mb4xgxrZbr0PLw4wvZ34qZIwCZriM4aXAjogNUqcpq5qBjYJLXiMQE36CEVgSrS5
Jd6616IrwQA/oM6BYRficx+M5rZKJ7pqSfwf9QJ85GWGwn3jyvrS1ZB9TXtxtuTM
oyK3QFzlMyS6XlU7bV5Cwdnlmonmimftf8TaQn9nU29Pq/lDfBKMGGbxWxhMV8HP
8HlsGmS3D0knWX3WSu5Bge7N79H7oF+p/+/u+Ds0ZI820h9QKI36K2GpokOeRNf/
05hXnAXQ9OSuw1avjwYGyWtXs2bsx3knGE67gtCb9uxuh/e78Xp7w2ZSxp9zD6tp
znyzW3Vy35h7XD9nLUPj4fZt8bi1MvA6T5KJ9lhelbBxhqiHHsrROt8j6aAROvwc
PvrKqisKAVIpg5hbLhIm2jqybRqSA/6Foz4USlfp20ZKr7/HUVAx5EvCgYYXCSRy
TLWMSkAFhQIMCXRa/RT4cm0i2h8cwTy1j0qrAFPOtuQ6DLKYcfeztweel/3dRyQQ
gASsQCv3LY6NBKrdzP4p/WkTuJpfBJT3GjIdDjiM5wYifHHT/3R0a/7K58FoM6l6
XLKp7LeGZ1AuZpsWnZO59CXlPTk0kqm+ySYV8wu2bvYFFoXS37HtXZrpVloUVWpe
5SWJcj1MlbvgJ7HfiwK5lTQ+p3fXeXUOasCbFE6fAua44ZVkOEwADoZBDLdJH4Vq
RHIoEMf4sE0IbvzuhNHorNEKQQPlfQIu3ZhqSys91H6eq2oJYBWBda+JFqwltRL4
anHRsQ0KNYYm5NBx6UKEwZ5WjAxs21Q3QStkC24VhBBk7BwwtOoRtRjf0mL2cCSY
J+/uULxPOoATN77pl4crb2XZN7dKFrsiioIZ/el+GcBEcYY+DqN6MTSfWcM8Atj/
HnAwPkK6GhJJ6eLbTNbr/9nu+ZjUKowDi6zCEKyvOVygAGAEZt/1uxxl9fQabiVp
w7xg4xIJPFFNVcPAgQSN3PETdwL3gtzPcWACc5fogzbdEIO1/Vg/yGLrX8mS/WqZ
HZEM7fQ11Q67NIbZjaWZLipgxNd2HvlvM2aJbZ8ry/B1sfolX+qf1TzKOF+NVBVW
yUc94HSyNeVl44U6TUx6/feuROEVAJtu7Nd8RAitRDblTGlsu4lDD0PeuD5dwdRB
Y12qF7WxXeegeCCAyyH13Fmm/0v1FoZoK7oySVBuwU/ql1wsZT+LlKz3pczg1wrW
KsaTg5/Xj5lwZlujuk7iX3E7/15aUkTUTUc3eWlsYbyH9LENMhK8GWnZ3QV+Na/B
yE9Q/A8E0Z7MyE+w4juvex9zmryrIdF4dlrAix7HtxH4QiiU4iubkn/R/yHTmvoE
JLDABg0Sab+XYL9IYuV2HIFwyrcpALhLmAUdtL22YOBlXmfwKho0UPieWG19GbA4
I8SrUi7wEI7F8aF9x2rnNXM7L/Y+jc11jLnX0xzP5X40wfqUBMTlT5sSSRSMy9Jo
9ACtKzKUoLjOJUz1o37DX7+k61KdJyw7HKNtCOMka8M9HLylEhl8IN7cGT/rogUt
CDJCV5yKl3tJvzaMLmj65axbQkLco5yM/M+GpSWzp/Y96K34Q93tAArHNlXCbJ2K
dpj24HeAsrdUCUObzZHqkF2ajz5QYC9Yhh1Fy7fBuLnYHWCSBjX38Gf5swNvOLW+
7bIeaT7Wc4ZOUg/wFpANOQJW/wyU70YtFXCzMNMx8jV4qTGckgClKuHn/kbCW4Gj
Dodf9CQvcjTcx2YJbljyWqblWPaJy2k8AvDA4tnm4iKlmEFBU7uyMEOecJYdKuuE
5Hh+eiqZ42T0yp5P7MDkPJ5BVTo/V/n0Rd8XgEUb8lFDnuZQ7FRuPXE2d1oR/LFA
VwF3FwK0+0LW0e9e1YVJAb7cu5D8B5Y811bv/HV7faCZ3j2NFvCoBH9Ju4xyv1Au
roGaW33Z+sktSKXrW0krrIEzp8vcYG/d9EKpLaJr5fqLBDY23asL/DMUF6KlFXT2
N0zluO+PUHGJ54BjonjiJN2j1nrmXa72ha3sOB7Ph4mZ8mDzKLCaabR9zCwEHDxP
hlVPvISmRFO52Ab/l3jNcqPGPJ6+Lf3dhs5dHxd6FXFV6cIBr5rALjy5kgjcuHC2
+a5yvcu5BZIVm1khp92jLQYQDhCRCyA4E6Av5n5WE6QsVtXrFiq2m5lSelcvZQOO
HBr7ohwSujn6XMKZGV/ZixbshF57A2qMpkWkhF+V+GSv4JZvmcdwgfJoIm/5UUvs
RC5U7FPGWr2AdRE7wiBIoFuHGG89EHPGQLC3EKchmYlk14W16wXIAl/0NR2m0pbX
91k8gK/V4UZBGoupagde5BOg/rvkdRKZXGUtMqNPvW+7a4GO6NiYA8LTTFduq3N6
4mfpBpES7hzez1+cHOFpbRLkGgksiO+GHtZkrXx3F7IzljnLh0kcXdbPAk7Xg6gu
y6U3UsDkugurVprNXAPX1MCU45b6rK1ruEFOhe9ZDosk4wQed8aDMa2g8jQMOXrg
u6INh+B/1beLFA36CkmpTckwl7AE0xLCV/fhVPO3aZQm+JyOCZ0BPAcrreqFtw0x
SJRx1iXTlpOvfcFAjt/eGUtD7wtSzJh+hGRfVkSz4LFZjbPxOgFZkj1yZ0MvjhyJ
OLlcc2WLHW34ZGopgSKgbBCULlBrS36C6+o9ytXQbNCPU7J871zKOQuZmMFORptD
7TkW1t5LZm2kIqTL882evbHNOcygywhHKr72cixtK4NCz+lcroWMxGNIeQNDDZhx
fPk7zEtJwBseEYBFLzWlnnuUdXLl8bbb6Ao6KUBdH8foPS3/MhfSQrGFkfzJS6CN
9KY/MzsGQqzBiBy6LIxxi/HWOSAWualPhkPjXEwdUbh4XB0b6F6GhV4wb5cHY/A/
DTXZov55q5HLSKg+RpgzIb1DrrOSZix3LYYAFMqCFlqrHqULSccZ3eCYj9bSwJk+
MEx8OPUw6t/zU0HQdu271S5Dtp2RBope/DRE36Fj7+Dnx0RoxhWMIzGUihlJlSYf
4zBnlBH/4d58QMePtll1gNN+NgO+K6F3fg0i73jvDFNizS+DAMaE1CIAE/EaNn7d
1YgEHSR6mtU58KOh+CYwT4Wje7pSm7r6+/Khl7wCKxjXZS20LMaFxayF8WEQmX7m
VW7dTevpWV6o3dChPaKtCSoWMnyxZ0kfldbW2f1fxmTY3xn4wWvqJbD6ehozMlOU
UBLJoisLhLzYkbQmHGnDMMda+XPXJOBtS79T7q0ZEzrLSOaT1epOuagHDT+R6ALs
IcQ+4JCj4TIIxkkMJsrFMyVbMeb4rDfR9QplW5flA2rtIhFoXHTOqzHeSSrKzp0y
P1eEG0MN194lPRFefVF/ulLW1NEUPpla+RZMn+UH+GmMwNhpZ06Tj58mjWJukPCJ
MiPC1iS2eZv3PSc/MMd/2mAfSFLnaBytFwY1gahLLJtMCODMqlww7J82V3CfG1Em
VhubiubqttmxxP2+kshJiMSFs02j4/NoknWIikI1W8YJZpYHKpaoPN9bbUpmMJbW
jOfhPveSaLNY9cyG/dqBCCpxVuPg2dLXrB+HzPPerEVA9LSJirnNqX9iraWIhZw4
h900YsXyexL6gNHLgnNfwYfPk7l6szVu7SIsBcmE8pBwFrbEhmL0FjP/1yfdDIo1
grODPn9OkGckOS9RUecDcTSzCuSLAhqv2XJPxomk3F+4jHH3DebMAaeJ2lhYDI7H
J6xQRYJrJt29KYNEMADAc00GdxCwy2NtCNwedriI7zdBBDdxNIJtJmWhpM6NwUdW
B0JIGdEA3VPZhaRj4LvVs1GLHgH1hBzNcHKw7//Sq7DBQkAfuU8dy3jLaNQ78RCg
noBZb6lc32mkBQlDUU1Z0CWonMIRX+WqMdZN2LkZYhaPD4PP5y+VcXv+HSukXL/n
ERsVeiUl1mRCpg8DBYmnM8lDIpxoUEyAVznZovONTq5Vk1Fa0H6MC3v4V6qyg7aR
edIJey7mS6Ywbdjd76MvagkhAKVtShRQRnhdblgAqOerR03iKbBHxWMEv83LHwr1
vfuu2VdpoKjEtGaki+alD0GjaprWkR9gM8tBVCRFUJCMjfr59yUPtBCqD3V4yywN
DTEOEYjUX8sq8rQlgJjQrv/sWazg44PpLv/DMSPkGw4WhaeD7ReJi6UNLEcdI7aS
ue3K2tjLIvUSuoZOaJ0u5DN0fzdoH7OUjUQYH5KZdKzv/G/crzzrbx2W8MroAMbR
QWKtBm3XZrdf0/f2jgYLmzn/PhB7lHpfUBP1VmhyUjm3jBClmMepA2a94rwWXjAq
IYfDplS8lAxQCFpv3mNPwmoAOi2BcxPhvvLwgl11/nCoDe6QGz6QE9o5sQI9uG8/
EmvvQKuVdiRTDjUEbR5UB5TGT+NQej3IRCC20v863BEpj0RwSKfPwa2OUWTvqlyl
7hZNAlTq/bT9Kq2Jgh4iP8APh6R8DbFx54x4tVuaccwnTmlLemGjZl/DQ/J6+U/V
yJfiUUqotAIsVWB5Vk7frnK3eEO6d8mlOPzUlKy7mSzVnifoZj/1N0CfoaX02BLa
5ecL/ek4DiC3oFuEHO3Ho47pJy1yei5dMEt3pyXo8WPC8iMN19w8VTu/6aP6tG7/
MD5uVy9hq74VbEiZGQJq9hr0olrda0UvQTRplySqXsFUyLa1i26gD13OxCEYAcQh
xtWR+8HTlWajpJCVPUE5rTqGCmU4Mqba5lSZDIEnqDO32Sy2dU5luKp3aSX97E6b
V5zIU4UDWkJTgxNIbRhdZVe+rcL7TY2wdh+URAj/OT5GHkSXdxsy89TaO7n5xOqs
sRzyqWZg2LFjsNqPUhPbPzOe+Jizc7DWFhhbZjRybz6De66+9fF3p8kZXvq1Wx7i
tJXm+M6EVj02UZbLUMhW69WfRUeQZJTttIg7fprTtlpBGd5rClRq5m3G/ZsHXAKA
amAFEvtv3pWBA62dUGVxogxuzWXf8AkEfIs2gsSSmFjXckW3Q0UUhxhSi6HpaVY0
LDgDSLSYCE+qSAk4Bj8FyhEXfIfpZf/RLX33ktqopnZlZVCDvnKP8vcQAEQdV9II
FO2UHGERGlblGxmT8ZsjAAxsl87RL8M7tBEKSUwK8zbRbMDTqTs6zQCp1QkKAwk6
ntXIPTOAIinxWuJaRE2jANdix35NJkrZwOQ0b9+D5m5zz8q0ggP1ixSUUfI9eArT
S/5zji/Kdy0dCfB3mcehvMjo+ZEpNIVcf+4eL2pmRUDmw/xoSiK+u30hI99CFS8H
fnbam7VUpv2wKpaGttUdvW1GWpoTuW6RyhmG195J4AJasB447O/AgQS1KsidJ6sm
EwK7FTtF3ogiMqfM7HAtqWnmImaJizsbScElZdycRcw5EQbtTCyykEMZ+7Qt52rF
dEYnhRZ7f8lBqsrLgB3pbj14tKBXkCb/AwoaP4KSAz3Qz6r410r+TjwoZHW6yp/J
YGNbQDT8W4cZgCoAwLqWWvuYOb0NXjrJmWw8ocRpc37z7RRR88ON8y4qB3PgFLSd
lxaxYchGb7eNiY6loU3XVKWd6MvixSWSQ7C2378yCqYQMrsjRmJvlknJhpHNBa/E
sW7FjbQ07skdlbbJj6kiDpkZS5kJaMMoW77m5aIOaoyrJAUHEiG2elHK0c7y6pd5
m1wobpU+7kXfhc0UmUOIe10aM4yxyL3YM0HZvl7cJPgc0BEvEUwaxRoYqAE1P7ov
cwmnaiVEM1kx7mQSLW2wwKplZ5jDi5LtxVgsU5Mgr3AIXAkQq//0FZVqKqz+F6pu
V0as56yxS0va8BPEOqT3L3P3Uk2s2oFSBVst3NRAA6o+wSgjpwrCZYsPOD1jDnnR
t98woefwjBHCi7EtueyuG8Ml7gX26T5VssyKIVhTUsFnlyNOSAajZUMH4LLSa0DI
HmDdXGgsbYxh9qPKN0hZVrDL6vqbMcz9fp++eWm0HTUTttVT+BYAl7CIY4ZIgpP+
FN5TNNj5T/+E1FAtL19VFNxYVZoud/QD1N6LLTSEkuemYxQe4orq2/8yQvfpQISM
xhXxgC2tjdw6SbSe0V05M1qx1X0UtomTymhfiTxgz4GzCTyb3ZrgZ8LrK8RsyXSd
NjTDk90OuJB4+P9flnEGCNfaODYIkHhiKXtfrrnJiOLL94kV/duUqhCFZvaxZuBN
/lCVXTABALC/Zi85S0kAv3ADguzaPI8c2n6PVT6wajXMvMkqwr0EZgLh3OVHoIe6
gW4DQq3GJ7wusfueMD66KcLFiEYgqXO3KWBc986mc3MXw0N7lGXOs9kCCUgy95JW
6Wnm8HuhcOk3Q/Inqst4IOJKE1AGgQBm1oNrsskW4EyhvfWv/APP4aiGXd5Lz3VW
pVw+27mulH4XnJSYd9XgXztHKW8q0AAPueUckBs4SWgUj38dzvSf3JPbHkyZx4yl
XAUMEIw4i3tF5WxcyLFtJqvr7lWlONmB0R8esJwWnubI110Z5pdHijHlgAz5Sepg
V/lSVHrejToFUwxMS68Ai1LpO3nqOQAB+URai9o0Pbo8QsvN1UpKT0/nn9l7Qb2j
2NAyH8JflxVQ2k+6ua2pVl+EkuQjWWc3/FEnRF0+vZZDgdBXjC9ALh9Z//L9mRJ+
3kx4EHij+br2OcCyPKHNvEGOTMbP7Zl/GXuWoevTFVam/vIevRo9ipnlK3qgpEou
NyeIxbsO+OmDYao9RwOkWKbDdjMykHwRONotLtJzATyDwtXtf6PpMZeWwSxEk7xE
HFSRleok+sW38+87TNtQ68mt3e1UtMxX1Z0xmpepECBniLCumulonP5ZdS5gZrts
3mWx7P34QqKKNb6W5L60VCaYY4HTWHqfS7yrbUVRw/Dp3+p5jEuWTwKtoVYqAzoP
dZhR5kbckRoqCEk88qRyvRjMrkGy7AfbGPOHlJ4Rc/hrOrd5blZoh25JYElvEnqj
2Vin2pP+fJl5Kl3xANJk4/hp0yQvO/EM6Sf/L2sLSLkubCScta40G1inaLHQAC53
Sig4DwjRZUaGulSEmR/nfp1j11LCqLgYFZ2mCnzBaVLDFepfJzFjrbRJfTISaJrj
h2rOts0g2tPaVhJm7xRYcutlVvmNzKbB8StmKgcNKRr+DiY3Sy0q9NqIt8gFXWko
vG2olR1rfJ6I6Wx7h3e7SxkCrCz6sMevLCi6gRtOovzh1YhYH3PfnwbTeTIZ5496
HKAMT7cOmoml8uZQDQ2QCg/jcYfP9DRs6Dz6su15OgAdxXgVshbMsTBcYrIqof/z
VE266IIw7wiUtIQiJAFDy0Zgw544cLtGp4qGhDyV01V95SbGiatv1qIPccU61uME
3JvXYZNCpxcvKM7SBE6c/kL4VH4teJegId2Y7rSHrCj2c/TJrVCjrKPyKq2XRuwc
YHgHenenwrnN03dqkVhh/SfF+60ERVi0VMXsTpR27ikMUcnz6lsz2ExqI7cczH0r
hehGcEF21Z1DwIIF5L/HRg8tEjzkDztdX7mm88OE5mui19Ja9kqyU8kRi4b2HJZX
NaG47woJstmMkQYfzMg/TuX0y/mXbi8iDE2f3cQibSH273sexr/W1JKDWRmgsrl2
EE0xJ8DuT8Gn8b00BKg0UoVC0KiTfRqAexNLi0/0rkJE2Pgy/1nYP/4tEQcU+Si9
IbS8ISlv+Xv54R2uU7uq5mPREKSIUfcxkSvvyfJRH8E7CuzMqKiiKsXsTc+/0w7D
tywPtHvMznK3I9/gie7M30EQG+LlgnwE8GUu1K9ZTVdKUFimu+yqL55dl8P8aZ3h
OUPNKKAn09bYP72C4+H3o0hQ1E73yGrZI5vEShFfCP8z+d75ce59DgSoMorszmUU
81VA1rGKVH91A8p0cEu6EGEy9TqIzqyL51Zmw/stmUpdWBMguB0ArFOS09CV2UNr
ikHbcHGyO6vx+TSrJlbtxvJPc2b4ZHVFI6TWuhu296qVpqWhOl425wYIWK0EuKzQ
23Mkqv7gdNQ6gL5ocSTUrVuDPZVtV3D+wtjL53ras08Y44PGMWb2dRwJEPJd0kTu
bR74OJ1u+h+VDAoudHZo4T2bZFmPPzymBaiqqVXMoPYlSw6oyfW2cjBdST0iNx05
M+nrcKT7kB9+M7IuLwz+0J2+arh2MaCSJoXUjf8WamX5Kt2i+ugdrVhMlFflsZBO
HsVzuIEAgrmku6JHZVSDkhN7xAnrOt9HWBthLVCqukyQnnLgGpPfq4yBJATcgoGZ
JC0Q6Ehb9AKZBmz/alp0kViT09nGnck5qDvtGCN4MrCoBYQ0vvWPT0yjsUInF0Wu
/6avj4a7b2Ghsc/4ieLuTllg01zKqhrtxN/g1XJO5F5YxdMP9AvxoDoQifQ+0b1u
Ks1inFuen3tCk/TKF54wZ3pCQHI1O8mDetaAAeyU5rqpyyyrr9dX6wYYiqCe/TYf
wrqNvqagpiuncxkfX3iMB4tt1rS9GWSFyGO/m2OyOc969MCmNqyPXmTT61Ie9Gnc
2vo7PHrgfyaCe97Pgwd4bBkBDXljjRr0Ye2w85tC4gti6+FlMUVa7A1yUOxq1mFL
vT2ASwu8zdWZ5HjEkNjO/ziT3brDQwQXQlb1uYGGvCp2FZBAzrr6x5drJx7bdbPh
FpwjJG15p6U8pL+CuZS8SRC5xM8ibTmQL7s0nqF5mC2f31d8/0zjslI6aaU4wpbF
CtJ1U5VHYZtR7s+2lonSTZSKdNdXzg6kDM0CGq04UDWDMw9EWa0srE2mbQo2wtKB
mxuJoS+5q9gWdSqVxlsZCB/H4FXtcJSFSVaHInpgKTL4riIhFutI0wbfSv8n7UZb
PTmIMphZIIPNDjSMAcfVxnMsQmEEbu1mEwmlP+30vQqfLR151d0qJl+U75Oe26c/
NBrskqzkyFwQk3N0wE+GkgfUtrBJiNkHiNr81f0ukQQylblKvisFvTBWqmNEQfVW
BBBO0DwYmrM9SZ/LtRTJ4GxUy5bLUfoIj69tVY27C+SNEebDiKPwc0KoqliL2dJ9
uANaSfQdRlkTJVbiFTMqm997y2icfQ3oWe4EIvuVsGf20cbLWGWawKHPkpGc3inc
mKq7Dww+0EXF9P/xhrn+tMNNLoqR3EDOatRLFH//G8/tLUwQUJfnhL7YuNBH3hvN
fF4t++f9diztsCvL69NfXhsaZq6e64xiMw/YRs2ZVu5ZDN4cxIMa9XXSMoppgVZA
DGzy7zifLKe23rR2c4Xs1kDlyshtvaF6lr/L/3DBIrpEe80EIcLd1yfnVKF5KGGY
9gqlIBMprCR1331bnkMy6M6fnOGlfGgGK1rxCSQ19ktnlmeyqvjrA/PedKrr+XwW
Bw/0BwlMWHVnc3G6ZuLMzVg1YxWamE65PMvP2WE6BVFwEdjjE652zm+PZj7Gespi
O01wWJ6xds9anA9Fw5FIJWM5dyuRMmUoYbNrlufLeR7FnzHQDRHjx1Siw5pYtC8o
q03oF1ffV6LiZtRpOEL21Ab9P+JtGD7Yp4OosVGtsYDFC7w6JO/9BJVl33TeUXeY
AHB3Wi6rPWK82RcZ4DinwvfskDzQ1qJgWKZXbZSb1e58Kd4Ik414kf/ciFSFO6co
dDVH58rOIe8EjfiD9FD0Q0DVlzBJ2V/AUZATgtrGGpR4I+93rm3P8Nqtoq9LaZvf
RjU+3K4jBnt0JFiqwg7V0vlKNDrdKV3UEOUI04Hb4FD125xwAZUGQ77IxVLKaC+A
g5MaDkZpWzYoV59eWu23Tf01r93VLbV5UZTzpQeQHJAqkObcOG7gN38cDuVofimB
RVJwdddzKSV/ik4iAaDzyt+oZc4YZyEz30HbKWRBY3eqVWhSdDILA0HiHdoWS7cO
DNa2DTAtn1+I1/xZSyEjleK8VSTAxqa8IWH+/3GE+1+8sfqdr0O7ibcfOI9205Wa
tdqAmw6TIlWZN8U4Sw6eR7vcYEwcEYm+RjgBPwomscAykIzUEznjAB0pJw6YkEEE
RHEYSWFQtDUuSriuKZRoimJ0POOAyNKnHBY9p79KMDYFSIyvDqFTMxVv/VdVcoUV
NbzVMzcxdgOpkUHPo6/P3eaQKvJrFfvG/Gu/cMBWhqJVjXQ4qY2T/FVxEeN/FRAb
kiPo4SEPmt/9kpcM2aseVwvqhY7BgVoOu95SX8Eq2ABrcREeYN/kyqK9V1y0oC9O
hovQ9/jEcj6gI4q2LddnVcmATlK6pbrPzOvfKTzNRdWcLZZe6CXBezJgMASVvr+m
3Th25n+wPNjWFX4e4sqC4N31R7TGtxLpV1Y30DhBTCfdN+zHu+h+IFvxtBjfBJxT
3dphOWUerKKMffsBzhu95BXweeh3ZnipjgewjY/WnI+GxWfhNTcLK8TRV0LCF7GO
T1fJv9Zefjwn+DpIPBMDEd0+uWN/obvnVyj3MG1h3cH1yiRTzOn4v1KXSRfHdExv
P0oWqCiG4KR3UuStvs81zFdrV3OFZmzb98dLghUFLqik1CX9iWkT5PjVQxU68j+y
HCMiGx0h42tEvtt1hizGyQmcqiPeNPtN6CAXXTU2boIMPKHW2DCkwRjC8uEmq/bZ
DzhPHksxa4r9abBaWXmJ/K+/pnlubqY5KsnpZavDwKVQ/gKw177MxQ3IwfdqXK1G
BFP8W2aXZB2fpCWajzxVc3+1GvHn6Tvlo7vVwFqHe1sf3iO+6FFqTH5PExZkCxGq
Lrb9NLM62ZGaRhMRWLdQFVmilrhkyEAtrZt3GnmXNrT3C4GXhA6Gykp6cuk3tK1n
zDVJ9pGq898t8bTXKDZMGRntcje5cH/JeqzA3Ubb8DFdP9TY8dMJPnikWuG7N/SB
ViYKYgQFx3Z2BIhpi6sYDn7DrQ1DLLiRJIUlIaUVFCVIgcjUZEPXL+UK6no2q1xc
A+VmqwIc72oSf0WcM9s2KU071IIeKNDUtPGtAoQDSjMvtrykw/xdnwo1aRAe7RwY
Vl36gAJJhAcvTFdIVZfH30jGkYF91rQdusBqmwtPRT6/dG+vocUCAGE92kC2N6a4
+TGflhl4vrDAMkbm70q2rA1gsMk1Lpo9BH39A/gPFgaOwThP747ihv7MhtHznn5J
M4XzkJPYd8KdlysI/E4t2sqeY5wrRNGbI4ba8IawvIlae5xQhjpoLXk0QK+dbLWR
985ZE9jPpBcUa4Rx6iG9J1/8ypsttArbPwDW+vLI4/S4X1rPdNqhMHaQyRDOiiI6
LnMARxoYFXbkV8k30hDDM3IOmtH6xVA8RWjahDN3ac0TlVfrivN4fswU+/MHfpTs
9FSI6F6cjlQejLCobLX9TY0sHhZvZSM9Awhyc/GmNlkwWoPC6ayPw9e4Ql/jrSO5
FB4OE5bIUVWNeV4mAWHqAI46DOkoeLGM2eYlHV0V+DoX1zQdFSw4FMvkgJVaxOYl
o/gTsnq+n1YeZ+47ouAGyWGz8OaQMHEJruL8M+M8OOLOs96c40a/UbXlO/HIqHqu
cStEWNyTyAnOJewv2kqtIRRRTzK3u7dWDEPpTpvUhhGnJeb6FJKluXeH8EC8q2Jp
3JwRZoHXbKtQIbUh1NpJbp5WAHeX0dEgl0+akygPE4FZLdiifafbZzFbmAIoOOnC
Az+diqPBBnn+cwvyjmBTCW6zMkFB53joDX3R9y+UWxMTJ5ejVWm21xjD/JHg92OO
5a5awXxhlWJeDFLXtBVfBzd/4S36oKqyxF7MgKB9NUmCAQh55DJ5nCb6pzbtDVMt
Nxx54VjPjawLqm+h+PESEy1WKQb5vNUfK/eFbyqmDYfLnq63sss/K905Y47W8Cdo
Y25LhZO6jaJqHlbKZEWEgn7gOvEZ+5XWnEkEQe/U8PT67n4VLTruXsJAga+X4hTE
12zdPzTIXs8GCIllq3WPJrUlJ2ehNBDh1GTS6D0thELULbkVv7xWErN3yGULszaV
8AoqHvJntVB7iaWH340Ko9SuJCtTVuZL3IPiU+nWhX/3ucTWR7HcDasf9kqb1Pg9
M7tpirIuSkqp/FvBcEB0ynec0uYOm10DzmweLAlqFfYyXU521GjNVHDFQf/P8+/6
ixR6rpSd54i8FQ+Vk76NC4rikG3/kWGHatyaEvXhCs2P0RuSa8a9DxeBycFpmq6P
upIukNqphMETbh/mq6YGcRwovQu0OKx+IgUmsbVd/QpwNZXpwXYRQnHojAYNbGJu
xHO7xd13/4L2pFaWoKOnH2ecUEO/QvltTRuV9zW8hzBN3GWKAFzBuXQXUOID1fzx
fJB5B3qC7nAqHmWhtj1DHgfkcLTA5YSIo/cjJVsJ4YcpRdxm0eaVyVpAUbum5O6j
pvRVRMRNPP5H1M9Xxq7tZxOOJJUgTj/q3IYQXuzKRhyZ3O1CHQP7Wvp5LWwaOPrH
voNuYWWThPOQg28vNrt1BPlox9GzMCAFbOSAfXAflKadMTwVyVJNwMHE/tNW7YZM
gqN3Bg/wo+rm9lT4ZmzyL5gXRWjBhfIwbOfYhzWgpeArTKmmFhNzPfN5jd0Qg/il
eYysHJmhu9fzXzWxdOowWno6/bJkXMOqW6c/GBuJHfKSuTVtL23RverosJTY+gOj
Lt9hAM6beMFRBJdyp9Rv9P4hVT3ak0q6QjG4UsMGAtbBLytvOZAoj3jlydRBotHO
q4RN30SA838L2G8zB+DrI2xIpjPIs/dRVIfWjCBDRV4riA+FIkxpgT39tkozfnfz
9p8X+YJHfIOO8GBI61hrBSxmRfpbNF3VwqNtkw69JBXAguciWfu0fAndyy1nDF7I
pSfwW3g1FDneMwDFSuOW7KVtBV4jw93xcTkxa9JdoipvDhWS8hr/dhWWb4U0zjzL
lrOMLG8ya9Q/YCgNVoygcAyOtb1anW+gWxmJfXjcufkb4aohJ57bwkRQJxiOCJ4C
G/Ly7anq1oNlJXW2f1xGtbcDhjhd7YdiogqI/I0yalxR3C1J/cm8GCP89aLts7EH
SRN/1Uwa+9gmj9QcchQAmKccI8sl8SQfdnF4t1JSYF3EVlxkcD/yKhh99pHocH1D
lLAnX8tczpegLykv3LclP4leizXAKFHN00kfyd3wKLQSgUS5ew/vWusA0p1A3t9F
Fac+FQr+IgpBhiMo2OsyyTBJgutk3cyHO5zWbNltXjjne+ZmZNwvRh1qk6qKL+Bu
7ERDizUNUxuOIGuZP1jS3UjNBhtT+KSKf/Hy9pa75VgpqVOEERrgymjobm6dDZtb
rtEuz/jQVNe5O2mi2o6RaI0YlNxSL24Q6+VFlVI2v9CRmWA6zffgh5sYwKOM8s8R
3rZRPfsiR/EdGwPViEsdQmejE233hdN2ZCaQxJ+orVwOfOe+Mupwo1SmYJKS7zWj
/63lRP/1YEfiUlE/Aku3ttfmEUSiyndWROoSOkov8HH4822ICJAkcvNb7qp8upYz
Pzc7L8x3hURQJlf0AT/BfKgS9E5trmZvvZOf+Dq5hD7wk9drAE/c9CJ5waiMOKZl
CuV9DgoQK+rngs4hfGWih8chBJpW7Q3wqB9PciDNSN77OQzy6t34n2t8I3zaixpV
iAsPx82zBX15boqFYe8tB0/C9qAAgghihkTGbqNQ5TNvIygqRnjtZhH2uZvSYoMU
NV7RHE6IIYLtxjvYuqtUq3UjKfD/njYwUqfJ+QNSEbCdcCq4kxMiq5Of4Qo+Sm2I
/IBH89S/5pOpdStjHKTOQDkr7wO2va82ZyFrOJ8AulU3mcgpxYl7sctWPRbWkkP6
1MD9EzY+bACgslCwZNqN7PWiTbsfApEot1chB4i41hjhkAHXKtGwEybh+RPfV7EJ
6fELBZegdIjH3bojKWsSexqoNPQGyX2bkb72sURVWA7cA1xX/82xLxy/cNxFfLoO
NQtvYEfqcnvpZkxe5EORlp3J0PKdaT+7JiaykkqaEJ7hs/ZChVRbivMd7Fyf6Wv1
EXujhTUL7U/Z0tznIJh0byPmsNxgFcAVg+qDldxoEJOlUX315TayHygB2wt6y4ki
YSRSPoM4+gebiuid/VeR7ikYSnVVOYTINhYaVughUTISdmHraWIJy8tN2zss+rb9
8nK8vZMR8dh752t5oNs+yvexAJLWDvRmMKU1BQXSlDpqygIKnI0WEkdrMzpIzqsb
qnwACumWfDGRUuchjOPWO8xB6tjdRDkGdyhVS00FMxzNpwGFeGYS+2KZ4FSAH60n
/JDAVg4d5H6SeMtV+d71xOyhhk1A4cIBT5X65iPlxLdNcMNqXQbfAuFkSswRSu3A
TErzM98T8+eV5c89liPBZt7Bn2SAhWZ6O2Qq8FsQe2dqo1KwtsQGZEC50+DykjBx
IQhOtern4Ppxk+gG/dc2jDuUe+DGkon5q6UfAvPTbFG+l8+MWOaHhU1c49/H8Vzq
RNV/MbZOVk2gBPYN1lPohjvVjkxdVV6oPtpA33eOcWiGdraZG7uSsTr+lGqXmo3N
54aovDRq5wv3J2nLJRioFtgWxtPo8MuHnzFdGTdsfaYK43ACFNyVlvjY4DS2s4/p
vtV7WP6CCBTmIfI/pmORiPJRllEAU5hpIk8LzjNaxvMEzGMsmBZd84K/4uvm5r5y
YRJzyzgysRI9+FHICWQf32i8sHvRVaT3OZ6PuuIvbj1NCmtQDiXinNIRVg+YC3tb
kj+HPzAvAPh2jJo4lvL7A4/aD9PL35DhyTmtrJVxCIQUTwhSCII+k9uTnNVA+I3I
aJ/9hMlrGkl5PsEf+cZWiWL6dBQ9YWeYZDGfhI8XabXewSmFcdNB2vOI4tSrhJGP
J6/580byJcUYR5iW5mu+lWejopTLr1GTIFEkngD2uSJSd02LvS63MAW2QPxMHcE7
ePAvuJil/FdA+NqT3DVkEH7Ond0D89/9NTwreL8ir9Ju6draHfT4JK0NCNoC+SJL
BCkwV9tnYMu5l2/c29/akSzwxjll+U8yJSzqDGS23yHRTmfRz1xoRaQyb9Cx2RJK
qj0uDbMpZoPXebcjabgaI3p3pr8ik83KwLdVuwUh6yHeASleLIKzhLnmBqvg8rzc
8MgUlLuJjz8ZbwRyvEgcjsjl4FEJUmBc+hJ+NqLh3LOW3PNqNj8qS/FANwowcmWr
Q40Z5y4q+u7kYztXhDPTI/zrs7FKj1oXTCxZIPskTtlzdGxmIcRhLAdMHYGOQg2F
c2fEbnGSuwyokU3NTaQfvUWvbmMy3RV1OIR3Rb9T9bvyG5BamlWfh6DBpxGnZYmB
O5WmoMViR8Gv/GMyiMfasfhVSreQ0gSYq3aN7kjV+AKjtxCaBF8VklfxJ4qZXbDh
1XCsKyM576diGDJZ6AKiFcwSj33UPLz0nhnzeji2BWpf7FZUSpC5hYTq14WLB/mp
ZfmQ8nH5TMq0naFeucdfTU+qn7g7g8KmtN9UtEAqQpc8J0DBvFcCpXUVDsbHoGdu
G2PInSZ3/yVgLs8SWufSZq5RG/fHXZwdcZ9VSQhMfGUYLKRw/14r+FhRbWWEBZ4u
+H4Ambo9ml1psqd0CL4Wqk7yMyoe1CoGRrA7q87/2+i3fAZX7aFjQ6vEj4BlgjHg
kW8rmdRxwQKNmPyBXFALqjxY+DOqm7QwWXWLrDiFFPwE601S/maDya2C6++f1Mrx
HWc9dP266hFS3n8jtVG7SlRyly0d19VsjZoOr9bUm3eE4Pp6hAk8uxBKoahDNBgQ
uuhrR0li0pxA6kx3q09v3fV3qxv6eyhquX0SlSXyP6CZAUW/94ZU6FSZZ92z3zKz
uxnLhBopYE7rj+JTzPEG0x0Ff4v8Nj8SmwsaQ4zSJF90/W60XLV2Ivpr3qmP06Gj
W8CvtJe2VTmqAvipjvE8DorjZwGSofqRam17XB7uQRxiE2hds4gMncwWzeHFR2SJ
jq5pYz5+Ylyo1Vz4YllU3tBixFGS64MJP3GhyimZhIrhi+/B5TYGDO1WaBYZMaJs
9rTIznxoAyyi+Qay1yw4SCQexUHXKFZKLp5TTWMDZSjrRP/uV3llsINuxhvMX5zA
aVmNNZPfNYd3BRdHyoZopLwMqKquBX6qqhkQpciv+0vlKAV/YMaHiHKfwWJqK5DW
bUC58fZMIbY1R8tnuUdy8YvLRH51RNO09s3ptFxniHuwAJ3JvtdDm7QglQUWSoWi
UiCjjGnppdUBqXPbLKa/J51xUfcaXRkWNX4vhVlFL/+EYEBoTvk9zdr0bdJLOVir
rvpAW22UUGGb66deWc0rCRQXbKcDFvCMRp16v+/StpgP9/8R4vvVCSNbMqCR7Kzp
7Hr/QUMLfDgMz80cxMoGzDggaB25jh8qs0PaPrV/VB+zr0s7OaOOqrigjFspq3IM
r4rOBZiSXGRGHda2tWKdczSGUhX/QIPpcCoGljSb9XTQe7FLqFiuJDfMEH2Vt72D
lwfYTzgR4w72XZPZbenE/UG8B+ObivcgSV1zXRqbhQKJvshRGk1JXAe7ciEL8xWz
z3npgeUU3G6C+iX0cvxMacEyLqkTGOgKRqkS9oWPRaQzjm4tCyv0AwwVMRP0OLUk
QOA/q2UgtUJtZedfwODjiVo6EbXHWM++23eoijUEefIEoTwRJH3LzsdQIjookJYj
N5pp9kBZuxyd9ppJBlm1A34gDfcXgnAU3WDQb3p8DzDCYLV1eXt3p2DO9boZMOco
Nbq6Z3kndaaruo7haxBVDTTWjsAfHIQ3kPwe9PdZT8YxXa7XTyyi6bbej0LzlzcC
jTU7DXpidFaOP2f2dqAzME9Vs0omotHZJkuJmRWI+g9p421mKRlBC8/X/g7LlZ+E
MVaD5bMQdkxnkpyeurm2YP6xLuYCoasmTfpl9dLJfC2ESGZC7wGKrWwd0abO8grT
2Mqbx7cNvJitissdipWS9otHr2dLXH5k06DeaVAVSKr9w1X6J/6CxXK+7Upf8tia
Q0PGBQZj/N0T+faBzPv6BMaEkS3SAAycvfTQ5Y1/K9Lr3TForLTtW2feky5W39yK
/dO1MduO00TchrM5MB4BofPCC7rWDZArcx+4XH9lOUNV5M65AbYxKNg5a4XCYr3O
G8B75IxyOvVLKfX5KyULMHrCvkw+Usti36vQIn+iY2qiBUiMbYiUZNbb/Sj5E+1k
VijdL39jUTamdy5ArZ2VJlIztbcGuIT6XELT2nJ6mKvx28awv7v0qdQMAMakcaf7
h0r0ffgAcZzVti/gLs5E1xFtThnk5MhM624i+XrjnZhkIrthZaruJ2F/TsBRINCT
nKI05D759YNMWjBdEmdrs5cxHvAOJK4aEja8jiTpMWGcDc0+srVgPPp9PDZRlZ8A
ol63vWbvbhkVEidBVvSkM7SCYz1JjP3+SU62e9GgzPEWymvIh8c2ZNjBdKr1AAqL
xiFjHEPYnxeYQtQ/7YahSipqUhfjznVakEscwfQ8JAFBdVBBJmOrCSbrM7Bz6MJG
qKgwJe5BB2VAGnqCu3bGs+WAgFm3n59qb8TwYdc260CSxZDtRL2s34Rvq6tYUKQ+
W1TKYe0va8X7oDGW7bsyaHYmJ4kkQlQzN1E7+3qKoamth6qQvYaQsq+NScQrtPqZ
Z7sHokmDV/UdApSY8uxNQSlF7JOai1JhXFGvRvFDV0nro7qlQdN6yt3oCFoLUUqb
1WAFoBGcF95e7+6z1T6KHXoSDRozx1AK8Ax681Qhyg5Z1hWys16yq2lSX8Fw6RSs
aXxffKR0q9mTErG101pMJQJr/+5DWh6K30257gLzkJUFKjCpKyMtO/fDxfejQIgy
83xSCkCQgk3yYH6to1NMkE79+6Bye6kG+RrHYZPY2AwtppAr0s7ZSzVqDTuPHMtU
0K4yL+Uh7Clwt2ypS0EevjIU+nc4E709Pw05y6z/I+DOmQH2mA0tUyBDA0voLZ1v
Xpq5V2uhSRwzspJT9/lXoce6GGVt2o3dYlvdGvbjrAZ6wwuSSidBrsKSOBtLfHBJ
SbAPCKHnmndkHX/ZwhinGb7gk/VLdU7Xo90gdK46y8XZjW2oqa53wE369donwrF6
eH0gh8Ryps6wOteo9vpjBr2PEWIyzr+3y1gsdYl4qbswU6UYKt3EOmSLIs9/GI2I
LRl+dxeTzkXkj1KUZjde820Mqqpe1jBOOe81rMC3cFHFgkKjM0GzPc0Lfg/fmz3S
BGk2SWNDPr0h84TWz0o2bx/M2yGkAWEBPCAwc14kHc/8Xjc3s73EFRBW8Pe4uaYP
Tb20/tCFEUAVRz21qB/Y+CL4D9mzNv60uwHDPA7fYNmjg8fM+6pDLUbV/Dzket9f
k9IIxv6QcRQKY6VrQblN5Y5Npu1bSUS7A2hEL4au3OBfywKUyuSR9VkhYKCCckoA
ldpmFIE4ynLLYNLzxM1jeB7jFJ+oLF/FkzV6aSQNFMd1AwVtriGFMF9zgmw1lo4r
Otfet/vIKVZt9WCQjz4fGrXY0d6RtqUwD7oc5vX+BmRXYDuGuL4mKazVCkxyjT2B
ZR46RC/3KS+hvag3mm85jAQJizPEHujHnDf21bqoufmTFL18RZ7CWCN6KGBJvuka
pg58/pVZapUIg2FBSmmNoICuZnUORplao6Llx/2cac4sD4rfGXwsKNBaVSlwI2Kg
rRS/nMUBFePhh4JX8mWiCAKeqIOxxzY57LiZSugv3gi4ObIjEsoY2xO3TVwX+bX0
98/N6pVdVkOG2sC5tCft7h0Kz+HZ/7cPQ+FZIib2OvtEi+p98OM8Zo+Y2rlO63Tu
8ATw9P0mWWUnf4mabxAZaEidjLl9hO+c/eV5c2qidTMN8YvX/uliv0W379AkvUf8
Wx5JyNvuv3DTppN91Zp3vTw8LvRfKdbOJk0HHcIqjPnu/ICSUsb2pxyrbbsX4hKh
KPoDpdYD/RLrajRSq5WtVCkI7d9482Co9WqqevoxQHw9MQZ8xnq2EMgwNNoDKLq2
z5MvvUbH+TWGBSXIkQyAVNFNO76lEw1sJ684RVG/exPZW7xv6TkDZHsG1L0i9g1i
cms2fwM3xPIY0yFpPAEUxEBxNbPjH9LMxNOPet0XuXdKYz6tkzUnyEG8c31lICkd
4+JM8aPbtOVI2wrfS+GfAr9jGFUqx/Ek9n+NntwPEwSe3CRXjycecvtCMsCNzf8C
FglckUUr+iXhNKzp56xbgqs/N6wv2HB39Nijs84dAMTWdi825QP+WIAGs6HFppMD
D2FsuxhktuvCaQNOnFMb9+MhlYVX3E3kpAZ+uhvug/Z/4m+nvAxT9jtE9amlJwyW
u8rIRGZaQNJEWIQ22RBaJvIbegmhU41dykI6+vljFu9+JWfjhnsWZppXMgVuAGGD
eKNp2yFZW+YA1vpPbPJqpV7TPQ9WGmR4U3xOYb53fnV4PTGEMfgozakIx92vlJuv
+6VSpzndpnu14akoW76IGI52DpiE8ZFrZX+/jo7lNlQy+N2XKB7J6hVxmv3i3K7W
Brg6kkp5m9Xeqb3It9DlTHE/9DTd3ZAp12YNbywyjA+AZCe1KCiBztBBQBLJrZft
s0lgmc0z5r7TM93I5RhgET88s4A8wfqrlLoBEdVCsuAq1ba2cyGZEMmiAK1Najxm
b7dNZs61YbPDkHL9LmN9j3mSX/L2pwvlV+PSWwjfQdB2XpkTTR7gOWrxd3xlCZ43
MDWQur/x09pghhur8Me3olExeI/ADgse0lfqBt4BGxYq+BjjWLsy2630yipGlrdQ
669PwVhMfZ7FDgGMQFBToIQHOtJTtOThTVFaIS80n9nxfIukKvV006/6acU6se49
/NMZsORqO3gm6fsyB/tqmvFpwqCcRA5tg98pJCQgSmgK9CHCPdzbRLdZtbZ0i5Rv
lk+wEh4F47FQkL8XErlaWxeiRH7BPLRl9TS66YXKOjehGONNY57KrQgYw+tlHcR7
jnE5voEAMZd5wHrZlLG3YmbBny1dPJPkfWAKC3mBysAHW1DzQLA76Z10gYpnkN9c
KI3J1UTfXRCZm153w3K6EEk6i4TRd+dURedtFq0zp3C1OD9QEzhAd9YPwb+q6dnU
YReQh19FQtgbDINLdnrzY8fQCmgBlhD+h89yjHzEx4oIxeg0AzsoBUcUlmBkwqxQ
PCwQK3zcVXoHb0ffDQIz1bzdGCFp1W2hf7nF8oCU4ZdB0FOXI4DFZO8FbFD2jW+c
1pUZnbmxDaXAn4z2k7sPtOnVxcIZeJo5O4ui942VPhH9EeRgryr00cf0jDNOyvgp
b4Wbz+JxHYAgFN4yZMpLnL1mV1X/JdJDkBxvMZaCAZpIM87vN8ubtvLy7OLGPsqY
+2l3UwJ3mo+2PQuKbxiT/CIOBnf1Yv2NbOPqjxu5FeDWvgep0AeparmSIDzxUv8D
VkE4b3ibZPT6UnJ8jwYuq/hZh7i4wxRY6/r1wmOQdpVwY8L1QyciNqCKc0VJtz4t
9Peh3N+t1/8p3BdrVRQVI8ll0bE3vV9loeskehYV+X0VInvsqXhdpsdfnQjDH8UC
CsvOcIs3FqsMUThbvYnVpQyPzKZuBRc09xVx9Y26DhhuM5cKh/KKnSt3E5+KyjQe
sdAKMZuNgFeYseXyiEl57puGD/jrO+N6im9oMhi4XZNP70KJNMdct4zgrOdVR1VP
+FK3e7HxPU1AckGCiM8HFDPOJIu9jy0ZWMSjpFZLYC5JQ+CbQNZj60mdLjrYt9eR
Q67TTwaUABufiXJiVYXhrLX9cB0c7iuu5BnkmGJwXSWnoYUi8AUZ/lf3JHJ/EqMG
5cHjZpQBagqbCxhE8axCTbJ9vQRrfzTgmfcnCfsYLV+YEooxb1tYJqJRaHk29ZB8
s8itr/cjG6P6UF1AmSsjcpJvr2t3jLk9mMztQpg18pe4keDwkfVJHeJVEQ5PZ4Fe
bNYrRAojBiDqHn0WMN4dLNct3SsE1PuqKLYIVVnkZwtxUiAzN2rRUypfqrXhKdH7
vNnrb1oHHTVCMO0mLcL2O8LrmiCkEBKvy4CavAe3cZXWv+UyZxyEm/kOl+N7bJLi
1ZYW00T2GdV9jVio/9SvApvBlQoRf/Z/UHe5GwBgHwLWji5yTpWanwNvsfbUrEZ6
yuP/5gaC6tWvHDEMGF1y+3WtRtDuIkVq+OrqEecnJfmWCZinpSC/XszOemM90e3K
+ithdpl5/i0PLOt5xvCXjY/ENw/t3B09WudZykpF5mRbcbOOSEVVvpKZQrawk6/L
k0d6o7kgjksLZUJN+gkoW624H1cJoU9ipCByEj1PXJUTrsD+y9p9SnW6h8W24QZF
d/9u/U2BDo/flo+LUzKUmUaa/7Ndxwn523U7qYdyTFzbv4iAHRlD3TI1u8aVT5g6
LeH2erFyraBSy02qD+YKrCg1FQt1juNakQ9IBCh0IuPBCJhHyaH8ef79szIj2s91
fFA1UO6TIaA5VaOTFlIKtn7P/tpUTeHzjcJHAzaz63iAnQot/2fb1tqJidAGycG1
fVEbFJGYq7rO3YpnIYnUcmxLZSv568V/lQ/X1cYrm9gd2S9fb0hA6Mbbp3RN5kIO
E7PMFTtq6m2DtWxQkYSyjmHUCvok72wNAnb8hKoQ6lPXMBARRzHlx5iGF5IVFVP7
rDuP2XPv+FgLwkPWE92upL0+ONWmxgxRXzZ/no0BHgKdX+LUorE8YGplgaIkxxkl
PQVo7FSMB1pHdq5JQswFyA==
`pragma protect end_protected
