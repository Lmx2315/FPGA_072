// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:37:05 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
RzB+ARRuIU51YNsYYAGDOpMOYnuoIV2KL6IXod4nTQnlhe5Ontuk6pCQuljWHFSe
6evbsZ1PxmTT+cxIeOPhi2wePWf0jhpHQo2mT+6WPsql4S/Bso/bKuFZXFKewWdM
FJHVOjmGt/RO5PV2Nn0y401JU+K68D0II4YoX939Zjc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 24512)
ez3JuUkv+h3RsORQObZ3A3UScECxA+kV0Q7pMX0PsV8s2zUqvWCHg9cZvuW/URr1
ptgGVDQ3VUmKKUfz9tQa4JF6zxZqFza3MaOYODyGRKSeKYdLa/8VA2Vt5qPVFeQJ
AGdRRKSsOTCja6k1IHdUNackhDZLkn7lWmBbeTsSkmeWIBX86DC2PpQZQK9Mywf8
OTpKzC+ei5/6hP0rDOxJ8iW+jZtuxalMg7h3l6Lq3f5YN/TN2WuLe9TaDSxqPKQu
rxSkFi2idp0pWpF32zBBEixJRtTn1ph/MAgaPSwz8qODzhS1/KOFOVujhSGYSsD7
X7ntPLUfHXxUlxlGCqVQ4y92+1KbbhR/FKIwzRbTnyW9RzEHmIKIlsVM6njOD2+a
JzKI+w+ESoxAQu9GPQyXOdM8XuoN6VbwVkSLDx8BpAX8cceFPDYM03ldNGGn8DpL
/HRvS9lUEuvM7YBcVUTAt7BZxw0AgcDg5Dj7bgK6gFz0OS8bKmKzmlbadMUR51Nd
M+jkpavPqwoucjIFpAjL1KawYR0SK6xlD/niMreBRuFIEqanXmXAAFVzIVxIr1vl
Dr88Fk0XEOrL88xNeW8ZrI+9Li9oieOCghApqtdsJREL2uTnF7Q56J1LwxXFdO/5
c4s7CxJUe1hS0aq6JbJ+gpX51IG9j+m9rgx0EHRRoi6BuXz/kcWQ9BMCJfSWVaV9
S1OgQEKn2l7jEJtueA1RFAorP9IL/i1JJVBC2jMgxsvbLzjitYAzbVvbUI1II7k4
q4iZywdb67kLYOb8TXdg/HFpPT+MQkDwdds7uTayEk23rh7m5AmDtx1mcmZoY4zv
raFuHQdOPIi0lekfpn07wYz/PGeM7zXmZnxgFxiEvGuoOvjaxsR42stec2kqOdFW
WqFR5g4UyMpQbwnJ0Un6Y/3Pa3tqzYMfMKvvwGnHne6nUd1cvT/NgfjAW6Nwiglu
RA2EU1KMsbm0Uk168QEgy3K7Z87Pu4bwWc/lyyXNAhUzK9rhnddWfu2+ozoB/nRc
eM5KwizyAlrMU+1cOsIlAdThQZm5TPno6qQGO1hK5+YUoWQyq//nwMOsfFDIJd7t
O7I6ysrCqlPXxwQtuCj7XvONEDCEJGs7Ab0i9UBTDbtN6mHgsfcljCP2AN4k2I6R
RGP4UAfzTCV3PF3BSGtQRzd/q2a9W3v1i3ym2ByGi/furX+BijOwDLSTP4diaB2j
ES2SFGg4QEew1XZXSAQGe9eqEDZ4BMgk4PR2G5H9QgD+ey49TKrZALhyvMpP3zic
nXxf4pqKGFOesr6Fz1D+rGGHoHqLKZ/9Wv0ClU5gpxuEcfIafXqf9hlPyQP+pYis
83v7UC/B1HwCjg28zGeizJhOdfV/3iiwC8n3uKLJEak4ClMRgs61kr9h3sb3tR4S
NJizdjOwUgkpnzBZ3Fsej50VQLVs2R7TFnfhUHVYZ63+k3WTXcFylDHxzxblQZhv
MZb0Pgf3oKUiB3J4mxDWCYzUnSdfC+sKVpssLr+A6uT5OcCIVNUikWqcmtFA/rjI
2JCaDcuEMaw6c9gLJzMXvUueXJmtswfOqtBikAsiRQq8Z2y8t2c3XeW+54Z6Ovpu
d2ME/GRzcUpXKL83Obvvr+zd2JgRJrXh4XTkw8AeJu2qp5aBfm/IBKkBSK9CH7GD
rzxyNb1KHoDVFHT4ILSor9ymwX8YpmmgE53Lqy2nxpZ+wZGzuIwVp8aXQKedpAa5
Q/V0gd2OBpJY5LfcmwKlObfrFYFWBNNNtmbRvoJSMITRCNr2hPFoTPfds4C7QFei
bUIYgsncN4uHtBrneUvt5VnbYwE00cew3bQ60BOQBPR9a1Sx/BQEY9ImkxFSSazN
7VMMhhUAUrs0Hvk6I3JLjBOC6zxZwPcR3H4ftYXW4h5uixjr4ELUKqf2pJcGB11D
JBPb8zoN+B6e8ZMTbhd37zSWkRmHozdb5nx9g2wdHsJiv55BOuHU3z9JvGHVOagY
RcPzKptKZJiWA+wLhJhLEwGJ2/Ko7PLaOfMqYzEi2DSKrZOLvv+n8OU3feak4kGw
ZZnXDqz8ukdCl7TRDLTj4mv97OkoVsPTI6+z99J9A+DFiGuB8i0PecOsRvhHBLZ1
HSMuLzEB9Wztk3g41O8w+3lTO8ZiSvsfE0CqOk3YraC9wJ68yxDWYIhUOnvnkHpF
N4AO+Qs5R3FQ7c/S3JLa85b2neaaHy/oj3ilmc8iwGp4n8PKGy212T2RkiaX68Nt
8fcdZW2FPlnD6bQ0MY+9PDPdA9hL8rglBQc193VbR7jym0pZW7RhfHPz2Gp23XbC
QTB7GB4kEEjQ5WO9Nx/bB2iaXjEVRs1TaSXU/ON9DbWuVd6xUeBWTbAgXT8HYgxU
Y+mVLyQtcpqUKDS0gl+4urexWuuMJ32IQTjzWtfai3/c1o/U0AsE7zubTVh+UWYi
730R57sPkzKC4uD8akydvSFn1h8hEqRxPUN0mzc97Gyy4qgmkHbXBUPOG56sT1Ys
YF8TTaR23GlZe3tNxlbuqZVuEfZXUqucCT8yWalds9yV/maT9fyK9WX2S31cShNj
kc4nQRCLc3vNXhH6OBATXBcAbCZVQXL8d790raMAB8flqUJ43kcHhr0otntnfSRG
SLp5AfBk0GgIrVu1ytsENOqZjqhrUQ4yFuLEl78eRB8B11tElYiRA7f8kGTxtkQA
amG3Zk+FL9wONvyV2wZ824Og7A94qOtCh9fmQ1ed0Q3X+LhAaQATVbpupZwj/KyO
NHoJqGi3Z/I8L5oh3S11Z1GRIdthVs29VbRBANU7nW0aivzCPnVlJm/ptBEWL/S+
oqjiwmzpFFJJCVVvElgJTbHW/SUxS6A9ISc5j/KPGl1I3BV41spT5QCZnAyWDk4+
w3dvyVZViP84V8mcMgXXYpjgBZgNFrJ/HIukGUBLwSw+OHrk2kIbIXzAVzaeYzLO
T53jqdVj9fdlLRPbGDrO5YsPMKxA1BA662tXRazgXeAUDoMXAbxKPaoKKwdk5DYY
JM3gUyzh/mPYwVIsVfag6iv4X0/F3UMUrnz6c5M9fOQ+V18G41zpIjUuxi1tRB8N
yhJ/aMSsZVLe5mhZj6/VM4q0IT9pWydnmwdGCpTBAvs0NEKzSJnqujKfv3utiY1E
uIzytUxR45lUF01iT7MUbQkwbkFswK7VW46E7VNJF1doUzTQ5Mk0G1wX1suWplTL
x+6hnLQO1GP2aSHubMe7MpF+MH6CgMRLm4YGRVQ8IgS2usnu6isyjwpiMsSi2AKa
d6t92LF0Q4Gnv5Vdu99XhX/7oPjKRqonTVVv+KPesmTu6iANg97YO9PoFfXb32bF
qYM/tZwGzNuf1YJShQ2DhQ4N4vEAJDcWSTsu0YDJsYOHCP8xRvyY9vIXO37kKZl7
dqLAFwt/L9xVR2NJwA7I01hUZAsvAnJuk5qjAT+bMTcDMI62lFO3Vz3rLYGcHFU6
sal1j4BKJuVVy3LYF6YrJsplEQw096TntvG+Bt7sQtzfKfvkjeRRaUmhG/cCj5BU
DxtBz+khrit9A8eRWg25D9XJ5f6+7ISpKrud+5xFTGRzOS8W5jONRqVClpOhq7FV
RAWSBNChYlIy+bYypliqrQqURvluMzqNbNeHLSPMC+tq6eTAoNp1s2zaGrH/Of5I
uv4EovexIMmsl6UbJq0FsVKTXfXQgv6vSbBItb6wcBX5hIJE8gO3MBdpihmA6XKk
YFq841YrK21P3PKnRrPL46wSMH2u2JUYavSrNLlxXSt46Y4BH/oU+w6v2cCioee0
UUTSNwV1jIWE4TGgG8+vA0RFcX9wPpOHWV66pECB+Z4JY5ZhDXdn3D8l3i7Kwofd
+u87g3Rjxm3Cs5y1YrncO3hF+oSpg+fNsXok8fWHr9dyF09xFKvo8azV8ldV6RxK
dA/ZDPPoDsaHla5xN2r0o/60n3kxssGyt4KrIYqafhj/QT+fgWDtlN9rwPji0+b+
DZzN7c64LR7xIUwesrUUMzWBUQppH/gSygZZMuFG5gXTOlBGTKMKxOoLvdFdHYv6
xKZRpChkLS3hdkW/OGtXJ3L1DZkBOUVkqqbDXkCXfWtYvV5IUFbscaoZf/l0wL/W
StPkPS+qQbNDqDlAkBGFc/eH+f4YZHcflDWCxPDcei8fTX2k5HTVJnkr9MF5Af+7
aMkzkDNgasje5m/3Y/BGMwJRHE70klxcBwo2hydvRYrblX7gnnlJ0nr/lg55unvH
VfLNkfTSpXHre7XPEYd+i3in4/GiNXpgI95xo/kf05G3o+c9VMdIo51XzSElObuJ
mH4oeseAwM+dhwU0vVDg3rYdTGzBMBBOgSHPvlkALf/Wvyjw8x/MNyozb/iSqZH9
+PszBAcX7KpPc+80Nz4pUgqs9oWdVMbfp4bCSxv9no35CEqrdtRftytmRzQmEgx9
qzPISFuIYzRgCz44vNd6gO/1Veecs5NJ8tMR879AALuQ4bRQVUZs8d0pY08eaWWZ
C2QJmkulW7WQ/PpMvZgtfKixsnjWWXZ+kT0Bg11MYrqyOGc4TgQB7umNLra2Q2aw
ubaX/0XJST2gWC9yXClSsS7Li/3C1Dcn8sIDJ0AFJ9nPhZ8lLxyVbK+8KqWEB/6C
mOh4xHe4VKF4ttw/zmYMIwiJxT3M5s/sJ/1R9Ri/3m6hZW3UxzaSIj26uGclQ+Ca
nWNYT7e7P/3LCRaE3iG5crajmXyeu09IE4bQSdGiYYIlQf6LD6Ifswe5h33qVmvA
7Ll3Ehx3a6B6uBtc0Lk6njWaYu32RNFWjSBbLR3sOU3XvD6vNk5YHwOkJlzFp1+I
irYCh8cx1gOEX8LlR6IPsRKv4V5TpE4GQ9Ls4qFIVU8F3vBcjgyZqJtOrnKC3mYV
fEzfeccHYH3+3VyGNw7sq/VNaTx0rk3Wseynv//aYZxFYQg2WA00XU+AENHK89XY
HlnCryclQHP/B1fKdoTtLDuSGlCiuT18kwwHFZJcjmfvNsamTUe7fSdn9WIqthCY
KBqqBAOI95q1Q6aGhGNo1m06YzeO+mbpSKdPKFMXeI/A9abj51GCf3FMqTMtS2lk
jdrb6VzRbz8luRHZwUo3tOyrRNVXIz0CzsGcK+yX174kt/9kOZmpCryOsrF+dS7I
8wkDCc8ezS18Bs4w5qgypQyLtgsCsvQhi/rdD0slQLwni84niKlKDfkh7CoAw8GB
qkWqhc9F1KZxdBI6g2gOELSP7kJfX0XFD0Ep7dZx8CuPy7tlGKHOIUEQfzbcH2/f
stpBhgjAnBdnc9xeWctHz9V55B1n3xE21gpsEDM0R+Z6cyOSTfOitUC/VyRn4UIg
npofRCawiQwFvmvePLrM5MWpQkLhIN3hQ/2+DBE2uu+dFsEibipQB7Xr7lGfEO3H
mvk16hkeaM+yZ/8lbFY0JjANOXRJ7b+kK7Zk2AqN/GoCJ90Dm7z8NPjMd/Z62dN1
O0HfX/Am2zhzo7NEZzUCPq7Hl2Ddkb2WZy8VWTyT0kgEZQASzKs0S/gH1r/cGcLb
uqZphkLnNtEhGeDcvh2fsyQztb/OqRlZ84/8ymEPq684InbByy0cj3VXrWuxxbyc
6Gj5fTInoKg7n+rnjNoEcptXn1a8hazwiOxwO0g7r+qPJXjEgk9QBixqbs4zxlbE
lq7/h0panTZZX2fd+of1Ap57kjQ2djI1DlEd8E9DbnXC2l1SaI0gqSnAG/+8Bjuw
1XMqoCKb5BRntlY4NtijBBxKfdXham6niHX5Wh9O9qw3ylovNNdRVvUKmfCn6QNy
T9pOF3huF3brw9DZCc7I45aYYZhSYDszZZhMzwDfktzLM2Ed2dJPfCBktKzH8M99
74tvhWpsNrjSuRZmAFSf9CaEq1w7SNFJ7smKD4JAoMVxUvanUIkqPZH7z+3LqmC2
ACAeWIVJ33JB6jhYoKCFiZwm7O/zfINnm/BGhWrhtyIpLWb74bguq7cPOsdAQqql
DJk9OrUS03I5is1vpQVHiw2kyej8nve7nbdATjFcjI8bjHxWV5r6D9xJydIuYrHO
AnYT583t7yuDuMmvB6jhKv1CQHxugHYehD23r4em9XRvqiZr13lrasZ3y7LJoaU5
OIN81TkZGc6v1jHX4VtFeByPYw/qAgySajvTLPkLln1M5r0TyOEm1RlX35FXxej9
XYojwpDCL91hp5EOLjWb9t5zCPqbz7sYEj3PBxOQDbuiSeXCKNSHYo483DAGm9vh
aO5coIB/s1tjsLyAUybzsU6S4fBsWnniFljOZKrP05wdMbi2I1iI2j9fK+Yi6ehF
Q49uIQDS2jRec7ipEDqSu5dmcBcpRvOYy0qib0ZS4TGF6DrYloeMInA5xckXzJiA
XK8foW3+XXcyBTJA53pUP9xmM/p2r6zBfVJrmFUk8CGw6SjDjTJeQmGLdjjBzHrR
61svft6oYFnusH9yXl9E2FpSDCWrMwtmECUi/nDvICBBqBtM72YVl5/TqmAkwHDg
Prq/srGsmKkvU3qX+NIOpynmVEk+XlPWx8hlR+gUNcrwQFwshNVI6ZEy1L+OkZl1
lZ3ODNXSiDRkeE6YavoC+IbAlHopnGsUANMYpimuNPrULpX2N2WeQPXrw/TUKVFB
WwQORCBzGUu1FvOwFUVBk2+C3++QWZz5KM2bq+EXkXgGOp8HVnuALwjcc4yLynrs
xvMpDijK0nwbx7Rq+r+70RzLQBDWI5qC/MNSLbvNIZy7FnmESO7ymAAZeWLUL7r0
3Hyz+/jqLQd8qa5VQd7A/RKKw/+M+xbU9N/S67acDEiZVONkZ42shZj2wMWiNdR6
d6m1q0eWv5Atyf3MQCahMTG1v1pIfB6fem14HR/MJptFSexzzLJf5pDdva1QMLKq
JRxgjTeEdh8tijwGrreP+sNELUmoY+Lc9bzKSCTCumRUC1Ey/duUKcfFXSDgFr7N
fpP3ysncVXXOm0mlQFKSKJqWK0eaObMVRKWzLgjiRsL4AeNlM2eYcdIu/q9aGU1q
HeOpvXm8zTKejZ1MNv5ixdvhxOGpS/U4oh2VhAD2dZMP5oqbG3jEV8JKy+j2zwIF
KBPq1tgnUE39tGOvD2ln2ZouePNAgB/5DBw2E7OH5zM2rGbdsfI79z0TjiFWpQY5
jiJGPaWkx2/VZ/T3mHJd0QUPe7bIH1IFEnpyWE2khgTIDjN61kIDOL8IXVplZNl/
Qe6bZSsu30W7M7z8pgWFPcNY9vj9wmn7UZ4Ebi+ypQmj4GbKYFDr0cJp2f2ljFzK
7i3xCE/Izn/+sL59+CsqMswrHKwtLnW+f/Udl7KxJ1oNmku4nE26bJ2bCnYQFJ9s
y9Z4SEm5X9HROdBgvO6HxH487WiiretKEe3lvUVrqbt18IQ+bPEl6izc5CkaHiLq
69F0tmDZWj1vhmoPhYU5RK2TjvckAQ7S/ui/9yzKPXPXpPL5KTZlePatO3mPNGmH
Olh9ow9my950B8ra9Y1vCXrJL4lwD1Dcyx0b4wlp0YyxCzdKUvHJA4nL4RQEaYhf
mN7rZRlQ69HFRralZ3MdHqBEdkJ2QTR2cUZX9Em659tt0CAQuxVOT7uHeD2QeljA
TDAFoiqZsM74A85ohQGA+69n58fVSK1ZQy/ziVJxx25UuAyfsTSmcvhMQv5KX3AI
RHywyRZOMod5i1uPGQcmEBEsHIY/B0vd0okFTWbyI+f0dK3xlVKgtPuf0PfgtEpR
bfP7h+AMRXYFrc0IF5pRZKBnLA0sThaO6CHMnSefnz03Q0xo34lhO2yPCxWXlnHy
eI5gfjGB14i1iKhpAQallkQCj6AB+OOoyCkoEmiXV8ld1AADSZqkFsf8wLSxvOok
l6jGCx69MENhQGWrf88aC/o9A/XFuVWsvs/7Z1+0kgmhn0zeBl+GvfFbMU+eBI2B
GJBsJ4Hzpm6C6iHJIBequl1M7V6cpQviPAMy2DoYr3XF4MT4GvOjucSyHs/QTMST
IAgCgapIrulRaHshmRLifhF/66fGEf68K2f/tf4cUyI7EORCL7uBHuXQ9SvTUqmt
zE6G6DW5gk8ZOVoEBqM2OTL9J0dfypd1k7z5PsQM53RajlvxKtDPohMZumXc4i4l
Tj91bddlbEgjKlMzcV8RS7PRwFVwOxGB0NzLqAoo9imSTWok0YTBjr2UtLbwEKut
e7hgcXMG7ROP/XXwXHJ2lD9H73NuzlizbN5RLY4jD9IulhisLUI60MCMyViHMEfR
MiAHgHPhE6/Hzl6rdKchbFPRVV0RgQIht5yzKUGjUCs2crs0FrFSqbCIh9FCXuSS
ZUb7RlnD2+w8NqpJloIVzmcowP05T0hANOUiBLrb7A4U5LDdtT+W5BrAiJHngIgQ
mrIJdMcI5+RWaKArEUAxsK/jkrlc1AR3KoUVafMR1G/itdrI3WgGriPbSw9+IJtF
zzUbVeEEvQ11bphn/bXTvBABAOU5lYR7HlfgS0SJ0or694J0rWBkobktJ/Np2oLF
lPgHYpBpv8g6EECgCzG0tZdrxMQ3uj09CXMJA1wivD0GkKNY0sbmzCvty+AMrlMj
az9zHvUf7ewgAQi+i5p4axEsengcftTXRNN50TFBHydFgEReQAjTi2CX5rbMCuWH
+B7NS5lrAfkI9+2iZWj02hGopvECdLlL390QXBNR89VjSi9NSoYBMZ3SI9M+VbUQ
3hq5OepzaCNHxRb7LAf4eXRyOpj8WG/r1wwkuFwpVaAKt/SB7EYVVpAiFkCCpM0R
VimKc1pPnJHtf8M0qvajRtWllIg6U9Kvdq4OzYIbpqNRQ0ut5DyzJ4p4ctKmFWoZ
ap3W5OxEOzntRBE+0tmnwWK8t4z1PyAXNBGkITFvb4Qyiyie4HoOAwUt62A5ITAr
6nT6r21EtKEbFucx/c2lDLQ4bsOAyzFlRduUV7W8xhWdBpNuGnhqBjO2nZgW/S4f
4xWdFGha4v20JoiUhTjj4c2PABJ98ngp7MaOKOqwHvb+UZeEw4Ap3DazIsLp87J0
PvR5/mmS2Cf8vLinxOIhmueq8Z6tzAaePZ7ods8zWw0S6nuotLCz9Gx8sJCmHeKv
KkseuChJ2LD4gCaf78vb5+r8M5MmS3p0/2DXZJTWf8NPC4UBr/5V2rt/N9ghXqcz
4RSbc2EVpGbsVks4NIsDM6rZBlUHLAP9ybeqCPamzdpABBwNkqITD/i4acHnfOT7
Kh0ZfIFKPlKoJYAaSatt4b4sBN6QOIXYxJ6pis4+fo2JaiR6UBkDNkxZWp0tTDks
Gt1bnm6AweTuigu7QuVBSREzZ4OTJUPrYlKz/ov5ZLg0sSL7EEoMtXWcA/wvjcF3
wrTdZjHfBzrBk3JYjzshwCF9oCdNMPRzxuqhbmWnQoFovDXpUanssk9iLsE45+Mj
Yw7YzRitvNa3vuj0Py13eENyoIqNIIm/x7JOsDXgnDfvMFXb7Dg+BChrdfMsSsGQ
clbbUZHTtc+JBdm65lMFeRMelcnsP1tNyfu11YlW4SnNUMyZ/WQgl8hVAZhNxu1W
Kxlfwuyt+LE+JQz+rsIG4BODRutKjqFF+Y5IjKtXzP1/sOExBcieQgk9k6KAIVv4
Sszz2Y2tuJ2IgXOXVefb6SU80QBgXrbw4VX0qAJrCLCCReKFGme/nmAYgEPgnVaF
OLlqB4sIhX+7oCgNuZ6xw4iRnFIYKqGvj9Y+U7uHGj/wo4paWf7pk91qmlDKtcvg
Dndnfm4C9AzlHmBCowOQNOUaNdK5ot2uxR1z1h/EzgHtflDZHPfuUFBullKUQ/a+
C3p1vWQchsHBoJHTIVTfCbL1cKimLKO4DPMlzDe94nbRx80M0mtnNGk8n7lzcgOw
4+H/yc+hwNUT4qgSFGh4uc0kkHPBX5uJtSYhInL3AUgVBg/LZipgA3wwN92pD/TF
en5BIPMx37aET7VROfCYmapwHvyhlCxCb+vgXlowGVcKEJuFdTMrOHcQK+DfIM4w
KiJV2HpFE4RgbE2wg0sLWC7g3+keRTbHQCHAyjLohJcEQh5f71UQvCCpL4lKwPyS
U5upTK6JEbeG0fEt2EsHq+rXuDRqlcu+PQQyto2+3bJyALBMtcZvsnT5ZSdyPH0a
EVxi2u9kH71Cvpr0FC5p0IOMadfGPvZEkAhhidqGwCQoA6AuvGCSEJoRFkYJXYgU
qvbnD/0Pf/c+MxbhJbE9jUt3XPHyg9Ilor3CjFPPHum4hLpRLAO4wMf7u/iADv3U
awh2A3Em17s95DJI4gnDYeF3LFlDEIBMs5aN99sXIdhhuHb6uLzXZrNrQyzZorvQ
N4Rqesaf0MI/JbIKQ4kySHU0aYk/DO6TLXVa9THCdC3vBF2s8Tl1CZ25X1NuS8cu
trPfw/dP9pGuBnCE1L6evB8HpAPjDWVaLVpH1bCnMyoQTDxSZNVEf05R6BJMiiMA
EkhEHH36JTDm25UI8B3dSznypXDAJWF3XTsYdKhevxt/eYICGAmRx4zOt0OmnfKh
UK6zUSx23O1ostmQKW2Yosj9UQfCRf3782vwV/7Q4jPskso4HdgdoVVzbYenr2cp
WKbebabt6JlyT5X1W1GHd3uU6Iixq1dPK3sldhgVW58/z3ZvEIJsxfvsI31HgUHM
sxv+V3OM+RC1ReI0qfRulhmyz7edrKtTqv/UJqwqwzwpuOG+AD9UrH1zU0nM8ePA
xF2aB0RMaU6jJAcUfQyW6aHf8dgiO5Q0Vay4LeYg/R497p0hg9+biw2XONnp/Fdi
R65UsHzuAzcRBrnxmt9wbp96+6sbbMLlxftKSYrJiPDKcMWSlvGFUjPeYVxp5n8g
pjRoIRr6dY/EwqGbz1tp5O1FNEW3NZw/zoMXA1XcRSejWusCkY0yUa35scp6/U6Q
S63TnCc1jgSoaV26SRSetiwNhNaOw8a/skyRKD78tvAwj6Skmcj1fyef/fm7tBO7
423gRzRZVT5RYjoBo6+l8McaVwigykwZGLjRQZeknO9T+hjs/vCkB4i98jv531yn
5QBgyyopChkLC3ni2UUycu/JR2jwNLdtXurZ/YHNv7auSwlxr5EaLCmv4pKSAP5r
o9/OGyo7BZCd1sT6TIh2tG15HebwDjocx0mmtzewMP8vZJzt9hjVdvm8Cf8LhVoB
MMPVpEWPiA5OCGFT10aCrruhYA4EpncZEaiA3sbmERpHhrHzQD9QBiIsCwad6xYS
TlPmHzMW7OfIyXOTzgO+ZILfJvihlg2N3j3r8kaLOQauLzmV0YxDgXD9NeYfqfc5
PEd8EUiLck05jadzg3YEZY/BJIgdgaw+y2bRH5dcqxD4mgWNkhn1uf8KHtpePt2D
eecuXjJtPCDe8Z/TthC97HLyWb3PXuGkBzImgDUwmd/qCNte2/w1iHBLBzMNBGzi
JvplEUI3kyXTOoA4oJ+H6A84Rc6YSEuyS94uk8HaeBITS048ieDS4mxV5Dyv9Y8+
l4f/LN/hh+fhNy0ZihMvA8mUBNExdWz1gNb4iq2s7cFoVkABxqcq3F+LZPiGJC28
MQm6J10igOUMlYSnNk4BSfYvowsesW59ymAwu20H2u+KS+kX2Gx6EL6pppw4rDzG
ITXBPFTZ021iY1RM3kuPNlNva68sPKScGKGL3ey+vkYy1K9sBaKiEMgqTN7YlQzL
z1RZAyjv9m+uxmRI/ReLxsxKA+eAMilXIvSMJCnqzgXlgWj4Fn6l/u9mdooAFjRE
XRQHN0V8R59306I7cTGqmJUs9r+tCBaGSjZSOgu2zxI3TMznL27bssOBfCItE7mx
Mco0OJuZzDlbXraXFzyyT+36VARWGCDGaTJdmhwMr91fz3+nOVKxahAOu3Ux8KZg
zBbXPRvuNLf+r7HasJN3i/eRwWyY3QQOX5Fug3Zm38RNXu+0zbVc1xkwTLA5/TTh
SBvo9e7d9hBV062Cq+fd1Unbgx02dR/11Ov2wusja2wuz8zW2WFnBO05fzUQfnzx
LdS9FsM1JwD1OXDJ5r0zZ6r8jXTTh/kW0f0h9gQUrYmqpr4qUdv6NVOqYOW9dOVc
07XIt4xq28p2IS7JnnADFFjbdzgurntcJX180/kmCyO1qnTUy6Fa6ydXN4tnA2lN
8i8rgulpyEznLUFvNA8gRaLtvS7z7AnovTYLvuQwn84CWYOa+7FjKBn6qzl0jbRC
+EdS5VgHqZstXSpxLDBo5Btaqc18eUvRyP4n9/MZHSn0DcQn4MN3bRdq8CuzjUDT
u3E4aievN7ECzgexkew8bW5Y7bEtGFLX6AUe3o+FJOq3tOTk6fQEU8/O25i2zSJe
4cMj1S+z+TAWAK+8j5ysKutBgsz8cR8gy3YskUObu1IxqnlBAKhKGJ1BL9NIb1d8
qbOwuqFsTcuxlPhjdfFqZawbRCEXmWHU+SMWTilWv/PQojdr34X/yE1bybGbzFrR
M0DtogqRuulybFFNXSW66bc0zvId/UiOT/Y5mmk9bDaauqlhyTKvoJDTDZIK2OrH
PK8LlQydf9gb8opwN451dylOEymt+jpKJlE2UdfO27ob/JESV7ah9ZcbA+rGRTO8
jxXxFkeJrv4vM49mr+jDWoNwl7Dm046YjsMI3NenGlS9exPpyKOQ+XRPl8pKCoUU
Z0y8FtlL9xOkMCII0j/1BIStVilOCvBEvfr91SeruE8xPb/DEkcjW7qkRsm86zuV
VaK6TTJRDMeMO8e5ggmfqVjji+EvnQxJ5VFs1JTi694j8VdHnzTgG+AXyJ08eZvO
wTAOq9GLZESWIjgkXpCNX6IKKi2LF2bMEdx1E8mxTNcH/DpeoChUXzyca/dDKSWx
TFiYacXaEdw2hB9t6gp8afdz3uw3Lwh0zuMffyNMPb7azkFOSFtEfBSRvIGo07uL
9nlNYcp9DelZNKk5ea6ND77ITRODFPEf7JgLoUes5jYsHxuLpIRum27uL3gCw7QK
s2jOaO5O53Qp8dQxIA6Q6BUrOBBUDfQgahAEgdo2pqUJCOwX0isVpV5hm3peQyDS
MJ6sbGYleZIwxnfOOjffvV13ykHVzSBbu+qmGGiGtJo5BjCDrFT0xm6HwUpQBwKS
digJycTCtrgdbhGVqXxWVK3aDXs9z2yjGrkd8+sPSfwdUoa/pDeBvNIAKn8vSzz0
DtfI4JFVVMtgstAHajad172Ucp3fXJVvnPkZ/Wq8l1+ncOP7vXpTvpqpKWwQAG+g
cQZYWcrsKJ+h/XI+stiEqFTuG+2vMHKtuQvy4TiJPlpK83x0yVXQDPKbLkrEulOS
x4xEIrQgAoXZ4BGXHUK1IilDm3CQ84aivj+5pPZfKn08j0w46nbBxBqxW8OZlGDq
78yHkjpTeTsNb89t0ysZTnL4svNYOp7rpOnXGJ3AhEW05fDZ78Y8vdd3pbo47KZO
nuWxYCg+5FCOwd+zkLN7nXgeDP0yn7eTEwD1r+QGf1Ycfln/QjvkJyhhntmUAq8W
AOG1BjwJbJN3eVyxTaYHVqvTOMz7ybnexK2cd8YprAptnI6Cug7Y5nswmDf/pOTW
jYQz89hzlYGxx2atfqB+PMag8eM1RzN52izBMT48RsvtImQlfN4Xnxw5VYPvNCLP
bs0vB66Xek/dYr3EQo1XzGpdAwciD09jgnimrjU2/E16MZmjQciSJXuwW/tWuGzO
3FpYu4TcDavZjwWEnb8qamYcqg7XsFdZiAkYJRiw56psN3Q8SECJ5rdQ/3wdjeZr
xlVnx9lXe3kK3mcLbRsM0mManwBskMqdHRt+jD5RtctR8LhygJxLndchk3ecd8EP
84ru/WPzPQUj7L6dM6ka12QcM56pB0bs5f/hkD3/tebq6U3sW2P2l1Nw309nBlgz
d/uoXNaVadmsWPBBkjotzSpZXayNS1faSHzdv2Lk7bZQAO0WaR0DnP3ETlcOwfQD
FZ7fezWluLYA7fTAR/TbWYIRiP9iC0zVGTrO7tCHsRzmR/XxNoifI5kNUbsuizr1
ds+JUgYhoHvPqU+q+eMoYaid8rF4eTHKcxwFzxzTEkP7cShjPssqEGCxFUfRWjzI
wxm9nokmlLcywFZkVr1hUfaF7p/C5KVjTI3pqgGv2l9nBwv8Kv6h8U2LFuFGY6JN
UVGGkBEteLOOgD/dfgrhyqVn0DQqUv7CxdvlEJLA6yeRwiOaNYrw4x+cnQ9uNQNt
caHJhtihYS2EOxpOqubbM4e1c+yjvua18D/J/FHkcXPkx/cIWR9FJXm5H5Nr75i5
dJiRI12QLsW6YnIfLMhFOBYI7FILpF9J8rmNea48WYcysh7ONJl7fyoWWPRacvC5
vSnG6lXnkNhMa90l6c47X+pFpD8exLvtRD7/jWmYVqTdHljDvXfadDhAML2T280l
/prcUT7YQ2auV94K5TEcvYrHZfLpDdecpsGEjqN4Mc85eX4AxlVJcAD8XfjanfBn
6wFjDcdSn7jrIry8oS0ZMIL4tpKAjoQJP2rINk5iBa0FZpolARvXa1wBLp17nKW8
wlQriYvcNEk+q0fvvK3dL4d4LN85al2Kul7lzKlmAk7RmSt62qlc+6J+oCpF2YIN
+tYW7brpAf8mXow0phcm7a+Ri6VXF+oU9+5SWYlPUNocnvmdumwrNIVkvCDOvi5b
tm/MY6sFnMGNBx9z02lxxnTOGDdiioFE7dDLHnfV6C+O+c2uiZ7ySNVudSw+IbPs
8MHINph8DdoyC27353gmvJP70GRvuj5qQsozawYHlIDUB1p0CMa7l914qtmLOltG
EHIJ0bM+OoOasHbXgo36A2vhoDDKurxTVNYeen/Ffi7vh1iMf745Xs7gsIXbpKhw
5bmhuhrvso1yMWFe36vD2AgHhWagrTqqlNHKbNlzDKkyIuXv3ee0FqST8Z3q/rwW
FdG+6mu636HYZzjRh1CTbUdpPjUa6xAIShdTTttR7JZk+CovsCnxr7kxKUu2OIrI
dxAtgtebudGL5ewoGkAh6Y4il/IvspAro6tM61HHWWRtgJiwXxo4DW9QvG4njCM5
XmVEY1Ge5MFovGn6GOnq9lv6g+4iaJP+c9d9NxCdO9nwUuTNwW7iC/55m1cSpiZ4
ei6/CRKBn7tg1fXvIlRBXvfcYnZlzMMSPIqSrdUleI3vm54jfBZTYEpQiLTSHw0v
KTWZUqNTf6+2w+pKApem2ya+oYK/SaIknF14HcSjyQ0LbNrZnAsFj2APICF8yWMp
jKvr5Lc93PwD6S2eSrIOGHgMiDs21I/R5I0LbjE83PM+8bvwaatzfyjsDRgkKZiW
uSeZmIIJkgBAVvMCDPoXPiUKTexj2KVcWtE/4tm9b5Zf0LhnfDXzlpZA1t00WE8B
r+ZF+jZwEueK9GiBrPcmactScRo+vTVL9gkB15QQruTQNQJpXfH8+4uKYg+m2SYC
F/zB/pblQQl1N+WjskU5v5wt9FlLl7Z0F4ZIwzWxIyXX1x8u45S58Hwq6bT5Vzbg
mi0l8tRWA/67st2Qx1WWR7JG69lJG1Pgw3MKPNP2S1GWkUM4upPjaql7rC8JJr0K
0o5H+Qe1T8eTlSz7v/Rnbii+Tf5V89FW9zYpEYp2+CsNA5NZAFU1IwI0dh59hZdX
7OATMppGoPA8z0kKM9DEObeLLFPDw3siMHmS5rXToCJbnqXxbKcg3EY5BE7Ul3Nf
t5ukxicxRX7KaRMSdmvb8NSqc/3Yow5amRkGmq04zsSV6qRtTj1UkcZAvMtaCTUO
GL15+YMlatn6AIxTENJ5kSIESr79IEOuiZLyw05Pda0HB/AyenMej1fCRErB9Ids
Lt3zOM9b6R58wbhlU7TioBvfFQmrUNs/WNdfJ8JedUHjoV7dhWXFwK5b5yo0D5R9
8G6tAzS0djhOBgKFd1cw1vqcsfN53mSmTUhh7sI1Vf79kX/4RaPNSBWXgqYS3wBK
zedpE01YKUDWnIoO9p3cEDy286cVVwQrYlTQSt6ZHhEulw8e0eE0WRjX/zwrCtIo
dkr9vqeHYUPZPd8sIY3JE4125I/JqzKi0WUrVuBxNurIb0z+gWnmEgkGLgwOYkHI
2o8waA27qLKCOhv6WwU6ohnDAeRhIHDM8d2XqxgjCwVx1dGfyPeDWh07N4uHHubf
AqluXW2zv61/eAqPuAg4InxLtGGnqMApNFezKPpHA3FIqHp6S/W7YkhXC248j9jo
fRq2M3O9x8Yq/aqgBuQZbhlC+b+W/Ua14TRwBRp39hzLijip1XHwYWmUkrG1WcVW
UNPpdubQK5Q03Wo4bMpIX8FV5WvxsuXzp12yHaFyBrHWl9XLkux8rrtP0kjbfQPE
gXq8SNGnVj8ubBvASKWvbneyLnanz6e/8sL0N3JQ1IGFE+Os1sFbLJvMItA0641m
eZ0LnyNDHJcyw/whIuZ/AKCXFuDXAOTF7QbOlQRRVvvYvNMw1nOZLo37snjiEwTa
JWki6CYydxl7WmKFDdF3jACyuB+sR+h9scxvxnffrgEZ0XGb45ZcRr4CIsNjLw0X
3JqtB2WDbuvezWtOM9ljTrBQSALltaISo+sSfUaRyti2dBQe4cJ2bM182HPWCbIB
Q+jRhtHS7Yh94p6jZNo0kaYHj1BPPVlf84XgyibdOno7a9Lt2SJwjoRSyhd2PQR2
iTSoeTJMEzyAJ02Footiw8CelVAVjN7eU2TSCa8ZGBX+8TQ82Si4x75yEufWR2ja
69Nf1pqjYRKGK2GbNBDuD0KSMWFhCq2lvWo9kLPENY7aIE6AQrHEAH6U9I/aZdTS
w802sbB4qpI6c9HscfI41cuz0pzIXqEuKy6bZ8b8K4qttYKGivNLnAf6BllKnvQ6
94NTaHGU5FQBRdY3pKaeDoR48uEzfsb7xDJD64UGx7PJETHGo0MMTOx6M2WQaXg/
+dful/dv8zfmCxNLP6OrAgIrFmnFsIvcStoOAcAHHApbgot+j2DiPY4xKugHhdTc
8qZFZFgMjDqseigVqFjmRRbm867ns9emEaZbaoL7BHNsKa+SVogDzvgvbyUUYoYK
nmzTJnKgy7dd0H1rwsVCGCW1i5FMRcNXhoxf6K+uB2V5fItyYNG3njrMiHuxak8L
KqaAdLqtjTfA0dOpSFcAXY+SquXvlKZ2Xn7QHzvy4gYCQ+Oi//I4FDbIycG6DXFU
Wfll7wB4K9WUtfQ67Xvk4qcAu29NG76N7dlb508HJcNjRNWJbdGBBN+ILNsdPPxt
CwjtA9AfqmcuPTn8L0Gx+Zmm+CO7zj0wf0crBiX7GJkyCyuVd5JK2cngYvGju9ug
0YSijNJbcVbTT5y7i9aFUUlS7O6EhFqmnhE5Fk76tQMe6WRyKxeAMfT559dJLy02
XzU/7pVhTxUwafNbcwNGo2Uf/+L9P/8T/cH+sW4zW4+dPp/a2TgUlSO1tjaHqQXn
Phk77vCQqldmmBQ2zzy1vXgCLXh5ck6uEqz6oB1WseyNUvQAP7RXfeeHSifOaaLZ
j2R5IiFupFGqIVEb6QPEzLqZgE3ysLiS7dHwAA10gejoGnmV+Rog48SAZh9KVhwc
2gxxgSGXuQuc29GjTRmYQOp5kgek634bw9uYgSZC6OGqRip2fskFFlXjfMM/KuMo
tRWq+6lWqR6uqRHtQ8AqieQrRtv41hIsAPHANAXWo074E9T3bVkZjLsvQM7/UPE6
6exMHv3J/20KtcW1UAHF9tI7phjkWuWJnIGBfDUqAB4u7dQmHomh90c5MVJh7Vgn
Akkl7omcI7eJy/MDGAg3OZjwGo9T18urT4uGAI1vCygfU7KquchqvCgmoMNmhdlj
DcJvRWZDUM+PC3wX4pNMUCkpCSr4fuKOMwe/B3NpPJp9l0kYH0PRnJo0UnXpFNxJ
F2jkEgMHGgDUgwUuQbruVp5rhnvWQz0+xoQSjemENhgm23zF6Yjl41ctlQ7jzEDz
N2smBRPt0GlIt6aZOK3G6tfq7RoTJ+XhzQTu2mKtTJKkhhbrDXiOWRie5kcp8lSo
AxSVkbwF7dq2ZBlVOqqoELi+VvpakcisN1K3NuYuCNoNNUGjQbae7dNxLDEtvSwC
1RiLBFU5JJCxUE2CEl7URGCBzUh55lIMli4OwNhYLlBBZyAM6zx8LiR0b9fQVjSZ
L0s4tclbMTd0fzV5pxuMUA6qlObvrg7RVtfeWRmPaV2hRf0rbfmHU7ASKnTHgxb7
/5XmjownhGx+f+xiwv/WQK17Kybrj2jSCJxBU3pSp8U/JymCNmz2rIVdZMEWjUZf
uzz+agfWpIk3HHW1HL4v98F9AAy3d78BNgPpxAG2ahe8SDQmo+eUxosMsyXAciwI
I+VuexDw0GW5mEYC1OFnbGRL3VtesEWv5/JSadqmpX41D/hKuaqTZTf52ffzDFub
YqHPHTFIwiqpXVc/tzjjFIvYUa7fQkvf7fgTixivgnciRUCsSaEjkVrP0Cqzoeex
anQ4qDXdEjKYJd3glGpDkcTNcjXOG/UDoY8v29qcHn82IvSCwwPtn8kZe6m559JC
LA/ylD6ALWeHTCxbmsNwh8YoUBXULz0cOUBC9w/qi4JpUIW9z/tN+eWMdkGAQAjA
KLDhl/cvJ9LeieJ0k78yOVZx/9gC780MVDflCWyzkxe+aKqDTXU7Xhc/zVcEk0H1
JwT5de2vB/RVij/aixMMRzK3GxATq13oOjkZIBVqtpxaFkPdWzE7tBZcDWLwlHpV
lX3tSDVer6B/PAs+HZ+RaCi3wxih0bl6/xHY13E6emTiINUR80GTZHCPxPWg5j5L
ZEADSQbWuTBuqCj7W80hQqIav9f1FM55Sm6F0/Y/OKkjsTm/K7vd2XO8zJK+FdgD
/A/EXYAQR7Tk8HIYhS9KhCl00On0EVsK+AKcm3JFw95FqbVu+2wgLkBk4ZP2BmXV
HGjPk0wCmhyT6+vaP8lz1HVIgdUvk2gFFm+HMUbvZmRTkusX8gYv53BAXlp8rCZk
HtEPM+w1LlJQXpuUTuLpDpMKRxAhi7tcpsPT3xe9srirAiY3ksTfOLWzVRTpRSDe
4U51qhs+ocMuOvIN1/JLDfw4DDQRj0UtQ7Zrv7nFHcd5T5MIRBFrwdlVvUcgqhwO
fBYDDLfP1V0hretj7PVzTMvZou2EuI/BmQzNn2PRk8EW0cpHN2HvOloaKwtKJ2WC
obi6/kE8Goq4cnTJs2x6+aewPBe7Oh4FqOoLSb/xkGHMCZYArVGJqdCKl81OKPmD
1QsZPT2F2bEI1HQleFCXxFn1sdLbXMPq7Q0O5xGMtE9zQEZmEcBKtREHy5AOImVu
GoGs07A/Q4kknHqCpI5nrsSYjZ4VSoFUbAJHj232wPbYnetGbSVLSfsIphc9UfjQ
ggNIjjO9RVljtw6aVuXdmOlByLSjZaDPZKoDJA0mrQejoSKmvwCed0UxtZZp4hm/
UjkGitqd0VtpM1F+ERkvD2+zNuMZ//BedeH9f8KvqzDRLvHoD3c47yDmPdxNe8HS
EqNv+Jgw0eXDxLdUm1/TKP7QB7JB2kGrB+looWgv3u/Prc//Ibv3kMC5d/YaCjCA
c5VkXr33OJS4QEpwX6mLf7CyPyjKfbcJaETZnz5nXmYT7FYe4E+y61ynyZILx8lB
mnK8QNzQxtwEMRFSGf7NDx3zKYXtUOcXLPrjaiqYj7GdqMojKnpEfZ1LVKXYDanj
uJg40pYp/jWu7/qoFZC9KHlIJX/JUSGmM6W01drwGEAtYhWW4ssb8oB6ZNweb8Y7
NqdP+lZJyFPweVjMI4UkiXTK5XnEB9Torve3XriShkswtOWub1yeCTMZumZG38IJ
dSbJGyin7U7i7uhj5msXrWywMtOL8eYUZ0Z4jb8vk7mREcobfFKCwhIst3IbEmrz
6NBAUR6JHfBYnnPxPUcsNhd2+gSURmLYPVJdgynXBEZHWed7Bob3OW2kzF9tpezN
cWDoIl2wWHwyPg+Wpy0BvklWnSzZIoc+qJgsiAeE0UnYQ8ILrFowOlpzcK3S1iZk
YpIWCBI/r7OkY352bo53nRCLczQ6//cZKdN4bX277Dh5af3SrZD1ztOteO1MsNAA
3XSOioQ3J8efUD+CvEnvLT+0MUVsNPHFxifgBp4cgZtsqDz5tmWb8+7qz+rl6DXB
CCzqh4xx9HX+acX5nliMkX8Bb8htmX2HQniF8kKAQ0Kr3+BxCxgkxtK39u5jsW/C
2xYXn53AG+EUd1t+5oNz2TRdsujejT/+xlrBbSw4m8CvDRA2oSoiPXV84amWTcil
ChQMb6uYT+l6YayT94IZz88G1wYGGHzkS7TVuNBbj/aQAVmt3B7kDnOe0AUAVLNb
4yjzuLbjOuqzpbuTAmHlGPACIBn0bl5kKBYkKUeoFv8fwfBLF5i030afNINigahg
aZ0pLroKcIN8jK67eUZjOjXX8Hxf/8CBjIY74bdV9Pp476CK0ssD6l+YMqVxdX4J
hrMXMSL3UCGHo/X+fXqPtnVMc9AxJcAAsnjWAUHa3IaG9twg7ZOaHT2sp7ySmo3r
TuzGNqWjfiqoATYpnj5GS+ZhuOfrQFTEfEdoolCnmAbnQzFy6ED1eyFSv7nbM36b
exoIc9rZUeII7gmQ3tUYOKjiX5BZ95L5aDMiKaIbRkQT3zTohGFS5WC8El4HaB3Z
1WqT5kWcWao5Fj3od00viIw4ZtpIsSFBZuvkF5YZNbeqinkLajQfjEYaKXpEFYrj
X9utlktocuL6O/jeyNtMx/yQ1Zpec+k2+fED3ia6hjsLQ8XBp/BExxT4wVZ7e03M
SWgHqsSsUJ5ulCoJiXRLVFTTYrXTOybmPiVYq8sLrGwpA7OBx2OtjLnN0aRkzhhf
ONDy+rYFCpli/DxxUB0Z4+AXTc+N5eLYK/9dZGzBuMFCyDvuIjzl1pEz2CGP6kC3
glVzfwmfwRTePe3WeasEAxS8Xi6XkJs0Iwkeyv+E+k11qqLIELNAi4SyrWMzXr6/
wsdc47itoaeyb4/rhCvnaTtPK8soGWTxl/mfJKkH98wSJGzdFAISoAvrA81T2D9x
c+nc+kQhsIEuLSyYWL0jSDwE1XJ3a9MM6KhIukjsYsziioma2DQpTkO7oCJ/U+26
hg46Y+8VPjIODMHKmxkxDfMIUMP8ojSjMdYme8YXZXveWopjx23vvkNEBGqOBwWz
TcfAHOFZWThRFDcWbsliQUPJ4/FmFEMG2dVKdZxUb5ZEZ+Y50iy+pPwTp3C0wHIA
3Cvp+Re7OfLYDTdSOdsyMOVqB9zZifenmISS/IYQGcMk9/bNK7fueymgTBKcaS4i
I3/r1Tl3mbod/Pr5lyWadX9TbJYZCcthnWInBfxp9TygsyJ3BGMMdCi3qRgIVNJx
xVXdPLpfw9+tXWjMs73ui9aDYa6x63HBI3xNrvu3b4D9mleJH6DTo48O/+txNujK
MawVwcxOU00WDC2uo90yNqLuL8e9RmJTtoWlve9SPssX6aOPWqAM03VLZxB7Wia3
ek8qzD+050uFIQlQhA9uMMdo7JPhPr+likP4fBOTGshqASf1ZaWKvRmd4qK6WIVd
VTnCta3yrvbIjNNXgXeyIJh3h89MUGW/s1tVtVOb/4jc1UVdNbw9ottLjGJ7bm0g
ltxuGdxHoacPgZjN+APEh41dwX5HUy/38WUGnMiIQmgeT5hfX4fmHVQ45JEUXAIG
qHXTIr0bhEojvAC9TEG0Skhr6TfB3W7BR4zKHFr3mo5ZSOmEbJs2kE4U2f9Q5a18
TA82T0k4gxz8mvpyW2Udb1NyzSl8VmocGaPoTfeol0SqzUCUzm5rxD0eESY4RLr4
o6SIqCeNbvIT8daMDTP1k5hircQuFADEj4YI5jU9QfHBADFwMonBzgCbSV+eGCF0
+Xg3hVzM+bzMn7dJsJXQ59XCVR3b6vTMAQ/cZWuq0fSOgnpsKsr5kRmzVb8C49gQ
BgH9SIL0+/SvcgFxkFPckZdRr4rkdR/I5xk6xpjIQZkxe5YO04A5rJEAfIvoicqh
n31D3XYXW546nSwOLvQhQyelQzX/Pw2Eew2saznOxdwS8eaA+eCOaXWjt9PEkHud
nSK4wLe8uCWItAFBZdCQqsSq4+QkKP+ez+6119ZEPMN+KLtX3RPeFwpnsqG3d//b
w8xcZS0vX6ZWn/ssKaB1LEAc57WUqXCGyrMdTbDtV6bnVti8UaA77cj02vu9CYsN
l0rAnwaTVejDgp3EdsZxMptPSwkXXDNBi+eEXW5r8vA7WYdAsMKUeoKOF6aNlr/2
5l1VBLfWIare8lz1hc8TWhvii9yYLtmPpD9bzKzvlHHAVWyWuuPpv/rDjnW1AjYU
x+bnpY3DaWoKk7gdCTExRc4g0ykBavKPULkDrAhvKWwvCT1oQ/aQqQv34XC+j6uF
Q72M3lDRT/XfbsVNcDa7RZIBmZ8IsSFDneDyMjJKcwXbZEjlsdHQpHWAdHuvEDPU
OxcFC1QplpkX4lAStyRVovJ1lZhqfipTw2qbla6c/V4TEM8ZEht3PAnoOuyqaOXT
UIpEKrlcfOuw03VT5yO1aTVh17wcRZA02DZfzs0H5KCAGdaPQDB7TgCz+eUCu13H
5po0H94lChPE1251BN82EZ6L1p7IGaIdyUGQaOIGr7iHPA0PZrKtcqqbt1QWvsHC
RKmJOi+gSv05SVmTpOAwPmvPVBsEhGwHDCbUiOUWXdUkTivW56OaXNmCQ+3N/GAR
98qILhRW9jagN9BDbeoSPDL/MGdvsA3OTIRpm7ene0z9hpvIpSa1O5mjP9sqZVVl
/sde7LQHBL1OAPlOwaxb33ntkAnfnc0HNjNxPMWyV2lHdqeezQkameN7iJg1aRJp
7j0EaV/3hlhDRpn8htFprJO5brP8c1gDr2xEwDf3iNes5bmt1Zc6Vxi2dZ0cZubc
5FHuxnqCtmEMGSgypcamkUDSUmHG5M57phqDT68q69Q2Xj2vWXQlhmWSw9EtkAM4
UYAeujTcpPaZ2dblPMOe9pvXAgsHJ+J+x1ubbllf4j8kt0sLUjmEAqgYe/OyMmTz
qDdFGctmXC+QWPFIyr6gQlaw5+No/OqE0qOm5nIQj3mz+HnHu+3Oap0vT2tBEDqK
+gruIac2TO9O1e0UgGNtoI6ZgcVP87i+mQWjtrrb1gKPEu1JBnfy9owEDdSGJQKd
naQY3MahHCL/go32sTSajHBcjIICzNLaw8JhtRFqTsp+ulJeHLlpR9nl0ChY4lXf
M0TooNhnQ7CsfrKzA1a+3yA0QJRdPbaM/QQRitSR1ky6EdeJD8eFE7N7hLKQXEir
8pnhZ2aZzvN/NSAdMFKe6f6kxK4KmV7KTNPrUcczKpX9tTr6DhkPc4/HiLGxghBM
ZkZ4i/Dh/uyNUsKKyRzygzDNbus7sr0PZ5rE8E/2y4NG0/HFLcqctIwKU33EhVOE
VgoV5pxEiPT2xx6zjGmrXlKf+fNqVj1Wb63XA6KCiDEtEeSPdNXpfTPTKycSnzOB
ziOtAgT972Yss5XuJpsHlwu6n7doBjqyCheUy//j/nLlGGrnPnE4DpAZ3Y52VlG5
fdAzr7Ie/AEiOAWHPTgAE98+xwkYxg82XgOL3foHkrcLgALXXBi+bv5HPmFZAzua
SRt3NsIQvvl2bFy8FWXvEx6c18uZ2llqKsrTHMt/93ZuMjIr5+3etJu0KBEBPOeB
pDloofQJOUCJ1jYumr3H695vdQycxecbuYQ/p7lx6VA1DsQ/7H43NZJsdm5hJlFa
xIQgKiZmh/LuS1PXtFe0yAzIwpT7dFKWTLfflcGkq5TRWlwrIfgUteFUFbVyXZXr
XCqoezgp+Aqojnp1mpAiNMv/4zoEIch9159TupuQLPqloqQ+0cqpM4/L94EpYOxs
zE6LNRWsrmSHZjgLj3Qe02euRwy+H+lIOm+LzgzGT48Zi1BWQErOoNOq12vRUsEr
qFbJOGa/kmZ5ccsiZfXU3Bad3iQvi3lzmFZEwB0D9/WjsT+eONHkE+pkThkSmn3A
DD27u+0ZSZSvPl1e6u200LDibducjGfrUoZ6DXPN6McMpwezTyF+Q1hNB33J0Ryu
seqGF4bsLF7j6WX8sZDprE2SFzNtFTKvpkt0Kb0ejUBW2IpSGOrgTRwNMUsJnSfu
Z/dr/p4ovV+OOQgbBhPodh3rflhSV/WyXNRtPXnFQSd6/L1yEVM2Qh0fmVN3sNZs
vNrWL9Bm4Sp1YlcYSVN3I3Xq/OlyMRXGmGgNcmD68hs58jl2GzVIsJfq+V9PJXv4
zOE/nQiryCIjlVMEOr0wfSl2PBw4LiwLLq54Y7AcgNIW38OvZR66celd0z1kX43h
OsyFVNBMt4DutReWr5SBwPd0d/eN4XhPf31Wqz3GOeUF+zQLAbqJBQHe/NnDOd1u
/iGM9qYxStnTU1NrMpJqdIPY5LlETt2Y559FPl1bneHqLBHAq+cqC+uZdg4eMOCt
T1Yw7vU86ujklfM+94laZtILpN07Uk8JyAsjwQ5REMxQPOY7mGZBxzdPVdo8Tj69
NIN+pxlfdGL/bgOVxVrig5S+7VLNJl/gUzD4mRCzi15FkQD34RhYvvVx/fi8CXYQ
5hgDPBFIndkrXxeIRsN9dWPSVEjQXVCD8HYa/ssv7LUGEVdEIV8Oy5xFhIXJqDRn
r97i0cwx7IK5mO0HKUO17xn5CzmockHh+EN+Y5KkhPjgVJoZfeTFrQcMPyoIbMXb
ZLhPluN5NxWH0ZvkWg4PUX0HvP+RU68TdAPP7lDsYjrGzvGPkSo4RjuGqDJxs6PC
7EcjY2pkJf2HssG3tNj/Rvu76VTKDl3numFhqnDvhJlO6YBZxFjv5pU+JnxVH+kv
oZxteFMf+vneA0JoLTXIeetSfa0ebF5vslGzMEqirQ17EhaRh5tf8oi7MciGN17o
VRW8zVtb/Vh/XsXxFaxCkZva8KUCebi1wwv57vt8x/Aa2B50B000Tf9eNh/bRmCL
CeHVT74aOiSmdR4jn6pdsx3wTNRMpzY76k0UrC1TpD7nHUK/MqN7z/dra9R5+h/h
FRTD+mWAR3Zt1oUGpDPAQ7Qol87+jdR49RVDdtNxRzG1wQLIa/ZkIKFQ8FcdERTo
Pen9NPVfAGgUd+ULpqRlepdb546ouGg77q60fIS+B46mDdJedQj1AMC9fqu+05OL
CgzTtXnM9cYtNUxMpPuEaz+dZCHCGMSRlQ8NKc2+rmUR+Uenot3BoFa2uabJgR5M
NNLnByL4ddAQfv3XRHH9/G8Gde3LuBr3BicpIlP5AEv/hX0uqMUT7+sZAq6wIxOZ
AwQSjOGY3wfkHz212MDxbeyBAq/APpLVeqYJbEaYuMElIMGfWCLGGeBPp80E+Cxq
tglKUaQ4bv7Ovi+kQF9DPlzro7Nm4379YwgT7lhODsBxq9WuwShCuryBIt5w44kA
rzG6J9HkJK+KCL3NvB9yD5l9z0YhHWBbTpiC5nV+A5yj0jTC6Ja53xMblzedt4jE
jYTiHiz9mqc5dwYkJfOWgMpIlhNYl/TGJZfBy5FNfjehzmsQ7JdvXSosPJ5AJSIl
XhWZk6yt4J98jS6LoZcgG4KQde9S7HAkku6U6sIQObaEYW16rEFySu7babezyRDH
txg1uYaVR2qxvT4rO4hTgbMk70L37bYKq2jUaiVqYoLkfsgg5B5QSDUB+FwWJAzu
jxvbvgO6tHZvhR1IMR8H68J/mZGpS863c79b22mfCCSSdaW4nNBpiAis5fJGtPFD
ZmxNWBShsES+bmykI9g53Eh1+3gDj9y61iV3vX8MwGom24JyddM7voFbOsU4O9Mw
7U2SDfzaBrKW7C1JZ4WKmui6pa6x0a/EeL0qi9lNJcCLhdZz/+t3mNRVpkxGFana
zfB20tiYCCgtOrSzR8IuxvSoR1rKmDA2c0Dsk9EjqsdlyeTqbVo31fnLEgYLI59F
XonNlgiD7xeTBegIgdfCjQdL+yVE341wADhiGn/JL6j+/OVmdsX78jYFHf/Qg76m
8vKQ9ZiTGXH4sNjZvTNOchCO+TtioS9784/qW9RqXO/+23WdAf/eFXLPXt4lupKU
30uGNYi/s+ku9QFoHI0hZpz1M2eGSOJcrv5W9hPJdQBX+3YyIb/qmNZA44xyexYT
f90VGkwpmnmdTrOD7xRc07gi+TTn4NOYLUWRb8/Q1GYKrKu0a1Feu61D3b6iG4UA
jsE8oVloQSfymTSEqfo+oQkUXDSpjBRmzYP8fTOMvAo7lZj1pQucbdfxT+V39rm1
/fWbzrkdTRBcIvZi2iJU2sawikGQUZoB3KGw6KzyYr8rqfEhwp0g/fcQBsUEEb5V
gGgurSvcSOibeaUpIzR/9nZcdxm5E+e8cohVIcBua7R8Kps22yJX6wGVCXYqBoRE
fBJXBjFSAcJ0BLb5D2nrHMq+gqwLFKG3IMr6lg1chb9FSdtiEw4rneaqUSrAIUSt
hu+H5SCr5ApmPjqlMKz12NtKrfudDDbjIG8eoPEeLxJc3VuAKxZDtpSB7q5SDUF1
396csgWjzc8suD2BR3ickPM+KbwzpWf9MgFc9Y1TcjAwz20u1/XpJiQig5K0GqTO
BcHOLsH+0kPcMAN7iI3SWYYnyS1Av2Fg5MnV+fOUripcwcZd2ghxVnUxPeztkFc3
b4rF5CDKDXJdDffrFADFwZXDq36FBAQ4tBpxBG4bIrf8KaeXZwzKMf5XtkENBlHi
aeoIASynVw3MuqZe55a/VvZkHvvlLC/0HhEU3PxbR7oEY0wRAExSSH80NBU8YM6O
hB/nR0wi9UTSrWAtsUPC1zCumY30ZBZbt/GmnqqQPKFE5ViX8Zhi7aMiq1d8MQ5q
AJVt1u/5QgiWo+hm2htmqA2kTeOFnf6v8I0AU1adMfBNt5BJqKSrVP+RZqdluFhb
9A/bjk0o2uKlZuBLxoVinn3OghCGlQjAwXp9ZKydwPIYYs5IRtTYyjEkULH3V1tc
UlyMnWoR0hJTE02hiwGAokp8r1Db5k2PsV2nDY2FFPoXEYk4ODHAFdpPmJigY9PT
0bJjqOswmVYOxanESSDQZ4wtjyMjNvTU1azqFX1mSz3XU4T1cVSZsD39ioE4TsHu
/nL0r0a3A8cVWVxZ6f/bqaUp6L3Jcgk08K4pH12ve5OwdI4WlzR6DTQybMil9yCp
omtzoV7isaWcjLDytUoWABZukWICZxGBC3AEM4AmF9MGs05isruv/BQlKC59LBOg
HwMbCFBIVB+osrB9QTmAQsI4PYkeUNPczbsSvuq7tPdVWaVLMRpQIYweuMhG+pcC
X8M8QwnZN8CG5pd1FNfEeJYW5WLNf0PKfM9qdgyvcNa9+4yaZ/axVRep2RgiLNJI
UZzF06JoJMoxO/CEuIZl2Saia9m3raA9uS100EFb0bHmmhF5f6P2ml9poNW5AsPC
eJNNb7RWHm6WZV1DqNXI2rRCm9/+pV/nD93d9CTCbPfmKYyREx22S4OjrCatqR+t
VPHEUR1p+CyW+IMLPQtcJsMpZadpZxdCWwrrjQW6+QaZxBUqvSyWaucWUyL1cU8T
cY+JxLN2fjLgpVX83toKSLn0d5py98YlvbGcjx9IcIAvQ4woCe4oVfcHRU7IhyeW
K8MAdt8aNQ1r5BGVaV/VcUpxS3Fiy1y/yKSX+KS8isqmellEnD8YlOvdpiEWa0OA
fB97CyJzGXVRGrqMsz9Ap8Ie18BiL5pEo21cKnbGJK0zF4jf7s0cDzniAA0uEo6x
nPOZMDZgmnw+/sfFdTd81HvywMvY2SCZaNQQCE8af+phHiXEwdgNMF20qdPorGtH
mFCDCO+cL3UYUP1dm1isKXkYfWKAk/v7qTn26Vj7+GJ9ZryZEtLgR0JRmv76AQie
3h7Wrn4gwn/xq2j5aysqzpF0RY0LhtYaY9u9OQDlhv4pbVIP2qInUBQ2dfGo7Gw7
zEUlEMlq+NA16dEKnRd7Ki/i+X3fDd2TSer5/kvUKiLgw7V9pdwWPsgXO9pa/oW2
/D4gTEeKKXCXMqQ4rMUYd+ObkwZ2X8JzoPBiW/3oBZtYJLRRMxFMXuQoIb7JXqnK
+FUx2K7LjbRGgVrmJjr3B9zNFuYMD13DnKPDzmAIGJghH7/18QUYW/aJ+zyLQJbs
WttFW+6jOjLIx9HQczcbcG+1qLysZ+nAG5+q7MPag9JFWfxn0sb/FNPPAM28+gsJ
Hx631tppLnz3RmOuLW0G8gsSvz0dFiKe+wtw9SoABvDibyTb07RvHvuEgarRjvzO
cXGimy7JHZoa7bEBlNZGNo6ypfiVUSHtWxDn6tqdMezIA3JOa+2Hb0zDFg3Rw15y
okmZ/SnYi/3Ca2jsFOvVSz7FVTik3QmM0mlBl1iLxKbbGxuVUVEcveYb2MkTajS9
Y3fEu07GeQgJpFAB8UabHeI0d6fOYG4LgWu3wIyzinxY2mWgTHYBMwsDNwcUf4AW
4NhbVvf9wi8smSSL8/4R1+ieBcogp7ZnX46zK23Wv6jBK3O04q8y3cYUJ05jn8Px
st8q2IJDGreCjX9/WHRYklXCuVo5UMTB4Nf9BJH0VvxDP/Z9l4EMp+BpzYRjNxq1
nYkyoDYyA67JYlpXRB60xT3TbekNC70QBhOGcnL1AY+tKwmRfcw5qW1uW+K+sDlu
GoSRifax5euP+jtQVKivHZ5aV0RfYEhjWq2dciiv9ew1l685rcJ3amoL6jw2zf6Q
AljDSYdNKnI34OgmdLpkTfCzin+9CSu93IjIOiLdAEWS6FuxZWcY3YQKz8fxPgIe
7ghBNU8gyRb7LTemaE7BYUm+Vy1EnareuKlN4vXqc719RngeTIv97nkOSlQnUJWN
m2MERTN4E/pvbco1Gl1nmjqgx+y28b1hFuMOjFybLVWOGdKIZ9WlmHhxIVquhEUj
d6g+XFNchfJxZzlHNF428BwC4Nnx/HxYQBxYmn2fAh7p0iv5O7BciqtEFOuK0EkP
LRHmw3QTbsdOPL29ouyBAmpZG+mHFQ+ooAWiOQWPQef1o9GabSdaTzeIN7j4/QwH
hjGFI1EFWS3gDKo/mW3pKm4B9RzkbjwQqEbBVR0WaUUG2d45cln7QAVaDVw+xzBX
XBIIN8CFe58AI07gf76YfOB4ns+kzRYA/4YKUgViKTVEC/U4Vy7ybKAm9GJekyfz
2W1BkO7x/sMo1U+IdEJNeRzbF+243KuO9Epvz2jPhlPKMwJACFfnatW7808KiLJc
2yi9RzzGEtVe5qjchiMkNh0A5Rwf72vGgnnfGvHrg+ymjNp7LIfvlDszVxuKdE0s
OXzuSlrMWQGkKBUMGO89Cft9D8hqESpXNJ5PLxtj91sjgS2YHQ1T583hengwBSgv
e7PSl64y1gwuDkMF0yvSCl5kOfy7I5w6I1FDRNXsx64dBW3gJXbfQfHgolzIw2yK
da79nTRxCtLjHKzZ05fW2uVy98bx2Stz1EIoO5c00pTYd0BlwbB+fbYxo1IkWPVg
HYgeakxQmjlXx74k69+cGqmCTxVCjE1pJW5TFZOggqWhDbpiIhJOd22x+MJoQz2P
aEnC0n31V+/vCnc5Kfr975UwfhAGqnador3nEV837ZC+rvKhp2SFtViP34vWG23H
HWJ/Phti/m+sthODSNx56QVOxKZBCU4wDp+/Z7VJGKSHsbnCH6Dw5R6DEWDg8Rt8
UKpAfj/7TxCylN3Gd6XXP7FEI5lqzqU3OR1QBp/zGwMLIOqHyXX2HRq4IOzq4l4e
lGbxlcuJqathXPUjV2oTfsIkFsf9AwoHzpcPZQOQMBhGYVCtraYZjjuzaBv3eAAd
YPuw4aGMD3004wgMREIn9K4LXRNmw1dHumDywPbIEPJDVpQ1tQUSW04rEJcL3o0H
8hkHqgOX8+UGwthcvSO7HBooEr4y4AwYdFmQbORHbhAvN85Ys+KRYGpbLGLou5VR
pY25A2uZ5bksxnq/udKeRrYN9aJJICElrFI3hivGbf7UQPPqAklRGY0lGreS9DPP
1/xIVxdwTqDl1GCHNJUgruAaiPatBJ3R2JsI4EE7jrp9RFNDnlnaaRoCyYXQOctD
fXn1NswIZlFtdoYhoCr91W/P9QOGHIs2HpEoB+KQcSfOhBjNkyZX7tzej/08Ilip
2x1KPJIiAvzjYyBuoMOynfsM+r4xNdt28qAednRxQRKc8aIf+L/lVp/2aUQt7x+s
gYKOk/KMplyz+KqEPw2ZrDPA/uSH53+yqdFA8vYIywF+WPjWcvsOmk2dFqUrl17p
pcBkxO0w1GpK97wwKOwNOw7S0u6vHRJtA2Z3fRetwSuVMMrpdhAyILq+uRjFizxT
v6qF0BMGZaMAz6KAI5ncRMdOBs09hdp66U7E7bVNhQ9NmXC+qI06YTw5MVj+uL7C
4jHLt1Z7SerhtN4oyXg5G4GDK4HuwN6TqeoFD/jVJFrFp6dMjG2IClbsj2Qq4hv3
LKQbMRjPhYqNy/C+Q8jXTrmlu9PTI5G94GB5LfyJAlZ+iHE12VNmm2USCMnvJxLg
1SOoNyOeLpM6T22hh6z8WszKSm/b3J6i7rNb1jIcFELWnOeUXkUNoxBqgyV3+6Xe
GK1Qi0yN6k8X8ZuLt/ysgRT4Im12ck0yGjwU1GsG9Rmd3XwnH3Lmz9F3QPp9cd1h
8H3vOXhAg+NkbjkHFphQw0bBxuyqKAWSc79JtvGAIpjPeX5+IrUk0ZXfmRqkaleJ
ANqcbxlT3egzcNjJNpMLTMOfYzhXyYjIwX/8/iNn+nNEAykedDiREWi8TIjL6m70
68vW96BE7gOwqFlePNTJwKKLyNZ5N7qr8BY6iBIWHJXNYoESuVLD/+MRuPDk8kCG
nqX1XcDnoSHKA12r22N9BbMUIlhWmtCE7ZvmYXIAmm78iT/4ztSaxL7oytK/zaTa
LeB6Q19Ut98RgrsyRpgZAJQddn4BLeGEVCZyDSKnyBmDiZemkUYhHaOjS1zXbkVo
dfkVU4B030FedQaNiFIFkPNaIbQ7L7MU7YDgAU8xmORKidldrl7MW/YPC4g0MfMp
q7jZGdwVeDIlTjOJcNpdwP2VzyMLkpTibYCQj2kiPE+Y82a/fXNyr3PJ/60PO402
yPoXz/ZQ/7si7YG8nlcBGJSXyGmQwX+LqFzQZYlUcjWnKKlvevnfaCFTQ8EZQz7G
UL2DPhTqBVaNVg5Ukmx6P73816qJMFjTUp61juStDXpkHyupMxcIqwymgyIvMHVu
I7HoGO6oC4kDdOFc8GitkRW7A4X1jqjQ3ZuJej4BLIuIWRLyWqUbpnrCSOz/gYUW
kZpwDgSVqRCAiTrZ3DdwvHAQdKRA7iMs23o2p1+eysGoEn8ZpZb7DglxZGnMKahm
mJBsLgsEkdY8DU/aPCPK6T4s69l0HPUkqE3oWEq90v2LUd1vMItBa+Qkr2Z7EUqs
gPFEAz/akdzgq85ZUvlFLBecnMtuEI0mSambCci/sVMn+X7i6wng1KHWCh69XUfs
5Rmnvwqv3uWKk85FOU1nPnCq2T45M1c174z53Hw8UrPyJTMKJHhE2pN+SYuCOya8
tSsXCdsLEA/48jyv6iSk50uws4QeVbmGAw4NVMdiJ8aaTilpRAkj8jb7madDdXo5
CWNawBm9EYnDH0dtpQgHpC7k9OzQByZQcywxDboRjPNM/Xjzjp+QcdFqdnc5wmmf
hstGpUG01fobi3EyEeVjB2H8kUFkz/cfBnWIfvSHCEvwBjyyCkW0A3JYxVBsMEtn
FekRwq0WRV/JGD5xzXuSWtX8LCjoLgz1Y2rGAwImdrOzo1ZkbC9oz/FLDXsZmSus
hid41Dt0ESKXNBsUfOzgiph9A1fV2dzpHZxFT4mMoWUvAWIbb4KJdtFyZrAMTOUD
ZBqK8oPaBMPPYePp+D1xcOnO4bTna3dNj720rDNROO4utnhT6Z1NDjffYliwGZU5
XlF5Lurd63cS56Q5UrTO9lLsV8HGT4oLc9y+0RN9zOJIowD6Tuig+c3hAE7h4rxg
BmgeifGFnEKzl0meO9lx0Ibbg2nYmuupAtw0OUPfB7HO2eVVww9+ShS2xrNORelX
RMREUfw8q7YoE2G3UBbf4lME2MMzPdkQ9HFv+Dqy4clkSAeWgDCYAjch7JQtRuKY
DEOPoqMJXcFxKBojoF5F6cCGhz0wVVb9YYaHF4wetgxjaVqyA2rp+HywqWHBwPtt
XQ6Ssd10fuZcHdUpxkpCBFh9QgxaqVEPgtnAO7+/X/NTpjGBvu4zRT5aG8I8w8iD
pkKYQSkOCQBof+vR12IrIgLWv5E8dMdOi5NE4wqQjZn9ltS4Auo/er80WxCQT3s2
pCubImCjE+FP6VHgTYHDV1bU9CPTsWiK31swlthUk7cdUQJKHv7VIa8Ohn1wZgxa
4QekFJFj6QSDziEH5KRtSyUOlcgS/8102lDM9H2M6jn3oIkfPJIj807cNlqunX/w
JqjILT+nU690cbtY+D7V+ArTL4LIUX8ymRmtFedJrfz211DCX1dsgEcATFps9uH2
EgzWl1un9y/XlpGVWQgcgaZSzMlBSB0731rnByZFwuOl6yyG2ErIxdgUZC4KHHkx
aaJaZ1RVDi29WrvMdKA5f1O3FnGWRaQXXuU6HVo/Mf5Rzd2yIuDhor4tu/Bch26D
HYnrhD7JE2Chxq0HSm6zHEbo0hLEOOjAUJKqFMtsYUWqkjfAAW4CSf6h1+DIOpZi
u5ZJFtS8pzMF9PCS5/kYG6YByy3CMCV4qnfUUVYUF3pZyakYRIPnc0Jtqo/e3Zao
Iiwh81h/R0iioHWXq8dyyNZTNitQkwR47gfZSS9Ck3UHHyAeIaGpUgUscIElxAER
JpZxn7TKqV1Z/oRfV+GUWRLnS3RJa1zwByFRMrhTiiOwarcKuXY2Yd14/Tff4JFX
/A6mdKt9D4+IncDNFkhbPYLHN/2N4srQ6Kf02Dc51xs=
`pragma protect end_protected
