// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:38:10 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
spiVyD6UHe6av5vYtgAykK7HfmgxtB/+HHmQO+/rMuo+TDWdPyUm5dSGHsowJ7fk
u0imkBs9mEOB58NaeaFq/KC5PqYUlW/cwFaxxY4Veppoly40dYgy5Xd2vCn7E3X3
GmNMx+QysAdDNaeck/cWOcvkYGq7nbaW7R7I6pQpUks=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11040)
ksOcrwtmAGaeDOAk2UrpLEIbKF+v/ilK7NzQVYLY+UhBs2xlAtvfBuY09ZThFkY4
N+Ctl3GcKChRjFQo0nBPz5OTBBZgGSllVKOx8i9CbbQiJJ1ENa+mLzZHOXsNE4Rw
NZ13ZzsrJlsFa9kUZwgQXHDgqwbmX8ZbRSQRCUvM3rb88v0sqwYeNl1vIBdZhMsY
2DDKZI0i0uD4Etro86fjn8qN8L3QRw63lHK11qw/A0r6dPPHHm+4yQNUstsYRPEk
qUAFOZgVFKPfSQC7AF5usxbzuHUcCKWgQjl12TtF7/F8qulqcojRBBgNog+0Q1n/
2RQefUVrh8UtKQ16B3Dzbge1EZnbFeOEW79nmeSTbMII9BApuaqP3WY/ukDCyP3o
n+nV2jxEsEB8rqT2zsxOA6jaVpCjQEzdhp9slPltvXp6P5YyjN/OUX1h4pg3evrt
CxEoJ3q4SSLAIp49EGCbmRw44y1tz9qypf/fySzviyO+Ee3LfP7DAlvzFAWo5wTl
WRcm4yZRuW9BnaKNml+j7BFeW0cBu+KTCUPQm1Jg+QKMyY77Jtio/t+vrdFOjbsP
2CnYtNZTPXso8oaJcYo38hBtdMZfyHIpOHR0oAGq+LqpvDDfVWJa3Oo5va8YmSlr
VpJOCPqt9/yoorje/ZXFbOXFPC6rVKBgsAyNdQUVQc+TLZcnlRsHf/KYk3PPuB4q
zvw5Bj1IZkV50P/kaZHpkgu/pEVjU2oZPv/fW+6n+wKKz2OspV1/uL2qDL6V7iD6
GbFm7bpki/ollAtwgsdLSeBfWPUb6uCLyukDjZnco7D1PIElUu6C+EIRNz2NYzJK
11QJ4kmlm8b2bypLU8p6pkxApThrsllgdPT8XzxhLhR4i2eYh0Y3yonnoTFuFbpt
3qMHY3rdUX7XeBQL8KBcdp15tNIZaiQdIU4qhiY9O89VlP5pv0okKIur3znD/CMh
vpt5qTHgHVeTOSh4af7evB49PdXPXjYpBVXjPI5IxgY/gIPa2C0PB9Ld4BtzsN6d
1U8dt8OyLZO9nmMeBj9TD/mZT+4/O2hdHBeDFaOZQvk0bJu0zxOFWoE74GllJcDH
0RbVVcGfDt/fSQbx/c0n2ehsuyOlwiroJmTN3JMQEOeFgVNBSLC6C/f7g2EDkSie
F1zwS79SPqZMB4fCg5NEmTGnUS5VM6a8KrdcRlRXiRSTHcGvRhZLPUZoKYQh5lGC
isnK9MffhaeldE60lcfDAR0iAF6JHsEtJjHmrGyaDoSj54nZ2um9pqntGBxENofd
YTT/uLc+81D6Q5HI/KeX6HiiV5Kqs7rvLW5eUxqgbBhAR1XUX/+an0/Pf0+hlT0c
5vvTv12qeXGUcRjgdL7PdcfU2s4ik4NI5qYkmhwz7IHN7mhCDffODmjJjCcOYmZ9
+tQqj4okTndL5FgGrQLHzrhykq/ehXRWDbZs4IFytjMIX9xzwwP7iDL6URnq0Qij
ZSZBBtOsCdat374ddKL2lw8Le0SPB58Y2tdusDn7uctkEFVDH2bAGKaTqUInCA2V
K81CNJ/sUS+6wiQ3YFu4tPxT/tf1UbDvXnVnAYuEdxpisMH5Ip6Edw+90TkDdRaa
UvoK6XS32brH6yaLDinMFJXN6MhMvr+RAe6Z8bIuR7NkYhfnC+tgxZswvwgchp8z
IS5dWDapFlnJsHDCvbTP3HtO/0kToz/D3r5bIw2pfSNlgLt44yv6ogv/2M/E2BCu
19S6dLyUhjjgXrBhLr0EWhDDGTZBjyr2U1wbiqDgnxn/WeLrEG0jWRr3ch1erCCV
1FpwBeVfhP+qtBk0DDYSh1Q6nVF3xEb44+v5d23pD1JRrHa7G1lKGyLyTKNjetTo
AO8M1019itblm5E8ap/40dxX8Lngjnwz+yG/wvrxOtn935NkEKGA4nCfn+1kxZLY
IWgOFtTKSAlBhmHIjT3D32uihJSX67q/xrRhbuaHeZOKk23AaU7Mu9Ky348qj0Jf
7TMLmvh8UdFcwC0CzB7MHRe0DhjQrb0bCbFcTpIwYv+I7sVB+B5m7PAWo+n77VK6
eDU10weR+OUL64aWurWXw95EOiMW4HHkNGMjBU6VPWGkXxexvD3wv+j95cJ4L2jr
JRErvqpZIj6G0MgRNP3ye9n1VG+IOphct3eAd9jtqjuxdaYgO6f2ByeFywW5QF/X
z0LbjIGP1wNC9IzLwy35w0B/HcHZmDALuOZJoiB+meU1ZfNAMSfLi1AIxs9fPFJS
q8MqhMSXLRB0OlnYRFjPmwFabVyya8a48WEEVcyH2nqfebSusxg+tDB1q5epXUGp
fenl7SdsAghH3iYcONYtVMc+3czM6EJcD6mALMG3nIgKmTlIhfnGGfCS6/6qAUcl
Ig03WKE7DW1nQJLwDVYbyJs4trgk3rdgPLSeZjUxvJQBIROv14A810wJ0ZhPFVmn
xIeRXh++fo3Y2E/AhFdseJg6yM1n+i+VGFN4Y0LhY/bEJzH0HrBHcUVwafSf8old
4no26t+Q7PX+TURUlTJr/7QPRZo0FJ8AoZgEQ+Cfxql6O0UVa7FvTWz7Ad4sjV7r
6IPmxKzwLIBVfmrOVnbEjaj82bwCtigD0jqd8goc4keZDQtdh9Y6vVS4/o0fEjsh
TrrxtR286X5JVw4B1JriowG5x9t5oCljjokQfFA6L4usAki4XAIa3+Uex26C1GF1
n8bqJNWK0Aj0AcSaqpRs2h8B4/4J9G3FTyWrXmcfFgK/n9bch5iwf1JPDnZfwyys
HEwfRZ4d4xLwW7d1CjXoALEzhHrFI4lA2ZMl51K4p7i1SksJPj1xbPaAR9UX/RSO
qip4RZ6VWwSXdTYP8yk695mufbjmcw6G8LCskotKAQV/uNelJE0jxJ/4su6uxM7R
pWn0blBu8lr/6jxpuicUqcN7GV16kfl+bM3T7ae4sJqh4by9Jlk6OEyl4dCZaOoK
r03TxjjDXjP+iWxgBm9hC1Up3zQ9pZtpV2O6ptBluf9r+hurYc4NhVNANc6IwSI1
gnuBwG78pFwGOIvw/fZ56+2gV3Bkz3PJ8s7LbcBDN9hDaHujL+/lUFB8kVIOREfq
PmqHSKitszASDq825PpRs8kZ0eO/3AYJUEu/Cz4E/HZST6sbe6mV+xWX1pcFB/yj
FsJEPRSGViYk5SsY9+0aCs7gH/DcV2kRRz5IHolvcJlbtby/+oTPe+xlSVPJDF6y
j4czvRKeXjSTBJFnjQVHC9yTIdWI9lPOtp9bQGyxdMXtxqy97vdkKshxsYdkt83a
XWrNbM2VfQpf90KcgSm5EeXFMRWdpu/SJzACUDD/v4tW62HX/ik3dOy+DSGo721W
5ruRq6eaH5hWK2lL4LqvIPFLtsz19BMyhXv2w8syt/CffG2Us4WdV8y+EfQR60/u
Vh3Du7MxqX92A42j3zn0aOE+Tzk8eXy4yGoVBCGp+uQd01VHiqI4kjPJQkuhPdKe
pRnN9+EqYXbnz6I9mxUxjNA/HyiIUCE8kyIQBe+iqoaUApwpEBGkzm7oCaXWgiUn
+DD9Mco1SjmAQRMhlnIGuuI7quJHETg0pMzrbfN+o4JvLM+W/7mmXsqjlq7OIHU9
cbgrocjYb5apmPDus3LdZOsrvU35n2Ciom1Clom7XC98S0Kld3tKAclPQUML2ATX
CJs3A1fsfOtlTczmXDeDiKn4vXAY0/E6b8zUXmlH5UpxPjGb4lvuivVetKIAhsmZ
b4IuQQiN8VvaaM3T4DLxxiIb0vk9sAWDn67/TnTSrICn5ko4j07/GHYYOtic4DYX
WmtqZnKikxYonq4iKHH2eYmcVytDaUsYYiC8NC6hG91yNxsy67Dderxp7pb/HqB9
KZBBSKYXmEoQwefy3QH38tmVezPZMmxDB1jO7pJXfwneVsKmSBWUVp+971X77gY8
MDHla/ZWm4cq3NxRQXRWxS24iqSU0q3+CCMrmul+AJyUGCidbJ8TrbMlcRts85lJ
kCk/2gYrwGuCsPxwTGKLNc3I4o3xYItEhoEvnDLiEmzwB8FqmZSfQPIpzPSTjxFl
Go/VU8XMc1FvjfGnTjmp8Zg/YkvIY+m9Ss7Avi8DifxiUD9WtaWK0kXXeak/9ViO
JOs2+li7iTF2qRsxA4AyzuLjvH6QLLR2yte2/PpPwolXJZqX4k6WllPLJXJK/AUb
BDahJcTzisJapnO5DG21pMZaur/qNhmMJ2T5apGUqG8DaD+hluAEBbVLp1Kbv/R/
Mg/4MFFOP7olzyu5faWz5zlpDJZK7RvNTuqVhGkDXuXlvynLWUq3QKh3+cruxNqp
q1bKBXiQ95qFbA3COLUqHlW3R5vQ2D83BgmeLrIPZb8PNx39PIn0xQuQTTDpPhmw
0Ed9voF8D0FgRhi4yHzSAJ5ZwdGIXZMJwWeurBeHxtejbZwvsPVkvQJqs8asBzeo
xCPMAfCwPj7Uot6vvxdhTRPCOni9/fsj09TOFp9oDNBSPJXDtyfhH/j/eFvSTcPD
49a9s0zzs+vqRIc08nA5OK+18Nf0Sz4McYaoKrgTxu5qjtMhLI0p5txPaSVrIk2h
s5q0EwRQkYAaH3ZByieZE7HDTmLptzK/XnCp8xhKBkKIP7tfXm640LQByXYnYkdO
wTvujywLLd7lMvFs/ZEJJqQbk/hCADhI32XNxzL6ir87TY6KjUhoguU6DfWa/hDW
x0M7k/esuFRO27TZm4MAqN/1jz9cvPD/3YDZDy6JVR7ASVAMdo+ROaI3QGNKaS4Z
M57xNHPqFcU0vbo8c2IQmZrSLlh86Vyo23JsD8pPQq9rDlNEoRijTrRZ3iEg+ipZ
aqo5hbjCZPOCOYAUn9hXpp/nCR+EkQhvNVCau8r9/B6NLggjplCUqaiBlrs/pawg
Clhzc1ATxMliWWyFn/a8NPlFh4d9sy7R+lrStRwKbiD1BUlvMs7MxUdQ3W8uS2lY
P9FaQrD4ENegWCjT0H0YN0tp3D9NNqa7Y9A8ywzQ1JNriui5YNGV7tQZMrY0S3Br
QdaCbMbZmax2QGbU3S+RMi1vg0SG8wPJglTaILpXgsE6sRpWfvF3CbroKGuUAZK9
nLuL4Lb+4UoKRz6aCtz01FbMucyjVOP0rIbxqErhxt0YBMgBMkH+dPQXxaM7J0pF
Dm9PM4q6Cyfogzlu5g2eP4msAb00bPnbuPD7G3hy6dpLxTrUL6AyX89lURYhrGBi
LbVE2i8Zx4iimdivw/YEejJkODTRC4VXLYGi9531/92Jf5ZqnrQYcaA0GCXgzLro
DHWOrETySAQNNnwjIvt/LL3k8H+WusREaTFk/xIWE0MWFnDoCJjPOu9nBsSWDGJu
ocQWgnVGo1DRl3XJLolYpJDasYsm40LeAjAQREnnt2rXlIxxAoXbF6gV2e26Q3Fy
Qhw0EaVDNb5nuIdYnVpWRUWg5N0jEU6zZiCQZuk7pyAAELYRITPUT207Ks5X2AJ/
njosue/YbSKYkr98Hf5RXGIAOTyFgFwd9jqvjtBhQWuD+wSxFtqKVdwPz8zh8Dj+
jVxw9ON4xPFtMLe+CqGmJJaK0grpbSUesP7bpDGFTu8R0ipT+HPpZmghegtXW20q
tCPJflDjTK10N+FsYzmzvKo3p2KWheScqd8wDR+pa1mVZJlQDRguWTqg3ntlTy5o
679kWZl0bT1mAgtlxffXRkssBpEZLVSUqoU1dy/EIEUjpD7wTwsvH2or4gEWKIMk
L1X4fkOCEItuLkMb2Ywbv985p2tkXGLX8WIsxa1wVDH1qNrzXzsrVuVugNFTazFw
zF/CBBPJOEBh5dA13bzAeAWO/YtH59T1bL/vqL4HJnjOl/Wa7O/xxwLb4PcCBIx9
X3gs4K0oZXx6yR+ZMcrCoASGo9u/+cSKQCiNQy1B0ElG5wzSX5FXYn2XjI68AgAf
1jktXJQtxUwc9dHWF69Sjrsbd6kzsJYuCMOlQ1MFZ/k3Ue93ogy62Hcb8EXAWcop
1NrVv7PtRniZcLsJkoqzJK64J57SrVJImJECGURBi2ZnBwcBkqrkAzXVnK3qYj1l
V+XOfdj1mqPQ3pHZW+Il2/3tIzN89PqCexh8ujg45q1Fh3jGDOgb9ausZKlzSuFO
ua5C19/7g8rZCAlI4xMcyTTdtRcxdCg2PHsI+Wlc9L0N6tl2+uBTDEKyVlSiWejK
t7eu+6L3amr1iKVuVW1yTRu0VbQijrcBUnscAEccEuI/GtzIFnuxMKJxYvyKRRaa
/MGNKLlzDkKBnZ92OiXXqJ3IYbFN3wPiB/AyYhffLABrEziAkptVt9+LXdEsb3mN
gSEVPGcWOiQaARfErZ3ZDj5FtZ6ideyTI6ofq28kVyYqLYJgDN9eCsgbW+/cO916
mZdp4rPAC7EDKBJhlhK3/9uCKXYlAJdFpKXo6un8RnU9JLcgL9bfcAZX+OFrj/3A
SFgBSRBUL3tzmguPPSYFvdo86vd0Xe+foD3JxaKvLUvAIpvFvhzL2uOJo2glzD6E
vYKWRrgR/SboGxMsIi4PbnS6DiuE7xNX6wVP60nN6W6dFTF15W+r1+jvUseYFGCv
TP4Xc2h+GN3pk2QsSS2mogsvAGI06B2tfhqBDEnCT8hJuR3CwAqA7HaL6gt+oAIU
JleieLesjG801PnaADlkuLAbtJc5ZgXQ+I+XJkn0jn/NTi3Y665SiLp6M470X3TF
GGuLoqjf50CbPZnBxRJsz1udqCobM8TXXcr7W9rl3Rl7y5QQuGi9PlCyYVyDmgAm
0UCmT4/WYwxYn/XiAZx6hsby2t0LwpzNSrTVMpufswYdcD28m8zeWcJ7mrJQj7x+
8NxG1nkEllv7e96yTPoplGAaf9Q1bfnOu6NKtoXIcif+6zXD7/WchnGeFtp/1eVI
pVqZE5A1sMvNa/PS/vw6yE5jVmyqny5snq+cGO8fiDKAKw/s2wDdKIIRxjb/103e
rj0n/YQId1DLtEa8CqLVl3lQpK7WsTA1DZnQrGEjAraHr/vBN8zCjevIGrq8STqo
c+T6XXYothP0GWErGuO1hZweD7kVjkqCVeYrJqhD3kjJ978BQACp0xDYgG04GbN2
5mW9kqh0E2hj9lABiL4Kv8blquXEmUQVWkVqkneH0H8j1UL6J6Y/SHtrl/Pv+SPy
kie1qCQCMUppcFoS0PnhWWMRB99EQhkI3zzsJ1aAftpfWYhqE4UI8Yjrs4JKlxxY
Gb4ihVe+b0B984HZhAPqB4uIqdnpIKHLEX6eXhm3zfxJORTrX/vLk+gZV8dlSzfV
hkhkdnm2oVQ6g9v1EC2KMLTFnyf9qnpUmHKdhKjoyLarzFnCXwyNIQEFIv7JZse6
oix8ccZbqeiyZWJQL4YNuIif91XWriSJSNtjOdih0UsECjPVkFfUu6tj6GLmUS7V
4/QaPIobnZXrfT+KeEdn5CxxkIBGxvW+S/I3L/e8unVI6L+Kkny1n2s3mzwAFN+S
1KXSDZvQiSamA1z0zqyvzyi0T9E8lmXnvUN7LSjwkONAidXbt24JsBnfkdju4/x6
oUU0Y/uofJc1h3B2YgxIa68xaWpuwSE2R0yFDX6KyPgGVZ9BuIE78KvqCRK4P3vF
x2ofIYDp6k5gaKaMM9XhvirI+euiTJ8Xq/+YDgNbqF5zODvIIk/h7gWX7ThSoVFU
f1k2TziGoIeKuMRLpF3taR3UNJowUbc49qx2Kil+NK7iS+x0rAJKvN7tnQ2ovPAo
ezq4BDFpvvhW5LS65b8aBXd9QgzCaY4OWcWm7DZYzD1y1uLyb8aaQNwfCIvHdU9y
vpy7s2oRIXDuFlI/T25EOH92rywBY059TEzJYP/pw/wOcb6jnscsqNvWmN4hpXFX
jUW4FvJdWnxbvr+N5q2YvJ9olZfWownZnsslQxM/z/0lBq/stBgSlISkFL+kQyAy
wB4pe9IP5sI/U2hLr8Age3ka+c/qoAhUsDuZ+CH2aUDE8Ruf8vEgSbmgKvzQ8xZu
nFt82IqI8HMhf2h5OqbXVpRBoTDRfvMKQoLUyhVYHvw0FZgDDU0KkNSai817hKsy
DJgiyS7qQbSGcuhLfVhvsezFOD041W/xBfBsKyWxVOQ+MJT1eKmJPhFVQHm70GdU
geunEWfKEuLTJ+ODK9uyMvWUKSzBFb8ZrmMinYftbE7wvBKCJ3uwffxYJ0jcbC3n
Echk0AoKcsU4cxq5GEF0D/tVcGBSoSqAi2UB51FxNYCAGwWq+bHSOet/6UuJFPkn
lGPxrPM11nvnkaSM6kkWpfO/ypR3X6KRV9oVEPLWztVYfP7YIEvBTIPuOp11CkaD
gc22hEWjxSgo8kVZS9RwIEqj+5l549Tr3/jr+j/pWMo3jiCrfq/DqFy7+ND3ciMQ
01QvGln4pc3rSFxKgkrBQ2T773R9sZaHXhJZhVHmBc5ptvh+TsDyJpQDakUDuf0T
bA/qS3RqxICjQAh+TXk39imqU2+ssgmhbFbdIGh7iTciztdWOuedQvIptmdilLTa
tNWAgu9JVkJWgv+ONPJcUmL9qgLIWUURFcE1IXdy6iKo8uVHMCRlygbtYX/UOXGk
uP8QCSjTEwyWGcicj8XJgnvmEVXRxlGJTLzFkWAYEH5zyvoFIZlZm6ZbZ20aO4D7
EAlC4x27ACt5Ea+ljeox4Daq3uf2sRBNtnRhWFkONYu8gkijWi/lM7nut/fGF6hg
uPG98kYZSqWLiOW3ccsHrkx4M3wperEb/LaPSFvuP6htcg/P5FyXSi/tzXQRdU9e
lZWPN/CyxO1v5xSuTIFAdyhXp50zuentSUg68lOwRwZ6qlzwfoZHsAwEETiVm/OK
9i/b9J7ToBSQT1jcBdlANl7VbFBAvnUCLdHLiKcKjEsBrvTyYBTrbMmrQUuSMKS1
U6e3eso8oJ+yQwUqVIgp5VD0V+GuCvXMvvRoAVVeL15Qp8F5snLWtrf6xbKm2P+w
3g8bZIGBBywC56YAl859vGWDVPmcYz+68SfIrwBlAGe1BafvrBZatIwEycaOj7Ia
X2WtjftdfBsmfDpPz0TLN687nlLna6ObXUONlt9TeFF5Ww4MTu/sB9gMcuWleWMB
oTKN1e/IXvdrqRWY5bpz552PifioPeascUx/Fo2VPIm476MypCL8CrKtlyau5+71
to0Wh69tWrYsoLQCKKOx5rghGwb0MxPz7K6HUh0jX2Jh+GTCzfXUpjrWDdJeS3e4
0goMpSSEzXjl61Odgek6W2tCqP2bD6KOYHVqP0mxJ9DBzUNEQ48qXf2OvqR3E1tO
hf6GxUnGferBhYPA1WRNGXgl3n0HlxPenceNe5Mnb7KgWvmQtymMwblpPMELG00/
1zqsLATWwv2HaSxHFiidaueQtUziPaU+aYlVkaKBplCklSfsFxBij6z350iGdoTk
7YFqF1CI4h3otBYnt9xMEUam1tlB0XEIYK4fbrhLixahFHBQmf3d/soQWQvzRw3U
XOS9MMh/k2Xw28sFaouuGW0IiGhl3uXO6l5/jIsPos4za93UF1sQW+XNOMiopxsV
m67qt4/5OY1ZLaYlafELSNzuy1ZIsJmOqfMv7+O8trtIZmPCO0PUuYaWFe5StWMD
DSsNmF6jQbu3T+TneDKuf1ak5YVjtszeX1Gf6lOemVYEu9bza/aODabQXfDB3Idb
8uqBCtG5B12m/IrLeJAEG2O99Qpy4lLY+gn+Edl+HZAPZDNXwt9r3K0LKV8vy+k7
fwTgUYbp8Z/Svf8FQrAH1RYAE6D7btd+3KUbt7wCL9+x6PYFiODl/zv4ZvDX99E3
DrwQuPJoOi2IOmU0PZXQGESproTrOmDH4S8xQgFFKKecy9WWBPDlAY8fhk3HdzXZ
0SrwZSYtRUzE0kSuoqNakrGqYprvkpf1YQTz2nrImXqgiXWSVqlV3Lg4EQPliEj6
45+XelI1BCSZxG6fTw0AR9A07zzIBMmhfDUvsfjYO5689ZvcKNYY796h5UV4YWnf
lmmrzk+WXdUYRRceyNHoc4hkpPGhzrkXvnTljJk6sMGcvD6KpRenWhx8MVSJujo0
mOt6LobgWXZ8LUdgc/8rAsMHQ7fK0x/im3JIbZ6DJL/qwfmJXEVGI/jpRGIrPRYC
ExQ8GcCQoU0p2/Vzjinz+geLFjkXaODmzpC+mFBum9XEyU8mvr6gZiaJmBLthwvi
rP1UGDKQJ7pzp5zce0yGctWvDqYLyNzlcxmGuJX71coP1J48rzoyd1rK3r9uCKm2
pE6GjhQk/Z4wmD3mLfG7y/NX2mIi1uki8aYsCABBh/B/oU9nUnRQgvKQy69d4r1u
ZfqItz/DdJ/5WCcYN0WV8sk3Z7HA2bOA8eNNzOmONDaE3OA2N18sazeGESWm+GCy
tuitZEQE25pj0nKZVEhSquCwuqtHHa4kxKBiYrUvkuYE4fmDOlMmlh71DXciegvP
kL9wf+M56WIUhANINcf97DDUaeMEdeX+WCco7fytMJYxuRVoqUkuDdI/fujtwcQB
5tE9fDVCs6IeOLW405iJJ8evi1Tw7B6DkSJBxSIt4yAwX6puWokKhDhGyeXMhA3t
+u3HGOWxB0Qq1sCRTmJzepT9xMqsUd45d5NxKHgRcvsf5me8X+H58cTHDuhi/eIJ
C4ZLc2eWKvxjlYshXUjbmzV8x2iMZfQ0HFVWPrseiiEoz1rptgvM/hDRsGry61/o
l+GvFuBOXUahZ+6+7Zj5o8yKuJBSlll5mVwo9JcXtaxHw3+D2uUEDn+WNdwf0C6D
I3rC4TDhYtEvkbTluID2XfDe2RidNPcBkLFjaMGb8mtR4iqKNQx/tbmtDtgNryG3
QJOzmubaHpsgDZdjiDazYjTirmuToCnAvDut/pgZbmyb0vR0O9Yq20kp61AZbGVJ
7Ll1mSQClMppTDr3EE9uH15Rfdep4PVrIJyIgiaLL6rFUqDnjsVRyYO8elhSVRJA
76VLcr8dk6i2firif3xVhIO+EunoAJgFSrBbXJSOrnEo4gCEgMV+Jx3Lc3I9A4WE
W/D0bcB/9HP+/vLl8JIL0m6dAIpYEwkXS2IUhNeAYphJIKOOsAIvRrjG6usnW9Uk
3VjAGFK5qhq/1YXhhVvIeOh6XlcgwieQsNAJgWAhWUNdemUl3OU1+KvY1faR9BYv
rcJPl5wcNwsbTrQn5jGx1+emdDqElf1TuoCv3C+DnK9huHJFHsQDxVQm/NF3An0F
6A2j7A+QAB8EwyFQRl47r9rEOxaR1KcsismrXcPIGggvXkjB9LE+HXDtNLpMZe8Z
5v73XICq/FDL+nyoD+HMv8dLkD5ea5EmUOMJIi9p0sDfk3jjSrrf23pSlAWO3LjZ
x0RxoUwVApaxCLe/03hEuE6Rlqz3Swl7LH7DhbXjbkz3muffqRd10RA3P6Wc7HUx
KvPuxR1iBBQIolK9XbJJz52py+oEpcj4Hp47W2JHpQz1++1Xm2W2I3wr2PI8QtBq
TfOOLWcY0kfmq4hk4hT2HFQ/Q52YtLdyfF5AcUsWV+7My4WyvH81nd/2UGLw3hLl
oE5FrJJ1F9JahVqxygiIWKMLP2A4l9nOzSc2NYxBmZUSMByV5pF51ARX53z416N3
CxZvBT0ZwiqPWmlbWtx73ofiDPHpXfkSAlGp1FoMBMYGJGroVr5a6fgh492MXZR9
IFGTU8mP0rhKMV4HBnl4a4aEaQKR8pTofbxMQFROJ2cQHOUEOKzM8oDN0FW30Aog
t/54q99MG1nbrPnW6lxp6jAzNmskSPvntacoYdL/m7q6O/bssAd7y0AsQ2IjB8qY
Le/t5g3Rfiovhwk9ppqSD96G8QWiLBFdD9ORB+Ynxt2hW7fHA1K7nJlpENUsdTaA
iXDVct367J3b2b/eXCCc4bvpl5n7TBhF81xJBDgfEWYSCHGCOymM7DB49xdO4Od2
9/Vgdhk/vzP+BCOUL8L9VyZv/oAg4VN5lB1EqP8RLSCkZzHJaTJGHSbg5PMuV2Zj
McV+REzHHA6VXywJsmPnMo1yK5otMf245Ocpsxvn7E9NJJDAa/g0n45pGjkLwtxi
5fEV57OIqXaeSq2flm7mfbbtpK3qM4Bq2CZUCj9Ce6XWJBfTAWBamsuGRiieE96O
F8He/QcSGnfmiZIdOy6dISVq3qNfYdfSdehkEgc9LF2hNJygc9wWASGJpq9Us+RE
X0M/OkwjfVWAsjOqAZ8S7hVq36P/lQuxsyRgs2+XKNHnzrDKuqQ6zkf09xhESPEL
LqNZGYusMe0q3ug//N7WynWT6rkaZtbzQb/mXeLjKCe8KvDHJlXmUxeY12mpGxrd
98zL+9HYJF+mGi5mm6RJUR6Tva1vT3H06kRuZixXJYrxOLtEOOAK508OGNzJ3knB
HWWE8T5lBly4YUaoDUkgbvWkOBInCXcoCbsDq8h3OcdH/gZ7in/UhruS1OwINWmV
IQiB34mGehpDoswssuwNsgFQ7iOifrhJEsMjk8VrNtaCrErejU20fOZ0jb/EHc+m
AsyJbPWsk/KXjh8lw0uoWndCVADqtizzfq8C6mQGa3p+n+AJNf3sl9MFRBXP61eg
tFpKIs+92up8nMG8p1gvzFkVnRStvj94d7AOPk09b+IKu6P4mM7cVJ/g1PYZa9cz
yDjNyz21GafzHq11S2JfOl/vouNIhTzbVOhEkDulQDNGIRPHVvWFvfiLDXUCA+i2
nr/WrP3271bzOUvXbEP4Ijf72/mNM4IzyxQ9T0c+l0c0bzIYq3nqi7UcHO3skPM5
1R5zbiQVUD+Ez4kecbhn0SpVrmpDCD6wEgYNIjZMS30pvhGe39GdZXAHVcXmUMBc
tjf9r2cH2k/CmOL28d/jr0VCf1Xv9vqd+SN8SolueJDpL07YXgpvv3bMhyBWPNjR
nQFMlpsCXUKDfjiaL2F9vxmspuZ8/ff7K1koVwCgwJ5btpQTCKm6pGiFV0qUh5XW
1Yih/J35QcREQbWBir1HmKuurd0cu9H5vHJhASSSpEATu5nPmVqaUhc8bTFbbDmk
iA49SgpjK+7+x/GPS7aZr0W3CKcCbxTf69QjaZYL2zUXunbBK5lLs67HxSSNUQ+E
UCSx718fGXuyRhO7PLBhHZTjUVS5YGNkHldINd3i2PGlQxxtgULVgXZ7H+04NVRJ
f0ZGcCN4HFxL0vGQWry0yY3AaM7Axt2Huw+qainYEeyGcgtBtxTiV7hoWacX0bJK
d/vEU5lxCshXV1c+i6bDpv40QLOYSYSDBogOoX6PHG0JgQlT27pt13rZOBkcgvSk
e0gV339Rjh68pJKr1CjZP5n1Y2tWdn7iz598EeNV6WXlQkgOKArBPXlEYiKdYoSP
1wnoJuls/nJMnxJJpIZ007dLmmMLuyGrUxeXpjAajMCVPkuk20uIDm7FI0x2jD1T
8cCyggLWJCqmbKAMx9uDejEQXxqhbc8wKcdOdqVPominySBf617+Wf1HgSIDOYT+
ovoGwK+JyrJxZS44ZXGXItsbXv+YeQyXstgX7VDqVnwM506bh7ldlWOkCtKkLXNL
wW/0sAGs/o3upiEf3fAsgPrs6a49TShkWm7A6dVsqgmMIr4tbKBvvrLfcSIZjBBp
3SqqRRT+5lLUjrpDIJaZ4HWixZvAxHtzrF7xA3f+utbR9Sr6Q08ZuDbgx3K++6fj
fca7OxcQeWEM39IuXXjS1qXG6rFxhnArSrxTw4CrAKHAWWwFImG8bs6R9sYi/PwH
zNecwytepZWlSqao1o98OluHBJ+DZat3c5wbZBca/WxoUHX+j+2rxEhVK7HHpgZC
4sOty7FkPiN0bGTSnbwjjjD+j/X5QEJPRtLIfYUqNHd06NDDLGZdFN6BzKHPhx7f
bl/I2j1Mi46/jYx4bf1timPA4eAnbhy9OTiR9L57dWqUgiJ+b5GXOVnyMefXrGho
OuYAIabFM+7xJgPgkaOcQFUTQdwYsMAMDaCGYTpVxH/FzxHzBFxUgzMgp2TGa2Fm
ei8zhMCP3BBw8ib9Tb8levv3f2Cu2S1MZL1v6PsHQUnw03tJ6LuY1Ta+YwOafOMx
W8cm5BFUdy1qsFoMgz0pYY5C67BYH1RDmiCcyiqwoV9IKdRmc5+g1h/T+2X6WLwo
4WEqRY7s/yzTsQOKPieyRVY0IjhzUV7IN8nNWPvixP2BFDoYaXIgSer5+bddnkxb
NICyk+pGQ/HtAvdg3xoifSY3XdiqAzDQjlCe7RFo5CDtrx0QBgris8LwRWNwuafn
MoZQkeqearEOFb8zwhGtmcCTZmIL6/80QEF7+hrC9/7KOJwkJr4Avyf/XqWmPOVM
kzW3/SBT/BivZmLt9Xl1GoFctRLPUMQ2Kv9Ik3w0xu+uUc/8hi6m3rINj+03Fgun
DxzUcL0DLL2+O7CtkxQ5Bz+qNI9hp5EiFJCBF9nJrzcR+WO8STuLHgnbPOEbBidr
dn8X+Ztllmjon6zBQyNoh/sQBkLum6n78UQf99ZKsGDssCBmvKhPTSKSSuSStd23
U2LMP8Pi97L9y+Iv0by4CtuRsImQJpdo0nvWFVHqbtg39PAKLmDYnaJChodZeVNT
TgBb8SuJm9FZfzpCx9lvZ7tduNk9D5XlYf6WsLL3gJEJsLduUfJwaSmm17iZQwRo
88OUTTd78zUyhcWqf5qqJ4xYwWj+bi/1x21imaxh/UsBw2oEKo2cl0ZcjGMDwXuz
d9LC7Pw3MlA+n7zcckWXSAwGd+VqkV+jgyXVslg2tVeKax6/hi8Yez69vC8OzF+/
riWsCqXZuWDvMi93Ogwwk8+O93wFiqbOR4uAGrUrJ7eG5wRHs6wkORETo1Ulbnb8
`pragma protect end_protected
