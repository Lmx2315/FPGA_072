// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.0std
// ALTERA_TIMESTAMP:Wed Apr 26 13:33:39 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
sxwhDtRMUD9DMrU+HXPMrt3vakF9vnqAS4utgXsGzLSPyNOjrDV0lXpxvMfQSOEJ
3sAM6Akh04Cf3jv0xRH3tUxB6sS8rDNq8ocNExOKHFMzpzUmyAWHTE1O8xIuq1u2
J20Kl/WZ5wyZG+SidmayjKv59CRgtOM4iTl1NieGDCQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 28016)
HUHNskYvxO1mSVG+J9LNzrPTICm4NeLVAh6Ks9HzXqPplnMpkYckqVR1N4SXK1NU
5pq9gVmpcqGPeJOJpoNgeiBzEND0Y/2CFWAA7xQOS0I+95jzlxBaiczlkB/RhbW+
QPTw6xVR/zhV07hr61UXLYYmVQAhCTBgl3RO1BLb0JhpJC1aGxGGXvDYWz/WTMAK
4m4IM8Hr0ENXI6L1h8D9GQjz+1oHcFO2iCzUOG/wYHzhQKqSTZRDP4rgwqF1UWcQ
mZ0myBiynzZofoi/jt/nMyGxYRK+tTY01EqM3w/qVUcVlpI3TdgvhybsI8jTwvYX
YGHpqxpP3ZVb4WiboQzMZbWjRz2+IIvISydi932c4uSShOraowqNwroihrmbnN9Z
4QvRBfaEYikWwVYkp7Rpyj047Pop0Jcc+fNIzFdRy5bOYKzA6n+894++JJWd3UIS
KOVjSCHWn8L3bzDRVnJNYGXufoNOSQ3m+F8CJqI+NxtF62XG9dOtQCnHXzJci6zf
CxG4kG6uzEumYMI5rF/H/inAjRC8bzqbd1lB9gHUTBJJ/6h/HVU9lKfHDsnnJwfE
4PDCUVxqXO2e76t63nCpzr0kKofT82iatpsJQDE71kZXPNespnQQjuQM5BuRrm6I
xatNONwGedmVfdIzKqR57HjU7h3m7CVk185G1Mh605O3lL+1xUrahiGOMPm+881w
1pPSNaOqtNq/9VBkhEVVfN8Wy7FjBZLvqeDAf+6P6Yj2I2xiq39OjlMt4+uL9zqx
LJHuZsCJp1sJ46vqI0egaG2V5kjNX4LFvFry7TcIFdZGcZrI4wPq+ZSPq1V6A6O6
iI+DO6up4+H7TV0hVV23YpYR7ov3GJe53zidC+h2Vw9J6d/7UfbGd4/rdP0PbUHR
V5JmW2m1RZO9NFoOz3aScbIBEMPYRB9H+SZIa9ljD+smua5xIfGQrh1SaCz2xA34
TZYSiSkisBwzj3sE70r98Aa8NJNbekkMaXoj/TPV5twsyAKkM6MbpQKXZzjvzUiV
nKKaoG05RB4CBAub/s9Q1fZMSryy5Qulh741Mq0j8W91IoPm7jF8wfBcZOELlseB
ENnk4IlHLu94bCo6ugsKEe0UjXCUFewcL3t1ykSGkeAn32k5NHEakvQgRlWnBhF1
VSGbuSTDk7g2fgyPyTUEdF69VQDvOZiDwO0uaq20FpfKZ/0d7+byUiyr1xOdNMBE
mhBM1DDlZ1sfWxUkCdDethjhNsgCdL2E9PTHc2fIp/qEUPKvCVV6KbI2atgH1d4X
2/IAQplRgj5Y7vJsV1evqISxxDQ3WJ+j91bVnLhw6XYJ2GjU++6nLxZNPUkSA9pl
3ZZfUJcCs96SSVtMuTGde2xi1taGik0LaXMV3qkmj6yaFLjHfcHXc/KqfcA2IxBm
6kHgRbDBYiaSz1Ruiz50y3gmUBzJS64w1lm5W55CuV9Vxc0MCQHshjs+qvg9e/Bg
TsAQh8V95FX/vUtrukvgQJqxKzCNcS/bm7MPXkmoaioUFckJC6BYMFdxyaRwvX/A
0WTz7N8Dqi/RqeuiIDDg8VfnMwG+7qnCQHhY4j9m9vdcw8QsIcWVPXZA3UklsFnU
syIqUDLd+JdzWdYJYqDDWnjzb1/mIlZLJZbVv8BKxGmYxsL0yb6oJvvNATmbqJIZ
5mWanJ/nyUMfw+FUJv51g3ISZFkRy+egQZkHM/NBt5QkswD3/HF0dhj7MG/CSjVv
tTQYdYCQobuvz8fQXfQDMYrNjvQbEpFEzeXMwAnR7UwkbVn79SH7stOKMu+eYHHT
b/lFVjgUGqeqNFsXrhKMjcgMkG2LQQTgh4vfqJ7b9sK4F7ISbbys4pzm71YvNq5E
JKRjxKGYgRxAVBoHnfdAXguZBauvN8KWLF8KCv9dHwWZZGllBQOgW1Galz9HPiF1
ELjbSmP9fq3vVe8I3Y8NHaiK9VANj9sWi0lW2dFt8GjtAIdbQJUBsfJju5OEHKte
bsy9kwwyOuXAF2cTL350Yxe1TI4WADRD/G1Jsb27uYf51wm0eLfPOA5ETxByOuKU
er3Ku6YIXsTXN9OPwn2mQhYzREatYWJu6Yl0HI6neXXQdmSXef1BA2WhRxYbVKNy
azfZ/tMfE8gJOWIqqTc8PZF47BX9SZcRTvBMkkiG83QSBaGUeZAWsw9Y0CSO1s4Z
FljsFxkc1FDiij5RR1AE3hFptsfq4DQ0LDbIwnTNKw2Jhl5QdwYzGkilHZ4E6ylY
qPVelZFOtT/PstIyA4QvJvfFcZ1o2SEPgHVKr6Havga5IadFzRW5zI7PqaILnhQd
yjIr53Ot0kzH9iGexernU5kyLoXhT1kOK6yhbK/zhjr2ILq6smQkRLrQkvcj1YpP
yDfFaX2B+b6MSgh0F8DUKXiV3fWxSHBhDCnzeXL1QCQ9E6HwKziukjd6tdU64RUS
xlPtYyau+s4NGi2bpP6PDT/qVYJEznutel16YFWdkPOntg0pQL+GzNHHAw3TvlGy
dsawjoZcYcoyCsa2YmzTEBnx9lXPEsLZw4eilqXOwhb5eu2yxeTiGhH7q+/xKlMK
rKoOX/LLoM7oytYDFfu+9vdLa28VLS0DJl8J5uUlQKTs5VxE0GEo5AKT4KbVRKdo
oTUeum/Jn5cmJv3j1Amg+u9qYqppEtEJdZMPhHqp7aupMth86F9KBU+y5COnORwB
CARrXb5RoMr1AFX4iq0OA6TjHndZv5F9u76irDO8KTwnOqTx73wWtlkhI+M7gHeJ
bfHn2v4l9R4b+mZUo3vw/WE2naVR25W7H1yKTq5Y+g3pxMYemkauEB9fcxp6faa0
Opv4+ABB9BDdVQzEIFkUe9dqUdCXb11VJxxZTq0VxD8noddEjfaaiHOPgnfyly8p
amT1ySUc42IxLLL8MH7es+gsDoGv+QPEb+bYDzMXqUjXMCpU/Ku9t0K4eh6UQNV3
DgOr/mEb7ktnKqNcN2qcJcOoWRMa/a0RlCFwCu7QxsKzZ9MMkTMz79KCCbyXPJyS
a7ni2kW0/6KZoeyidVh6e+4RI9DXyn8OVMpMd2V4MJ1dmOOt+Kzlayq/8S++A60E
xdGg+Cm8mFeQHDdYz97dmL0varqhgZl/pjt8TE0LUWAdLkcjvdj32sCYX0vx5yZ4
jbH0/0pC1uoG86c+NJ5KH1EH9yEKvdi0pnrP+utwFAT9dv4u9592gdhQwVBYLDiU
5n/YnCBasc4Z8DGfRJ1+7dgloOQDlUGIibm7hmbwdYlJEnqkDu47iEUZHT5TabNN
9tY4ei5cn9NzBDb9tbg4ANj8v5prfwXM9LH7qYDKYRRGXS9mfx//JeVKrgATAJVu
yOa1+c1MkFzEzB0h879BobU1U92S6ojoKCpHh03PYTjjb5HRilq+v1/fovJGIs1k
Qm1zKQ18fMMc+v3y8NNQ0D8/2k+FycLAIGGhcbygN0qOEujTkanYGt/cKcAoBm5M
e6ztxc9g7apBVk7tiMix8VUdXM7kQQRWPoqb7miT4HIE5pMPITHPhe9hJv7E7sOP
KT8RI5FrrNrwKSkDzvldSfn1GOeUvNazmYxDEY6Bzs7krhJOComQcpDPLCmZv22P
xy/JYwq46o3vpKC7Ukv3oRXz6iwd/KB480QERd9MImvOW0ZcVb6QRNvbxPgRankP
/v65e4f27EBjMWwRIiISlO1fZuVFklqOAqPMBd/lQh9yb8AX3BKjfQLFnckirrhc
xbPgT1wTBJMJ9jj2W8V7QN8E5tZ/O8Mi5zRj4Jg5PhtgIa4jMV0j8wwLGvngYWHT
KaFaGSjjdcOzxblIYN6Z4ZpFbWYxqx2tHjd2vg1Ps8LAgrR23INQFtBwHjEqOebT
MyKct9EZRiiCvVSJ+bIgzAmkR5QzYVqV4ZTrnwdZqkNGLXZuTimmn2YP+7UflEYq
WgmuXy64uTdoYqR2NEOXiDALrEOexg2I7fezn2kfG7PH2ojD2uGrgBr1Y2BU6AWg
/wxDX5dOKnMdjFRlv4c5jF4KCsFaGw5GLKLzVVJOh8+UEewrbQYnIDwF3YBaCYvH
cpcReGoG27WFzFe+l9aZzppDvigwtoInR6ewTbLOOjZVirxHKUVXNYbv5hQHCQOp
w1eACaG1eiPlPoFtcGiHiYbwMv4LnpNBBG+h8mYO7EbFQVxW3E0r2ROwdJvohrds
G0X5I/z9TN+pfEIPloJM2CLz6SORXHAgqcFivDUm4EW2Z7DvsUTM+jfAEsgePTNc
et2hjWlxvgzIqT5xIEUT3G3HQeVnjJmh9UtQ0uva3icGudhCY5idqW8MGEOcl5no
6np4Akd4/+rqIwFFfzPKBCedc9l63qdmTGoP08TSbVQVnhjtZay5o2u10+l8NPeD
fKoj2nOQBUC/bxwXyu5iEliMqHDvt5M+d0zzvCXuY6jdi4MDbsXp7IEBomezjzr/
2t8A9g9nAakJQl2IjRPDMj5RuCcQwz8zCUiAJ6082FisqsTVgE/9Xlnv6tKejVPb
UdfDnDoCk0rxEEj43ZNNbMFiubtc0mWWLE43zb8mBB9Zdgx3XO/7gjhSvFNYyqk/
Ji0T9YZl0n3sLeNi4vRiTt/QEGpMs81DO7eM6waGNXNPUIPQgFuJUl+6zgrVukMZ
kAaDmvaMlwV0++HWrnvVEBsN+GOzYtxSJ44tSvxURjbwtj0bcmYCxh7Igqn9b+dV
ixBW5HYsTaqj4Sw/itkjRo6Yhr8QYi29JnzrAvvqfxzuiYF/3xjc8munARa6RQj2
JKdCnLuTw8nABBx1Bqmv+Atg/kbZszW7Xa2bxG9mAKjN+Ec9ukOBTy8Eird83jwB
3Q7yWuqcfun1y8ek9OdWtabxG9gOOgxjSurH2NESza55Zwha/NdG0gMmBtEN633o
+BSu0Tdg7lmpXYEQfw/Vkjdju9MvgFC+9eNRIg6tlmd9sWX5VK1eSqZ7KGTpD5ua
k/DFJz+EqeaiKJ1IbWsE2LUsyiKvRqYdRmAQr6aMCrB8Vu1+k+K4j/cF+g86DJAy
2lna+RsDewEZD60m5U6/eG4B/yXUuw6VuWrbwJGBuS3qNe56ZBlRe4l5nlUgBwfs
swtBT96Ni3Erhv7Jjnv5LHImOBSefmOaLnfwu+Hxgz8F4GAe7XVD+agGxwsl8mnN
6fqZQPPr4j4b2fT86mrWg5DWecxR/Jio70nc+g8T4nTpyVzSWVzNZcDVUO8tZTJH
Xk63bsZTzmOLd6mPhEXRZZsixNLiBTTjo32ftrLpe/oOa5r9ZThM9fTI2hcDuFBc
m/c7D/5BdAJBYIcpIJiyp478kPa41iwjpv74SSyeMl0ACU8UlMIaI0HhBV68UV4J
K+rG665RoSxsa1BfrH18B4chgpgb+7xdMwI2IDrnj+Jx/QsjERpbfzUwLlVUlGtf
a7Ww29FPjQj4V6oJHrFXhHtM4MHOjHmg8jpw8dBP7TVhM/nghb2oBwW8lWa4B/jX
f56fdfzJoahwj03q3G8NS5Vl1Poz5AgSQKQGXyLkvUxGOXl01HJ206Nni5/UDCPj
dAxJvWOD1gtOpNRPfWL9POiHRb9zfTWZgcIHaM4gRBlawwWpHxZXyej+RBGeajB7
F+rjNJprUnqgNkwZOt4SqEub08n51c7vMA8SmZ4030DOMssnj7ENlAl98rYY9vGz
HrKvh6zqKYSUQxGc4657dXq21zOhp0oj0MKtkexOwL86+Bh+2FpWOFyewc7zr0mj
f+YtQyHUAcNLlff8B9afTkH5UhkkLRKyNkDxJLVSVOlTlKHqbYlIDSMR4qXsjFUu
hFH2O60YmTC85O1FdsKRUHt6tja9m25vbHV5VtccDQNzwbpFXUWi4lEZYdidT9ku
ZGdu5ePTnD/GPJL/8UOhoPg70pGgxbpKapiN+6jiRrZKo2hlAxD2e/ugGue8oDP6
NkIdAXGNma9Puz9hITVs53pdQenQeKSof/HIr2bQo/fL9wz3+ZmKbLfmkS/hUBEE
oofr3xyUHeQdcUc/Q4USVSMgOQqWcIifJUdpAQrCNTTsWUTezrMUnACM8krPCQIW
meSfDXP+/Qr6NHwiIQx32kKW+/kIXyBlSYM+UVMQeAGJP3d22XvjVvHlVOtlktTJ
UR7iMJipFmQAZ/tjxsW/CKrcUf6h9mAnm7yJtpV+OQPkhVpRT5swiPjfsViCEBg/
dBS75o/mMMLoVhEJIDGWlEq6quT2z6y+M1Xy4GiCDcsa9HpsOkNykIuyOvBByNW5
guSeRwVKtsnXLf4pM8tluxdH7j3BeBAk97NSJjO/CjV6FWRiy+rhSQGEr2r6oo8G
4aLVOkRCakPsOnn1uaQVqsUMKCxmFG54rcCmzWJBtu3Ml5+aTIaqnXW3oRy55BDg
NcN4PZt6ppVUGnr0VPCcM1hV0YlPY69ueX6g2qu3IBAUCPL9iXl+GtrgSR4t6EiJ
oNdRBxWNrJwkrXaNYVJzu8CvB+YBYLknwsD1OVE/wzm8v4X5X0bfBpOP/ezxPaD5
SM041SJIDHHZfWTK62vyAnH3lcRuxwAUV+OuclSljDirf7I0r7NEAsaZpx5xc8f1
J1ORuYmztEVNoRXtybp07XU896WSbKn/D0cPsOYrbObhKp/bjbI4Ziyf4IX68xyy
cft/V/73S2jpCr67lNaM+4/1KA2gFTiQkWiudZ3L7SwsT69XyQ7whdw1NNAjJhdP
WkoqhvcY0NxJm2rL4BfE36c6uXrgKLJAnISOzthD9BZLkxfIqbDMvhUgOBM4YlOs
115cK2zC++1t0Xkmf5mDo3gTe47dG/t3udG732x1eU2AfkVr9T+JPAj5y4iIVrWC
L73y4v2Fma26LZB6LKeTtEMGM6z8RHcCMSRSpfwSCUrhjuu+HmkadFotrGWKNMXb
mQ6efzK9alP8lPTAxk1A2g+oX+UeYXwzpyUvF4q1EhNmCZMjWv72H9J3HAWWe+Vh
G5zEma1JLx1xUoJtUbofm7IK9DaBcOFj4cLfEXPkj7JTdr7VvetIfr6L1HnU5GkV
NukamCUNr47X9Mg0bU4CMkO2iWJZAi9QDQG4AusIfQ8ThMs59dFRmYpQ2F/8fsmj
z0u5mxNUsQxBNfVYC/aTn5d6RjCG4PsC6NEQCbmNIKtsqEf7tWtYJXHFLzDkuuFR
Bn+207q3NUpz38ttM4YQxkAKau6ZDIf0u7eBgGeLhMioGpixd28iHXcJvG2n0XLc
b06dB7vbxxeUG15oQ9EmWb24aL6sLggiZ+tcFjr/Ilir+U1rFddqso/PW2ehfz4g
a7ks+/IHqGn3TbUapwB9TQD6GqhB2OTOw45zbR9BmalE/NPfC9WMTM9oMqPjXF9w
0xYaqCNYFHjbZ6t/q5LfCTcI6F4L+iz/hV+DJViPoaX/zmrZQ4GSq7hB08nlfAjK
H+VBKhC/THk6KqlDf1rPyYTYPAgw9nPZwFc5c2vNsn2WlKP6NQZ6qLq+FEtP5BPK
rUour4hqo5AouXhzFiuDYEBN3x54DDHr8uJ77TnUwFxgByznPdWuG/cOncbf/dVM
hrTqKdnAKIkzCFoPahNOx3bxLn0JmyBEZgFf/3rYvk8BjrVBmjMSzM1A5TWD39BW
8y3QfRXVjLPsOuzJyjPbh6OQTodQVV3GQXgvrQY4B12Kh7ICD54/Y7VZgNCaVOKC
R5EdrILEaUF6EQ4RsAebEUXL3JfnLYwU8vGEt55yMfl5q6nDT7caCGVihnJJixvZ
JnUJnO3W/jfJQVbTLJyz0cwc2vGCruqZGZNDOOmFJtsaoVrm04TmdOQFL5Xj/qjp
Ak0zSk796pjEPBOx3IBQAXfsSnVanT2xmZadQXPw/CSclNX0+AO001WihbwRLp8J
FAq4SekjOy3ql8xyV56aLmhIkHVB1Ki6iz0mjrux+ue5hOAA5PSSu2H+jdEUewfo
u2lwV2vK0BALnpgWOSXPQbM63ihLdCq5L8lCJIxt2PE6s7j4CvKhEaLBWybZKM7+
Vxy1XQ/20NcppGcPzx6pJtvROfbQVzQvZFgVgqrQKAt7J9MhsQN7N5Xof4UgZA52
nJlWRUaXNl/hSV/1Jy+hvpjAMWUALc5Vc9I7FG+wbpbFrKvquOWnJJavIpJ271ix
fHjHNTLeSzp2QKLRGpaBsxFru3zQEUh5/U3hfjADtcky21KnbJrSlk3PonuGjvEV
33QGF1f2sUL6g8X8oxNXStlEIUuWDdmjdud3KONNCzUAY1Ic/05qbU1cao50+gpj
52wz1VE1+V/6285wtOfZT7/dmdHE2dG83PFoW6UGUqn1ka42NnrlWlwgycooI+A+
XX+j5UAbYyyi6KJ0l32gotdv7klOQA5wZ9ii52FVJEP9HrIRHF+ePrTaCaz4cArU
brZKll3270thc2+TrWRMQWguWtGJnBSRRDOc8KCupwOEovaLuIBf4+J16AF4NfG0
OUv/HFegUoeFfn/i2KN5aof3Z1fzOPPK5OLb3Wgu5s/AJ/zy63RDj/jC9J1mb0i2
o0nu9YF7rV0ocQ5W6YPakEX2ihXkQdujUkm0jqMZZfwBU0fjO7yAQMiuVkPouodN
YJ9EWYg4+pOj5G/pESsces3NFnDJCx1pkl+zQfyOkLHiLmsCTgSP05B02w/OM4VV
JmzZPmHMJ2+RhmHd9NC2D6YWbNBbClg6JBSxp2CnISUYxyiIGj14OqRnmZ+VhVak
jxIGABJKLosgKkNiG5UadEWxQqcXrCRIrYKWaJHFbDEm4cVSrE1pqtHo6okgDF3s
HvZSQLIOXEGeEBLyVHPKrZ7YYZYPsUo8py6B1sNxZKi/QONVCK0a3BuDSQWx0qEj
fJJj3QTuL415H4iOascoBA7DZMlUPkpJpIARXssbxYPpsPpQeIDQTtRso1/VJOK5
Vd2P0EfikW6gCODbUPZjVIB1c6r4uK7fbrxKuCrvHCKMw/Qs3kEq9k3jLg9EIRL9
yckqiHzmvVHnMVKlei7Of4Te5eLbePhDSkN3x3T9o9VswjLBiN2fMRexezx+o+Z9
hSeQTwwmm4lmOgS1RZ+yLd6nnQR6LQ4qESZf4WSSOBxpbi1GyDxAJ27SFKHyIOb5
0rzRVKsvCo4dtKiRaI1+T/M8ARRHaJtjW7+u/QPOR3p3l518vL9WOgfn1kLaTTIQ
iKqOgR8SiyyIVRPUudq0OubbaWjahGDMyxQmWneNxGJB45n0df85RBamPB5t0rQW
jOMUQ9xGnptNKEfUXZIshJObo17eQOVARTnXXD2Gppn52E0p+3ICEvXJp05DyX2l
nKmgYDBkLXdCOQQ1DhULRxjk7BgfRdwnQHK8B6QFeoFDcChYi2P+kjZ0WAZW4Dxe
1UgreJ4zL1T/NPA2fLnWOQ5l+xHxZigeWA9N6n3OOehV44Zqe/HoQHNsdyH03EJg
qj307BgaKmP7s0I1/Zl5w7VX2tJIdEuqz+8yvNJmqMHe3uoRLGktZBrUf/ebz5ZF
fafWuRgXXmSucsVYWDUBPsEt7OPiJLFFOUGOAHJBRRw69oMyPASb1VWSkbBCpFpm
+hSXM6QzdyYR2X6uYJj6s6OBN4tyzuDCWabttiDKgj/jEjWyvjFZWOyTQKKlWgpU
pVlZBT5sbKFVMjwSaIHOE17nRqrJ6sHScPMtmQtbg6/ZVdc94eEXscBBEv2K6ZJo
WphdLC206/u4o4/rEwjwikIL43IDdiiir+WTTiIfKLrolw/EoAgh0//1cOKF1TZt
b4BoKf9zfiEvJrhKVuvBRkUL8QEDiW1xjJOBpQruvncNFsf3WfUKqdmlriZXFXf0
orWbUsLPMCg6ItXbKGj6A3QmdUsnlh3N1w8YaGZ1SmrDQeKB+NcK72UCMNHqLFcQ
xdPd3BdeSbSgjFzM2AllnT57vAOocyv3qHOHK/8nuzOJwXkt3fTfIy3vQxIM4Z42
ByIIo8Lq7KJmWOIevg7g85zmDrYHZuQkXJwehK7cyU0bBJSLe1cudZ+gat58cceR
xKq0749DAvcEH8qcZB+UZ8/ivuNB/mBXjyUqjLmxxDm6PjKGAFncZQpf5mUp4bRw
iGvKO2C4o0fiZwunMRUW9yH+dUbOO9Mp5ltNLNTVOcrlVbo+xg+sQUXlMasB5mm2
W0Gzpm0NCdVEEJX3acnCm3w5trEaq5dlWc73DPUahk9gw+kcFsQcW7YHS7QlmClq
IH/ol7goTbrjJoIHn5csT8UPPUYWrlXM1ymetSGVXScSFx46nFCMVLKEaW7XZpb0
371HxIBFWwvvfYcQ6kii1K2eycQn+8ZtdUYPJzY0+juD9OzmJPYYXYY5DpTZqizr
suqx6ghUJGXwcMBQUdS2QztoriqndnSR7Iq/LLXwTJr58peyUQKPvk265Gtkyg8F
YfTzLpNHwU2WrwpAV7blhks1oBc5W2eMJ/mbDgDaJa4oQSVjw7AfJA+LCWP0UzW5
D8FsK/vFe/IsDqgO2iOkjbm2eeaOwm63i4dnU42HBVtd+7G+Y5ls6RiRSh6ZIFqC
a2tzJ40KaTM5RrJ70alNLY4uRrrEJKtHin/TN8yZHdyKUFMmL/TSciTZ9rTCI+YW
Nhd8uWj2kGLkqIuON5nWz4BpenN7hROPz0SESGccZMRO/KHP2g/orYzAmqc1WUyb
7y5MD1wCukkRFSqyldOGOwXuSQEmFliAvPxdMTjrm91FInWWRbMx/OJHJpZVp/JD
0WKa3u/d0V7OUHVG8RycBJO+TvdNeekCXobk4q7enD6tJ9fQZVfaAPpjXTtk/HLe
OUh+vBosj/kW26h90OE+Pv3k3ggLOIwBm3Rr5fjuTs6sEH4afGRY080rj7Uf2yMh
vBk2UbqkBDSj+eQr6tQgOV9AFcgNQObw1dljvqtQkR7AbSo1LXmv0IoRtP4zeSOd
XMweMZSLBpa6iu1yTYAxxjZvi5HXaa9De0mh4GcDUmKsL3kV6ZRRG+CXgjVFb39/
SFqdz6bSPtjcZVDSuk1H73/ym6Mt05QOSIvt/USENGcJykXZ/MeAashEUm5qlXbJ
q+kflT7g0NLjPyJoJIJtx6QrQ9ZNY7+jGkxyoo8RPaJxDvzCOVHUFOU1CaB4Lyyj
fgTQ12frHyGy66IegAr/+ouu2LlQkQI5J4AsvdRL32kFUP1cdS5XMeV8NGquRx13
VAzoF5gu8f4Hc/zyts4c7m0ha+rSMLRVLCwFnbw/PRgCwfjJ0UylP7XdWJYKExZd
C2nzlOeHTJs1KtfepgiloM7sln4E/VdDy7IMkkFc1DEEdPEcckux12Dlrb/AMj1q
OuqcDHhMHLe5gYsCMdcoerlKRPor41uy+eQfN58GPMeua88iA4msWK9F7OlGg721
gmbW5qIeVmaeX0YJ5/AcgM7PDBjVscEsBqPKmZPgEuBOzuUgOlx3Pp7b5q5SBB2M
3idZCXfk0GfBxZOS9zIC7tkdhFrmmBVhdYMH2he6XGnkzHn52Xeo6mE+/mNMET0R
Ku3Ee1RyK/jn6Uv5cjc4NoKtbSmE0ihspaYu2I05/qfB2/63rqH4zUfqDJqNXgvL
Tq4zd5EijdhdpsaICAgwlbb8LzX7JMC0pUXO3fc9GX4kcHm3/VLsBDvhuEXuMtKR
3pOc0r3w7R1pT7k5yAcbJnDn9BlTKf4TgT7SxSveuhdbqFd8F5b3U2D0ayQADdCG
8fW34IB9lW2ZfaGQVhyU7iKvzBHwn5xTXjXrDFeAKtdk3yzHEQ/ZLN3Bd7OAQH5q
JBZ+0BXrXyoXbDSnZPY4m1EiKsOaWGmWGxXIuyF4AOzCe5Sw5PwgJs4LhVbDtmhb
SuPRnWKgv0f5/69U4uQDurAiCOhcymS1JFpmyaXTohPdsHGLlvv1N+rZTyP4IyKr
JlIoo+QqngdP3jxo8O7u26qb6ggeLlO0RHXw5ITzbUj3QGBE6S/Z/SLzdAvPx1xC
FxTUcqtDhQqQFH4uT21HzhsrLKG5tJsBBBFxEv9/XFEeX3wcGKVpYYzYLYwqJDRy
S9G8yeGK29Ip9XXVwaOZXIu81r4d0k1t8H/JfSgncuYvp0v9goBkWLaX1gMTzqbu
dtif/CN9bbjC3FPvxA8de5kd1o0mdIDSsq1jGAGG1RlehBNi8abr0SceGVY+b8lX
k3JOIz2fsUw8ph6BDC+QJB8XHqUrA3qGRWwS8plUcBEJ1HqBZf25Hv0DQiE3N96A
17t3a+PRpAayULFfXQHpFeMkfkSeMbzBTyrLC1UT+0s3sd00KtOASa10Bd0oo0L+
fq2ROA5It8FQldy8I5/kQHcuYldXE4KGThnG13+ewI89mOOMb/V2UTqSdcbKNXB6
OBhtrzTM2g6zP8PKaPN/zuTiv0OhoOF6606TigkK2o2+TB3S/OIi8EXjM5hxNrKg
Pgmqk1mM/PWdJ0owQEi9MS7LS2XOPQdjzX1ueQGUX5Fm2h+/opWKMbZFWKd2PmY0
FETDniicgfZYKlcViIyQSm9NJr1RPx2tv8nH6UBVRoPPv3gxpfYYvuu97/6kbPfQ
GU/2QkLjBr/Jh2qvZ6wIvgtx4b0++ziSlEDMN1yhVlScrmRnqnQulGBJSN0EOZac
iDdsScKM1x8mcNfbms4B4kclPwDI86sbsL3tR9H+5xW0DlesUoJgEvyWQRpkrUyv
Oh6MTHYpFUJny2DB3cQGJFfwj1vlSVtBayPmsU//dsZ/2rLL4/0c6yxgXhTgZ604
t3vIjVEjrT1qj2QQ1hcJyh2PsSbM8hDYV0+hz20AYu8p3gXpcyHzXQzxPmVIBuDL
FzsDpqgR2pKjezb2TZj9zubjIn4V4WbtHuH6qxqtRUiixPCB4CepyTUs7weGyShG
x1C2cJNDaL0OhzTjzwy8xQRjWaW1DtzG4ILigUZXJdDw06qt10ufhpJWFLKu93D5
3bUwPvLsFHniRoZil9tP5+jRPL7xodM4UzUoKTi+nwMaHg762u0eePXDzfrLl5hB
YNdY6gNkwnEK2/3Pd9kN6w2tjCp1PtaDhlsiNJiiAowS2b4wg3AHzCbx9o/sQSxT
M9EQhDOmnhf1fUi0ImZ0s2fsxiF6mUkhgH8YCRM83BmGUi3aUiQqfNyyb9sD+1c8
tsGzocMZOTnSp6vV4N41KH3Gbp8tLbEijjDaRnTUfsQl+jNs38fbGiVWZRzzYQrj
TBpBjlLixeiih5T0J9NyzCOHZX4f7kiHSN9mLwPN7fTWk8496yT5HMYc+wC2nlen
pkmYTNzrkvSFJMbxP5yoQtGDdg+6lrhUZ4TBkKjgVwObzYJMPJkkDvs3ALCcy2jp
wzlNjtuwz7OmY1kfGn/aRPTtU4XcaPSmPnkTlfm90WmS83ivujAI/8lcpzaeRLss
HGcdlV1k4HVELdpJsgByh7Z5MJN/0bfkmzjdylGNgIcS0AKq4JcgB1iEygDlF5Oa
1Lz9YiOy+yJQnPzYhXmPXZYhE7Jo3/r0hq7fbJnO6zJZoGrVCvfQ++8nxHiup5qy
TwJzJshL5nsSpQ+Qo7arAys80AmksxchHlxIYguIssV97e8SxXlSu7PklTS422FD
HrGLszC64jPvai8VvgpJGE7agtm2PMIOIdVvi3Tsue3iuOFUjU0TBzIj7OEX8Lli
68F1UN81yYb+gTF6RWoE4aDdBCJ0I8C/e6XtZVXPRAzOMYbjovs3ylcK/COmlICa
SnuCR00Iu1rDQkQYlfHRrmcVUPN/I9YigUhBnWf1ltcDieVfa/fS1QJWglJSfMwO
jhz0A02GcwSAWieGPIDgDhUuFZfiHLDJXF5P9kpKUwWg8/yhjKiBv1dp7yi6b2X6
768FZ5/UsHadVod12pXKqxR1yydFgfvY1G3yXcn0qTVqjZz318uzGiT5cQtp5Ec/
ntFJi02twvyT8Q8zVrVsJwbupu2GEjPGCpTcQmCatNyKi/RzKqzCCgPIWFXsvMQ5
oRXTkjhEFjiTjRnasyDJjy52W7uwV19X8j0w302XyxBp/rS9U2BuEycQDGEvJykL
Zl3u5Ooujt5Wtb/KE6Zy89+tXhHOEe4ovO/ln97zfiR3nW18WfJkjGmbXwbBXQ7H
vshONbVTaVQNID6zV0SLSugAScsgbDIWvq4CFkQ30rRFftWQvNo22EvBBCfvv8Q0
RZQ6UyFGaqZx9HM6o1A4iQcc/NhfQM/7ZXv3LlB21E4adNdiLLghtmO0YV3Czh6t
MzdM9sWW/awEXDrRNPclwYDQSUi+Z/zdUmbmBya4Ua7qIjELzljHNiLGN7B1Tu1s
yWCVYoIUwlW3kKb/hUcMRjUBs1gUzojNl15u7uuBRcvqd4a8VAS3n69/Aq9WLHV8
RRfu989c5r6sWBXpMuxEF1H3QE9zx/FFO2J8ia8cihReOrS/7i34uJ9cDb3A7alA
h2g8DNN9820/kcPXZNAJFrPSRTQmUX3Nehnz/2rKi5YtSTzC1NQKPr/OvRyBXh4X
lmh596uqSsTUxqM/+JDA4+YVb5CU7M0xS7jFp70NiYDx+MBQXpvf5mJx0TNh3wwr
qkn78lNx9g6QevU+h9FyU7du2IQs4STuDY1r7VBIOm6SLD7begfaSzHV5vlNmkPK
8/Y5Hi6E9oevj0oWu6jpfjNkrHocmvfUKb09Xq7mqLtfmYj1otyFomkPRm9rbxdf
Jj0W4ojjbXjL5MkPcuRArYev/LU3UJqCkLOebh2ZtgeUtGpcDfubnMPW6+rokYfO
xOUTjWad6J3AHEhfzQB4r2BS8qx8A9g0i2MQU+ZVtrJj4mUIMcv9QBm8rXNNkhki
TlE3fVlSi1OJs8Htia2cxoNJSrqi+7T1yWfJrExrCBstvqR9mIDHgSvvVMT3ko9P
b+xXFa9hqQjiVH9xllfdXLHJPS7alV5H3hQUZxOUS2sONOC/5228w1KPnRbxKlYM
B7/rtSL02vU5Ii8+RbuXpcEbfun6zDfdw8yJc4S0/sHS1xmmGYQqja7rAsqy2kSh
CYP+b+RyMPiVSjTegCn1mdAIzD1P5TL34YJ/7iPOAwlX1HutCdADJ7pN3gvOOapi
XR+bWOS0ySLLznfYxjgGB8+BbJ0wf0/fKfJjexxUFy4vrVsseP+LZXaAh3XE7J0I
9DBxJi3vZLMvZOuqMXoIJbJwghE9vmWGB7QDUschWjmQcv3Rk7777jgG7TXL63ir
lVttPiQvi04XDR5ztWsCcoiVzGWMJk3QnPjbZlD7Lw/6BQQALIga+csgfLeM87lC
ufzZi6KuprSF913vwOYMCy85BTnCdTsy9xGR3e1GZQ6pmS1xHB8/AjqasTLYTY2g
8mykM71Md4TFeyJVIh0S7gxi0b1oQ0wp7qD1Cb6XLmXJHIXwNHcIfjUsbtwyrRka
Bu/cwhg/WPW8ixsYSV3Rl+NNtoEHS0YmMBnR+eSzYxvTq/dDWeqAElrjRncBMZN0
a5mrtGlVixFYbdXXpqpHSUpSNZzq38+ed0ES9d0Ocs+SFvNVaOq5nw+aQUNDpYjQ
S9YLv9IozFRBAt7WPQfyRHhT8PJ9jCMS2Iye8Zsob304nt1TiVjYdyhYgEw02U/I
wrDW3mhYhtxosr4pLTRulj6DGn6/mb5nXC7SGTkWD3eClA+XFRmgwXsrnlazmO1I
gcuIeUCh+3UQlJuXT0JONiq+qPaE5pZsGxqFGg0PxFzq6fc/fEFKp7pu3pAWcVJD
SFlINrsgQixt6YIQy1RyFWq6t/WDWeMVPMX8FpChAKqboKk08VxiTCDY3AJjO00j
9BNbetAyWcY0aPDCqvKz1TVIL/ZJCy7ekCa3RCHqG1Uf2h7GA8lcYORyCHtWJvt1
zutYqcLDh10EIqdVJliPhF0VZlWBLifHCUHVTAUMd86kCLOUhwNILcKXdN4SQDai
Qolew5p+58gofeY3Y32f+f9Pv0zJmtDtNiFjjZcwx0z2Ytqq0kJm3M3ah29jXgYk
Pr+jV0S/Tk+DlvfFxTWIK7h6Y1OwTBVAyW8nAVsX1BQLqn7PEMTqJggr4wqzU1Za
XfE6oSHrgAkQyA1ysmiuTcesBfYoRgBB0GbcjfRfgn3PXVEHQW7HrjrwHjFQkUNQ
WGm83JTHesR7lSzM6Tsd2uQVLT8wQwewjYImk0cZmIKDN0Vq37gGTCKlnnXH3EyC
mTJfkMhVOFOdU2x5M9ydmAlZ7AGV20TkFRH42LDm6ZSwT8TRi+y5XTGijNybJA3x
yFbHi48dAI+FwtW1W072Cdu05R5WVaLiOBb4HxuJ25KdNILxFJYMzwjwI91d2Lnz
nUssaaoFFzXx4StA6pu8hMe8qY09lNrqtH1EBSZ9fgk++xNt1CCZRQlCL2Lbolht
6Fx26osV9QtRLr/XU+0D6JwkoFp11lBkoGhILO0Nl9a/lm+Lzd21xxMuQA/42Ecl
/1FHBYusOmUA2STmzYeH+R14DTgZP0agQ9FhZ0yZihk7dYEhL9/4OemnjtTAdA+c
yzutYoXFisvI+2FQUvD+Vo3ACE5U33I/CeWQ5bqYtFXL+XQjUSzRxf6Omqd9vjcE
V5sj/s7hjRFLvMw30wym+qqx+psnhn4pMVS/aVfKqgBzOQq1494RkM1T70KovQ4v
/M+Wyu3eXBYoAKuE6tCpzhhu+W6TrNhqtuRGgSeDC4XCc9TiwmEYZN3gctmlrxkh
NH8Sg3biTPlRGJ8VBcRuQJPaYBwAAwdT1CYik+vAciu+NMPWfNZkkcaDTU6RGWOn
w1287MsNTB/phvKi4UKfBnrohLVM/vVSltIFJ5/zPH45fNZZVnUIVkLaHOisWe9z
fpnAZe545Ulmky7uM3GdJNX48BYsqRqOKet58QUNkBpjjqTnL3dDjvnJq4MhpAIV
9qW5UserjEenyl9yaHY1SUDx3fPAfW1olNMvpmf7yfJFEONNQtfDvNGSZ+/9/3pS
bD01pHG/BUVMo9+9Lfbn5uLZ379m4jH6dWYLdFdWI6rPD0gGUGNyOEfe1JoOXDTP
wOnALglYF5nnH3q9DarSUqzZp5pzFXt04+3Clu24ohfxzYV/mW9H70O/LXLHTyWw
OVhesbFQMwu+vBQP/+67A9T3H1tx1Y3s/dXErO0E97Y4SPFFk4IS66jiQUdcsdNZ
2VgZhsTrBLTCU0p050O6PI1lNye99rtAsEUPTE8nkH0FwMcEBWnLhSNjsBNkI/3C
CF3H4fWNBMXqa9b7n8uEex5rmmLRugS7Gmu0zG8dJzy3Yw0HMbEOdhGZDjRuAhih
AKmh+LsTVVvmjS0/zK4+4euTqlRGvVudRrRchwFh0e0wF5FmrmcJv9EMMeUUjg89
bWfHMLtalUqSaZF6I4hVbuz7Do0HugaZE8YPzr/YuKcVD6SZQTaoBYqyqj0qssb8
M6J+11MMezJmfgIdtS637zT848ptJU2VOn4EpVvRKc0voqqOhH8r1uR26lHu5Dfr
FIkTboeyLXG37s0vLWzkXJuKGSKl8XwvDVoc146dnpyiwR4jEwKiK3njANd1Oh4x
DPfRYGmyN/uGSWaYSh3aJ3YvtjiMaPSv8IF+W7tdNs3FfOL4cBroTDN96XqAJAT1
rLZxwNB7A0i8wW0wltnjgoMCZGPaoh2aoX8VtCVTNrbEVnxeRzz6wJ467ZSGMUMB
YcPrGIP8ZfVOAK34yiJEA1QiTwA6h7HTxWOxMxOplyBsysrpEwq6sXSIrbJ5YKRC
5pU2MrIKk5M60qjD1UbiPwMu0ymwGDTwE17LfwGuYcaUSdEYPOE9ek7xuV3pYxUu
rpuX4MVrGej7CQkjJmFs5nMTWSEyyiT+b9b7MUX6hIIhmC3ri2jOXqDYrpKs0Ufg
wk80Jnvc6lBQBaAcoMpnAn2FHPUaLJC6PVLZ0gP0yY65r5dDIEJvELKbNLbZ4suh
ExT28UshiIZWWtkjF/ssGb1vh020Lpqu5G4SMdpIy+MN+iLkB4tmiQ+uE09dyfsp
2QkhP1EHgpMGL7o8Q8hx9qNNXfWKWQtmpMhclpd6RWX5obfrSmvoYj2uOlDB6yGK
+LUWIyO1FR4YiqcVEStGRcb3o1IBe3FMMotyQSnSvhrR2YZtjA1QPDJYX9+V1pTM
tPVGpeD8Z2N61k6a4USr85q9ueudMLR7+cNdw3rjRKHFaYgtrWObMdUusadmsOln
U6lNvpZ2YPiucz1XRqQycordAYOwxDHVHrH+Re+MP+NGMDPY58Bc9ElCDlkXiCEU
Axb89RqoS+bWVFR/WNYjyOaXN45Xk1tpLQHHqwsJ42vgHaa/lZKQWrPcRqbTLI2N
4rj4z2AY02lwSzhM7YEp4kYnuqEAtgEPrNCx3UMvb4W2dJ1Nz1e3vYOtBV4f6yGn
eplRbn7pgRT4TLCn/9WYeeiMt7RIVGSKD69y6yc2vGUfiRakiDz+Tiyt/iiTXmCM
wG8eiH/vbBD2yj4gnC1a7c0OvStufvpG2+zgkKINg2gEAhR7oAIHFQpjTYDFDmHr
PP2V/ZevWiYcutyQHhAIDhSWRoMnpwS83v3Z/g1JJ/uJg2iJS3xrduLULY5hPQ39
xiESvXwUam+b14D8ECv2KIwx6TTwdacNMXoHsF9J9wq62zyaeELjBl5R1KO3tVV4
hSGbNrn9/QlXq9bP9/mVSHfH3TKfhp360tGOXsuc5dDBi2uxi4T03aZlOaX2LJFK
3cu0S8n/NSMOxjRcCGgjO7kj7lC7Iksd86SgqMpx/6hyu2kSLzzzd6+oz70BuAFu
SJNP/KuVL/3C0JgDDPfMz2ZbbcJRtW5SjsKUM2Uqc2li+EJojv9Mtu43M6xifJGv
+oa4QH6oONseC+uDKYLR3V/ZOF966rb0gd1leBrLJoR7bTVV6nOtEYNwnoyT/StR
YNpQXXc2HOKn+T4EExrfSpHrIOzsQ6bluojSVgn2CVIIysB7nyY/xx0i+F1YvWBa
3/ZqU1k3Nqgdh5tuurYa32Oj/501s8UI6fVivkUAKA34mmwOTe8zoGVR4Sbkd9XX
Dyssy3Vaeg0DeUhMcFTjTM5b3RReftQTp0/g2FLNwfVdjE1IPjcY6QpKk0v5bqF2
u/v7SDMTzE8cj7E3TJ+/HOGhtcio/feCx9GKrTVn+tB82O7bTLSdIKFdSTGiJj+j
aGJpVFHaMyi5VMgtno3Pc/xdE5czqDrNmAToPYb/ldLfPyAEgGiCddRm+5vPlbFs
9p9AhjHxCzhQqbV/eU57tQyS8Q0QQG8Ib/5d1QMDBiC8rAhqkh9gfZg0+Yc54cSs
iUPNMaNup/MjlH9EYTqGt47i3pPG+aHc2RUJmYTLHNy2ehoOV7AfxCqUQBeNuW5y
RGmwhntWdKUY7M4wSujZY3BXuS4hgVxxHC64bfBqkSg4xNp9KG2t4Dga5VEFTFF7
tqdwpgsBCdQID6EsBjd3KV0X8MKyk+zgU+ACSiaFHt24gJXn8e7655YvFrTuTffu
oSOAQPRiukoNPsJBXDHqg+lJCrR2tXtFaLhCvL71Gz0b1pNwXKJJfVyiWH3Cf7nk
XVM4JgIiWRF5x5Df/F9mLgKz60BZZ82eGWToDcnvyNy/lF5lOmJXI9CNurQeOagp
L1CR0XG+vq/cxhCxHqYth0JUh7F7JxlzHucJsWkSPN+AAU7wUyqJ0zeM/H3HBLD9
o1owtQ0m4CxZ/ywePSHFhWC2Eyj9qRnST0S8Oe/ARs+BM7ilFXVxav5Ld+SVSAUZ
Wdq4pjdG1FA1DkI90LB4hQO1saIH058Z5aEoTAAYq/lTNrLkWnXCSHxx/NUg8iH8
7fILglawfuP24Rj4HxIda1HGZD3R2plZKYTNit35uADV1tbgjotksOYPtdA1XgKX
BazK5yUCDPCWcF4z2flMGsF+W6tMfG6IvKWrWnJ6bVntZvRSKjezdGxVCOK7tkd2
rmMaIP2IWUvGEz8HaTl4KiiqP3zPiXJHD/vJVyg9xhta2zAU/PEUX7wIJPBIy2UD
K+OubBhbYmA7h4hVNFf+VkpfOs8A6SKtDCSy1/mkzu+RHjS6C2ejSV5wce4tjRG8
Myrq+CI0HVSOCNHKsfKFEVqe55V1VDoDMsFLXfPBI1SnPUbWN0NdcRdeGqgm0ySJ
vLwk3zwIaPYpIRo3BfOtpYAV4xQawV5/zJs4yLrqR5GW1ObBvsYx2WqD+Numx7Zs
gV00qtVyiitkG2VnyNO4Ls1K4RB5ZN3fN6DHSkj1XeTMtrEgRcNx9nqLxKl6IKvl
mbXTtLp0RH0/JmAAvl1rx4KNj6GKhiSWWwsA601KS3zFoHrivmPiV4AqBMHAJzFL
UNjawgGwi7oTBo5/KTZQa/yrXozkhBGBS379hmy5Bld163pt/15WZLQVPhka7kxw
uDulxzZ/nZHPVaL2fPJVJL31uCfo0H6j/lCw2v+tf+d97UjTzJtFdE/LT+87Ey5P
duY+dUbFMttq6cKILUmKXbGilkMdckcacB72YECccJeJXN6dC7mSOZUtNkT8nJfM
fIhlR36qo6epu2MoA34AQcXeKjNzhmwuxMADWLDDbNDhzN0A72H26SHiTW7Blmt3
WSGArvW2Uk5HSxyyq1daZzLofs2WWFD69ajPeQm4boLcvm2JZ71pAM8F288fT77Q
J1AeJhgr5WeiuLXXHFDwSREOiDrRTOOL6lFcWMmBlxdThOoKL4+/e0tGO+0SXzYb
5JOtr4HRAya4p3xAW1pu72qxK7aaWSvnycapNGvM1bY+xJTySrAM1Aj2z8+b7mVE
hxc779xjNwyLMqtfpZJUUlF/e6OtY4t1Y8Ylg8T6/ocAUmDN2QLLtXSi9QEq0/0/
B7ah6Tm0JXRrDSPOQn+cXyvz3fYwLfk6l6qG/GOcYP8F541lbNi8qM/zaZhva0dq
iDLIWOEOqqkqFvipqlvOXqMnKD/uALvRfgObiLoX+gJuEEPl68L6EVskiYQItdbR
DUQWN1bv/RmrdaxAz7fXDyWac4oRGu6nt1+Iq/P/rw2asrNiE7dW90TPth8QxZ4d
S8KwwWylZVPLJ1NJQfVRmRpETkefLwh87h52xbQQJZBsBEJU+VqpwNUj9o/BZjZ+
JwxyGQ4tlhrq30lLRYB/crXv2n/aImBujVloQPaUzOM//BXS7cfGnbdFXmOK4yFw
Y/2oePuvTSqjPj9bDbQyVXOHLzgkS4cs++06rqhh4y3xYSiM7d4zRkUOyZZr5pVh
FtdxL3Zy/UZsDXXsleYPb5aYcyMZCQRJB2S0sbSde7wcHiJcxvd5RhxGAMEfoWpF
/gAWQCIfi6wAk8GuU0S35Uz5mP9q1rhNOJewm+/6YyeaE6KQQ/HrEPu430dYErKc
gmfRTfY1Y8vgqhcqpmaB3+sAlX3W0gOhAxSv7U5Jji5VLCNFc7pxyfBUrZ6vDrD8
kBbUeEEVh6sEXqs9u0hd2mQmVvY5c1vMXbF1ZOVe+lhrCEDV2x/+YwMEP7EE9KrZ
pI7f1m5PdPnRACmyjFRqP9flgC54hEf2RDsfWo7JJ91z4aguc3EGnis9dAhjr/Qo
E07HFFwPD1LKUucdlI/wvnL80DKNI6N+P+rmnxM5BQnt8etQWB2KV3K3+bsA8BQJ
FvK9qRiIPd68g00AeO6gfzdeqyAGu2IDDgpwAfqSmtd0d9CKx3pERFid6/0qWCJh
rjtHRQHviV/05GipS0uZLOQVLZICMCm36TiBSIHtcjmoOgweflMHOOeNW05RyU2d
+VSrcHpMHwfych9Y55lscAUlglpdRkxuyWbybxvg+CHGmMn8aSt+9s7Q+AdR/nnK
yRYfVb73vzpACFYO6sxuu/B9DclklDBMHR2iX9O9bmaSzJui3LfOPMsiTqWm9W0x
0EK2vxo7rhoS7zEfVXf/PKZsAUwkaohWKX6doZZzhVv9SwFPF/gZ+MoBepnQPMG7
aq7o5lSszXZD45koBKW9Qhf9Obr1gJ2wCRu9kylquEivXQnQkjpyC8gPjGAVWoTr
aw4UbpYHv4vIikEipz4eXNAGfUvuy0QUt3wcpm/cufy/wB4rkfeQBunZx/snaZ84
/B5kCvCLdZcA+oLibFRrXoWxO0pqBUCpQy+zWqVYV6xEcWVtjnaS6T5qes1qocc6
jYCkRB0oI4OfxcDL8ymY/xR7EDG9uxRjfF3D0V9jj3GAOL9IiprL8fe5/8QZnwuy
5joje8hICelUQcAvbenrXahCtGGQxl81kBByn8Yc1M4uRgDMnQ1jNhehXB1380z9
28fSfsOyqqU7/9akuer14RljKO+a4N5TPPqqJp+EOcpOWkA35j99CNFKOxS2/rgZ
mLYGmxYHEmJ0f5+sGbLAflIFuUl3CIfZ/N6Wu1DOmdmfa4NigSCg0mRZgQ68DZ8w
CB17J5gILW06XzCfhaVJJdD/VovAl1vViNLUg4Jdq/GtEiI+WOUGIhN33vNVE79y
8piPcVsNtMEQkYAIdrvVsIqIrXTf5DG0wIlrPStCw64xboxq7IuWXhqwhe9FdcDi
pq6YNKCmDwqTzUqQTwyHrYnNoKY4icC3nAIa9DqiSwqY30/x0JSTR3eymv57xjqk
zFUj1yasTUAtHpPmQDFY8aZ1PmtcDWJbglC3Hi2RE0E3Dg/mhG/7NqkEuwOPh0/C
qqtf75CoJ+72Pwy9FZHFZUUZp177eKJVfxiNIlCIuzJyBeNbskU6YXa9RR2Esogv
VIh9ufi4V7iB6PC06aV39gW2G/0Obtgov8UXRZnr8/5aSX4YGActggjx7+SFabMF
DPTcqBPRmDD7B4sXEi2smD1a+bFvtTCs99h7KRxIroeAqST61eEAg/YOUv7pvTlW
Yxz8XAqbYxTaYQAfcfuScRp1yG7X6q1P+FVG4AUG6DxAdYe/4WJ2jP/c9XTu1iT6
wx6zDE/rCkiieOo9CMHV4BGN3bf5+wTqVJC0JLg1ABeRO+4gfGWXWQU7l0F4t7S4
fMyYhEUjk8G/aV5i7kKKQleT8dj0MfU/Qav2X0Ur9SKUqHa0YyAw4DRN7lYfg3Bn
dCApU4l9y4BSZggjl8g6peXB10OW98/Iqqng8TOukxarb1hH86ItCqh/y3sMj1xY
y8lm3Hm2yFI1BsdwKyY17yPMVYEBT309XEnNQ2FJjcvHfEMZ+4sxx0JDW5OKEo2E
mBvcSY0Qv2v181lcEvwNEk2Dq8+1AycsaQzvvacpXt03kD43zrbCDXiyk1K3UD7P
z+/+Nguz9VqQmoIVxkbzQqBPph1AEermM1wI8ivyNyKdF69bMy94hmOeOEdJh8ZP
ARj5n0sODlVtghNHOvbKfR8FjRawA1qy1ZoFyAvPykG6Bn4NAYs/OI1j3+TpkOk/
hpbmf2R0wmkVfbQ9jenpBbONEzhS4WoRShJ8dYdPv7tL3HDycTwWkmoO+WtEqmw6
9zAwbcrPR74LdxIh35oUvS2XIVa+zr9Mxq1HrdGAeqkQ4MTKSe3OfDbyz0I0t7pP
sO4UvagjntEhYlpBP3kj5geC0QMG4+CRSmVnyEDIp61jteyTqh5jJv0B/cwLeQvA
z0ZB6nAd9K0LWC+6DYB7hd7rQ7Z0+zkcPNEwPUgJZbk8ltbm8wNOuyu4qEG7Tm5Y
OOzCk1L9lqxcnL7KZ+QQSVOLWsOXajtXWERGNgonkKJxq0Ec2wHuoqlXvqjNxldB
Win6G3yABtP0OkS4NzhkEbp6NJsdU4n7IGimbGkRoY2D26h2xFIHZebP24dU7qdr
n+CpQDB+7HOJFeM64G0ZYPh8rlNAz51ZM6zlXZN0S6Bo7nVtoKdp5lpMnmsO9ERG
NcHaq+8BN32Hv9TvgnLChz8VSD+6Q15Nsojz/Rsu6+8i+2quF+oPNuLXjuhivIBj
bqxC1f0EoAufX7uCFk1eTZhbUPLnk6qppiJVINLMaSpQRcrptEiiwWnD5FXtWEeF
cy6C3PKc1ljTcbI9D4SUGCWH/KNSPKfK9FVCE6saqY5Tx6b8NhaTFWZenGocw1vG
WFfS9dvbpAniHiQWfm9v6Qn++I8kKoPaByA/6EqGxV3xtHJD5wmmjtnEXXx2WIkn
c4woi5Lf1R8U0vyZLCXjqTtdEdvA5w479QnkN9uEBwG3DaJpP2efEKucmuyQFEWI
rsJSgB9f55DVtbv6tST2DpuNkEOFez3rZs69z2l2kdC4dhSFNYTfRWmrUKhFhxY3
ni7wLzlLIp1ffasfOn3E+v0VdT8lXBU01YJP2bu5CFD+mBisXhWwGtpoaOzbVIAd
8hlFGpGBxNDd/t7/o0hld8L/7TmpTMQhr+mY4d9KN6XSc2IyR2+XWIEN+S16enG9
egpL7WBQlUHQO7TtW5g9nSIsl9dDIZ8ow7BFf+Z1AF8tGcZ6Ubor3e2fL9mvPzpa
obZcjElj06grDyiO4WvBzAcArsbcNieZ+MMGMfmtxmMDW6J9mxBWXSCuOgjpHaxx
97OMmFZXRS2ldXuAsVBsBQLNixiy0pLnoUNQkXgsrfUPWJD0V9QnVe3SZ8OxfWKQ
vy7wXqbFj411Z2M+kM1f4uKSzFeTALWQl96CaDAu8i/u2OAxI5sMvbNAMr60zHqE
cByx9fy5klmXApCVjdoTY5BtDu79GJTPxq++k6bmtE0zwJZQjvdXWbH75uN2M0Bx
NnuuxpjXM2bMey/k5zFbUN9ACZJhTlIUC0MVSmZo2jlH84EDQjiUhO6b0M9tMp6H
0IxUCm4CRGCAfU9CmtcjhLRrwfJtazeovD/UEWgQlGx2GIdlEuX6+wjO0DBgNQGR
d+dbUmB595U7vShV28mA8uiWXOz7wHhpuMt01ag4RKkvbsjpUlfU48lAeSaD0yvz
ZQNasR4VHaVtb2NsSCfUVuEwCQR8kbZqvQAKq79LEDSSarxrcprWgBjqXdE7Hx2N
LPeqPsC989jxokHs8i27Cc6IQ/2+LYV6ie/xER9IMxrNSSmM4iuG9XmAuRRNtcAz
Zi/Bj7vkUBuae7iLK8V63UrdoZGMpqmrga1NQd0sfV2C6DqPwcVkV25yiIf9D7eu
CWhejtzhADIeR1Y5Aqh5wIfU5FC4P5MXsl1CthadfwF5InuC5g2AvTzjjDiAsiJI
I7VEyzls1aQ4ECjZF8PW4HrrZRxQ/Oi3HE4MtSBEChFeSgK1iBU5wOXYKIckztUR
TJeIzZOaI1FK5DnTpX1cEsPAvYPMUH15PfX9V8UlloNM681mu2yRHwgaasHi68Vc
xKnMpvtZxu+5VULV9Eq0fs4QnYV6L3zeYZCqFTdyMYUc54UCufGQ1rcFobynAtZp
tXyvYpK7bTrN6XTKoQp+qHgG6s6Xdktt1CWNoXmZdZi/gThLqFNQcdPOhLFIR7WT
c/8Y23BpC82YM6NX1sXK1b7YGSkjSW0FXclPA2RN3uoJaxolKMFLO0b2eirTPOKQ
VrUqd4SxC5mKSmey9MwuJE1ltISxNafO3Wo5lZdki1eJJRFbQVYpi6obE40IW7gr
LsF2iFaQcl9tTEILTJMluo3exzCTOKSVQieNBDDvCFHfsYcBV2okVfFHaarumu4Q
cRXLUp8Vh0Xl5osZy7PRNPbU4sfpqljiIJLbRlXO74H1CFVU2/AQ8EccswTl/jld
U2D1KiBnkcE5Nsgx2GyHEhULS6LfRBzJvxaNcGT2WDbN0OpN0XZAxYSjz1op5OcL
G8oTsClxB/1mjrM0NkfArDfgdKhIkfIOudI7EgXyOlu1GGut+Gn5rVkVehSJyIhA
0s3UsYUvMKId4R+OiAnDxb3hd5p7SiM70LZ/jG3WV4mPqVzu5uFLdOuJlostLqED
9EEpzpStsOvknjSZcTzpeaKSssN2yoGSSk1gqDve15MQ5VfV9HZMM3aexnCUJHgT
FJqGC1rwc4mNIQpU7HpsRs6NnzZICURsFUfPH5jhl18Fiq3Cb2VKtOkBfU58U2MZ
lLGUSHPtSYO1kJPx+4OxhjT4/fOUvSKBRrgkHqAzoD6Ml/MAyw7wBrWECk2k/A+Q
hoH4DpqgH+25X0gvpEBBGkafwgb2oXP535UMxXlx3NKWUvwhb3b+KTJgDZa7VAAk
k62OJzRl0+57ZlpOQfQqOyLsm1mZ/nY19UsdWB/hqhQ+N7C3cvfxxyr5nhDrUWmz
U63kFt2RVcA7AvaBAuLR+AyGA4kEejH00Gae0zPG7CYsHws6jtFr+VLYZJU21QN5
2tM7tEYDmZ1pBAl7PZnw4yygPqqrfAOvHveEUBSZiWPCU/QHPe0glpVA7MDq3SPd
ed4PqK1FYgRIU4zLoIDmKzFEctl7dcKkXWwANrV7DUa7c4MH0/uBFRT3YUK9XFJ3
2TwbZ3yhX5jTvMK5syB9Yz0QD+rSiWg3LiRy0SJQpFyOKQgYttWf7ePeeuRNer26
c1NW3nfTUK1dwfL7zgurwmTqp6FVxT9RkgskPwD8uxBWQeLG8eDZMwYUgl5y2uFs
IM/dMfgyVe0HNO5AyeXQh//H8Kq5VJL+D8D4OrthjlC9LJ7rXlYwGsOYl3LFlnW2
ijq9mm6S3OSJU/tA7loq7eiGntXQzWpV8ue39Y+CMCLX7XeQMAE5jFSPFpBZdiC1
H/0fcnR7uyhbGzlW8R6Ce6zJ0j7glEyEeJ+EoL7oFM4J8VsBFJ000ObjXA3R1zf7
1u4Lrg3iiQg9dR10lOUrtp5KUirG9eEeTwBikAkyzVJ1tyNJJAi9ZfD2r1IrHKfJ
t6Gvwwdq0GuOu8tkm9s+qkQvFpkHa4ztvte3EhlPk95rBPxdJv7INI6HeF2Y7JHp
IFy0niFCANt2NVHdx/ad38gPipRE2XlX5lIFUN01D3tcU9+DNMODE4JBfYGq5CT8
xEwnsC6+8W2XcT3/1HbvRNiP25rqAkp2iWD4ZqQTw4gs7Y1BBV4cgH7J/8DHSSP1
YhbAvhyf5lVXX5IJmezwEm+n0dJvADYQsnHKh+742vySH3iXfjpmBS02kHJBGMMn
C32KJsyqPjdKnX7Je2TwDSXZMYxI6Ka6waoz0u4C1cv3zyM9LtkzP3Pqd1m8f9F5
oQl8cNkByEr5XUdXhmK1aypKg+a3qHVqkR1tXCt0lgV4h/B+57iTpkU3PDWTib/B
b+hY4xetVBRI0u03lbamXrJoQXbJwCF39E1fpyrY86IKw9iFhFsgb8zojpYbYM3w
a8MII4wJbHzkg9VAjEqz2JkyrMVsXPIEQjLWCxqqipKJDJ3hBr6/66V30273jrm8
h4ubB01zXIOTTUDqlxGZkFo80NDO34Fp4DAks2subkBIvomnDttNeeDML36VGNps
neiZKV90GeQDjDpIbGqm2QqqwAHB2N5mt+0C0pT6Qaf0DVoukVOe9fyJxSFgckGX
HdbEs62rvuQ8lTAJoC9Jr1MuHDhnblwQDeC/bJ7yhL07Sk+998JYKIDmDv4E1Df0
4gOMiGL1BOWkMoTa6PTdXrSsTe6HYHYWXpCm2/01Mz2/yA3KH4koCTcN6JhPrHiY
0L7bY3lTu+SSeb7U6gLOzrVKi2N/7i3p9YGFYXHVzV6YF/lcHqfxZeOOgzdGgdf+
W/6aU+lHFTMDWPW2MC71AWp8sPxIODlSvgNozSvcYhi4If45NPCXIoDOYNj8obQK
t49N1eigycVWNTtlg+jprCOo2veq07pD6bnNsCJ6OM5oI/3h9WG+gAqy27EGwVD7
s1zVoyOk122FJwjWIKtRnzQgAxVxJQi29mFnft8VRPLSZCtGQKboG1EyL0Cd0pMl
KXD6JeYvgDUD9Onozz8xCQOfywOnMkqOgwbaP8il0s7ezrpEqm0Nn2TV9lSNxaG4
7XbpiP4htH5wW8z5E0OR85R+7oReotm3O+0C1Trw2BkWzRBAOgedVYakCn12JpJ5
L3YfXBkmz81gSp3HJ9EPO5jVke4TdmU/hOIjhXFEkeS5c9oxah1beEeH3XqFXUGx
ryQhZ9arxSdhtHcxl8kFmQb9mETT0iU40yC++L/MqjLczUjr/JUHjoQMp9Ico1Ne
h/boXtOYjJsT7xQWEdBw7wtXOJJsK4dJACOHNi0K81g+z5tFd4onfNFB7IGDelRy
7hEoWo4E1ZrKGDs6qpWHg+g5cbd5h/GK9jLshLFk17SQVu0/sKkisBnc1NqcCl+Q
BLso8GC6sRfthOGQvU7B1FzJoNXYr6Vw/THm86OMcSkHVbXBhr+b36lgjGJQA12X
eO1hyzgr8t5DzErc0QMxraXJsCngFl+SraHWaP2JsY32jziE+T7EZ27QOdV/bju4
56WSKaiyyyvV61i549/3ttwXM2Y0h4H9AcXFOQlAs/gAsCn18feYYrvwkrrIsPZF
9Vszf5pFVNh+17oUOATclhcdTO1DJAOkcfngM4FWlnuPwNgjuOuJzAmoIpwsF/Gv
ZSHRIHxyuK5TrQDz3zyda5e3imlPIH+SL9ccBAYh78h4vRnaitHzPyv00lZI7NSP
REt1n1/FPfHGOQJ7oNnK7SthAjvX+8gC4INrpXYBy5xsfj2G1W+JpADHHh7Js+d5
FpkozTVEy24xRYxZjvGeELgbxweMoJhQzz/lwwJgq2w8ecA1OsEMdB8zgojXvhV9
wJ9UAma2w7tfs5xqExgWgIQM6nRP9macTzGB/7UnQI60D0/yuFzG+Qmd3TTOo5El
0al+n9HK8q7j+cJ1Gd6rGSSMO7xyXDW4AK3ydgoOQ12tKKIOr5RUbu13LHb8emYG
1vSZ9lEJ3LWmBiNSv0KIHiYHEJNspHrT0P1uE+dNLtnyVxgoxLwpfjX4ye5qNlkG
sOXONNvW3iVTxYwBdkE5tyWyUCpa/vKGaE/x1ZyM3NackbL4tCOk6g7a60mcg6yu
Rj+SGfkityayjOl7INkGfR7qplYIYOiFJkSJb6egNsebHR/iDMS2qzriewxvKSC1
5lamjTOyK1iqAqcXLPL49eHfAx4qnTSN5jlcHMv1qzl1eMWOGFvRaYsAMOnqrFyV
p37FzfBEIOklKeiXjZpDIt1ezEiq133AgXadAaTsUeiK3VtidjPfgbcMyVMgWVtd
rG/idKaZ93AAGYJSPsVN4VevhweBRKPdIU0NYkfTjyuADoENl80PmmBHo9d0FgxH
6ZIDhhO06u0KyPZKLsMo3spfrlC2cfxEhwEJkTEugTu9l61LE5JH0BOLx79641Sn
IKaGRerwnzH5O8zlRIN+fIy7j+OikUbn1b6Fxxdli7AM7uIYqMYxZxu5VskiLW1a
dujCdb8vJMhz3qbGaOWSbXtaVfpism3hGanT45t3UgubXHAksV9IopFOIwfmxmC7
dl5x9Xur9ebkNbjys5I7kkm5Fn/BOTHvcIbgncDkyaEQjtylAZFUWV9EM6ZSjsjU
0ywdACzj0FWGPXCZrAB8aH3Y7qI9Y31Io6BwUdRyUkHGMmxMN8EVG/nwgWiKWGr8
INysbZy9I/jwe02xpBNts55G3dAT/D3BKpIJoM2XGjW+Eo5Lv/Ztxepl+BTK6adl
fB/QnoCdODHeKHhf4whJbusnv56LHDh1wK8WLwlEIxy5jCw8I2qvfBDeoVaw0kdJ
ZjE+mdIXqXCGZUKYbZKuwOHEgbVLWBBBEi+TAXN8IlPPMDZkuPnT8etQwfQ72pg1
+kEx6a1dj6hl1mIg/NyO31COOKQC27Fl8yeyncyg0reAnLmKlJwJBskK/VuIrkum
ywyPihfvqD0JXuPFLYSXOAy93tl7iK9Hhgj/i85RtcGpP9iPHglTXfLkTk+rZc+0
xufzjiEcws6GO813Lwh44ErjigfTfVrbqFiqrrmF8IvQvxQOrNUwXO+SmU5SlZy8
g741Xgk5FEnHtQLtlv4islDatFQVeQehqeIjTMICtvIyx3+Mno0OfD+PSqffw756
mdhwrMu56paKRpmPA6/hfKhuXbIwCQwXi6PRH0VZpbZvurxEj3Jrh5FXmYE9S0ay
euH44x72ScSguS3UE6tUjtBR4Co8fmhw2P/kXQKNYhqk4QKIBibZRJRltNE+awh2
k2M9lVkmJEUPMkKiqYK1uKytphd8rTUtmJc/b3U6Zo6Rt6pd4+Bnn8PWekrt65OU
CQqDZQgPEHNVHDO5ZKyg66ziatMMSAh5J4FyRFLEhYEi9T+5EiuWtHPHtXu0acLR
DHSsK7eMUXyLRHt7cvUqNeK6JZaE35OthXXzTSOkxeEk0hcyJkx7VcXpuA6Aow2d
h4/y9wGOUGI+LBE6Xiz/VusKcfkzwu3Tap48x7tsB23wAYz1PU3+XkPoge9v8Uv5
uGOXlGHWOPTGQkmDF4zuaT/kRyoYPXzjULFpA6CePhKBapRKeQNLUjV6X5YvlF7D
NRGGo/G7VhgHWylniWeLMT4A78+5lX+btu8rA7s74CMfgJkitlpGDpi9/K9oIWkN
YTRXZ4pJCPSKgY8+u/85XTFk/+57YGMOuWKKZSsMN5TzzvN8zeF42XPTPfaAfSS+
odaERxLzwcfjm0lsBFhUlIjJsTopnlHV0c2V9NXaoDlws4IOAAvFXbPI6c4EbJCz
SE1vrIC3+0rwqwOrTvedsIsAGXroLAtFOMucr10Pa6jxYUQ4xVYw/NzWr/59GuIJ
0QSV/Vxnp9uPrbCI5aRiHOqvIuJrYlOiQnSvXCa3WgGBr48j5aOuWWSjNNQ/sIvE
GTSmoBwPFa2B/bApFmzWb+sCLk6x7FoFGqLyN7pW2OwvHf4a0kqs0X0zeuzyAjOb
OJePXf98wWDtfEkybP5L0tx/bGMHO6i8fg9M4hk5UAPoljN7cDOx0r5+bx0JOjYx
fEcjVTqQLJLOjJrBm+aK2Jk30xzz7r0ZPHqZsliawphT2r3HSExsVyL0ftRwRTDF
2WxrfZwfv9Mn7Sw64yrectCv6gLClcoGnnMRTl8Qoa1YgTEwwk/m+AiG2WGQV/us
J8RTy5de3gbdSjEjfAGrglPN38MU7kY1N3aJ2a8cQMqZoa7u0GeWdu4ESEb7STr2
FfJx29x6SjZgbDSPrrHN2XWZjFKwIto7Px3YR9b3kb0XEKLraJ8hlif7CwwTYS9T
b3SeFbVvSBNE9oLsUbOE5SVfpeGwIqbr3xAq6IBpS0wmwF66/IMfB0rcZox+ipnE
TuL7mL/7D9E6b11XvEdBl9r2wLl1pN0372oQuxPqCm77pTahKo5AhHDnQTGWqkaU
Wi/n3vxmPEQhrG/hyWwOabokwagUwXx7YKyOo8xicvjakSxIPbYADm6Y9xR3N0B1
gXHzQx5RTBfH9lmW1lNKMa37rQbKKZ25dPAgQj1Zuqk/Smnqqo5gw2/f5rdCxbu9
ZObaIMZvCg/6UzLGIME3RwECD1p4N2gBH3gY9hVtBgkPNH+n25PDTwc1smDHNBzs
YaNBI7TOLJyzNEPNe7c/ObwShM2TiV1Gj2osG+sO2Je6KcK2GonFL6IoNtCm6lmq
HvtOHsfm0sqGIDuYhSy+ALaIL9gMFSPNJ0ryWNWEYA1o8AN9XIyE+G/z5jKVk67w
CtcpjuUBkXPmepYNpUR2+33TMr6pNkXe8Z/u9lbZvus1mxY0GBDat29COcCrUDZD
3c1q1T71IaJp7JFVf/hAU7OZA9f2ceHiaXL2PVP7e/O0hGiBTFei6HHlssdrNETW
02w/yox5Dk3r656EE8DTqGVp8C8uDhLq6byIaQRlsz3r7ErmhFfdeLWE4diqeiKy
vp8BeARyPFV2avoNm/vtE8/WpOGPJUWDcnw+pPMsGXKhpXMX5NyuxqkDofXmMqZh
A3J5TpKONS5Q0AoQEwXo5ukPKbdvLTLFr+LFaLnucvlPjbYvol3syjwe+BLbzVe1
7XU/Tszs/rOGF8FfRXZlDqxPXEivXoz4UQ22QU2hzQaWdCUqKIBLaLMhBtuR9y2z
tsJufabERNp41xXRRa8e1kc5OvIdE9ZqhU2tOZxoNKAswODkHB8nuCiuiWKzcYqa
IlNHgYTqZkaQ9RHGML2ENFE/gFCBQfMB2sccJ8vldIrGbdZSmyKffVOYnqiTq5pa
erQOAqsAopJrq/E8vpm68gArLgQW1Cm9squvTeRk9hzyAVxTmOBAmo/O/469KRGK
Ma0MBSd8uPpUSUNd/G7r9R4RAGO6qRpfPDi5IQ3DmJ0FC0dWZioMQoAFn772l1u6
mIqu0taEV4b62OALVxC8ecfl54TxuGTlw+VgwDRL6xnPV9BaJK/RzbuH8Tm0s2IE
7DGD9b++Kap6pOXIwcGO1tx0yffLQPSsCNKxh/cmNMVuhumvpwX66mJskCHcXhTj
Sa9bajnxZBXipl+nqH+fsPhhgXEPigFJysXC0x6gxauhI8p9/A9G4CAuG01aQ3DF
FZ2r/rCOtidufZJDMsodoJcYgA5OYxYqjueX/0kxm5iyKkFgWgnRsldelNyRZnX6
Pq1kmaPIu4CvmscAnx0BzvrjUnC01ficyJToP5jv/QJZr0fTbzb1IPpfgnEhp534
rKTCBtgQI8EjmGShIUgg+B2uLBiTBVKQh3h28OtiQaxRs36o5g1i+ECpawVKOHpr
kwMQkBEo62SsYnn4Mnm01OJt7Gs3gvtUTXhvRpGywj9DOR2iMvDu3V7Jso1eOYqd
SqYFjfSXmtcXg6F8sZFS7v46Mcd8l9H8foYEWwz6WFzlFfdgIZP/okwux07rn341
VO2eVJJ1YuHuXlHdr6zHVPKJqo2zKq54I70XEv0MyYaEN1CtC5o0pKJar0Cr5VSu
0ExgiWTU304ilXI0JdfCLGMEOEh2UxuDut9dBm6Y7h4Gek5qvJ0swZVzU+ckdy65
aPYSjyul3IbgesHvknGaYrGwG4ahNa2tUTa4VAOb8A9J/gdi9l7p4N77skfFZHoP
ln3YT6oqAKrfYKENxyMWRit24nh5Vt2OcNLJIrj5HXEppdEd+A4u7wUOLyPZ4bO0
e2DaMydXPcu/hZkwuyv2NeIt5F+79yaR6kRFBdW7BnASDocIle6csI5UxIMUn1FF
JnzltgWvC14iEQY8nuZzDOaFakRg9K9VKig+xJoP8AXI5gtmKhSAJwjjLaDH1v0C
dXnh/slQSYrOc0xQU2d+5xqHVGSpOKLl8baKvHhLE39NCPPkE30Zlxfhk9qkpvN3
1LAe1TJnhrWU887YK1uoVbGaZI/lBv489a0ZER6GG287uGA9Th8c/C9IXyaRrXGg
S7Ie8YR0LipEdMZotL2xqQxB+NCBFgR6b1DH/fXT8BEDiKr5dMil9HaptKYuNDis
qyI5tk1YJUrLWtyGY4uaMNo96ob3HElUGL9PeRiGWnLtuQKgf/CgeBaUgUugWGUP
SND2CmbL2zRBsT8SHl/SD8/8GJxIYwQPZEEboayawHKo1JUmp71ElWCzlXSbdyug
xMIQtjMuRj0r+SNsa8MbTRg7sdGkxd1vlA9CYaGjscybzD5XRxX6vVJ8Enf8nHPH
iZqEFdCcXHiB+zx94fGStZNdE4gVu5kLtDPBw0gv8yS0Cr2ljTPohlL4qAYCfnSJ
+nJhU+D8/krVGih8urwP/VasiDvqPSrItfapxirlDNKi8zx5aZxJ/DpA1LLYgakt
AZbEXHvMVQ6Ix5hFrlA0MhAKX3Db/i9qy6+4BqugHATFh3cr20EEpHYKq3/yAjlG
QPHMi9LsBnuNVSSSZWA8Kc/b6pewOpUa86szbgaWl2WLz1Z+G4udedYJRCzkk0FG
mnRyi9Ih7KsR6U2Zew1vHYG3t2tIOHn4cxHlL3N2y6LfTpCslnA7lcZdjliuVU/H
6ExKlCskadUwJwn7f85UTsDX/j8Mm72U+qbNbr/IDWvJBgk2nMCUr0HlojDLW/ge
wwr4/AlbvO5ex2d2laUL/q2QajaYUeaV+WLJZJLRLeMMUDQ0QIO/48/RBOeP/jjC
+TEr3cexXELKIptMT/XOdmc6rOYAm3ChwQEzaVi6xL1PVt8KWG/s8jLDolkMijuA
HSzsLo65CUuERLsW68RbULaJcdh+hi5uc44pVHsd5vfWDdnmFxIJARNko39lvFPF
LwIVmBbGVb5L5JAeMr7hQBLpsMxUp922nXhgr0CiFy0nMvaNmdBFdQNJPTmr46lo
eqOZNiPoGPtgg74mDTkdHVg142+pDAJbdn4hg4BLhIuZu7LeIvzMHcEgAKcfpMVS
PcQfTF7PffxGkNjvVY3z2ztUh8wPAJFe2wCsyCkhgkg1nLtQKI5soxDDj56LzkgO
Tv2DFaC0zB4keWmCwlIiyMrs3RI6o8LAt+LxlQ4vr6t2NuUhPvY+4Thc4kwK8DS+
syCgQ3h5o8X5x+lNyQ0da+RgoqOJe5YtworeJIA1f1s3weTmkyC0C+NBzARZaHlf
Wd25/UmpBDmb7c1KtjPVa4exjZxmTY7ua3HlRh0CscGkboMg3rm2QTpRv813bExB
a6WACK1FvjAYxLN3lsuxZLGKUQiaTm5iylf/DqJ0zNvhS1Q/+Zo4hRAUjpKo01pE
A5hL0X2y41bgaHj9a1KD9zPgxnYdZqLKbOEjL2Cq0ZE/XNJszxPMWXnkb7Ze0+ib
X3q7GpxZYAM2wlWDG73H4UlMyMF+uGb3sk3oDkeN9IPFmHM7dEBm0Dju+dfVKPZV
BkP3QwZM1LXiSPXoavhdeQsx9/Yh4yuauthoXy3Eek+s2IeeGxtqymrVoGV2x1YO
iJsO29z7Vt8NM//fGwhIzJvCsYoH1sV5zmgx/cibauH6fqk5oUdz6Oy2lg3Y9UYp
Pc1aO0rA0DsFltqGk5NKVravezwYz8cBTchffMh4qH9SJJT5g/YtSN9l1bTkbn3e
HoyvTOat8Ha34u7JZfbOXMl/epEhk0fUoyIFR30I39KtOvDOd0wD81rs8nxFVYlk
GqxSmJrumvO+PqOQzgU/YThyfcaeAK6wJQ0psjNa+Bi18tL+mlbvqQjIgY93tTM2
HiNoNGyNDwA/wQo/383YoJHJkLDsvGZL65oh/bT1q1v7X1Y3XiMegOd2wdvXmV75
Fhgz06+UBEvapQt/TukAVlJoBVXuuJTRMjKSH63zHB7fSxOlcEBzYgTcnxfY0Tu9
GM4tuWoicU6oNt9IrLWOpSxSS0sCeG2WKddAzekrRP0fDVk/Bl3oL+JSFZTbuUzn
8Ft610kr5y/xX1EQA4ilwASzRwOx3ddapU+piVe7RPxT1YlDM3Gizq84JJ3ZQhPo
TxH4WTVwcBD6O1r+xiCoFOdPXfx4xHxX/HvjYZHygGisolpmHkSL5m9Gniy5Vgt7
wPyhd8O5IY22L5atNtsjeTrTaJYxDjwv/nNyGhk5qkEuLEvkYEg6ACoFhXduab6D
3UjwMOog+/RBue89OdpuoAlzU3fHXYaNwfRITMCfiRlxQBEBb5r5ZZzPBlF2jEYq
byO99VUqkMmb6kpID5/KmiNCA1BjuKdf+HORA/pkYS+SdMSqM2rYgc0Z07p4D5wm
zB9bDnNTjRKp5Kb8xHTpiNx9mmhQAxOAlQMWofwM7GnzoqyMrQq3gQ/GsSx5H0gt
nhEUA0amuk7aXMi9Ylw6ZTbmLINLT3KmJINseSBRuP90vj7aJ9UZC78NUd5c9qf+
CX3x3yQLfuREpPDAe1T22Er3t+dNhqBjJnSDr6G1BYtoGFrm8PmnGHobLmT98gN4
wjC7M+3Dh7OnARxxuZQuPEDKjj4EeE2/bK5A27/oLo347Y/nKeATVqYpHbrmrF7M
hH7VJSsFO8jhlD7Yc0wDrzPvdD008JjcAztbJEXpBuuo7A5RxqPPWsbUHh3cesOk
7FJM7vFCQErGAnLwkDntdfW27TKGF2At414voHRZCHeBNuNeNw1w5tlJRdQvtL73
9AR6PqkdoHkxEA54jrDfed6NrdeT1+m/Tldrgtht+JywpSvw2sNKrgGl/buPm9Bk
3qJGiEgeeimGfoQ7BmfqoAx/V5MJEJAce4fazc3TIZp/JWaAkoQ/SR8F6x8W2g9Y
kA1XiMfh48CHTtkTtb5bgGPPwSx95ShNJdKVS6p4UxF67oSZf9SUC7YSC77expmr
R1N/HWK+FD09V2jBYNpD4WgzSfb3Km5eJjjLbeolNlS57zC82Uye+mCNJjByWyTv
vVEkNjoCbkNIPpB83hQChLM60FjCeDsL0Ivgi8vZ1Yz/ALVr9yWWWm0zH0UaDToB
eFDEXIq5WDh7K8ZOEX0rewkC5ZlLdoGGQV04uMzuXfLzfi66gngXv2jUT9k+6pE3
jHcGc7ouVpLDW4QmwVop72kjfext1xJlvnDZ/i3DAl5eIKP/QTcVhKMWRv342RSP
NsHICipBy8LgPqRVE/pm/1qAc1Auab9BZfsENYkSEU9YqzbnMA1FbejBJKFx7XWR
2ypfTASy9NpiCJVXIY+tm1+ltds/gSX93lO67uotp2VqaZQa4v1anPditAtEyCKM
c/3HEWOr628PsaFjjD/neHg2xZLretWfX2gIGVt1cQJOBc365R5DbwlYes+tNV+N
hfAbDyM93zAToQjYXFJUDJcNeKVYR+EYN3pIzhjOot7W0u2uOYFwynKPF3es1lOa
kJGNRqpZ17YGEpO/5gnESknmPm2sx0RdB5z8Km3Pr86l2VG3MzgXqaHLVZoCVZOf
YsN7ZPdpMwkBz59wwb5pfu+R3khg/URZCIrCwTmAAF9aCA/CJX+ixDqW4RlJH/3M
BdDNtJdpDyftBhERHxZJtFk/5vkraFwOfwC43gZM5x+iegQJ/ps9kzoc9p3VjCwc
pf/3Q9HxhYrt7EW+jZ6Cl/7lZAn3SvPmRMUew1+qMGHOJBf/HdEdglIPg8PUS94q
rW3ehOQCx0eOjnEWGwOxs2A5HxApuK++1nBItnMezjg1gygVdnEd2izkMmbWviAG
thJXwRu5Iat4eIcrckijUaSikbl3DcZAFQ20DYit8OptkZDUApmjmXymrbPRM+5V
dhHbSF2Xk4xAVpcheAtfR3ivI9WoSlmtCLhWJ9UnUGKQgEmS3UqwWUPFXEZJGoGx
C5glzhD8INjCFkFG6w/sc/9ON2oMYqLHqkFFIpcvEvN+zVtw8CJuHRlk1Ao0BHQh
WcVyme+t06i2WVn5QZLNnhEIvykQmocbSKJpx7ZIS62t03Tos6PNObh9CyddwM6P
ZeQP7/lj6r61hApiZsAwZw1Efm31a8hN3aVYajCbrHl2eagcHkC2/11HuQlQdGkE
Wqc3mHFw83wHDoq/NXxWxQzwLUn+0F9P+CTkH987kV/SRjIj8xZN+pxXjG9hO3dh
7B5zbC8UG8zDPlwxjDTOdz6EoaDGJnhh+ba43nH6ySXvXNj4f5+11vY2l0OdPRPB
iQN6svUcj/i/DkFr8xn/yV+0fh6qBdACrLw6MjJQzghsqgq1790NCy+zZtRffC1q
Y0UnC5Vqy350DhTmnowe1R6WyBXy9HW0H9i/b8pH7f1aHDt/cHSuKHAmKG69t9ea
hWbp2K1uBMSjYwOU9vMtQ/54mVTabZAUzs/xWxUQ+reVUEAE3egGB4GemcXHqRtl
YYrW1UAcitLtUWnnW/P5hOdWpuATawL/1oEPdvMHWR7yZ020D8fOF2EFv/uPUjcG
utuobKSXv670C9QuzXrwz0Wbh+3ozn0GHiEpDpHc3wmt7bDQaB0PKttn+AcNd0g3
GvFsqO4i+QvUmuzc/7J0RmpR/6lZoaSqZZcgshYubKOUJPY86mVRF6niMoi+5Kvj
dxavkytVbD1F1hqK+61AtsfJUiLimEgN+w4TaDBgu+8=
`pragma protect end_protected
