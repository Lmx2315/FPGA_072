// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:36:44 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ElIOlmKvseS+lTV1hAtLsN0c+ZcCjArDDW77N9P/gwimjSG2j4xOsNf//JkKPFwn
6l6dXNhhbEKxdoQ5mT4gvJqAofVS4c6rakf0Jf3CeXi9uttFr2kTjiRmpvkhpSKD
VqBYx9qz2v4JUP4rcURWsiiXwX3GW5ZcLhEOnk0kDOM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5792)
pWvxmB1QikU7Lyu0kguJSWWsdyiEj7rVppUYNe+P1yrZPlz7xuoy9zm77zFo9orz
7tJm4v4X0GD/skalmu5bZIkGHPlIz1qPs3mw0QTvPYZwn+JoESBDQrJ9t3t4IhJb
1Fl+W5zmnth1qDMXrxC94l7yMvach92BxCJa5APsg6zgMLuOaW5u4WU7ODqsYCcu
y3SQVRx7IrBGHAgwSaShynW4gkcJysTRzfytcDxFAc0IiI9vJqMIJvDAWMkw1jd4
mgMVYTdHORIsnMU0iNqXPxvG8ugofjp9ISMQ1asct/282Tvp5hfgd3NAzkjXUigE
MmvKhh+9NMMdel0qsFPDh9VPXvtl87+APgTUkp3OjdeKsZYPqVxz2AP6KNl5+c/R
3hxSdNsSIq/QFpUlJyctffPIFbvf/MAFyy6WkAV2A4rWLVd9gzRdxxBTK/H6ODNO
kdvmPkp/jAXIHNlXMaF/CE3hs/CK+4BwLKd4SshAkY0O72WaIxdZGkT+aO4c123d
YpYVRQPMV7Lq8pNuycoTgY2sNkLDQThkyzEQPudhh2N5BT6t7mDYVPFy0i0DFH9p
jpS8NSR0Y/3RHKaIPzJ/AM1ys5BUk9p6mlQL1CXjD5IVFaHHSMCKidNrKGbyErsG
PKVdf8ucyun6m1tczBBZEBvstPuySt51+X5xbWKsQE/bLHTZX/v7JXzf1SRmwCpz
7/OjOBnhI/3YxOMr09+ZKYtW5cSEoBemN+4sWkDai7VI50E20BswWDrw6//kLepP
t6CBeG1y0tXjzOAmfYUi16geQpy1hY//jXBvX3FL6HRTl0SfSnM9SUBpmTEfEXIG
7AxF8AbjvDPsVlF+LCvDhx+ZmcJewg3NI834cPSkWnlbZhzkNEiw5/K6hKknBBGS
SGxEl9jb/c1EZsmLc1ldxUc2ULrXlUPDq3GRH6qF0AHjrmrhZg8axTp1IkkqxI3s
MEmXFmYTl5aQwaSJKDZGiWyd6AahP29N/PJuu7zqa6PQvhjTb/NWGfHEySMeUAQW
Dj6Gmc45/q2jKIlmS3iFZy/XXrKN4/gMVlSLWGIlJQ56bmO7sBU2FN+N0xecUfG7
ibjFEkuhQlw1vrVJORBMbil9QS3rdlNpKIJENATsm90cvWUsgtGatEfxcILzSjLd
sjnrPx9pfkIwFn8LkN/mM6+e1PUrO58Yjgi+gsHIxxfuXL1SpfR7qL22Om2HNDV6
FWMivHlDHTZFBs0bZFpxX+5P06FtnUNUiwHl60kuQfj633/eQ18OmWo5oLoeO1OB
l8SLvpKksa+fUmnWS4a2/ZaBJCp+GJq8N6TrI1TLIrE3WAnIfs898GaTuKXeiupT
BjSGapD3djCE3LkbZKIRGkF3fYMwm4RocwRqWfBm1ZjPc59OHUkMjY+KVY5OIErI
dnzhdPVfRfl6yFNb+YWpECuYP0f98j5u/bjv1DjeNiJYMq/cp40XgLRcvVGSwDJ3
a0+y/17aW6kE+3j15tpKOjO1oduNzieZ8Tw2kK4248c+MKdGKEqxjD3CpaoudB6h
UUs8Sqx4MRyeWi09/9tRsJt6wPm2Rpyuh3qRTYQDc+HSZrKWuBCY4H+nQpnf/uHi
ZXfRWzRVwO5vdLeJypxgqK3ixe36B3N/9LOA/c8Ievx/QBi8SDfPbBvT494gRuue
hemaAa17l9hZCVZ1YDC8Imhbpt3Y0TVO04aipafcqxOyADi1hVoswIU+9sWmKBGd
cC5IAFXCB9RdPfZ8CSdUnI0rGWHK2FI9alnAStNLuBEeWhVL2/ODH7+t6m0HQW4d
mGT4OLOfmwIPieeEinFHxq2ISmkBBY4QHGsNCQ6AU7UDny2sXYXDUXQpswJxqS5a
vUMcOgWITrwaqiBpnTiYMbFg7x9H3tIVXAnGqWPa8v0xbLCRyhZiUKlCKbr5rbFx
5yTPEJzLHEKI2UYv+gQ7G0DupxgobCZ5/lbmW+Yrb6L6n1E/TGDtgul7PAMCw31l
xvLMKz3SobUriwkXtRCofeHL9kQ00Ems0DC1h80MQhHwi36FBHYx3oVsiCMD+CL2
iq2eLkd/FHZaxA2Tq+CNg71qeTdz8dpGBakQePP2ogG+OKRVUyHB7nDYfOIh4oOI
3uQyLm4ZYer37xtf9KOhqWgA85j/pcBR2ZSlDGCZ+C8ygq17clvlDWdZuKHiOO58
vZDZ8oOn/qFoTFxplNhMEHVZIQTP17ICgvxJNomgg51wetaXMT2NsGQOOUd5Ssw7
rxhamDuOEmNB9I+5h9mvcxisr+rwLSSpYQS4C+Pre/dKn/PJ+bDrS1erBDq/I5iW
LJv6fEEoakvFLbSgKBKZwBsaaX1eSYvDKmXnPiBcl297TOk0GEwdwAfdZ8UUx34d
hvrMqZsYpKdFYuwIDMMKqxQ/pKTu+mFDbgoU4pj+DOOVtofUm7HXaImdVaBN/Ko6
WToSk/SpyPaE1laLygL/jr8MW906RTZOxzFKm75agmn1x+7nOD6AkN98qGvRCcf6
noNJuXIjsIABhFhnTTIfTAl/C1G61Jdc8mzXTwES3+qdOGZ8p58LD2XMFrQ2i2XW
Rz3dAz1wFby7a5dYcs+ToxekiuebbgplOBMUMXELCAUHpUInzliXjiHNA7z9EpvK
8WDqTYehlbpi8bIH0gltekXQiPvu1R/lObidZ6HG3ggHEFMBAtarabeR4i0gPh7i
tdCsvjBhgY1MJ5q0zXO8DmgP6PA3Gp6JdW7c3t3PQbtlOknYufx0kFyTMjT35US5
lbMA/LVi1Mu6ih8TF4lnGC9d1pW4MUJ/Apy3iYuUDgIbhNCh3PX4VGWB0NzDVBay
u9vjVFJ94dS6BbD/EGWBfmT9AVsFBaTD9X3oAymsUWyrX5Cj69FvQz/Ssv20Yb1h
PgvwmnKxxfYzcDHf0rTzje+9vfF+FdhbMXHMb6lZ1Yf1f++0fLbMnd9A4PSkvCS5
UBdXY+vS3/tAbRNHZmLPcTj6xn5iC3gZHUttGqnPlT9a1CzX8vfbt2e7fD/REFTk
fIqdsv+0GbslzlyiSDHECc3vkTCF7kY6z+8Gg3eCtykkKwfsgISZ80EBwppmXgbL
ypG6rbgjMk5mQAk0O8BUytbZvNFuQ9zgT8Yy9xcVU+OCBBxSnwLRVRcLq+nCF/gJ
hkks+4tjmtKdu1mj0DrOvtkP0Xn9LC1FhpyBZERCrFAt2R8KMipv3GvIpun7fa+p
J4TqMDLEEILWHfNS9pqV24KX/ZG/1XkrF/zVpNmHO8R+qqowPi7tGIOskVzWVFT2
yY14SzHZ8JpqlonD5HRJJ+FM9+yOzCMnxVoGnAePUUGDk4YymnJJV+CJu5/MUFJg
Cb8g5zSh4uMrMyPvmhGwLcLCusC6Sa7FnjucWarKxyrd1QLd7FG7ZX3xX+/It3K3
9OD2FgZE502L2Zyz/x9rdj4tG+HStwXZHnmvOEnM0jKafYw5T8Gn8hL+lfazVZao
0Kxq7740/KrEDSFcUEPw93KeIqeeZNprvFaX46kp0/FQCSYaLd74k9bC9rmdBo89
xGm3pE4Bf9fhM7JMtHoEY88B6SHfaq3vxfeLE/utlHaWG80hKohaUNDRe04cV5Ph
t8p7R+csWuXV0tkQbcsuaMNOSz3ggSn+MMhmsp1ctsO82aKqQq8K8h2NzOTasTqH
VccAgG9tWJXHNyGO2Bt2mDMfrVNE0lyYPuYfKPr6MmXc2IQUM+FTdVlt+czOEqPC
8Htke3BsSG2cW1+9IEBeEeWQCsPPuLOwyEwEGREnqkc8wh3Rh4zmg+O9+J4N6A4j
nnv2O9czdzAbwV8EW/UdExxnP3NxifNBSBjlKp6fhkVsh2ZlWxpWUYnXK9RZG9iZ
wepyWWL3lDz567UXYVig3RnIcTZSnjYeguhjz+TcjueyJZ40qPmSEB4tWPZdnJKe
Ne15wO9FYzxX/7ZS8z6lqNSjGiPePNxMpwT9A3YMUrrKaLSglTMmgv4sa5yNi0kE
AWlQDB0Evb9VfMSxTbiMmMskpkgxbQ9e1s3ejtsZS4Mm0ZErMd2Pa0pAgc4u2KDi
Iau7E2BM0XCs4hbJnDJVIZB1nNznlxz0CvVEgbBSA6NoMmN4MEmsCtlzXDWd5PBk
CsUKqfflmVMAWNV8enEQ2u/UOgP1/OGJkWQuk15oRqUYya4SA1U1IVCur0krt552
cC9H2y7Q+QswZNHXoBIFdcfkLxvrbVA4Ef0CGShs4kBtUN8pxUnYDRNGxJnbOwwF
2+KKgOuyJG/tEJgck1ACj03UyEGo5wvCp+AuK8qKPjmopwerYhWVieoABuWdcW+7
YedftqcUbB/UyvDXf7Obm1DZkjv7+8PRGHqoLckb3VhkuZI8ViDp8tDNcMFvL4v4
dNWfKkxwXp5PNtoXIHLptaYXoSRgIvatwSeb0MD7pkpG2Vwa1hPD96nGVsHAEJeM
yWkl6M38AUK8UoeSjTOqWagFOhn/qSNdvU1jChPOIIuK4Pm3iXJke5AgN9vD0Sfc
7h2SC4yAaKy1+npSKS62wbwsZc4lrlN6JDc1t1cxh5PrwwzlAEwffT8qxxlZRKyO
q4wY0PvBmFYPGNpBNIh2vokldo3nVM84dnGHngVm9bJ/9sy9FCmG4Nuopcrzx7OX
eFTZfkT5ZlXEojs2xQ4wihVScqcQNfXDV2w0jhFqJxxNsb0l9EAurXRn0quhoH1H
OYdM8frf2YSPmZBB+CzBG2OFUYtCPzb2mGRlouD/RBbe2hFgqVgDX+GdzRkZ8ymu
iZjH9NMzIEBAMiTExpOXz3QSrpKrr56k/pUgMp4V6nRj253A7U0ZDPgjj09zRd2y
67wAJOOfo6xQ/xfPWraDlXFOhUpvD7Kz/60svEVE+zfPvdnWn/+M2ySX1ylZjZAk
80u+yKKiaqy9XnfCRxtPJlaoU6ggnHZhFNxsiGADPgwPWbuo9u3QG3g7y4E7ZqND
XpZaPgsjgv8KFLEK1gTZ/Pkj98wFZFHLr3vjURW+n+PUadKg6IcTTZpkX9WQkaal
LXcVFrGvvFW2o6UY601ISjwUR77+qD1EZx1ebROV7ZmPOhne7dpOGmjLl0mVA45Z
tYQY8QuXMhbF3u9f7HbHUxx5mQuE1pptAMhH0AWEkWGM7a5moK3L3VBBhvLEeCSY
2PPX4jeSN7/kzNlBdtzdC0xkLKDr0QWi00G6TTyT/67QC6znADlf/DZ0XmBQFcC2
RsDXNV8IYEADzYzfu92al8yW3E323nR9D3hWyXmxw0dMuXRly8Q6WGleSSQeHHgq
WXoD/4brgLFKR2N5O4pilNtMIIyfJYr+I1ebROadaEUuyWgk8xKxjsKf8npAXBEg
1ITtGm7IjlxFeyLoeI3xNaetNUhm4sugadyxp5N9c5lnbRlPFEB/Cc3BTH4VWSek
1GM0dx2aId8vAVlaIaxb29zUiw0+UhmwLL2cnGBz+xrBq/xvpdp23aHsqF0L5LGP
MBW4vKPaA8yiTSJnVqT4N3b+RkqOquPVz4ucyacnn3Gv9ZCDJMm/BBWD58PE3RKu
sHaq1L/SWzz0QVe9sTm87vLidjgpuC9KfzbarIXkv34h1Iak5lUNDPjbAK74cux+
UT2xvhk5DQO3+bvxI2IIFrHTrmsBmP6Q3LeH667jV169VBPuB0Qioc+jyON/HR27
8qVMXQPpfAOfaMkKdgZi3JdaU6LKgV94GCvx+IsqGxgfFs1XC0owX47BW8N9a3bT
oq2K48klzVKYIptIri/hTETY41U+xLb8ire3bmwHmDfpsIFPZv9f1soVuuZXmWsG
S5WesVVb+0bD7lbAw2EhqAoOXZm9ec7D/bpeZ145Lzm9h4OjlmxvlkZOIsFhriFe
I2TEAbr5EeqibaPQSJYH0qsI6OITzZWywYF73r+Jn/aPjyylWEZzecTW99egyGBi
UCvTYrbfV1UcA8A2d2lasqGt1Yr7mIrjt6j7HS8oFlSC02s5q6GqZVFwYyB+VCl6
xBcXGPhfICxF4QC2jTnVJd7xa5vjCgCZ9C+DgX3xCEsSMRq7Wz5tXnuEu4uW08LL
SjkanGZhTysWxI5nPPNc+TkzkBkVOtv1Tbtvv5S7nt5jDQnKSNs6h/zD7a17QKcX
KTipwGl9e4j7ATIsjzTJ2kjgCUXSb5rAWl5crKTU3gaWu0HCGTGg+D32hbsurkTE
Bgw7ZlJxk5Slvq2hIK8rVXg/Bp7zYkTSXHTiQER7+yXU8oe6yh9VeWtqMf3w3tB6
rD1dQzAZqeYi50LsqEv73YNcScEDgZxHQ/uHSlLV84jMadOyjBX8eYMpJaAgpWZv
PNCiTneH98Qju4F6NOYCn3Jyf3XCLzDcDl91zcA8UxeCONpdvoI/22UUPaO6glvD
O2mup1/Pg1XPLIcf/HHFtK2EG1o/cs4SWnspczt1TtksPbKtRzOFzN6ngE2n/f6p
S9JCfkcfYRAJBN6Jr/DFb9qfB49a0TgLcfXt5nf1thkHchIkgTvewq6xgW9IEInq
50FGygqF/qP7k49ZuTIefOYgAP6DPzWRPlBbASRA/AQcUgdDOzHwbfBzOKul48Ha
sqVz/K1NvX1d6KdmuppdNMbtvsQh0bPxn/L1QfrH2nQMj7O3SawnASnJqnoHW6bo
uJ8gmYM3VfjHWJWsliC4J1s07j0tc2CYag0rCDkWzPzMllvKfNdSRI1gHKz4LMlA
0Ai9eAGorN/Zbjoo7934EQTaQMZGckzz1XHLL7zKGaZ3k8rJ9qsHBu9XxNg/jrog
dfPG+UhMHO8v4Wcs2twE84nmnSrp4bJc0uB62ReshBiA138Lqf2Eq7AW+E58u8B3
8/2h6ibVhdAy7GECfs0Rcigv0b1iq2px481J//i2JG9tDC8Pmx3Tw52g1HUPmdF+
ArqNI3J6dE43rTIprtd6bJOlKjxf2b9WTz6IgUGA1DLL7yGVL7iz6ZkDKuMTP3+s
Bw8G+28DK5J1a8r/3vlT4TRqkbLvIWXMRQ1/zghmNgmtCcMmuTDq+CWc8xtaulCM
Y0be5RVt6RugksM4AiEbKsN3imy0lY1qdirGzH49UXlzoHQI7l4NHDrLAQApGvlu
N7lSf+TQBDT5KhjJjGeAZU4IRFBFPDnLtmICzmiBDmNLXM/pMuWQQM1qEJifqAFM
NqwbTOlBmVIxPgPFxC5htNIxR9WoiNMZqIE1+nvl+uRm7eUwTET8HCUsDgPkgok4
F4bn0jPHvsQnj0psIcDms3IxCLMWlgxNI1R0yTW4W6AU14jjeUhUDn0q4Xbge36i
jtZBiFdQiQepGbzNRPej4XDI2MLUvhnz2I7XK9Wr3HZuu4c833g+DPyuExH2ylVy
ClayyJ6+o4WmUygfNKfP8Mv4GKSyAA6YLPygPfDJHyz4+VUooKLH3Sf56IwOQ20M
vOAQfvisfDiTLJkxes6veRB6DKuCxW3/HKjstxMUCPEETK9P0Ow6VgPdIHo46cmH
GlmKcM327guniNvR4ZxIXSkvQCoGDNtVdduM1uEBmh9MGGeIYrImxH/qVb5R1TDy
eZu7bWutAS8/+10bcVPyt4QZvqLcBD0C97OUj9OO5o8Y+uT3976R1Mg54rjX+lGI
f42gETveI0xILizWuRhmTJZOtZX3wyCR/mE4RBnnTBzar4meepJvVTuGj2fK02nC
j1vf5Vzz42zM2AGsESYTJRG7vwgIWecCjqNHNOaYmuT9EMSbWr24wG4dbrpL2E5y
QGVGbhp9NOfSKCEoCVsJ2kGWbr6iM1yCZ5tJheVq8Zg=
`pragma protect end_protected
