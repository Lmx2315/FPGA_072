// Copyright (C) 2018  Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License 
// Subscription Agreement, the Intel Quartus Prime License Agreement,
// the Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is for
// the sole purpose of programming logic devices manufactured by
// Intel and sold by Intel or its authorized distributors.  Please
// refer to the applicable agreement for further details.

// VENDOR "Altera"
// PROGRAM "Quartus Prime"
// VERSION "Version 18.1.0 Build 625 09/12/2018 SJ Standard Edition"

// DATE "04/30/2020 13:56:40"

// 
// Device: Altera 5AGXMA7G4F31C4 Package FBGA896
// 

// 
// This greybox netlist file is for third party Synthesis Tools
// for timing and resource estimation only.
// 


module DDS_48_v1 (
	clk,
	clken,
	phi_inc_i,
	freq_mod_i,
	phase_mod_i,
	fsin_o,
	fcos_o,
	out_valid,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	clk;
input 	clken;
input 	[47:0] phi_inc_i;
input 	[31:0] freq_mod_i;
input 	[15:0] phase_mod_i;
output 	[15:0] fsin_o;
output 	[15:0] fcos_o;
output 	out_valid;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \nco_ii_0|ux122|data_out[0]~q ;
wire \nco_ii_0|ux122|data_out[1]~q ;
wire \nco_ii_0|ux122|data_out[2]~q ;
wire \nco_ii_0|ux122|data_out[3]~q ;
wire \nco_ii_0|ux122|data_out[4]~q ;
wire \nco_ii_0|ux122|data_out[5]~q ;
wire \nco_ii_0|ux122|data_out[6]~q ;
wire \nco_ii_0|ux122|data_out[7]~q ;
wire \nco_ii_0|ux122|data_out[8]~q ;
wire \nco_ii_0|ux122|data_out[9]~q ;
wire \nco_ii_0|ux122|data_out[10]~q ;
wire \nco_ii_0|ux122|data_out[11]~q ;
wire \nco_ii_0|ux122|data_out[12]~q ;
wire \nco_ii_0|ux122|data_out[13]~q ;
wire \nco_ii_0|ux122|data_out[14]~q ;
wire \nco_ii_0|ux122|data_out[15]~q ;
wire \nco_ii_0|ux123|data_out[0]~q ;
wire \nco_ii_0|ux123|data_out[1]~q ;
wire \nco_ii_0|ux123|data_out[2]~q ;
wire \nco_ii_0|ux123|data_out[3]~q ;
wire \nco_ii_0|ux123|data_out[4]~q ;
wire \nco_ii_0|ux123|data_out[5]~q ;
wire \nco_ii_0|ux123|data_out[6]~q ;
wire \nco_ii_0|ux123|data_out[7]~q ;
wire \nco_ii_0|ux123|data_out[8]~q ;
wire \nco_ii_0|ux123|data_out[9]~q ;
wire \nco_ii_0|ux123|data_out[10]~q ;
wire \nco_ii_0|ux123|data_out[11]~q ;
wire \nco_ii_0|ux123|data_out[12]~q ;
wire \nco_ii_0|ux123|data_out[13]~q ;
wire \nco_ii_0|ux123|data_out[14]~q ;
wire \nco_ii_0|ux123|data_out[15]~q ;
wire \nco_ii_0|ux710isdr|data_ready~q ;
wire \clk~input_o ;
wire \reset_n~input_o ;
wire \clken~input_o ;
wire \phase_mod_i[0]~input_o ;
wire \phase_mod_i[1]~input_o ;
wire \phase_mod_i[2]~input_o ;
wire \phase_mod_i[3]~input_o ;
wire \phase_mod_i[4]~input_o ;
wire \phase_mod_i[5]~input_o ;
wire \phase_mod_i[6]~input_o ;
wire \phase_mod_i[7]~input_o ;
wire \phase_mod_i[8]~input_o ;
wire \phase_mod_i[9]~input_o ;
wire \phase_mod_i[10]~input_o ;
wire \phase_mod_i[11]~input_o ;
wire \phase_mod_i[12]~input_o ;
wire \phase_mod_i[15]~input_o ;
wire \phase_mod_i[13]~input_o ;
wire \phase_mod_i[14]~input_o ;
wire \freq_mod_i[31]~input_o ;
wire \phi_inc_i[32]~input_o ;
wire \phi_inc_i[33]~input_o ;
wire \phi_inc_i[34]~input_o ;
wire \phi_inc_i[35]~input_o ;
wire \phi_inc_i[36]~input_o ;
wire \phi_inc_i[37]~input_o ;
wire \phi_inc_i[38]~input_o ;
wire \phi_inc_i[39]~input_o ;
wire \phi_inc_i[40]~input_o ;
wire \phi_inc_i[41]~input_o ;
wire \phi_inc_i[42]~input_o ;
wire \phi_inc_i[43]~input_o ;
wire \phi_inc_i[44]~input_o ;
wire \phi_inc_i[47]~input_o ;
wire \phi_inc_i[31]~input_o ;
wire \phi_inc_i[45]~input_o ;
wire \phi_inc_i[46]~input_o ;
wire \freq_mod_i[30]~input_o ;
wire \phi_inc_i[30]~input_o ;
wire \freq_mod_i[29]~input_o ;
wire \phi_inc_i[29]~input_o ;
wire \freq_mod_i[28]~input_o ;
wire \phi_inc_i[28]~input_o ;
wire \freq_mod_i[27]~input_o ;
wire \phi_inc_i[27]~input_o ;
wire \freq_mod_i[26]~input_o ;
wire \phi_inc_i[26]~input_o ;
wire \freq_mod_i[25]~input_o ;
wire \phi_inc_i[25]~input_o ;
wire \freq_mod_i[24]~input_o ;
wire \phi_inc_i[24]~input_o ;
wire \freq_mod_i[23]~input_o ;
wire \phi_inc_i[23]~input_o ;
wire \freq_mod_i[22]~input_o ;
wire \phi_inc_i[22]~input_o ;
wire \freq_mod_i[21]~input_o ;
wire \phi_inc_i[21]~input_o ;
wire \freq_mod_i[20]~input_o ;
wire \phi_inc_i[20]~input_o ;
wire \freq_mod_i[19]~input_o ;
wire \phi_inc_i[19]~input_o ;
wire \freq_mod_i[18]~input_o ;
wire \phi_inc_i[18]~input_o ;
wire \freq_mod_i[17]~input_o ;
wire \phi_inc_i[17]~input_o ;
wire \freq_mod_i[16]~input_o ;
wire \phi_inc_i[16]~input_o ;
wire \freq_mod_i[15]~input_o ;
wire \phi_inc_i[15]~input_o ;
wire \freq_mod_i[14]~input_o ;
wire \phi_inc_i[14]~input_o ;
wire \freq_mod_i[13]~input_o ;
wire \phi_inc_i[13]~input_o ;
wire \freq_mod_i[12]~input_o ;
wire \phi_inc_i[12]~input_o ;
wire \freq_mod_i[11]~input_o ;
wire \phi_inc_i[11]~input_o ;
wire \freq_mod_i[10]~input_o ;
wire \phi_inc_i[10]~input_o ;
wire \freq_mod_i[9]~input_o ;
wire \phi_inc_i[9]~input_o ;
wire \freq_mod_i[8]~input_o ;
wire \phi_inc_i[8]~input_o ;
wire \freq_mod_i[7]~input_o ;
wire \phi_inc_i[7]~input_o ;
wire \freq_mod_i[6]~input_o ;
wire \phi_inc_i[6]~input_o ;
wire \freq_mod_i[5]~input_o ;
wire \phi_inc_i[5]~input_o ;
wire \freq_mod_i[4]~input_o ;
wire \phi_inc_i[4]~input_o ;
wire \freq_mod_i[3]~input_o ;
wire \phi_inc_i[3]~input_o ;
wire \freq_mod_i[2]~input_o ;
wire \phi_inc_i[2]~input_o ;
wire \freq_mod_i[1]~input_o ;
wire \phi_inc_i[1]~input_o ;
wire \freq_mod_i[0]~input_o ;
wire \phi_inc_i[0]~input_o ;


DDS_48_v1_DDS_48_v1_nco_ii_0 nco_ii_0(
	.data_out_0(\nco_ii_0|ux122|data_out[0]~q ),
	.data_out_1(\nco_ii_0|ux122|data_out[1]~q ),
	.data_out_2(\nco_ii_0|ux122|data_out[2]~q ),
	.data_out_3(\nco_ii_0|ux122|data_out[3]~q ),
	.data_out_4(\nco_ii_0|ux122|data_out[4]~q ),
	.data_out_5(\nco_ii_0|ux122|data_out[5]~q ),
	.data_out_6(\nco_ii_0|ux122|data_out[6]~q ),
	.data_out_7(\nco_ii_0|ux122|data_out[7]~q ),
	.data_out_8(\nco_ii_0|ux122|data_out[8]~q ),
	.data_out_9(\nco_ii_0|ux122|data_out[9]~q ),
	.data_out_10(\nco_ii_0|ux122|data_out[10]~q ),
	.data_out_11(\nco_ii_0|ux122|data_out[11]~q ),
	.data_out_12(\nco_ii_0|ux122|data_out[12]~q ),
	.data_out_13(\nco_ii_0|ux122|data_out[13]~q ),
	.data_out_14(\nco_ii_0|ux122|data_out[14]~q ),
	.data_out_15(\nco_ii_0|ux122|data_out[15]~q ),
	.data_out_01(\nco_ii_0|ux123|data_out[0]~q ),
	.data_out_16(\nco_ii_0|ux123|data_out[1]~q ),
	.data_out_21(\nco_ii_0|ux123|data_out[2]~q ),
	.data_out_31(\nco_ii_0|ux123|data_out[3]~q ),
	.data_out_41(\nco_ii_0|ux123|data_out[4]~q ),
	.data_out_51(\nco_ii_0|ux123|data_out[5]~q ),
	.data_out_61(\nco_ii_0|ux123|data_out[6]~q ),
	.data_out_71(\nco_ii_0|ux123|data_out[7]~q ),
	.data_out_81(\nco_ii_0|ux123|data_out[8]~q ),
	.data_out_91(\nco_ii_0|ux123|data_out[9]~q ),
	.data_out_101(\nco_ii_0|ux123|data_out[10]~q ),
	.data_out_111(\nco_ii_0|ux123|data_out[11]~q ),
	.data_out_121(\nco_ii_0|ux123|data_out[12]~q ),
	.data_out_131(\nco_ii_0|ux123|data_out[13]~q ),
	.data_out_141(\nco_ii_0|ux123|data_out[14]~q ),
	.data_out_151(\nco_ii_0|ux123|data_out[15]~q ),
	.data_ready(\nco_ii_0|ux710isdr|data_ready~q ),
	.clk(\clk~input_o ),
	.reset_n(\reset_n~input_o ),
	.clken(\clken~input_o ),
	.phase_mod_i_0(\phase_mod_i[0]~input_o ),
	.phase_mod_i_1(\phase_mod_i[1]~input_o ),
	.phase_mod_i_2(\phase_mod_i[2]~input_o ),
	.phase_mod_i_3(\phase_mod_i[3]~input_o ),
	.phase_mod_i_4(\phase_mod_i[4]~input_o ),
	.phase_mod_i_5(\phase_mod_i[5]~input_o ),
	.phase_mod_i_6(\phase_mod_i[6]~input_o ),
	.phase_mod_i_7(\phase_mod_i[7]~input_o ),
	.phase_mod_i_8(\phase_mod_i[8]~input_o ),
	.phase_mod_i_9(\phase_mod_i[9]~input_o ),
	.phase_mod_i_10(\phase_mod_i[10]~input_o ),
	.phase_mod_i_11(\phase_mod_i[11]~input_o ),
	.phase_mod_i_12(\phase_mod_i[12]~input_o ),
	.phase_mod_i_15(\phase_mod_i[15]~input_o ),
	.phase_mod_i_13(\phase_mod_i[13]~input_o ),
	.phase_mod_i_14(\phase_mod_i[14]~input_o ),
	.freq_mod_i_31(\freq_mod_i[31]~input_o ),
	.phi_inc_i_32(\phi_inc_i[32]~input_o ),
	.phi_inc_i_33(\phi_inc_i[33]~input_o ),
	.phi_inc_i_34(\phi_inc_i[34]~input_o ),
	.phi_inc_i_35(\phi_inc_i[35]~input_o ),
	.phi_inc_i_36(\phi_inc_i[36]~input_o ),
	.phi_inc_i_37(\phi_inc_i[37]~input_o ),
	.phi_inc_i_38(\phi_inc_i[38]~input_o ),
	.phi_inc_i_39(\phi_inc_i[39]~input_o ),
	.phi_inc_i_40(\phi_inc_i[40]~input_o ),
	.phi_inc_i_41(\phi_inc_i[41]~input_o ),
	.phi_inc_i_42(\phi_inc_i[42]~input_o ),
	.phi_inc_i_43(\phi_inc_i[43]~input_o ),
	.phi_inc_i_44(\phi_inc_i[44]~input_o ),
	.phi_inc_i_47(\phi_inc_i[47]~input_o ),
	.phi_inc_i_31(\phi_inc_i[31]~input_o ),
	.phi_inc_i_45(\phi_inc_i[45]~input_o ),
	.phi_inc_i_46(\phi_inc_i[46]~input_o ),
	.freq_mod_i_30(\freq_mod_i[30]~input_o ),
	.phi_inc_i_30(\phi_inc_i[30]~input_o ),
	.freq_mod_i_29(\freq_mod_i[29]~input_o ),
	.phi_inc_i_29(\phi_inc_i[29]~input_o ),
	.freq_mod_i_28(\freq_mod_i[28]~input_o ),
	.phi_inc_i_28(\phi_inc_i[28]~input_o ),
	.freq_mod_i_27(\freq_mod_i[27]~input_o ),
	.phi_inc_i_27(\phi_inc_i[27]~input_o ),
	.freq_mod_i_26(\freq_mod_i[26]~input_o ),
	.phi_inc_i_26(\phi_inc_i[26]~input_o ),
	.freq_mod_i_25(\freq_mod_i[25]~input_o ),
	.phi_inc_i_25(\phi_inc_i[25]~input_o ),
	.freq_mod_i_24(\freq_mod_i[24]~input_o ),
	.phi_inc_i_24(\phi_inc_i[24]~input_o ),
	.freq_mod_i_23(\freq_mod_i[23]~input_o ),
	.phi_inc_i_23(\phi_inc_i[23]~input_o ),
	.freq_mod_i_22(\freq_mod_i[22]~input_o ),
	.phi_inc_i_22(\phi_inc_i[22]~input_o ),
	.freq_mod_i_21(\freq_mod_i[21]~input_o ),
	.phi_inc_i_21(\phi_inc_i[21]~input_o ),
	.freq_mod_i_20(\freq_mod_i[20]~input_o ),
	.phi_inc_i_20(\phi_inc_i[20]~input_o ),
	.freq_mod_i_19(\freq_mod_i[19]~input_o ),
	.phi_inc_i_19(\phi_inc_i[19]~input_o ),
	.freq_mod_i_18(\freq_mod_i[18]~input_o ),
	.phi_inc_i_18(\phi_inc_i[18]~input_o ),
	.freq_mod_i_17(\freq_mod_i[17]~input_o ),
	.phi_inc_i_17(\phi_inc_i[17]~input_o ),
	.freq_mod_i_16(\freq_mod_i[16]~input_o ),
	.phi_inc_i_16(\phi_inc_i[16]~input_o ),
	.freq_mod_i_15(\freq_mod_i[15]~input_o ),
	.phi_inc_i_15(\phi_inc_i[15]~input_o ),
	.freq_mod_i_14(\freq_mod_i[14]~input_o ),
	.phi_inc_i_14(\phi_inc_i[14]~input_o ),
	.freq_mod_i_13(\freq_mod_i[13]~input_o ),
	.phi_inc_i_13(\phi_inc_i[13]~input_o ),
	.freq_mod_i_12(\freq_mod_i[12]~input_o ),
	.phi_inc_i_12(\phi_inc_i[12]~input_o ),
	.freq_mod_i_11(\freq_mod_i[11]~input_o ),
	.phi_inc_i_11(\phi_inc_i[11]~input_o ),
	.freq_mod_i_10(\freq_mod_i[10]~input_o ),
	.phi_inc_i_10(\phi_inc_i[10]~input_o ),
	.freq_mod_i_9(\freq_mod_i[9]~input_o ),
	.phi_inc_i_9(\phi_inc_i[9]~input_o ),
	.freq_mod_i_8(\freq_mod_i[8]~input_o ),
	.phi_inc_i_8(\phi_inc_i[8]~input_o ),
	.freq_mod_i_7(\freq_mod_i[7]~input_o ),
	.phi_inc_i_7(\phi_inc_i[7]~input_o ),
	.freq_mod_i_6(\freq_mod_i[6]~input_o ),
	.phi_inc_i_6(\phi_inc_i[6]~input_o ),
	.freq_mod_i_5(\freq_mod_i[5]~input_o ),
	.phi_inc_i_5(\phi_inc_i[5]~input_o ),
	.freq_mod_i_4(\freq_mod_i[4]~input_o ),
	.phi_inc_i_4(\phi_inc_i[4]~input_o ),
	.freq_mod_i_3(\freq_mod_i[3]~input_o ),
	.phi_inc_i_3(\phi_inc_i[3]~input_o ),
	.freq_mod_i_2(\freq_mod_i[2]~input_o ),
	.phi_inc_i_2(\phi_inc_i[2]~input_o ),
	.freq_mod_i_1(\freq_mod_i[1]~input_o ),
	.phi_inc_i_1(\phi_inc_i[1]~input_o ),
	.freq_mod_i_0(\freq_mod_i[0]~input_o ),
	.phi_inc_i_0(\phi_inc_i[0]~input_o ));

assign \clk~input_o  = clk;

assign \reset_n~input_o  = reset_n;

assign \clken~input_o  = clken;

assign \phase_mod_i[0]~input_o  = phase_mod_i[0];

assign \phase_mod_i[1]~input_o  = phase_mod_i[1];

assign \phase_mod_i[2]~input_o  = phase_mod_i[2];

assign \phase_mod_i[3]~input_o  = phase_mod_i[3];

assign \phase_mod_i[4]~input_o  = phase_mod_i[4];

assign \phase_mod_i[5]~input_o  = phase_mod_i[5];

assign \phase_mod_i[6]~input_o  = phase_mod_i[6];

assign \phase_mod_i[7]~input_o  = phase_mod_i[7];

assign \phase_mod_i[8]~input_o  = phase_mod_i[8];

assign \phase_mod_i[9]~input_o  = phase_mod_i[9];

assign \phase_mod_i[10]~input_o  = phase_mod_i[10];

assign \phase_mod_i[11]~input_o  = phase_mod_i[11];

assign \phase_mod_i[12]~input_o  = phase_mod_i[12];

assign \phase_mod_i[15]~input_o  = phase_mod_i[15];

assign \phase_mod_i[13]~input_o  = phase_mod_i[13];

assign \phase_mod_i[14]~input_o  = phase_mod_i[14];

assign \freq_mod_i[31]~input_o  = freq_mod_i[31];

assign \phi_inc_i[32]~input_o  = phi_inc_i[32];

assign \phi_inc_i[33]~input_o  = phi_inc_i[33];

assign \phi_inc_i[34]~input_o  = phi_inc_i[34];

assign \phi_inc_i[35]~input_o  = phi_inc_i[35];

assign \phi_inc_i[36]~input_o  = phi_inc_i[36];

assign \phi_inc_i[37]~input_o  = phi_inc_i[37];

assign \phi_inc_i[38]~input_o  = phi_inc_i[38];

assign \phi_inc_i[39]~input_o  = phi_inc_i[39];

assign \phi_inc_i[40]~input_o  = phi_inc_i[40];

assign \phi_inc_i[41]~input_o  = phi_inc_i[41];

assign \phi_inc_i[42]~input_o  = phi_inc_i[42];

assign \phi_inc_i[43]~input_o  = phi_inc_i[43];

assign \phi_inc_i[44]~input_o  = phi_inc_i[44];

assign \phi_inc_i[47]~input_o  = phi_inc_i[47];

assign \phi_inc_i[31]~input_o  = phi_inc_i[31];

assign \phi_inc_i[45]~input_o  = phi_inc_i[45];

assign \phi_inc_i[46]~input_o  = phi_inc_i[46];

assign \freq_mod_i[30]~input_o  = freq_mod_i[30];

assign \phi_inc_i[30]~input_o  = phi_inc_i[30];

assign \freq_mod_i[29]~input_o  = freq_mod_i[29];

assign \phi_inc_i[29]~input_o  = phi_inc_i[29];

assign \freq_mod_i[28]~input_o  = freq_mod_i[28];

assign \phi_inc_i[28]~input_o  = phi_inc_i[28];

assign \freq_mod_i[27]~input_o  = freq_mod_i[27];

assign \phi_inc_i[27]~input_o  = phi_inc_i[27];

assign \freq_mod_i[26]~input_o  = freq_mod_i[26];

assign \phi_inc_i[26]~input_o  = phi_inc_i[26];

assign \freq_mod_i[25]~input_o  = freq_mod_i[25];

assign \phi_inc_i[25]~input_o  = phi_inc_i[25];

assign \freq_mod_i[24]~input_o  = freq_mod_i[24];

assign \phi_inc_i[24]~input_o  = phi_inc_i[24];

assign \freq_mod_i[23]~input_o  = freq_mod_i[23];

assign \phi_inc_i[23]~input_o  = phi_inc_i[23];

assign \freq_mod_i[22]~input_o  = freq_mod_i[22];

assign \phi_inc_i[22]~input_o  = phi_inc_i[22];

assign \freq_mod_i[21]~input_o  = freq_mod_i[21];

assign \phi_inc_i[21]~input_o  = phi_inc_i[21];

assign \freq_mod_i[20]~input_o  = freq_mod_i[20];

assign \phi_inc_i[20]~input_o  = phi_inc_i[20];

assign \freq_mod_i[19]~input_o  = freq_mod_i[19];

assign \phi_inc_i[19]~input_o  = phi_inc_i[19];

assign \freq_mod_i[18]~input_o  = freq_mod_i[18];

assign \phi_inc_i[18]~input_o  = phi_inc_i[18];

assign \freq_mod_i[17]~input_o  = freq_mod_i[17];

assign \phi_inc_i[17]~input_o  = phi_inc_i[17];

assign \freq_mod_i[16]~input_o  = freq_mod_i[16];

assign \phi_inc_i[16]~input_o  = phi_inc_i[16];

assign \freq_mod_i[15]~input_o  = freq_mod_i[15];

assign \phi_inc_i[15]~input_o  = phi_inc_i[15];

assign \freq_mod_i[14]~input_o  = freq_mod_i[14];

assign \phi_inc_i[14]~input_o  = phi_inc_i[14];

assign \freq_mod_i[13]~input_o  = freq_mod_i[13];

assign \phi_inc_i[13]~input_o  = phi_inc_i[13];

assign \freq_mod_i[12]~input_o  = freq_mod_i[12];

assign \phi_inc_i[12]~input_o  = phi_inc_i[12];

assign \freq_mod_i[11]~input_o  = freq_mod_i[11];

assign \phi_inc_i[11]~input_o  = phi_inc_i[11];

assign \freq_mod_i[10]~input_o  = freq_mod_i[10];

assign \phi_inc_i[10]~input_o  = phi_inc_i[10];

assign \freq_mod_i[9]~input_o  = freq_mod_i[9];

assign \phi_inc_i[9]~input_o  = phi_inc_i[9];

assign \freq_mod_i[8]~input_o  = freq_mod_i[8];

assign \phi_inc_i[8]~input_o  = phi_inc_i[8];

assign \freq_mod_i[7]~input_o  = freq_mod_i[7];

assign \phi_inc_i[7]~input_o  = phi_inc_i[7];

assign \freq_mod_i[6]~input_o  = freq_mod_i[6];

assign \phi_inc_i[6]~input_o  = phi_inc_i[6];

assign \freq_mod_i[5]~input_o  = freq_mod_i[5];

assign \phi_inc_i[5]~input_o  = phi_inc_i[5];

assign \freq_mod_i[4]~input_o  = freq_mod_i[4];

assign \phi_inc_i[4]~input_o  = phi_inc_i[4];

assign \freq_mod_i[3]~input_o  = freq_mod_i[3];

assign \phi_inc_i[3]~input_o  = phi_inc_i[3];

assign \freq_mod_i[2]~input_o  = freq_mod_i[2];

assign \phi_inc_i[2]~input_o  = phi_inc_i[2];

assign \freq_mod_i[1]~input_o  = freq_mod_i[1];

assign \phi_inc_i[1]~input_o  = phi_inc_i[1];

assign \freq_mod_i[0]~input_o  = freq_mod_i[0];

assign \phi_inc_i[0]~input_o  = phi_inc_i[0];

assign fsin_o[0] = \nco_ii_0|ux122|data_out[0]~q ;

assign fsin_o[1] = \nco_ii_0|ux122|data_out[1]~q ;

assign fsin_o[2] = \nco_ii_0|ux122|data_out[2]~q ;

assign fsin_o[3] = \nco_ii_0|ux122|data_out[3]~q ;

assign fsin_o[4] = \nco_ii_0|ux122|data_out[4]~q ;

assign fsin_o[5] = \nco_ii_0|ux122|data_out[5]~q ;

assign fsin_o[6] = \nco_ii_0|ux122|data_out[6]~q ;

assign fsin_o[7] = \nco_ii_0|ux122|data_out[7]~q ;

assign fsin_o[8] = \nco_ii_0|ux122|data_out[8]~q ;

assign fsin_o[9] = \nco_ii_0|ux122|data_out[9]~q ;

assign fsin_o[10] = \nco_ii_0|ux122|data_out[10]~q ;

assign fsin_o[11] = \nco_ii_0|ux122|data_out[11]~q ;

assign fsin_o[12] = \nco_ii_0|ux122|data_out[12]~q ;

assign fsin_o[13] = \nco_ii_0|ux122|data_out[13]~q ;

assign fsin_o[14] = \nco_ii_0|ux122|data_out[14]~q ;

assign fsin_o[15] = \nco_ii_0|ux122|data_out[15]~q ;

assign fcos_o[0] = \nco_ii_0|ux123|data_out[0]~q ;

assign fcos_o[1] = \nco_ii_0|ux123|data_out[1]~q ;

assign fcos_o[2] = \nco_ii_0|ux123|data_out[2]~q ;

assign fcos_o[3] = \nco_ii_0|ux123|data_out[3]~q ;

assign fcos_o[4] = \nco_ii_0|ux123|data_out[4]~q ;

assign fcos_o[5] = \nco_ii_0|ux123|data_out[5]~q ;

assign fcos_o[6] = \nco_ii_0|ux123|data_out[6]~q ;

assign fcos_o[7] = \nco_ii_0|ux123|data_out[7]~q ;

assign fcos_o[8] = \nco_ii_0|ux123|data_out[8]~q ;

assign fcos_o[9] = \nco_ii_0|ux123|data_out[9]~q ;

assign fcos_o[10] = \nco_ii_0|ux123|data_out[10]~q ;

assign fcos_o[11] = \nco_ii_0|ux123|data_out[11]~q ;

assign fcos_o[12] = \nco_ii_0|ux123|data_out[12]~q ;

assign fcos_o[13] = \nco_ii_0|ux123|data_out[13]~q ;

assign fcos_o[14] = \nco_ii_0|ux123|data_out[14]~q ;

assign fcos_o[15] = \nco_ii_0|ux123|data_out[15]~q ;

assign out_valid = \nco_ii_0|ux710isdr|data_ready~q ;

endmodule

module DDS_48_v1_DDS_48_v1_nco_ii_0 (
	data_out_0,
	data_out_1,
	data_out_2,
	data_out_3,
	data_out_4,
	data_out_5,
	data_out_6,
	data_out_7,
	data_out_8,
	data_out_9,
	data_out_10,
	data_out_11,
	data_out_12,
	data_out_13,
	data_out_14,
	data_out_15,
	data_out_01,
	data_out_16,
	data_out_21,
	data_out_31,
	data_out_41,
	data_out_51,
	data_out_61,
	data_out_71,
	data_out_81,
	data_out_91,
	data_out_101,
	data_out_111,
	data_out_121,
	data_out_131,
	data_out_141,
	data_out_151,
	data_ready,
	clk,
	reset_n,
	clken,
	phase_mod_i_0,
	phase_mod_i_1,
	phase_mod_i_2,
	phase_mod_i_3,
	phase_mod_i_4,
	phase_mod_i_5,
	phase_mod_i_6,
	phase_mod_i_7,
	phase_mod_i_8,
	phase_mod_i_9,
	phase_mod_i_10,
	phase_mod_i_11,
	phase_mod_i_12,
	phase_mod_i_15,
	phase_mod_i_13,
	phase_mod_i_14,
	freq_mod_i_31,
	phi_inc_i_32,
	phi_inc_i_33,
	phi_inc_i_34,
	phi_inc_i_35,
	phi_inc_i_36,
	phi_inc_i_37,
	phi_inc_i_38,
	phi_inc_i_39,
	phi_inc_i_40,
	phi_inc_i_41,
	phi_inc_i_42,
	phi_inc_i_43,
	phi_inc_i_44,
	phi_inc_i_47,
	phi_inc_i_31,
	phi_inc_i_45,
	phi_inc_i_46,
	freq_mod_i_30,
	phi_inc_i_30,
	freq_mod_i_29,
	phi_inc_i_29,
	freq_mod_i_28,
	phi_inc_i_28,
	freq_mod_i_27,
	phi_inc_i_27,
	freq_mod_i_26,
	phi_inc_i_26,
	freq_mod_i_25,
	phi_inc_i_25,
	freq_mod_i_24,
	phi_inc_i_24,
	freq_mod_i_23,
	phi_inc_i_23,
	freq_mod_i_22,
	phi_inc_i_22,
	freq_mod_i_21,
	phi_inc_i_21,
	freq_mod_i_20,
	phi_inc_i_20,
	freq_mod_i_19,
	phi_inc_i_19,
	freq_mod_i_18,
	phi_inc_i_18,
	freq_mod_i_17,
	phi_inc_i_17,
	freq_mod_i_16,
	phi_inc_i_16,
	freq_mod_i_15,
	phi_inc_i_15,
	freq_mod_i_14,
	phi_inc_i_14,
	freq_mod_i_13,
	phi_inc_i_13,
	freq_mod_i_12,
	phi_inc_i_12,
	freq_mod_i_11,
	phi_inc_i_11,
	freq_mod_i_10,
	phi_inc_i_10,
	freq_mod_i_9,
	phi_inc_i_9,
	freq_mod_i_8,
	phi_inc_i_8,
	freq_mod_i_7,
	phi_inc_i_7,
	freq_mod_i_6,
	phi_inc_i_6,
	freq_mod_i_5,
	phi_inc_i_5,
	freq_mod_i_4,
	phi_inc_i_4,
	freq_mod_i_3,
	phi_inc_i_3,
	freq_mod_i_2,
	phi_inc_i_2,
	freq_mod_i_1,
	phi_inc_i_1,
	freq_mod_i_0,
	phi_inc_i_0)/* synthesis synthesis_greybox=1 */;
output 	data_out_0;
output 	data_out_1;
output 	data_out_2;
output 	data_out_3;
output 	data_out_4;
output 	data_out_5;
output 	data_out_6;
output 	data_out_7;
output 	data_out_8;
output 	data_out_9;
output 	data_out_10;
output 	data_out_11;
output 	data_out_12;
output 	data_out_13;
output 	data_out_14;
output 	data_out_15;
output 	data_out_01;
output 	data_out_16;
output 	data_out_21;
output 	data_out_31;
output 	data_out_41;
output 	data_out_51;
output 	data_out_61;
output 	data_out_71;
output 	data_out_81;
output 	data_out_91;
output 	data_out_101;
output 	data_out_111;
output 	data_out_121;
output 	data_out_131;
output 	data_out_141;
output 	data_out_151;
output 	data_ready;
input 	clk;
input 	reset_n;
input 	clken;
input 	phase_mod_i_0;
input 	phase_mod_i_1;
input 	phase_mod_i_2;
input 	phase_mod_i_3;
input 	phase_mod_i_4;
input 	phase_mod_i_5;
input 	phase_mod_i_6;
input 	phase_mod_i_7;
input 	phase_mod_i_8;
input 	phase_mod_i_9;
input 	phase_mod_i_10;
input 	phase_mod_i_11;
input 	phase_mod_i_12;
input 	phase_mod_i_15;
input 	phase_mod_i_13;
input 	phase_mod_i_14;
input 	freq_mod_i_31;
input 	phi_inc_i_32;
input 	phi_inc_i_33;
input 	phi_inc_i_34;
input 	phi_inc_i_35;
input 	phi_inc_i_36;
input 	phi_inc_i_37;
input 	phi_inc_i_38;
input 	phi_inc_i_39;
input 	phi_inc_i_40;
input 	phi_inc_i_41;
input 	phi_inc_i_42;
input 	phi_inc_i_43;
input 	phi_inc_i_44;
input 	phi_inc_i_47;
input 	phi_inc_i_31;
input 	phi_inc_i_45;
input 	phi_inc_i_46;
input 	freq_mod_i_30;
input 	phi_inc_i_30;
input 	freq_mod_i_29;
input 	phi_inc_i_29;
input 	freq_mod_i_28;
input 	phi_inc_i_28;
input 	freq_mod_i_27;
input 	phi_inc_i_27;
input 	freq_mod_i_26;
input 	phi_inc_i_26;
input 	freq_mod_i_25;
input 	phi_inc_i_25;
input 	freq_mod_i_24;
input 	phi_inc_i_24;
input 	freq_mod_i_23;
input 	phi_inc_i_23;
input 	freq_mod_i_22;
input 	phi_inc_i_22;
input 	freq_mod_i_21;
input 	phi_inc_i_21;
input 	freq_mod_i_20;
input 	phi_inc_i_20;
input 	freq_mod_i_19;
input 	phi_inc_i_19;
input 	freq_mod_i_18;
input 	phi_inc_i_18;
input 	freq_mod_i_17;
input 	phi_inc_i_17;
input 	freq_mod_i_16;
input 	phi_inc_i_16;
input 	freq_mod_i_15;
input 	phi_inc_i_15;
input 	freq_mod_i_14;
input 	phi_inc_i_14;
input 	freq_mod_i_13;
input 	phi_inc_i_13;
input 	freq_mod_i_12;
input 	phi_inc_i_12;
input 	freq_mod_i_11;
input 	phi_inc_i_11;
input 	freq_mod_i_10;
input 	phi_inc_i_10;
input 	freq_mod_i_9;
input 	phi_inc_i_9;
input 	freq_mod_i_8;
input 	phi_inc_i_8;
input 	freq_mod_i_7;
input 	phi_inc_i_7;
input 	freq_mod_i_6;
input 	phi_inc_i_6;
input 	freq_mod_i_5;
input 	phi_inc_i_5;
input 	freq_mod_i_4;
input 	phi_inc_i_4;
input 	freq_mod_i_3;
input 	phi_inc_i_3;
input 	freq_mod_i_2;
input 	phi_inc_i_2;
input 	freq_mod_i_1;
input 	phi_inc_i_1;
input 	freq_mod_i_0;
input 	phi_inc_i_0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \ux0120|altsyncram_component0|auto_generated|ram_block1a64~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a80~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a96~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a112~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a32~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a48~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a0~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a16~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a65~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a81~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a97~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a113~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a33~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a49~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a1~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a17~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a66~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a82~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a98~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a114~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a34~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a50~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a2~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a18~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a67~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a83~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a99~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a115~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a35~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a51~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a3~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a19~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a68~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a84~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a100~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a116~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a36~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a52~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a4~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a20~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a69~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a85~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a101~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a117~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a37~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a53~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a5~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a21~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a70~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a86~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a102~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a118~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a38~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a54~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a6~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a22~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a71~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a87~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a103~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a119~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a39~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a55~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a7~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a23~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a72~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a88~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a104~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a120~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a40~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a56~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a8~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a24~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a73~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a89~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a105~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a121~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a41~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a57~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a9~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a25~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a74~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a90~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a106~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a122~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a42~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a58~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a10~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a26~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a75~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a91~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a107~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a123~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a43~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a59~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a11~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a27~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a76~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a92~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a108~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a124~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a44~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a60~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a12~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a28~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a77~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a93~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a109~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a125~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a45~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a61~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a13~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a29~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a78~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a94~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a110~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a126~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a46~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a62~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a14~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a30~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a79~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a95~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a111~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a127~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a47~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a63~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a15~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a31~portadataout ;
wire \ux0121|altsyncram_component0|auto_generated|ram_block1a64~portadataout ;
wire \ux0121|altsyncram_component0|auto_generated|ram_block1a80~portadataout ;
wire \ux0121|altsyncram_component0|auto_generated|ram_block1a96~portadataout ;
wire \ux0121|altsyncram_component0|auto_generated|ram_block1a112~portadataout ;
wire \ux0121|altsyncram_component0|auto_generated|ram_block1a32~portadataout ;
wire \ux0121|altsyncram_component0|auto_generated|ram_block1a48~portadataout ;
wire \ux0121|altsyncram_component0|auto_generated|ram_block1a0~portadataout ;
wire \ux0121|altsyncram_component0|auto_generated|ram_block1a16~portadataout ;
wire \ux0121|altsyncram_component0|auto_generated|ram_block1a65~portadataout ;
wire \ux0121|altsyncram_component0|auto_generated|ram_block1a81~portadataout ;
wire \ux0121|altsyncram_component0|auto_generated|ram_block1a97~portadataout ;
wire \ux0121|altsyncram_component0|auto_generated|ram_block1a113~portadataout ;
wire \ux0121|altsyncram_component0|auto_generated|ram_block1a33~portadataout ;
wire \ux0121|altsyncram_component0|auto_generated|ram_block1a49~portadataout ;
wire \ux0121|altsyncram_component0|auto_generated|ram_block1a1~portadataout ;
wire \ux0121|altsyncram_component0|auto_generated|ram_block1a17~portadataout ;
wire \ux0121|altsyncram_component0|auto_generated|ram_block1a66~portadataout ;
wire \ux0121|altsyncram_component0|auto_generated|ram_block1a82~portadataout ;
wire \ux0121|altsyncram_component0|auto_generated|ram_block1a98~portadataout ;
wire \ux0121|altsyncram_component0|auto_generated|ram_block1a114~portadataout ;
wire \ux0121|altsyncram_component0|auto_generated|ram_block1a34~portadataout ;
wire \ux0121|altsyncram_component0|auto_generated|ram_block1a50~portadataout ;
wire \ux0121|altsyncram_component0|auto_generated|ram_block1a2~portadataout ;
wire \ux0121|altsyncram_component0|auto_generated|ram_block1a18~portadataout ;
wire \ux0121|altsyncram_component0|auto_generated|ram_block1a67~portadataout ;
wire \ux0121|altsyncram_component0|auto_generated|ram_block1a83~portadataout ;
wire \ux0121|altsyncram_component0|auto_generated|ram_block1a99~portadataout ;
wire \ux0121|altsyncram_component0|auto_generated|ram_block1a115~portadataout ;
wire \ux0121|altsyncram_component0|auto_generated|ram_block1a35~portadataout ;
wire \ux0121|altsyncram_component0|auto_generated|ram_block1a51~portadataout ;
wire \ux0121|altsyncram_component0|auto_generated|ram_block1a3~portadataout ;
wire \ux0121|altsyncram_component0|auto_generated|ram_block1a19~portadataout ;
wire \ux0121|altsyncram_component0|auto_generated|ram_block1a68~portadataout ;
wire \ux0121|altsyncram_component0|auto_generated|ram_block1a84~portadataout ;
wire \ux0121|altsyncram_component0|auto_generated|ram_block1a100~portadataout ;
wire \ux0121|altsyncram_component0|auto_generated|ram_block1a116~portadataout ;
wire \ux0121|altsyncram_component0|auto_generated|ram_block1a36~portadataout ;
wire \ux0121|altsyncram_component0|auto_generated|ram_block1a52~portadataout ;
wire \ux0121|altsyncram_component0|auto_generated|ram_block1a4~portadataout ;
wire \ux0121|altsyncram_component0|auto_generated|ram_block1a20~portadataout ;
wire \ux0121|altsyncram_component0|auto_generated|ram_block1a69~portadataout ;
wire \ux0121|altsyncram_component0|auto_generated|ram_block1a85~portadataout ;
wire \ux0121|altsyncram_component0|auto_generated|ram_block1a101~portadataout ;
wire \ux0121|altsyncram_component0|auto_generated|ram_block1a117~portadataout ;
wire \ux0121|altsyncram_component0|auto_generated|ram_block1a37~portadataout ;
wire \ux0121|altsyncram_component0|auto_generated|ram_block1a53~portadataout ;
wire \ux0121|altsyncram_component0|auto_generated|ram_block1a5~portadataout ;
wire \ux0121|altsyncram_component0|auto_generated|ram_block1a21~portadataout ;
wire \ux0121|altsyncram_component0|auto_generated|ram_block1a70~portadataout ;
wire \ux0121|altsyncram_component0|auto_generated|ram_block1a86~portadataout ;
wire \ux0121|altsyncram_component0|auto_generated|ram_block1a102~portadataout ;
wire \ux0121|altsyncram_component0|auto_generated|ram_block1a118~portadataout ;
wire \ux0121|altsyncram_component0|auto_generated|ram_block1a38~portadataout ;
wire \ux0121|altsyncram_component0|auto_generated|ram_block1a54~portadataout ;
wire \ux0121|altsyncram_component0|auto_generated|ram_block1a6~portadataout ;
wire \ux0121|altsyncram_component0|auto_generated|ram_block1a22~portadataout ;
wire \ux0121|altsyncram_component0|auto_generated|ram_block1a71~portadataout ;
wire \ux0121|altsyncram_component0|auto_generated|ram_block1a87~portadataout ;
wire \ux0121|altsyncram_component0|auto_generated|ram_block1a103~portadataout ;
wire \ux0121|altsyncram_component0|auto_generated|ram_block1a119~portadataout ;
wire \ux0121|altsyncram_component0|auto_generated|ram_block1a39~portadataout ;
wire \ux0121|altsyncram_component0|auto_generated|ram_block1a55~portadataout ;
wire \ux0121|altsyncram_component0|auto_generated|ram_block1a7~portadataout ;
wire \ux0121|altsyncram_component0|auto_generated|ram_block1a23~portadataout ;
wire \ux0121|altsyncram_component0|auto_generated|ram_block1a72~portadataout ;
wire \ux0121|altsyncram_component0|auto_generated|ram_block1a88~portadataout ;
wire \ux0121|altsyncram_component0|auto_generated|ram_block1a104~portadataout ;
wire \ux0121|altsyncram_component0|auto_generated|ram_block1a120~portadataout ;
wire \ux0121|altsyncram_component0|auto_generated|ram_block1a40~portadataout ;
wire \ux0121|altsyncram_component0|auto_generated|ram_block1a56~portadataout ;
wire \ux0121|altsyncram_component0|auto_generated|ram_block1a8~portadataout ;
wire \ux0121|altsyncram_component0|auto_generated|ram_block1a24~portadataout ;
wire \ux0121|altsyncram_component0|auto_generated|ram_block1a73~portadataout ;
wire \ux0121|altsyncram_component0|auto_generated|ram_block1a89~portadataout ;
wire \ux0121|altsyncram_component0|auto_generated|ram_block1a105~portadataout ;
wire \ux0121|altsyncram_component0|auto_generated|ram_block1a121~portadataout ;
wire \ux0121|altsyncram_component0|auto_generated|ram_block1a41~portadataout ;
wire \ux0121|altsyncram_component0|auto_generated|ram_block1a57~portadataout ;
wire \ux0121|altsyncram_component0|auto_generated|ram_block1a9~portadataout ;
wire \ux0121|altsyncram_component0|auto_generated|ram_block1a25~portadataout ;
wire \ux0121|altsyncram_component0|auto_generated|ram_block1a74~portadataout ;
wire \ux0121|altsyncram_component0|auto_generated|ram_block1a90~portadataout ;
wire \ux0121|altsyncram_component0|auto_generated|ram_block1a106~portadataout ;
wire \ux0121|altsyncram_component0|auto_generated|ram_block1a122~portadataout ;
wire \ux0121|altsyncram_component0|auto_generated|ram_block1a42~portadataout ;
wire \ux0121|altsyncram_component0|auto_generated|ram_block1a58~portadataout ;
wire \ux0121|altsyncram_component0|auto_generated|ram_block1a10~portadataout ;
wire \ux0121|altsyncram_component0|auto_generated|ram_block1a26~portadataout ;
wire \ux0121|altsyncram_component0|auto_generated|ram_block1a75~portadataout ;
wire \ux0121|altsyncram_component0|auto_generated|ram_block1a91~portadataout ;
wire \ux0121|altsyncram_component0|auto_generated|ram_block1a107~portadataout ;
wire \ux0121|altsyncram_component0|auto_generated|ram_block1a123~portadataout ;
wire \ux0121|altsyncram_component0|auto_generated|ram_block1a43~portadataout ;
wire \ux0121|altsyncram_component0|auto_generated|ram_block1a59~portadataout ;
wire \ux0121|altsyncram_component0|auto_generated|ram_block1a11~portadataout ;
wire \ux0121|altsyncram_component0|auto_generated|ram_block1a27~portadataout ;
wire \ux0121|altsyncram_component0|auto_generated|ram_block1a76~portadataout ;
wire \ux0121|altsyncram_component0|auto_generated|ram_block1a92~portadataout ;
wire \ux0121|altsyncram_component0|auto_generated|ram_block1a108~portadataout ;
wire \ux0121|altsyncram_component0|auto_generated|ram_block1a124~portadataout ;
wire \ux0121|altsyncram_component0|auto_generated|ram_block1a44~portadataout ;
wire \ux0121|altsyncram_component0|auto_generated|ram_block1a60~portadataout ;
wire \ux0121|altsyncram_component0|auto_generated|ram_block1a12~portadataout ;
wire \ux0121|altsyncram_component0|auto_generated|ram_block1a28~portadataout ;
wire \ux0121|altsyncram_component0|auto_generated|ram_block1a77~portadataout ;
wire \ux0121|altsyncram_component0|auto_generated|ram_block1a93~portadataout ;
wire \ux0121|altsyncram_component0|auto_generated|ram_block1a109~portadataout ;
wire \ux0121|altsyncram_component0|auto_generated|ram_block1a125~portadataout ;
wire \ux0121|altsyncram_component0|auto_generated|ram_block1a45~portadataout ;
wire \ux0121|altsyncram_component0|auto_generated|ram_block1a61~portadataout ;
wire \ux0121|altsyncram_component0|auto_generated|ram_block1a13~portadataout ;
wire \ux0121|altsyncram_component0|auto_generated|ram_block1a29~portadataout ;
wire \ux0121|altsyncram_component0|auto_generated|ram_block1a78~portadataout ;
wire \ux0121|altsyncram_component0|auto_generated|ram_block1a94~portadataout ;
wire \ux0121|altsyncram_component0|auto_generated|ram_block1a110~portadataout ;
wire \ux0121|altsyncram_component0|auto_generated|ram_block1a126~portadataout ;
wire \ux0121|altsyncram_component0|auto_generated|ram_block1a46~portadataout ;
wire \ux0121|altsyncram_component0|auto_generated|ram_block1a62~portadataout ;
wire \ux0121|altsyncram_component0|auto_generated|ram_block1a14~portadataout ;
wire \ux0121|altsyncram_component0|auto_generated|ram_block1a30~portadataout ;
wire \ux0121|altsyncram_component0|auto_generated|ram_block1a79~portadataout ;
wire \ux0121|altsyncram_component0|auto_generated|ram_block1a95~portadataout ;
wire \ux0121|altsyncram_component0|auto_generated|ram_block1a111~portadataout ;
wire \ux0121|altsyncram_component0|auto_generated|ram_block1a127~portadataout ;
wire \ux0121|altsyncram_component0|auto_generated|ram_block1a47~portadataout ;
wire \ux0121|altsyncram_component0|auto_generated|ram_block1a63~portadataout ;
wire \ux0121|altsyncram_component0|auto_generated|ram_block1a15~portadataout ;
wire \ux0121|altsyncram_component0|auto_generated|ram_block1a31~portadataout ;
wire \ux009|rom_add[0]~q ;
wire \ux009|rom_add[1]~q ;
wire \ux009|rom_add[2]~q ;
wire \ux009|rom_add[3]~q ;
wire \ux009|rom_add[4]~q ;
wire \ux009|rom_add[5]~q ;
wire \ux009|rom_add[6]~q ;
wire \ux009|rom_add[7]~q ;
wire \ux009|rom_add[8]~q ;
wire \ux009|rom_add[9]~q ;
wire \ux009|rom_add[10]~q ;
wire \ux009|rom_add[11]~q ;
wire \ux009|rom_add[12]~q ;
wire \ux009|rom_add[15]~q ;
wire \ux009|rom_add[13]~q ;
wire \ux009|rom_add[14]~q ;
wire \ux002|dxxpdo[5]~q ;
wire \ux002|dxxpdo[6]~q ;
wire \ux002|dxxpdo[7]~q ;
wire \ux002|dxxpdo[8]~q ;
wire \ux002|dxxpdo[9]~q ;
wire \ux002|dxxpdo[10]~q ;
wire \ux002|dxxpdo[11]~q ;
wire \ux002|dxxpdo[12]~q ;
wire \ux002|dxxpdo[13]~q ;
wire \ux002|dxxpdo[14]~q ;
wire \ux002|dxxpdo[15]~q ;
wire \ux002|dxxpdo[16]~q ;
wire \ux002|dxxpdo[17]~q ;
wire \ux002|dxxpdo[20]~q ;
wire \ux002|dxxpdo[18]~q ;
wire \ux002|dxxpdo[19]~q ;
wire \ux001|dxxrv[5]~q ;
wire \ux001|dxxrv[6]~q ;
wire \ux001|dxxrv[7]~q ;
wire \ux001|dxxrv[8]~q ;
wire \ux001|dxxrv[9]~q ;
wire \ux001|dxxrv[4]~q ;
wire \ux001|dxxrv[3]~q ;
wire \ux001|dxxrv[2]~q ;
wire \ux001|dxxrv[1]~q ;
wire \ux001|dxxrv[0]~q ;
wire \ux0120|altsyncram_component0|auto_generated|out_address_reg_a[2]~q ;
wire \ux0120|altsyncram_component0|auto_generated|out_address_reg_a[0]~q ;
wire \ux0120|altsyncram_component0|auto_generated|out_address_reg_a[1]~q ;
wire \ux122|data_out[12]~3_combout ;
wire \ux004|acc|auto_generated|pipeline_dffe[0]~q ;
wire \ux004|acc|auto_generated|pipeline_dffe[1]~q ;
wire \ux004|acc|auto_generated|pipeline_dffe[2]~q ;
wire \ux004|acc|auto_generated|pipeline_dffe[3]~q ;
wire \ux004|acc|auto_generated|pipeline_dffe[4]~q ;
wire \ux004|acc|auto_generated|pipeline_dffe[5]~q ;
wire \ux004|acc|auto_generated|pipeline_dffe[6]~q ;
wire \ux004|acc|auto_generated|pipeline_dffe[7]~q ;
wire \ux004|acc|auto_generated|pipeline_dffe[8]~q ;
wire \ux004|acc|auto_generated|pipeline_dffe[9]~q ;
wire \ux004|acc|auto_generated|pipeline_dffe[10]~q ;
wire \ux004|acc|auto_generated|pipeline_dffe[11]~q ;
wire \ux004|acc|auto_generated|pipeline_dffe[12]~q ;
wire \ux004|acc|auto_generated|pipeline_dffe[15]~q ;
wire \ux004|acc|auto_generated|pipeline_dffe[13]~q ;
wire \ux004|acc|auto_generated|pipeline_dffe[14]~q ;
wire \ux000|acc|auto_generated|pipeline_dffe[32]~q ;
wire \ux000|acc|auto_generated|pipeline_dffe[33]~q ;
wire \ux000|acc|auto_generated|pipeline_dffe[34]~q ;
wire \ux000|acc|auto_generated|pipeline_dffe[35]~q ;
wire \ux000|acc|auto_generated|pipeline_dffe[36]~q ;
wire \ux000|acc|auto_generated|pipeline_dffe[37]~q ;
wire \ux000|acc|auto_generated|pipeline_dffe[38]~q ;
wire \ux000|acc|auto_generated|pipeline_dffe[39]~q ;
wire \ux000|acc|auto_generated|pipeline_dffe[40]~q ;
wire \ux000|acc|auto_generated|pipeline_dffe[41]~q ;
wire \ux000|acc|auto_generated|pipeline_dffe[42]~q ;
wire \ux000|acc|auto_generated|pipeline_dffe[43]~q ;
wire \ux000|acc|auto_generated|pipeline_dffe[44]~q ;
wire \ux000|acc|auto_generated|pipeline_dffe[47]~q ;
wire \ux000|acc|auto_generated|pipeline_dffe[31]~q ;
wire \ux000|acc|auto_generated|pipeline_dffe[45]~q ;
wire \ux000|acc|auto_generated|pipeline_dffe[46]~q ;
wire \ux000|acc|auto_generated|pipeline_dffe[30]~q ;
wire \ux003|acc|auto_generated|pipeline_dffe[32]~q ;
wire \ux000|acc|auto_generated|pipeline_dffe[29]~q ;
wire \ux003|acc|auto_generated|pipeline_dffe[33]~q ;
wire \ux003|acc|auto_generated|pipeline_dffe[34]~q ;
wire \ux003|acc|auto_generated|pipeline_dffe[35]~q ;
wire \ux003|acc|auto_generated|pipeline_dffe[36]~q ;
wire \ux003|acc|auto_generated|pipeline_dffe[37]~q ;
wire \ux003|acc|auto_generated|pipeline_dffe[38]~q ;
wire \ux003|acc|auto_generated|pipeline_dffe[39]~q ;
wire \ux003|acc|auto_generated|pipeline_dffe[40]~q ;
wire \ux003|acc|auto_generated|pipeline_dffe[41]~q ;
wire \ux003|acc|auto_generated|pipeline_dffe[42]~q ;
wire \ux003|acc|auto_generated|pipeline_dffe[43]~q ;
wire \ux003|acc|auto_generated|pipeline_dffe[44]~q ;
wire \ux003|acc|auto_generated|pipeline_dffe[47]~q ;
wire \ux003|acc|auto_generated|pipeline_dffe[31]~q ;
wire \ux000|acc|auto_generated|pipeline_dffe[28]~q ;
wire \ux003|acc|auto_generated|pipeline_dffe[45]~q ;
wire \ux003|acc|auto_generated|pipeline_dffe[46]~q ;
wire \ux003|acc|auto_generated|pipeline_dffe[30]~q ;
wire \ux000|acc|auto_generated|pipeline_dffe[27]~q ;
wire \ux003|acc|auto_generated|pipeline_dffe[29]~q ;
wire \ux003|acc|auto_generated|pipeline_dffe[28]~q ;
wire \ux003|acc|auto_generated|pipeline_dffe[27]~q ;
wire \ux003|acc|auto_generated|pipeline_dffe[26]~q ;
wire \ux003|acc|auto_generated|pipeline_dffe[25]~q ;
wire \ux003|acc|auto_generated|pipeline_dffe[24]~q ;
wire \ux003|acc|auto_generated|pipeline_dffe[23]~q ;
wire \ux003|acc|auto_generated|pipeline_dffe[22]~q ;
wire \ux003|acc|auto_generated|pipeline_dffe[21]~q ;
wire \ux003|acc|auto_generated|pipeline_dffe[20]~q ;
wire \ux003|acc|auto_generated|pipeline_dffe[19]~q ;
wire \ux003|acc|auto_generated|pipeline_dffe[18]~q ;
wire \ux003|acc|auto_generated|pipeline_dffe[17]~q ;
wire \ux003|acc|auto_generated|pipeline_dffe[16]~q ;
wire \ux003|acc|auto_generated|pipeline_dffe[15]~q ;
wire \ux003|acc|auto_generated|pipeline_dffe[14]~q ;
wire \ux003|acc|auto_generated|pipeline_dffe[13]~q ;
wire \ux003|acc|auto_generated|pipeline_dffe[12]~q ;
wire \ux003|acc|auto_generated|pipeline_dffe[11]~q ;
wire \ux003|acc|auto_generated|pipeline_dffe[10]~q ;
wire \ux003|acc|auto_generated|pipeline_dffe[9]~q ;
wire \ux003|acc|auto_generated|pipeline_dffe[8]~q ;
wire \ux003|acc|auto_generated|pipeline_dffe[7]~q ;
wire \ux003|acc|auto_generated|pipeline_dffe[6]~q ;
wire \ux003|acc|auto_generated|pipeline_dffe[5]~q ;
wire \ux003|acc|auto_generated|pipeline_dffe[4]~q ;
wire \ux003|acc|auto_generated|pipeline_dffe[3]~q ;
wire \ux003|acc|auto_generated|pipeline_dffe[2]~q ;
wire \ux003|acc|auto_generated|pipeline_dffe[1]~q ;
wire \ux003|acc|auto_generated|pipeline_dffe[0]~q ;


DDS_48_v1_asj_nco_fxx ux003(
	.pipeline_dffe_32(\ux003|acc|auto_generated|pipeline_dffe[32]~q ),
	.pipeline_dffe_33(\ux003|acc|auto_generated|pipeline_dffe[33]~q ),
	.pipeline_dffe_34(\ux003|acc|auto_generated|pipeline_dffe[34]~q ),
	.pipeline_dffe_35(\ux003|acc|auto_generated|pipeline_dffe[35]~q ),
	.pipeline_dffe_36(\ux003|acc|auto_generated|pipeline_dffe[36]~q ),
	.pipeline_dffe_37(\ux003|acc|auto_generated|pipeline_dffe[37]~q ),
	.pipeline_dffe_38(\ux003|acc|auto_generated|pipeline_dffe[38]~q ),
	.pipeline_dffe_39(\ux003|acc|auto_generated|pipeline_dffe[39]~q ),
	.pipeline_dffe_40(\ux003|acc|auto_generated|pipeline_dffe[40]~q ),
	.pipeline_dffe_41(\ux003|acc|auto_generated|pipeline_dffe[41]~q ),
	.pipeline_dffe_42(\ux003|acc|auto_generated|pipeline_dffe[42]~q ),
	.pipeline_dffe_43(\ux003|acc|auto_generated|pipeline_dffe[43]~q ),
	.pipeline_dffe_44(\ux003|acc|auto_generated|pipeline_dffe[44]~q ),
	.pipeline_dffe_47(\ux003|acc|auto_generated|pipeline_dffe[47]~q ),
	.pipeline_dffe_31(\ux003|acc|auto_generated|pipeline_dffe[31]~q ),
	.pipeline_dffe_45(\ux003|acc|auto_generated|pipeline_dffe[45]~q ),
	.pipeline_dffe_46(\ux003|acc|auto_generated|pipeline_dffe[46]~q ),
	.pipeline_dffe_30(\ux003|acc|auto_generated|pipeline_dffe[30]~q ),
	.pipeline_dffe_29(\ux003|acc|auto_generated|pipeline_dffe[29]~q ),
	.pipeline_dffe_28(\ux003|acc|auto_generated|pipeline_dffe[28]~q ),
	.pipeline_dffe_27(\ux003|acc|auto_generated|pipeline_dffe[27]~q ),
	.pipeline_dffe_26(\ux003|acc|auto_generated|pipeline_dffe[26]~q ),
	.pipeline_dffe_25(\ux003|acc|auto_generated|pipeline_dffe[25]~q ),
	.pipeline_dffe_24(\ux003|acc|auto_generated|pipeline_dffe[24]~q ),
	.pipeline_dffe_23(\ux003|acc|auto_generated|pipeline_dffe[23]~q ),
	.pipeline_dffe_22(\ux003|acc|auto_generated|pipeline_dffe[22]~q ),
	.pipeline_dffe_21(\ux003|acc|auto_generated|pipeline_dffe[21]~q ),
	.pipeline_dffe_20(\ux003|acc|auto_generated|pipeline_dffe[20]~q ),
	.pipeline_dffe_19(\ux003|acc|auto_generated|pipeline_dffe[19]~q ),
	.pipeline_dffe_18(\ux003|acc|auto_generated|pipeline_dffe[18]~q ),
	.pipeline_dffe_17(\ux003|acc|auto_generated|pipeline_dffe[17]~q ),
	.pipeline_dffe_16(\ux003|acc|auto_generated|pipeline_dffe[16]~q ),
	.pipeline_dffe_15(\ux003|acc|auto_generated|pipeline_dffe[15]~q ),
	.pipeline_dffe_14(\ux003|acc|auto_generated|pipeline_dffe[14]~q ),
	.pipeline_dffe_13(\ux003|acc|auto_generated|pipeline_dffe[13]~q ),
	.pipeline_dffe_12(\ux003|acc|auto_generated|pipeline_dffe[12]~q ),
	.pipeline_dffe_11(\ux003|acc|auto_generated|pipeline_dffe[11]~q ),
	.pipeline_dffe_10(\ux003|acc|auto_generated|pipeline_dffe[10]~q ),
	.pipeline_dffe_9(\ux003|acc|auto_generated|pipeline_dffe[9]~q ),
	.pipeline_dffe_8(\ux003|acc|auto_generated|pipeline_dffe[8]~q ),
	.pipeline_dffe_7(\ux003|acc|auto_generated|pipeline_dffe[7]~q ),
	.pipeline_dffe_6(\ux003|acc|auto_generated|pipeline_dffe[6]~q ),
	.pipeline_dffe_5(\ux003|acc|auto_generated|pipeline_dffe[5]~q ),
	.pipeline_dffe_4(\ux003|acc|auto_generated|pipeline_dffe[4]~q ),
	.pipeline_dffe_3(\ux003|acc|auto_generated|pipeline_dffe[3]~q ),
	.pipeline_dffe_2(\ux003|acc|auto_generated|pipeline_dffe[2]~q ),
	.pipeline_dffe_1(\ux003|acc|auto_generated|pipeline_dffe[1]~q ),
	.pipeline_dffe_0(\ux003|acc|auto_generated|pipeline_dffe[0]~q ),
	.clk(clk),
	.reset_n(reset_n),
	.clken(clken),
	.freq_mod_i_31(freq_mod_i_31),
	.phi_inc_i_32(phi_inc_i_32),
	.phi_inc_i_33(phi_inc_i_33),
	.phi_inc_i_34(phi_inc_i_34),
	.phi_inc_i_35(phi_inc_i_35),
	.phi_inc_i_36(phi_inc_i_36),
	.phi_inc_i_37(phi_inc_i_37),
	.phi_inc_i_38(phi_inc_i_38),
	.phi_inc_i_39(phi_inc_i_39),
	.phi_inc_i_40(phi_inc_i_40),
	.phi_inc_i_41(phi_inc_i_41),
	.phi_inc_i_42(phi_inc_i_42),
	.phi_inc_i_43(phi_inc_i_43),
	.phi_inc_i_44(phi_inc_i_44),
	.phi_inc_i_47(phi_inc_i_47),
	.phi_inc_i_31(phi_inc_i_31),
	.phi_inc_i_45(phi_inc_i_45),
	.phi_inc_i_46(phi_inc_i_46),
	.freq_mod_i_30(freq_mod_i_30),
	.phi_inc_i_30(phi_inc_i_30),
	.freq_mod_i_29(freq_mod_i_29),
	.phi_inc_i_29(phi_inc_i_29),
	.freq_mod_i_28(freq_mod_i_28),
	.phi_inc_i_28(phi_inc_i_28),
	.freq_mod_i_27(freq_mod_i_27),
	.phi_inc_i_27(phi_inc_i_27),
	.freq_mod_i_26(freq_mod_i_26),
	.phi_inc_i_26(phi_inc_i_26),
	.freq_mod_i_25(freq_mod_i_25),
	.phi_inc_i_25(phi_inc_i_25),
	.freq_mod_i_24(freq_mod_i_24),
	.phi_inc_i_24(phi_inc_i_24),
	.freq_mod_i_23(freq_mod_i_23),
	.phi_inc_i_23(phi_inc_i_23),
	.freq_mod_i_22(freq_mod_i_22),
	.phi_inc_i_22(phi_inc_i_22),
	.freq_mod_i_21(freq_mod_i_21),
	.phi_inc_i_21(phi_inc_i_21),
	.freq_mod_i_20(freq_mod_i_20),
	.phi_inc_i_20(phi_inc_i_20),
	.freq_mod_i_19(freq_mod_i_19),
	.phi_inc_i_19(phi_inc_i_19),
	.freq_mod_i_18(freq_mod_i_18),
	.phi_inc_i_18(phi_inc_i_18),
	.freq_mod_i_17(freq_mod_i_17),
	.phi_inc_i_17(phi_inc_i_17),
	.freq_mod_i_16(freq_mod_i_16),
	.phi_inc_i_16(phi_inc_i_16),
	.freq_mod_i_15(freq_mod_i_15),
	.phi_inc_i_15(phi_inc_i_15),
	.freq_mod_i_14(freq_mod_i_14),
	.phi_inc_i_14(phi_inc_i_14),
	.freq_mod_i_13(freq_mod_i_13),
	.phi_inc_i_13(phi_inc_i_13),
	.freq_mod_i_12(freq_mod_i_12),
	.phi_inc_i_12(phi_inc_i_12),
	.freq_mod_i_11(freq_mod_i_11),
	.phi_inc_i_11(phi_inc_i_11),
	.freq_mod_i_10(freq_mod_i_10),
	.phi_inc_i_10(phi_inc_i_10),
	.freq_mod_i_9(freq_mod_i_9),
	.phi_inc_i_9(phi_inc_i_9),
	.freq_mod_i_8(freq_mod_i_8),
	.phi_inc_i_8(phi_inc_i_8),
	.freq_mod_i_7(freq_mod_i_7),
	.phi_inc_i_7(phi_inc_i_7),
	.freq_mod_i_6(freq_mod_i_6),
	.phi_inc_i_6(phi_inc_i_6),
	.freq_mod_i_5(freq_mod_i_5),
	.phi_inc_i_5(phi_inc_i_5),
	.freq_mod_i_4(freq_mod_i_4),
	.phi_inc_i_4(phi_inc_i_4),
	.freq_mod_i_3(freq_mod_i_3),
	.phi_inc_i_3(phi_inc_i_3),
	.freq_mod_i_2(freq_mod_i_2),
	.phi_inc_i_2(phi_inc_i_2),
	.freq_mod_i_1(freq_mod_i_1),
	.phi_inc_i_1(phi_inc_i_1),
	.freq_mod_i_0(freq_mod_i_0),
	.phi_inc_i_0(phi_inc_i_0));

DDS_48_v1_asj_nco_isdr ux710isdr(
	.data_ready1(data_ready),
	.clk(clk),
	.reset_n(reset_n),
	.clken(clken));

DDS_48_v1_asj_nco_mob_rw_1 ux123(
	.data_out_0(data_out_01),
	.data_out_1(data_out_16),
	.data_out_2(data_out_21),
	.data_out_3(data_out_31),
	.data_out_4(data_out_41),
	.data_out_5(data_out_51),
	.data_out_6(data_out_61),
	.data_out_7(data_out_71),
	.data_out_8(data_out_81),
	.data_out_9(data_out_91),
	.data_out_10(data_out_101),
	.data_out_11(data_out_111),
	.data_out_12(data_out_121),
	.data_out_13(data_out_131),
	.data_out_14(data_out_141),
	.data_out_15(data_out_151),
	.ram_block1a64(\ux0121|altsyncram_component0|auto_generated|ram_block1a64~portadataout ),
	.ram_block1a80(\ux0121|altsyncram_component0|auto_generated|ram_block1a80~portadataout ),
	.ram_block1a96(\ux0121|altsyncram_component0|auto_generated|ram_block1a96~portadataout ),
	.ram_block1a112(\ux0121|altsyncram_component0|auto_generated|ram_block1a112~portadataout ),
	.ram_block1a32(\ux0121|altsyncram_component0|auto_generated|ram_block1a32~portadataout ),
	.ram_block1a48(\ux0121|altsyncram_component0|auto_generated|ram_block1a48~portadataout ),
	.ram_block1a0(\ux0121|altsyncram_component0|auto_generated|ram_block1a0~portadataout ),
	.ram_block1a16(\ux0121|altsyncram_component0|auto_generated|ram_block1a16~portadataout ),
	.ram_block1a65(\ux0121|altsyncram_component0|auto_generated|ram_block1a65~portadataout ),
	.ram_block1a81(\ux0121|altsyncram_component0|auto_generated|ram_block1a81~portadataout ),
	.ram_block1a97(\ux0121|altsyncram_component0|auto_generated|ram_block1a97~portadataout ),
	.ram_block1a113(\ux0121|altsyncram_component0|auto_generated|ram_block1a113~portadataout ),
	.ram_block1a33(\ux0121|altsyncram_component0|auto_generated|ram_block1a33~portadataout ),
	.ram_block1a49(\ux0121|altsyncram_component0|auto_generated|ram_block1a49~portadataout ),
	.ram_block1a1(\ux0121|altsyncram_component0|auto_generated|ram_block1a1~portadataout ),
	.ram_block1a17(\ux0121|altsyncram_component0|auto_generated|ram_block1a17~portadataout ),
	.ram_block1a66(\ux0121|altsyncram_component0|auto_generated|ram_block1a66~portadataout ),
	.ram_block1a82(\ux0121|altsyncram_component0|auto_generated|ram_block1a82~portadataout ),
	.ram_block1a98(\ux0121|altsyncram_component0|auto_generated|ram_block1a98~portadataout ),
	.ram_block1a114(\ux0121|altsyncram_component0|auto_generated|ram_block1a114~portadataout ),
	.ram_block1a34(\ux0121|altsyncram_component0|auto_generated|ram_block1a34~portadataout ),
	.ram_block1a50(\ux0121|altsyncram_component0|auto_generated|ram_block1a50~portadataout ),
	.ram_block1a2(\ux0121|altsyncram_component0|auto_generated|ram_block1a2~portadataout ),
	.ram_block1a18(\ux0121|altsyncram_component0|auto_generated|ram_block1a18~portadataout ),
	.ram_block1a67(\ux0121|altsyncram_component0|auto_generated|ram_block1a67~portadataout ),
	.ram_block1a83(\ux0121|altsyncram_component0|auto_generated|ram_block1a83~portadataout ),
	.ram_block1a99(\ux0121|altsyncram_component0|auto_generated|ram_block1a99~portadataout ),
	.ram_block1a115(\ux0121|altsyncram_component0|auto_generated|ram_block1a115~portadataout ),
	.ram_block1a35(\ux0121|altsyncram_component0|auto_generated|ram_block1a35~portadataout ),
	.ram_block1a51(\ux0121|altsyncram_component0|auto_generated|ram_block1a51~portadataout ),
	.ram_block1a3(\ux0121|altsyncram_component0|auto_generated|ram_block1a3~portadataout ),
	.ram_block1a19(\ux0121|altsyncram_component0|auto_generated|ram_block1a19~portadataout ),
	.ram_block1a68(\ux0121|altsyncram_component0|auto_generated|ram_block1a68~portadataout ),
	.ram_block1a84(\ux0121|altsyncram_component0|auto_generated|ram_block1a84~portadataout ),
	.ram_block1a100(\ux0121|altsyncram_component0|auto_generated|ram_block1a100~portadataout ),
	.ram_block1a116(\ux0121|altsyncram_component0|auto_generated|ram_block1a116~portadataout ),
	.ram_block1a36(\ux0121|altsyncram_component0|auto_generated|ram_block1a36~portadataout ),
	.ram_block1a52(\ux0121|altsyncram_component0|auto_generated|ram_block1a52~portadataout ),
	.ram_block1a4(\ux0121|altsyncram_component0|auto_generated|ram_block1a4~portadataout ),
	.ram_block1a20(\ux0121|altsyncram_component0|auto_generated|ram_block1a20~portadataout ),
	.ram_block1a69(\ux0121|altsyncram_component0|auto_generated|ram_block1a69~portadataout ),
	.ram_block1a85(\ux0121|altsyncram_component0|auto_generated|ram_block1a85~portadataout ),
	.ram_block1a101(\ux0121|altsyncram_component0|auto_generated|ram_block1a101~portadataout ),
	.ram_block1a117(\ux0121|altsyncram_component0|auto_generated|ram_block1a117~portadataout ),
	.ram_block1a37(\ux0121|altsyncram_component0|auto_generated|ram_block1a37~portadataout ),
	.ram_block1a53(\ux0121|altsyncram_component0|auto_generated|ram_block1a53~portadataout ),
	.ram_block1a5(\ux0121|altsyncram_component0|auto_generated|ram_block1a5~portadataout ),
	.ram_block1a21(\ux0121|altsyncram_component0|auto_generated|ram_block1a21~portadataout ),
	.ram_block1a70(\ux0121|altsyncram_component0|auto_generated|ram_block1a70~portadataout ),
	.ram_block1a86(\ux0121|altsyncram_component0|auto_generated|ram_block1a86~portadataout ),
	.ram_block1a102(\ux0121|altsyncram_component0|auto_generated|ram_block1a102~portadataout ),
	.ram_block1a118(\ux0121|altsyncram_component0|auto_generated|ram_block1a118~portadataout ),
	.ram_block1a38(\ux0121|altsyncram_component0|auto_generated|ram_block1a38~portadataout ),
	.ram_block1a54(\ux0121|altsyncram_component0|auto_generated|ram_block1a54~portadataout ),
	.ram_block1a6(\ux0121|altsyncram_component0|auto_generated|ram_block1a6~portadataout ),
	.ram_block1a22(\ux0121|altsyncram_component0|auto_generated|ram_block1a22~portadataout ),
	.ram_block1a71(\ux0121|altsyncram_component0|auto_generated|ram_block1a71~portadataout ),
	.ram_block1a87(\ux0121|altsyncram_component0|auto_generated|ram_block1a87~portadataout ),
	.ram_block1a103(\ux0121|altsyncram_component0|auto_generated|ram_block1a103~portadataout ),
	.ram_block1a119(\ux0121|altsyncram_component0|auto_generated|ram_block1a119~portadataout ),
	.ram_block1a39(\ux0121|altsyncram_component0|auto_generated|ram_block1a39~portadataout ),
	.ram_block1a55(\ux0121|altsyncram_component0|auto_generated|ram_block1a55~portadataout ),
	.ram_block1a7(\ux0121|altsyncram_component0|auto_generated|ram_block1a7~portadataout ),
	.ram_block1a23(\ux0121|altsyncram_component0|auto_generated|ram_block1a23~portadataout ),
	.ram_block1a72(\ux0121|altsyncram_component0|auto_generated|ram_block1a72~portadataout ),
	.ram_block1a88(\ux0121|altsyncram_component0|auto_generated|ram_block1a88~portadataout ),
	.ram_block1a104(\ux0121|altsyncram_component0|auto_generated|ram_block1a104~portadataout ),
	.ram_block1a120(\ux0121|altsyncram_component0|auto_generated|ram_block1a120~portadataout ),
	.ram_block1a40(\ux0121|altsyncram_component0|auto_generated|ram_block1a40~portadataout ),
	.ram_block1a56(\ux0121|altsyncram_component0|auto_generated|ram_block1a56~portadataout ),
	.ram_block1a8(\ux0121|altsyncram_component0|auto_generated|ram_block1a8~portadataout ),
	.ram_block1a24(\ux0121|altsyncram_component0|auto_generated|ram_block1a24~portadataout ),
	.ram_block1a73(\ux0121|altsyncram_component0|auto_generated|ram_block1a73~portadataout ),
	.ram_block1a89(\ux0121|altsyncram_component0|auto_generated|ram_block1a89~portadataout ),
	.ram_block1a105(\ux0121|altsyncram_component0|auto_generated|ram_block1a105~portadataout ),
	.ram_block1a121(\ux0121|altsyncram_component0|auto_generated|ram_block1a121~portadataout ),
	.ram_block1a41(\ux0121|altsyncram_component0|auto_generated|ram_block1a41~portadataout ),
	.ram_block1a57(\ux0121|altsyncram_component0|auto_generated|ram_block1a57~portadataout ),
	.ram_block1a9(\ux0121|altsyncram_component0|auto_generated|ram_block1a9~portadataout ),
	.ram_block1a25(\ux0121|altsyncram_component0|auto_generated|ram_block1a25~portadataout ),
	.ram_block1a74(\ux0121|altsyncram_component0|auto_generated|ram_block1a74~portadataout ),
	.ram_block1a90(\ux0121|altsyncram_component0|auto_generated|ram_block1a90~portadataout ),
	.ram_block1a106(\ux0121|altsyncram_component0|auto_generated|ram_block1a106~portadataout ),
	.ram_block1a122(\ux0121|altsyncram_component0|auto_generated|ram_block1a122~portadataout ),
	.ram_block1a42(\ux0121|altsyncram_component0|auto_generated|ram_block1a42~portadataout ),
	.ram_block1a58(\ux0121|altsyncram_component0|auto_generated|ram_block1a58~portadataout ),
	.ram_block1a10(\ux0121|altsyncram_component0|auto_generated|ram_block1a10~portadataout ),
	.ram_block1a26(\ux0121|altsyncram_component0|auto_generated|ram_block1a26~portadataout ),
	.ram_block1a75(\ux0121|altsyncram_component0|auto_generated|ram_block1a75~portadataout ),
	.ram_block1a91(\ux0121|altsyncram_component0|auto_generated|ram_block1a91~portadataout ),
	.ram_block1a107(\ux0121|altsyncram_component0|auto_generated|ram_block1a107~portadataout ),
	.ram_block1a123(\ux0121|altsyncram_component0|auto_generated|ram_block1a123~portadataout ),
	.ram_block1a43(\ux0121|altsyncram_component0|auto_generated|ram_block1a43~portadataout ),
	.ram_block1a59(\ux0121|altsyncram_component0|auto_generated|ram_block1a59~portadataout ),
	.ram_block1a11(\ux0121|altsyncram_component0|auto_generated|ram_block1a11~portadataout ),
	.ram_block1a27(\ux0121|altsyncram_component0|auto_generated|ram_block1a27~portadataout ),
	.ram_block1a76(\ux0121|altsyncram_component0|auto_generated|ram_block1a76~portadataout ),
	.ram_block1a92(\ux0121|altsyncram_component0|auto_generated|ram_block1a92~portadataout ),
	.ram_block1a108(\ux0121|altsyncram_component0|auto_generated|ram_block1a108~portadataout ),
	.ram_block1a124(\ux0121|altsyncram_component0|auto_generated|ram_block1a124~portadataout ),
	.ram_block1a44(\ux0121|altsyncram_component0|auto_generated|ram_block1a44~portadataout ),
	.ram_block1a60(\ux0121|altsyncram_component0|auto_generated|ram_block1a60~portadataout ),
	.ram_block1a12(\ux0121|altsyncram_component0|auto_generated|ram_block1a12~portadataout ),
	.ram_block1a28(\ux0121|altsyncram_component0|auto_generated|ram_block1a28~portadataout ),
	.ram_block1a77(\ux0121|altsyncram_component0|auto_generated|ram_block1a77~portadataout ),
	.ram_block1a93(\ux0121|altsyncram_component0|auto_generated|ram_block1a93~portadataout ),
	.ram_block1a109(\ux0121|altsyncram_component0|auto_generated|ram_block1a109~portadataout ),
	.ram_block1a125(\ux0121|altsyncram_component0|auto_generated|ram_block1a125~portadataout ),
	.ram_block1a45(\ux0121|altsyncram_component0|auto_generated|ram_block1a45~portadataout ),
	.ram_block1a61(\ux0121|altsyncram_component0|auto_generated|ram_block1a61~portadataout ),
	.ram_block1a13(\ux0121|altsyncram_component0|auto_generated|ram_block1a13~portadataout ),
	.ram_block1a29(\ux0121|altsyncram_component0|auto_generated|ram_block1a29~portadataout ),
	.ram_block1a78(\ux0121|altsyncram_component0|auto_generated|ram_block1a78~portadataout ),
	.ram_block1a94(\ux0121|altsyncram_component0|auto_generated|ram_block1a94~portadataout ),
	.ram_block1a110(\ux0121|altsyncram_component0|auto_generated|ram_block1a110~portadataout ),
	.ram_block1a126(\ux0121|altsyncram_component0|auto_generated|ram_block1a126~portadataout ),
	.ram_block1a46(\ux0121|altsyncram_component0|auto_generated|ram_block1a46~portadataout ),
	.ram_block1a62(\ux0121|altsyncram_component0|auto_generated|ram_block1a62~portadataout ),
	.ram_block1a14(\ux0121|altsyncram_component0|auto_generated|ram_block1a14~portadataout ),
	.ram_block1a30(\ux0121|altsyncram_component0|auto_generated|ram_block1a30~portadataout ),
	.ram_block1a79(\ux0121|altsyncram_component0|auto_generated|ram_block1a79~portadataout ),
	.ram_block1a95(\ux0121|altsyncram_component0|auto_generated|ram_block1a95~portadataout ),
	.ram_block1a111(\ux0121|altsyncram_component0|auto_generated|ram_block1a111~portadataout ),
	.ram_block1a127(\ux0121|altsyncram_component0|auto_generated|ram_block1a127~portadataout ),
	.ram_block1a47(\ux0121|altsyncram_component0|auto_generated|ram_block1a47~portadataout ),
	.ram_block1a63(\ux0121|altsyncram_component0|auto_generated|ram_block1a63~portadataout ),
	.ram_block1a15(\ux0121|altsyncram_component0|auto_generated|ram_block1a15~portadataout ),
	.ram_block1a31(\ux0121|altsyncram_component0|auto_generated|ram_block1a31~portadataout ),
	.out_address_reg_a_2(\ux0120|altsyncram_component0|auto_generated|out_address_reg_a[2]~q ),
	.out_address_reg_a_0(\ux0120|altsyncram_component0|auto_generated|out_address_reg_a[0]~q ),
	.out_address_reg_a_1(\ux0120|altsyncram_component0|auto_generated|out_address_reg_a[1]~q ),
	.data_out_121(\ux122|data_out[12]~3_combout ),
	.clk(clk),
	.reset_n(reset_n));

DDS_48_v1_asj_nco_mob_rw ux122(
	.data_out_0(data_out_0),
	.data_out_1(data_out_1),
	.data_out_2(data_out_2),
	.data_out_3(data_out_3),
	.data_out_4(data_out_4),
	.data_out_5(data_out_5),
	.data_out_6(data_out_6),
	.data_out_7(data_out_7),
	.data_out_8(data_out_8),
	.data_out_9(data_out_9),
	.data_out_10(data_out_10),
	.data_out_11(data_out_11),
	.data_out_12(data_out_12),
	.data_out_13(data_out_13),
	.data_out_14(data_out_14),
	.data_out_15(data_out_15),
	.ram_block1a64(\ux0120|altsyncram_component0|auto_generated|ram_block1a64~portadataout ),
	.ram_block1a80(\ux0120|altsyncram_component0|auto_generated|ram_block1a80~portadataout ),
	.ram_block1a96(\ux0120|altsyncram_component0|auto_generated|ram_block1a96~portadataout ),
	.ram_block1a112(\ux0120|altsyncram_component0|auto_generated|ram_block1a112~portadataout ),
	.ram_block1a32(\ux0120|altsyncram_component0|auto_generated|ram_block1a32~portadataout ),
	.ram_block1a48(\ux0120|altsyncram_component0|auto_generated|ram_block1a48~portadataout ),
	.ram_block1a0(\ux0120|altsyncram_component0|auto_generated|ram_block1a0~portadataout ),
	.ram_block1a16(\ux0120|altsyncram_component0|auto_generated|ram_block1a16~portadataout ),
	.ram_block1a65(\ux0120|altsyncram_component0|auto_generated|ram_block1a65~portadataout ),
	.ram_block1a81(\ux0120|altsyncram_component0|auto_generated|ram_block1a81~portadataout ),
	.ram_block1a97(\ux0120|altsyncram_component0|auto_generated|ram_block1a97~portadataout ),
	.ram_block1a113(\ux0120|altsyncram_component0|auto_generated|ram_block1a113~portadataout ),
	.ram_block1a33(\ux0120|altsyncram_component0|auto_generated|ram_block1a33~portadataout ),
	.ram_block1a49(\ux0120|altsyncram_component0|auto_generated|ram_block1a49~portadataout ),
	.ram_block1a1(\ux0120|altsyncram_component0|auto_generated|ram_block1a1~portadataout ),
	.ram_block1a17(\ux0120|altsyncram_component0|auto_generated|ram_block1a17~portadataout ),
	.ram_block1a66(\ux0120|altsyncram_component0|auto_generated|ram_block1a66~portadataout ),
	.ram_block1a82(\ux0120|altsyncram_component0|auto_generated|ram_block1a82~portadataout ),
	.ram_block1a98(\ux0120|altsyncram_component0|auto_generated|ram_block1a98~portadataout ),
	.ram_block1a114(\ux0120|altsyncram_component0|auto_generated|ram_block1a114~portadataout ),
	.ram_block1a34(\ux0120|altsyncram_component0|auto_generated|ram_block1a34~portadataout ),
	.ram_block1a50(\ux0120|altsyncram_component0|auto_generated|ram_block1a50~portadataout ),
	.ram_block1a2(\ux0120|altsyncram_component0|auto_generated|ram_block1a2~portadataout ),
	.ram_block1a18(\ux0120|altsyncram_component0|auto_generated|ram_block1a18~portadataout ),
	.ram_block1a67(\ux0120|altsyncram_component0|auto_generated|ram_block1a67~portadataout ),
	.ram_block1a83(\ux0120|altsyncram_component0|auto_generated|ram_block1a83~portadataout ),
	.ram_block1a99(\ux0120|altsyncram_component0|auto_generated|ram_block1a99~portadataout ),
	.ram_block1a115(\ux0120|altsyncram_component0|auto_generated|ram_block1a115~portadataout ),
	.ram_block1a35(\ux0120|altsyncram_component0|auto_generated|ram_block1a35~portadataout ),
	.ram_block1a51(\ux0120|altsyncram_component0|auto_generated|ram_block1a51~portadataout ),
	.ram_block1a3(\ux0120|altsyncram_component0|auto_generated|ram_block1a3~portadataout ),
	.ram_block1a19(\ux0120|altsyncram_component0|auto_generated|ram_block1a19~portadataout ),
	.ram_block1a68(\ux0120|altsyncram_component0|auto_generated|ram_block1a68~portadataout ),
	.ram_block1a84(\ux0120|altsyncram_component0|auto_generated|ram_block1a84~portadataout ),
	.ram_block1a100(\ux0120|altsyncram_component0|auto_generated|ram_block1a100~portadataout ),
	.ram_block1a116(\ux0120|altsyncram_component0|auto_generated|ram_block1a116~portadataout ),
	.ram_block1a36(\ux0120|altsyncram_component0|auto_generated|ram_block1a36~portadataout ),
	.ram_block1a52(\ux0120|altsyncram_component0|auto_generated|ram_block1a52~portadataout ),
	.ram_block1a4(\ux0120|altsyncram_component0|auto_generated|ram_block1a4~portadataout ),
	.ram_block1a20(\ux0120|altsyncram_component0|auto_generated|ram_block1a20~portadataout ),
	.ram_block1a69(\ux0120|altsyncram_component0|auto_generated|ram_block1a69~portadataout ),
	.ram_block1a85(\ux0120|altsyncram_component0|auto_generated|ram_block1a85~portadataout ),
	.ram_block1a101(\ux0120|altsyncram_component0|auto_generated|ram_block1a101~portadataout ),
	.ram_block1a117(\ux0120|altsyncram_component0|auto_generated|ram_block1a117~portadataout ),
	.ram_block1a37(\ux0120|altsyncram_component0|auto_generated|ram_block1a37~portadataout ),
	.ram_block1a53(\ux0120|altsyncram_component0|auto_generated|ram_block1a53~portadataout ),
	.ram_block1a5(\ux0120|altsyncram_component0|auto_generated|ram_block1a5~portadataout ),
	.ram_block1a21(\ux0120|altsyncram_component0|auto_generated|ram_block1a21~portadataout ),
	.ram_block1a70(\ux0120|altsyncram_component0|auto_generated|ram_block1a70~portadataout ),
	.ram_block1a86(\ux0120|altsyncram_component0|auto_generated|ram_block1a86~portadataout ),
	.ram_block1a102(\ux0120|altsyncram_component0|auto_generated|ram_block1a102~portadataout ),
	.ram_block1a118(\ux0120|altsyncram_component0|auto_generated|ram_block1a118~portadataout ),
	.ram_block1a38(\ux0120|altsyncram_component0|auto_generated|ram_block1a38~portadataout ),
	.ram_block1a54(\ux0120|altsyncram_component0|auto_generated|ram_block1a54~portadataout ),
	.ram_block1a6(\ux0120|altsyncram_component0|auto_generated|ram_block1a6~portadataout ),
	.ram_block1a22(\ux0120|altsyncram_component0|auto_generated|ram_block1a22~portadataout ),
	.ram_block1a71(\ux0120|altsyncram_component0|auto_generated|ram_block1a71~portadataout ),
	.ram_block1a87(\ux0120|altsyncram_component0|auto_generated|ram_block1a87~portadataout ),
	.ram_block1a103(\ux0120|altsyncram_component0|auto_generated|ram_block1a103~portadataout ),
	.ram_block1a119(\ux0120|altsyncram_component0|auto_generated|ram_block1a119~portadataout ),
	.ram_block1a39(\ux0120|altsyncram_component0|auto_generated|ram_block1a39~portadataout ),
	.ram_block1a55(\ux0120|altsyncram_component0|auto_generated|ram_block1a55~portadataout ),
	.ram_block1a7(\ux0120|altsyncram_component0|auto_generated|ram_block1a7~portadataout ),
	.ram_block1a23(\ux0120|altsyncram_component0|auto_generated|ram_block1a23~portadataout ),
	.ram_block1a72(\ux0120|altsyncram_component0|auto_generated|ram_block1a72~portadataout ),
	.ram_block1a88(\ux0120|altsyncram_component0|auto_generated|ram_block1a88~portadataout ),
	.ram_block1a104(\ux0120|altsyncram_component0|auto_generated|ram_block1a104~portadataout ),
	.ram_block1a120(\ux0120|altsyncram_component0|auto_generated|ram_block1a120~portadataout ),
	.ram_block1a40(\ux0120|altsyncram_component0|auto_generated|ram_block1a40~portadataout ),
	.ram_block1a56(\ux0120|altsyncram_component0|auto_generated|ram_block1a56~portadataout ),
	.ram_block1a8(\ux0120|altsyncram_component0|auto_generated|ram_block1a8~portadataout ),
	.ram_block1a24(\ux0120|altsyncram_component0|auto_generated|ram_block1a24~portadataout ),
	.ram_block1a73(\ux0120|altsyncram_component0|auto_generated|ram_block1a73~portadataout ),
	.ram_block1a89(\ux0120|altsyncram_component0|auto_generated|ram_block1a89~portadataout ),
	.ram_block1a105(\ux0120|altsyncram_component0|auto_generated|ram_block1a105~portadataout ),
	.ram_block1a121(\ux0120|altsyncram_component0|auto_generated|ram_block1a121~portadataout ),
	.ram_block1a41(\ux0120|altsyncram_component0|auto_generated|ram_block1a41~portadataout ),
	.ram_block1a57(\ux0120|altsyncram_component0|auto_generated|ram_block1a57~portadataout ),
	.ram_block1a9(\ux0120|altsyncram_component0|auto_generated|ram_block1a9~portadataout ),
	.ram_block1a25(\ux0120|altsyncram_component0|auto_generated|ram_block1a25~portadataout ),
	.ram_block1a74(\ux0120|altsyncram_component0|auto_generated|ram_block1a74~portadataout ),
	.ram_block1a90(\ux0120|altsyncram_component0|auto_generated|ram_block1a90~portadataout ),
	.ram_block1a106(\ux0120|altsyncram_component0|auto_generated|ram_block1a106~portadataout ),
	.ram_block1a122(\ux0120|altsyncram_component0|auto_generated|ram_block1a122~portadataout ),
	.ram_block1a42(\ux0120|altsyncram_component0|auto_generated|ram_block1a42~portadataout ),
	.ram_block1a58(\ux0120|altsyncram_component0|auto_generated|ram_block1a58~portadataout ),
	.ram_block1a10(\ux0120|altsyncram_component0|auto_generated|ram_block1a10~portadataout ),
	.ram_block1a26(\ux0120|altsyncram_component0|auto_generated|ram_block1a26~portadataout ),
	.ram_block1a75(\ux0120|altsyncram_component0|auto_generated|ram_block1a75~portadataout ),
	.ram_block1a91(\ux0120|altsyncram_component0|auto_generated|ram_block1a91~portadataout ),
	.ram_block1a107(\ux0120|altsyncram_component0|auto_generated|ram_block1a107~portadataout ),
	.ram_block1a123(\ux0120|altsyncram_component0|auto_generated|ram_block1a123~portadataout ),
	.ram_block1a43(\ux0120|altsyncram_component0|auto_generated|ram_block1a43~portadataout ),
	.ram_block1a59(\ux0120|altsyncram_component0|auto_generated|ram_block1a59~portadataout ),
	.ram_block1a11(\ux0120|altsyncram_component0|auto_generated|ram_block1a11~portadataout ),
	.ram_block1a27(\ux0120|altsyncram_component0|auto_generated|ram_block1a27~portadataout ),
	.ram_block1a76(\ux0120|altsyncram_component0|auto_generated|ram_block1a76~portadataout ),
	.ram_block1a92(\ux0120|altsyncram_component0|auto_generated|ram_block1a92~portadataout ),
	.ram_block1a108(\ux0120|altsyncram_component0|auto_generated|ram_block1a108~portadataout ),
	.ram_block1a124(\ux0120|altsyncram_component0|auto_generated|ram_block1a124~portadataout ),
	.ram_block1a44(\ux0120|altsyncram_component0|auto_generated|ram_block1a44~portadataout ),
	.ram_block1a60(\ux0120|altsyncram_component0|auto_generated|ram_block1a60~portadataout ),
	.ram_block1a12(\ux0120|altsyncram_component0|auto_generated|ram_block1a12~portadataout ),
	.ram_block1a28(\ux0120|altsyncram_component0|auto_generated|ram_block1a28~portadataout ),
	.ram_block1a77(\ux0120|altsyncram_component0|auto_generated|ram_block1a77~portadataout ),
	.ram_block1a93(\ux0120|altsyncram_component0|auto_generated|ram_block1a93~portadataout ),
	.ram_block1a109(\ux0120|altsyncram_component0|auto_generated|ram_block1a109~portadataout ),
	.ram_block1a125(\ux0120|altsyncram_component0|auto_generated|ram_block1a125~portadataout ),
	.ram_block1a45(\ux0120|altsyncram_component0|auto_generated|ram_block1a45~portadataout ),
	.ram_block1a61(\ux0120|altsyncram_component0|auto_generated|ram_block1a61~portadataout ),
	.ram_block1a13(\ux0120|altsyncram_component0|auto_generated|ram_block1a13~portadataout ),
	.ram_block1a29(\ux0120|altsyncram_component0|auto_generated|ram_block1a29~portadataout ),
	.ram_block1a78(\ux0120|altsyncram_component0|auto_generated|ram_block1a78~portadataout ),
	.ram_block1a94(\ux0120|altsyncram_component0|auto_generated|ram_block1a94~portadataout ),
	.ram_block1a110(\ux0120|altsyncram_component0|auto_generated|ram_block1a110~portadataout ),
	.ram_block1a126(\ux0120|altsyncram_component0|auto_generated|ram_block1a126~portadataout ),
	.ram_block1a46(\ux0120|altsyncram_component0|auto_generated|ram_block1a46~portadataout ),
	.ram_block1a62(\ux0120|altsyncram_component0|auto_generated|ram_block1a62~portadataout ),
	.ram_block1a14(\ux0120|altsyncram_component0|auto_generated|ram_block1a14~portadataout ),
	.ram_block1a30(\ux0120|altsyncram_component0|auto_generated|ram_block1a30~portadataout ),
	.ram_block1a79(\ux0120|altsyncram_component0|auto_generated|ram_block1a79~portadataout ),
	.ram_block1a95(\ux0120|altsyncram_component0|auto_generated|ram_block1a95~portadataout ),
	.ram_block1a111(\ux0120|altsyncram_component0|auto_generated|ram_block1a111~portadataout ),
	.ram_block1a127(\ux0120|altsyncram_component0|auto_generated|ram_block1a127~portadataout ),
	.ram_block1a47(\ux0120|altsyncram_component0|auto_generated|ram_block1a47~portadataout ),
	.ram_block1a63(\ux0120|altsyncram_component0|auto_generated|ram_block1a63~portadataout ),
	.ram_block1a15(\ux0120|altsyncram_component0|auto_generated|ram_block1a15~portadataout ),
	.ram_block1a31(\ux0120|altsyncram_component0|auto_generated|ram_block1a31~portadataout ),
	.out_address_reg_a_2(\ux0120|altsyncram_component0|auto_generated|out_address_reg_a[2]~q ),
	.out_address_reg_a_0(\ux0120|altsyncram_component0|auto_generated|out_address_reg_a[0]~q ),
	.out_address_reg_a_1(\ux0120|altsyncram_component0|auto_generated|out_address_reg_a[1]~q ),
	.data_out_121(\ux122|data_out[12]~3_combout ),
	.clk(clk),
	.reset_n(reset_n),
	.clken(clken));

DDS_48_v1_asj_dxx ux002(
	.dxxpdo_5(\ux002|dxxpdo[5]~q ),
	.dxxpdo_6(\ux002|dxxpdo[6]~q ),
	.dxxpdo_7(\ux002|dxxpdo[7]~q ),
	.dxxpdo_8(\ux002|dxxpdo[8]~q ),
	.dxxpdo_9(\ux002|dxxpdo[9]~q ),
	.dxxpdo_10(\ux002|dxxpdo[10]~q ),
	.dxxpdo_11(\ux002|dxxpdo[11]~q ),
	.dxxpdo_12(\ux002|dxxpdo[12]~q ),
	.dxxpdo_13(\ux002|dxxpdo[13]~q ),
	.dxxpdo_14(\ux002|dxxpdo[14]~q ),
	.dxxpdo_15(\ux002|dxxpdo[15]~q ),
	.dxxpdo_16(\ux002|dxxpdo[16]~q ),
	.dxxpdo_17(\ux002|dxxpdo[17]~q ),
	.dxxpdo_20(\ux002|dxxpdo[20]~q ),
	.dxxpdo_18(\ux002|dxxpdo[18]~q ),
	.dxxpdo_19(\ux002|dxxpdo[19]~q ),
	.dxxrv_5(\ux001|dxxrv[5]~q ),
	.dxxrv_6(\ux001|dxxrv[6]~q ),
	.dxxrv_7(\ux001|dxxrv[7]~q ),
	.dxxrv_8(\ux001|dxxrv[8]~q ),
	.dxxrv_9(\ux001|dxxrv[9]~q ),
	.dxxrv_4(\ux001|dxxrv[4]~q ),
	.dxxrv_3(\ux001|dxxrv[3]~q ),
	.dxxrv_2(\ux001|dxxrv[2]~q ),
	.dxxrv_1(\ux001|dxxrv[1]~q ),
	.dxxrv_0(\ux001|dxxrv[0]~q ),
	.data_out_12(\ux122|data_out[12]~3_combout ),
	.pipeline_dffe_32(\ux000|acc|auto_generated|pipeline_dffe[32]~q ),
	.pipeline_dffe_33(\ux000|acc|auto_generated|pipeline_dffe[33]~q ),
	.pipeline_dffe_34(\ux000|acc|auto_generated|pipeline_dffe[34]~q ),
	.pipeline_dffe_35(\ux000|acc|auto_generated|pipeline_dffe[35]~q ),
	.pipeline_dffe_36(\ux000|acc|auto_generated|pipeline_dffe[36]~q ),
	.pipeline_dffe_37(\ux000|acc|auto_generated|pipeline_dffe[37]~q ),
	.pipeline_dffe_38(\ux000|acc|auto_generated|pipeline_dffe[38]~q ),
	.pipeline_dffe_39(\ux000|acc|auto_generated|pipeline_dffe[39]~q ),
	.pipeline_dffe_40(\ux000|acc|auto_generated|pipeline_dffe[40]~q ),
	.pipeline_dffe_41(\ux000|acc|auto_generated|pipeline_dffe[41]~q ),
	.pipeline_dffe_42(\ux000|acc|auto_generated|pipeline_dffe[42]~q ),
	.pipeline_dffe_43(\ux000|acc|auto_generated|pipeline_dffe[43]~q ),
	.pipeline_dffe_44(\ux000|acc|auto_generated|pipeline_dffe[44]~q ),
	.pipeline_dffe_47(\ux000|acc|auto_generated|pipeline_dffe[47]~q ),
	.pipeline_dffe_31(\ux000|acc|auto_generated|pipeline_dffe[31]~q ),
	.pipeline_dffe_45(\ux000|acc|auto_generated|pipeline_dffe[45]~q ),
	.pipeline_dffe_46(\ux000|acc|auto_generated|pipeline_dffe[46]~q ),
	.pipeline_dffe_30(\ux000|acc|auto_generated|pipeline_dffe[30]~q ),
	.pipeline_dffe_29(\ux000|acc|auto_generated|pipeline_dffe[29]~q ),
	.pipeline_dffe_28(\ux000|acc|auto_generated|pipeline_dffe[28]~q ),
	.pipeline_dffe_27(\ux000|acc|auto_generated|pipeline_dffe[27]~q ),
	.clk(clk),
	.reset_n(reset_n));

DDS_48_v1_asj_dxx_g ux001(
	.dxxrv_5(\ux001|dxxrv[5]~q ),
	.dxxrv_6(\ux001|dxxrv[6]~q ),
	.dxxrv_7(\ux001|dxxrv[7]~q ),
	.dxxrv_8(\ux001|dxxrv[8]~q ),
	.dxxrv_9(\ux001|dxxrv[9]~q ),
	.dxxrv_4(\ux001|dxxrv[4]~q ),
	.dxxrv_3(\ux001|dxxrv[3]~q ),
	.dxxrv_2(\ux001|dxxrv[2]~q ),
	.dxxrv_1(\ux001|dxxrv[1]~q ),
	.dxxrv_0(\ux001|dxxrv[0]~q ),
	.data_out_12(\ux122|data_out[12]~3_combout ),
	.clk(clk),
	.reset_n(reset_n));

DDS_48_v1_asj_altqmcpipe ux000(
	.data_out_12(\ux122|data_out[12]~3_combout ),
	.pipeline_dffe_32(\ux000|acc|auto_generated|pipeline_dffe[32]~q ),
	.pipeline_dffe_33(\ux000|acc|auto_generated|pipeline_dffe[33]~q ),
	.pipeline_dffe_34(\ux000|acc|auto_generated|pipeline_dffe[34]~q ),
	.pipeline_dffe_35(\ux000|acc|auto_generated|pipeline_dffe[35]~q ),
	.pipeline_dffe_36(\ux000|acc|auto_generated|pipeline_dffe[36]~q ),
	.pipeline_dffe_37(\ux000|acc|auto_generated|pipeline_dffe[37]~q ),
	.pipeline_dffe_38(\ux000|acc|auto_generated|pipeline_dffe[38]~q ),
	.pipeline_dffe_39(\ux000|acc|auto_generated|pipeline_dffe[39]~q ),
	.pipeline_dffe_40(\ux000|acc|auto_generated|pipeline_dffe[40]~q ),
	.pipeline_dffe_41(\ux000|acc|auto_generated|pipeline_dffe[41]~q ),
	.pipeline_dffe_42(\ux000|acc|auto_generated|pipeline_dffe[42]~q ),
	.pipeline_dffe_43(\ux000|acc|auto_generated|pipeline_dffe[43]~q ),
	.pipeline_dffe_44(\ux000|acc|auto_generated|pipeline_dffe[44]~q ),
	.pipeline_dffe_47(\ux000|acc|auto_generated|pipeline_dffe[47]~q ),
	.pipeline_dffe_31(\ux000|acc|auto_generated|pipeline_dffe[31]~q ),
	.pipeline_dffe_45(\ux000|acc|auto_generated|pipeline_dffe[45]~q ),
	.pipeline_dffe_46(\ux000|acc|auto_generated|pipeline_dffe[46]~q ),
	.pipeline_dffe_30(\ux000|acc|auto_generated|pipeline_dffe[30]~q ),
	.pipeline_dffe_321(\ux003|acc|auto_generated|pipeline_dffe[32]~q ),
	.pipeline_dffe_29(\ux000|acc|auto_generated|pipeline_dffe[29]~q ),
	.pipeline_dffe_331(\ux003|acc|auto_generated|pipeline_dffe[33]~q ),
	.pipeline_dffe_341(\ux003|acc|auto_generated|pipeline_dffe[34]~q ),
	.pipeline_dffe_351(\ux003|acc|auto_generated|pipeline_dffe[35]~q ),
	.pipeline_dffe_361(\ux003|acc|auto_generated|pipeline_dffe[36]~q ),
	.pipeline_dffe_371(\ux003|acc|auto_generated|pipeline_dffe[37]~q ),
	.pipeline_dffe_381(\ux003|acc|auto_generated|pipeline_dffe[38]~q ),
	.pipeline_dffe_391(\ux003|acc|auto_generated|pipeline_dffe[39]~q ),
	.pipeline_dffe_401(\ux003|acc|auto_generated|pipeline_dffe[40]~q ),
	.pipeline_dffe_411(\ux003|acc|auto_generated|pipeline_dffe[41]~q ),
	.pipeline_dffe_421(\ux003|acc|auto_generated|pipeline_dffe[42]~q ),
	.pipeline_dffe_431(\ux003|acc|auto_generated|pipeline_dffe[43]~q ),
	.pipeline_dffe_441(\ux003|acc|auto_generated|pipeline_dffe[44]~q ),
	.pipeline_dffe_471(\ux003|acc|auto_generated|pipeline_dffe[47]~q ),
	.pipeline_dffe_311(\ux003|acc|auto_generated|pipeline_dffe[31]~q ),
	.pipeline_dffe_28(\ux000|acc|auto_generated|pipeline_dffe[28]~q ),
	.pipeline_dffe_451(\ux003|acc|auto_generated|pipeline_dffe[45]~q ),
	.pipeline_dffe_461(\ux003|acc|auto_generated|pipeline_dffe[46]~q ),
	.pipeline_dffe_301(\ux003|acc|auto_generated|pipeline_dffe[30]~q ),
	.pipeline_dffe_27(\ux000|acc|auto_generated|pipeline_dffe[27]~q ),
	.pipeline_dffe_291(\ux003|acc|auto_generated|pipeline_dffe[29]~q ),
	.pipeline_dffe_281(\ux003|acc|auto_generated|pipeline_dffe[28]~q ),
	.pipeline_dffe_271(\ux003|acc|auto_generated|pipeline_dffe[27]~q ),
	.pipeline_dffe_26(\ux003|acc|auto_generated|pipeline_dffe[26]~q ),
	.pipeline_dffe_25(\ux003|acc|auto_generated|pipeline_dffe[25]~q ),
	.pipeline_dffe_24(\ux003|acc|auto_generated|pipeline_dffe[24]~q ),
	.pipeline_dffe_23(\ux003|acc|auto_generated|pipeline_dffe[23]~q ),
	.pipeline_dffe_22(\ux003|acc|auto_generated|pipeline_dffe[22]~q ),
	.pipeline_dffe_21(\ux003|acc|auto_generated|pipeline_dffe[21]~q ),
	.pipeline_dffe_20(\ux003|acc|auto_generated|pipeline_dffe[20]~q ),
	.pipeline_dffe_19(\ux003|acc|auto_generated|pipeline_dffe[19]~q ),
	.pipeline_dffe_18(\ux003|acc|auto_generated|pipeline_dffe[18]~q ),
	.pipeline_dffe_17(\ux003|acc|auto_generated|pipeline_dffe[17]~q ),
	.pipeline_dffe_16(\ux003|acc|auto_generated|pipeline_dffe[16]~q ),
	.pipeline_dffe_15(\ux003|acc|auto_generated|pipeline_dffe[15]~q ),
	.pipeline_dffe_14(\ux003|acc|auto_generated|pipeline_dffe[14]~q ),
	.pipeline_dffe_13(\ux003|acc|auto_generated|pipeline_dffe[13]~q ),
	.pipeline_dffe_12(\ux003|acc|auto_generated|pipeline_dffe[12]~q ),
	.pipeline_dffe_11(\ux003|acc|auto_generated|pipeline_dffe[11]~q ),
	.pipeline_dffe_10(\ux003|acc|auto_generated|pipeline_dffe[10]~q ),
	.pipeline_dffe_9(\ux003|acc|auto_generated|pipeline_dffe[9]~q ),
	.pipeline_dffe_8(\ux003|acc|auto_generated|pipeline_dffe[8]~q ),
	.pipeline_dffe_7(\ux003|acc|auto_generated|pipeline_dffe[7]~q ),
	.pipeline_dffe_6(\ux003|acc|auto_generated|pipeline_dffe[6]~q ),
	.pipeline_dffe_5(\ux003|acc|auto_generated|pipeline_dffe[5]~q ),
	.pipeline_dffe_4(\ux003|acc|auto_generated|pipeline_dffe[4]~q ),
	.pipeline_dffe_3(\ux003|acc|auto_generated|pipeline_dffe[3]~q ),
	.pipeline_dffe_2(\ux003|acc|auto_generated|pipeline_dffe[2]~q ),
	.pipeline_dffe_1(\ux003|acc|auto_generated|pipeline_dffe[1]~q ),
	.pipeline_dffe_0(\ux003|acc|auto_generated|pipeline_dffe[0]~q ),
	.clk(clk),
	.reset_n(reset_n),
	.clken(clken));

DDS_48_v1_asj_gal ux009(
	.rom_add_0(\ux009|rom_add[0]~q ),
	.rom_add_1(\ux009|rom_add[1]~q ),
	.rom_add_2(\ux009|rom_add[2]~q ),
	.rom_add_3(\ux009|rom_add[3]~q ),
	.rom_add_4(\ux009|rom_add[4]~q ),
	.rom_add_5(\ux009|rom_add[5]~q ),
	.rom_add_6(\ux009|rom_add[6]~q ),
	.rom_add_7(\ux009|rom_add[7]~q ),
	.rom_add_8(\ux009|rom_add[8]~q ),
	.rom_add_9(\ux009|rom_add[9]~q ),
	.rom_add_10(\ux009|rom_add[10]~q ),
	.rom_add_11(\ux009|rom_add[11]~q ),
	.rom_add_12(\ux009|rom_add[12]~q ),
	.rom_add_15(\ux009|rom_add[15]~q ),
	.rom_add_13(\ux009|rom_add[13]~q ),
	.rom_add_14(\ux009|rom_add[14]~q ),
	.data_out_12(\ux122|data_out[12]~3_combout ),
	.pipeline_dffe_0(\ux004|acc|auto_generated|pipeline_dffe[0]~q ),
	.pipeline_dffe_1(\ux004|acc|auto_generated|pipeline_dffe[1]~q ),
	.pipeline_dffe_2(\ux004|acc|auto_generated|pipeline_dffe[2]~q ),
	.pipeline_dffe_3(\ux004|acc|auto_generated|pipeline_dffe[3]~q ),
	.pipeline_dffe_4(\ux004|acc|auto_generated|pipeline_dffe[4]~q ),
	.pipeline_dffe_5(\ux004|acc|auto_generated|pipeline_dffe[5]~q ),
	.pipeline_dffe_6(\ux004|acc|auto_generated|pipeline_dffe[6]~q ),
	.pipeline_dffe_7(\ux004|acc|auto_generated|pipeline_dffe[7]~q ),
	.pipeline_dffe_8(\ux004|acc|auto_generated|pipeline_dffe[8]~q ),
	.pipeline_dffe_9(\ux004|acc|auto_generated|pipeline_dffe[9]~q ),
	.pipeline_dffe_10(\ux004|acc|auto_generated|pipeline_dffe[10]~q ),
	.pipeline_dffe_11(\ux004|acc|auto_generated|pipeline_dffe[11]~q ),
	.pipeline_dffe_12(\ux004|acc|auto_generated|pipeline_dffe[12]~q ),
	.pipeline_dffe_15(\ux004|acc|auto_generated|pipeline_dffe[15]~q ),
	.pipeline_dffe_13(\ux004|acc|auto_generated|pipeline_dffe[13]~q ),
	.pipeline_dffe_14(\ux004|acc|auto_generated|pipeline_dffe[14]~q ),
	.clk(clk),
	.reset_n(reset_n));

DDS_48_v1_asj_nco_pxx ux004(
	.dxxpdo_5(\ux002|dxxpdo[5]~q ),
	.dxxpdo_6(\ux002|dxxpdo[6]~q ),
	.dxxpdo_7(\ux002|dxxpdo[7]~q ),
	.dxxpdo_8(\ux002|dxxpdo[8]~q ),
	.dxxpdo_9(\ux002|dxxpdo[9]~q ),
	.dxxpdo_10(\ux002|dxxpdo[10]~q ),
	.dxxpdo_11(\ux002|dxxpdo[11]~q ),
	.dxxpdo_12(\ux002|dxxpdo[12]~q ),
	.dxxpdo_13(\ux002|dxxpdo[13]~q ),
	.dxxpdo_14(\ux002|dxxpdo[14]~q ),
	.dxxpdo_15(\ux002|dxxpdo[15]~q ),
	.dxxpdo_16(\ux002|dxxpdo[16]~q ),
	.dxxpdo_17(\ux002|dxxpdo[17]~q ),
	.dxxpdo_20(\ux002|dxxpdo[20]~q ),
	.dxxpdo_18(\ux002|dxxpdo[18]~q ),
	.dxxpdo_19(\ux002|dxxpdo[19]~q ),
	.data_out_12(\ux122|data_out[12]~3_combout ),
	.pipeline_dffe_0(\ux004|acc|auto_generated|pipeline_dffe[0]~q ),
	.pipeline_dffe_1(\ux004|acc|auto_generated|pipeline_dffe[1]~q ),
	.pipeline_dffe_2(\ux004|acc|auto_generated|pipeline_dffe[2]~q ),
	.pipeline_dffe_3(\ux004|acc|auto_generated|pipeline_dffe[3]~q ),
	.pipeline_dffe_4(\ux004|acc|auto_generated|pipeline_dffe[4]~q ),
	.pipeline_dffe_5(\ux004|acc|auto_generated|pipeline_dffe[5]~q ),
	.pipeline_dffe_6(\ux004|acc|auto_generated|pipeline_dffe[6]~q ),
	.pipeline_dffe_7(\ux004|acc|auto_generated|pipeline_dffe[7]~q ),
	.pipeline_dffe_8(\ux004|acc|auto_generated|pipeline_dffe[8]~q ),
	.pipeline_dffe_9(\ux004|acc|auto_generated|pipeline_dffe[9]~q ),
	.pipeline_dffe_10(\ux004|acc|auto_generated|pipeline_dffe[10]~q ),
	.pipeline_dffe_11(\ux004|acc|auto_generated|pipeline_dffe[11]~q ),
	.pipeline_dffe_12(\ux004|acc|auto_generated|pipeline_dffe[12]~q ),
	.pipeline_dffe_15(\ux004|acc|auto_generated|pipeline_dffe[15]~q ),
	.pipeline_dffe_13(\ux004|acc|auto_generated|pipeline_dffe[13]~q ),
	.pipeline_dffe_14(\ux004|acc|auto_generated|pipeline_dffe[14]~q ),
	.clk(clk),
	.reset_n(reset_n),
	.clken(clken),
	.phase_mod_i_0(phase_mod_i_0),
	.phase_mod_i_1(phase_mod_i_1),
	.phase_mod_i_2(phase_mod_i_2),
	.phase_mod_i_3(phase_mod_i_3),
	.phase_mod_i_4(phase_mod_i_4),
	.phase_mod_i_5(phase_mod_i_5),
	.phase_mod_i_6(phase_mod_i_6),
	.phase_mod_i_7(phase_mod_i_7),
	.phase_mod_i_8(phase_mod_i_8),
	.phase_mod_i_9(phase_mod_i_9),
	.phase_mod_i_10(phase_mod_i_10),
	.phase_mod_i_11(phase_mod_i_11),
	.phase_mod_i_12(phase_mod_i_12),
	.phase_mod_i_15(phase_mod_i_15),
	.phase_mod_i_13(phase_mod_i_13),
	.phase_mod_i_14(phase_mod_i_14));

DDS_48_v1_asj_nco_as_m_cen_1 ux0121(
	.ram_block1a64(\ux0121|altsyncram_component0|auto_generated|ram_block1a64~portadataout ),
	.ram_block1a80(\ux0121|altsyncram_component0|auto_generated|ram_block1a80~portadataout ),
	.ram_block1a96(\ux0121|altsyncram_component0|auto_generated|ram_block1a96~portadataout ),
	.ram_block1a112(\ux0121|altsyncram_component0|auto_generated|ram_block1a112~portadataout ),
	.ram_block1a32(\ux0121|altsyncram_component0|auto_generated|ram_block1a32~portadataout ),
	.ram_block1a48(\ux0121|altsyncram_component0|auto_generated|ram_block1a48~portadataout ),
	.ram_block1a0(\ux0121|altsyncram_component0|auto_generated|ram_block1a0~portadataout ),
	.ram_block1a16(\ux0121|altsyncram_component0|auto_generated|ram_block1a16~portadataout ),
	.ram_block1a65(\ux0121|altsyncram_component0|auto_generated|ram_block1a65~portadataout ),
	.ram_block1a81(\ux0121|altsyncram_component0|auto_generated|ram_block1a81~portadataout ),
	.ram_block1a97(\ux0121|altsyncram_component0|auto_generated|ram_block1a97~portadataout ),
	.ram_block1a113(\ux0121|altsyncram_component0|auto_generated|ram_block1a113~portadataout ),
	.ram_block1a33(\ux0121|altsyncram_component0|auto_generated|ram_block1a33~portadataout ),
	.ram_block1a49(\ux0121|altsyncram_component0|auto_generated|ram_block1a49~portadataout ),
	.ram_block1a1(\ux0121|altsyncram_component0|auto_generated|ram_block1a1~portadataout ),
	.ram_block1a17(\ux0121|altsyncram_component0|auto_generated|ram_block1a17~portadataout ),
	.ram_block1a66(\ux0121|altsyncram_component0|auto_generated|ram_block1a66~portadataout ),
	.ram_block1a82(\ux0121|altsyncram_component0|auto_generated|ram_block1a82~portadataout ),
	.ram_block1a98(\ux0121|altsyncram_component0|auto_generated|ram_block1a98~portadataout ),
	.ram_block1a114(\ux0121|altsyncram_component0|auto_generated|ram_block1a114~portadataout ),
	.ram_block1a34(\ux0121|altsyncram_component0|auto_generated|ram_block1a34~portadataout ),
	.ram_block1a50(\ux0121|altsyncram_component0|auto_generated|ram_block1a50~portadataout ),
	.ram_block1a2(\ux0121|altsyncram_component0|auto_generated|ram_block1a2~portadataout ),
	.ram_block1a18(\ux0121|altsyncram_component0|auto_generated|ram_block1a18~portadataout ),
	.ram_block1a67(\ux0121|altsyncram_component0|auto_generated|ram_block1a67~portadataout ),
	.ram_block1a83(\ux0121|altsyncram_component0|auto_generated|ram_block1a83~portadataout ),
	.ram_block1a99(\ux0121|altsyncram_component0|auto_generated|ram_block1a99~portadataout ),
	.ram_block1a115(\ux0121|altsyncram_component0|auto_generated|ram_block1a115~portadataout ),
	.ram_block1a35(\ux0121|altsyncram_component0|auto_generated|ram_block1a35~portadataout ),
	.ram_block1a51(\ux0121|altsyncram_component0|auto_generated|ram_block1a51~portadataout ),
	.ram_block1a3(\ux0121|altsyncram_component0|auto_generated|ram_block1a3~portadataout ),
	.ram_block1a19(\ux0121|altsyncram_component0|auto_generated|ram_block1a19~portadataout ),
	.ram_block1a68(\ux0121|altsyncram_component0|auto_generated|ram_block1a68~portadataout ),
	.ram_block1a84(\ux0121|altsyncram_component0|auto_generated|ram_block1a84~portadataout ),
	.ram_block1a100(\ux0121|altsyncram_component0|auto_generated|ram_block1a100~portadataout ),
	.ram_block1a116(\ux0121|altsyncram_component0|auto_generated|ram_block1a116~portadataout ),
	.ram_block1a36(\ux0121|altsyncram_component0|auto_generated|ram_block1a36~portadataout ),
	.ram_block1a52(\ux0121|altsyncram_component0|auto_generated|ram_block1a52~portadataout ),
	.ram_block1a4(\ux0121|altsyncram_component0|auto_generated|ram_block1a4~portadataout ),
	.ram_block1a20(\ux0121|altsyncram_component0|auto_generated|ram_block1a20~portadataout ),
	.ram_block1a69(\ux0121|altsyncram_component0|auto_generated|ram_block1a69~portadataout ),
	.ram_block1a85(\ux0121|altsyncram_component0|auto_generated|ram_block1a85~portadataout ),
	.ram_block1a101(\ux0121|altsyncram_component0|auto_generated|ram_block1a101~portadataout ),
	.ram_block1a117(\ux0121|altsyncram_component0|auto_generated|ram_block1a117~portadataout ),
	.ram_block1a37(\ux0121|altsyncram_component0|auto_generated|ram_block1a37~portadataout ),
	.ram_block1a53(\ux0121|altsyncram_component0|auto_generated|ram_block1a53~portadataout ),
	.ram_block1a5(\ux0121|altsyncram_component0|auto_generated|ram_block1a5~portadataout ),
	.ram_block1a21(\ux0121|altsyncram_component0|auto_generated|ram_block1a21~portadataout ),
	.ram_block1a70(\ux0121|altsyncram_component0|auto_generated|ram_block1a70~portadataout ),
	.ram_block1a86(\ux0121|altsyncram_component0|auto_generated|ram_block1a86~portadataout ),
	.ram_block1a102(\ux0121|altsyncram_component0|auto_generated|ram_block1a102~portadataout ),
	.ram_block1a118(\ux0121|altsyncram_component0|auto_generated|ram_block1a118~portadataout ),
	.ram_block1a38(\ux0121|altsyncram_component0|auto_generated|ram_block1a38~portadataout ),
	.ram_block1a54(\ux0121|altsyncram_component0|auto_generated|ram_block1a54~portadataout ),
	.ram_block1a6(\ux0121|altsyncram_component0|auto_generated|ram_block1a6~portadataout ),
	.ram_block1a22(\ux0121|altsyncram_component0|auto_generated|ram_block1a22~portadataout ),
	.ram_block1a71(\ux0121|altsyncram_component0|auto_generated|ram_block1a71~portadataout ),
	.ram_block1a87(\ux0121|altsyncram_component0|auto_generated|ram_block1a87~portadataout ),
	.ram_block1a103(\ux0121|altsyncram_component0|auto_generated|ram_block1a103~portadataout ),
	.ram_block1a119(\ux0121|altsyncram_component0|auto_generated|ram_block1a119~portadataout ),
	.ram_block1a39(\ux0121|altsyncram_component0|auto_generated|ram_block1a39~portadataout ),
	.ram_block1a55(\ux0121|altsyncram_component0|auto_generated|ram_block1a55~portadataout ),
	.ram_block1a7(\ux0121|altsyncram_component0|auto_generated|ram_block1a7~portadataout ),
	.ram_block1a23(\ux0121|altsyncram_component0|auto_generated|ram_block1a23~portadataout ),
	.ram_block1a72(\ux0121|altsyncram_component0|auto_generated|ram_block1a72~portadataout ),
	.ram_block1a88(\ux0121|altsyncram_component0|auto_generated|ram_block1a88~portadataout ),
	.ram_block1a104(\ux0121|altsyncram_component0|auto_generated|ram_block1a104~portadataout ),
	.ram_block1a120(\ux0121|altsyncram_component0|auto_generated|ram_block1a120~portadataout ),
	.ram_block1a40(\ux0121|altsyncram_component0|auto_generated|ram_block1a40~portadataout ),
	.ram_block1a56(\ux0121|altsyncram_component0|auto_generated|ram_block1a56~portadataout ),
	.ram_block1a8(\ux0121|altsyncram_component0|auto_generated|ram_block1a8~portadataout ),
	.ram_block1a24(\ux0121|altsyncram_component0|auto_generated|ram_block1a24~portadataout ),
	.ram_block1a73(\ux0121|altsyncram_component0|auto_generated|ram_block1a73~portadataout ),
	.ram_block1a89(\ux0121|altsyncram_component0|auto_generated|ram_block1a89~portadataout ),
	.ram_block1a105(\ux0121|altsyncram_component0|auto_generated|ram_block1a105~portadataout ),
	.ram_block1a121(\ux0121|altsyncram_component0|auto_generated|ram_block1a121~portadataout ),
	.ram_block1a41(\ux0121|altsyncram_component0|auto_generated|ram_block1a41~portadataout ),
	.ram_block1a57(\ux0121|altsyncram_component0|auto_generated|ram_block1a57~portadataout ),
	.ram_block1a9(\ux0121|altsyncram_component0|auto_generated|ram_block1a9~portadataout ),
	.ram_block1a25(\ux0121|altsyncram_component0|auto_generated|ram_block1a25~portadataout ),
	.ram_block1a74(\ux0121|altsyncram_component0|auto_generated|ram_block1a74~portadataout ),
	.ram_block1a90(\ux0121|altsyncram_component0|auto_generated|ram_block1a90~portadataout ),
	.ram_block1a106(\ux0121|altsyncram_component0|auto_generated|ram_block1a106~portadataout ),
	.ram_block1a122(\ux0121|altsyncram_component0|auto_generated|ram_block1a122~portadataout ),
	.ram_block1a42(\ux0121|altsyncram_component0|auto_generated|ram_block1a42~portadataout ),
	.ram_block1a58(\ux0121|altsyncram_component0|auto_generated|ram_block1a58~portadataout ),
	.ram_block1a10(\ux0121|altsyncram_component0|auto_generated|ram_block1a10~portadataout ),
	.ram_block1a26(\ux0121|altsyncram_component0|auto_generated|ram_block1a26~portadataout ),
	.ram_block1a75(\ux0121|altsyncram_component0|auto_generated|ram_block1a75~portadataout ),
	.ram_block1a91(\ux0121|altsyncram_component0|auto_generated|ram_block1a91~portadataout ),
	.ram_block1a107(\ux0121|altsyncram_component0|auto_generated|ram_block1a107~portadataout ),
	.ram_block1a123(\ux0121|altsyncram_component0|auto_generated|ram_block1a123~portadataout ),
	.ram_block1a43(\ux0121|altsyncram_component0|auto_generated|ram_block1a43~portadataout ),
	.ram_block1a59(\ux0121|altsyncram_component0|auto_generated|ram_block1a59~portadataout ),
	.ram_block1a11(\ux0121|altsyncram_component0|auto_generated|ram_block1a11~portadataout ),
	.ram_block1a27(\ux0121|altsyncram_component0|auto_generated|ram_block1a27~portadataout ),
	.ram_block1a76(\ux0121|altsyncram_component0|auto_generated|ram_block1a76~portadataout ),
	.ram_block1a92(\ux0121|altsyncram_component0|auto_generated|ram_block1a92~portadataout ),
	.ram_block1a108(\ux0121|altsyncram_component0|auto_generated|ram_block1a108~portadataout ),
	.ram_block1a124(\ux0121|altsyncram_component0|auto_generated|ram_block1a124~portadataout ),
	.ram_block1a44(\ux0121|altsyncram_component0|auto_generated|ram_block1a44~portadataout ),
	.ram_block1a60(\ux0121|altsyncram_component0|auto_generated|ram_block1a60~portadataout ),
	.ram_block1a12(\ux0121|altsyncram_component0|auto_generated|ram_block1a12~portadataout ),
	.ram_block1a28(\ux0121|altsyncram_component0|auto_generated|ram_block1a28~portadataout ),
	.ram_block1a77(\ux0121|altsyncram_component0|auto_generated|ram_block1a77~portadataout ),
	.ram_block1a93(\ux0121|altsyncram_component0|auto_generated|ram_block1a93~portadataout ),
	.ram_block1a109(\ux0121|altsyncram_component0|auto_generated|ram_block1a109~portadataout ),
	.ram_block1a125(\ux0121|altsyncram_component0|auto_generated|ram_block1a125~portadataout ),
	.ram_block1a45(\ux0121|altsyncram_component0|auto_generated|ram_block1a45~portadataout ),
	.ram_block1a61(\ux0121|altsyncram_component0|auto_generated|ram_block1a61~portadataout ),
	.ram_block1a13(\ux0121|altsyncram_component0|auto_generated|ram_block1a13~portadataout ),
	.ram_block1a29(\ux0121|altsyncram_component0|auto_generated|ram_block1a29~portadataout ),
	.ram_block1a78(\ux0121|altsyncram_component0|auto_generated|ram_block1a78~portadataout ),
	.ram_block1a94(\ux0121|altsyncram_component0|auto_generated|ram_block1a94~portadataout ),
	.ram_block1a110(\ux0121|altsyncram_component0|auto_generated|ram_block1a110~portadataout ),
	.ram_block1a126(\ux0121|altsyncram_component0|auto_generated|ram_block1a126~portadataout ),
	.ram_block1a46(\ux0121|altsyncram_component0|auto_generated|ram_block1a46~portadataout ),
	.ram_block1a62(\ux0121|altsyncram_component0|auto_generated|ram_block1a62~portadataout ),
	.ram_block1a14(\ux0121|altsyncram_component0|auto_generated|ram_block1a14~portadataout ),
	.ram_block1a30(\ux0121|altsyncram_component0|auto_generated|ram_block1a30~portadataout ),
	.ram_block1a79(\ux0121|altsyncram_component0|auto_generated|ram_block1a79~portadataout ),
	.ram_block1a95(\ux0121|altsyncram_component0|auto_generated|ram_block1a95~portadataout ),
	.ram_block1a111(\ux0121|altsyncram_component0|auto_generated|ram_block1a111~portadataout ),
	.ram_block1a127(\ux0121|altsyncram_component0|auto_generated|ram_block1a127~portadataout ),
	.ram_block1a47(\ux0121|altsyncram_component0|auto_generated|ram_block1a47~portadataout ),
	.ram_block1a63(\ux0121|altsyncram_component0|auto_generated|ram_block1a63~portadataout ),
	.ram_block1a15(\ux0121|altsyncram_component0|auto_generated|ram_block1a15~portadataout ),
	.ram_block1a31(\ux0121|altsyncram_component0|auto_generated|ram_block1a31~portadataout ),
	.rom_add_0(\ux009|rom_add[0]~q ),
	.rom_add_1(\ux009|rom_add[1]~q ),
	.rom_add_2(\ux009|rom_add[2]~q ),
	.rom_add_3(\ux009|rom_add[3]~q ),
	.rom_add_4(\ux009|rom_add[4]~q ),
	.rom_add_5(\ux009|rom_add[5]~q ),
	.rom_add_6(\ux009|rom_add[6]~q ),
	.rom_add_7(\ux009|rom_add[7]~q ),
	.rom_add_8(\ux009|rom_add[8]~q ),
	.rom_add_9(\ux009|rom_add[9]~q ),
	.rom_add_10(\ux009|rom_add[10]~q ),
	.rom_add_11(\ux009|rom_add[11]~q ),
	.rom_add_12(\ux009|rom_add[12]~q ),
	.clk(clk),
	.clken(clken));

DDS_48_v1_asj_nco_as_m_cen ux0120(
	.ram_block1a64(\ux0120|altsyncram_component0|auto_generated|ram_block1a64~portadataout ),
	.ram_block1a80(\ux0120|altsyncram_component0|auto_generated|ram_block1a80~portadataout ),
	.ram_block1a96(\ux0120|altsyncram_component0|auto_generated|ram_block1a96~portadataout ),
	.ram_block1a112(\ux0120|altsyncram_component0|auto_generated|ram_block1a112~portadataout ),
	.ram_block1a32(\ux0120|altsyncram_component0|auto_generated|ram_block1a32~portadataout ),
	.ram_block1a48(\ux0120|altsyncram_component0|auto_generated|ram_block1a48~portadataout ),
	.ram_block1a0(\ux0120|altsyncram_component0|auto_generated|ram_block1a0~portadataout ),
	.ram_block1a16(\ux0120|altsyncram_component0|auto_generated|ram_block1a16~portadataout ),
	.ram_block1a65(\ux0120|altsyncram_component0|auto_generated|ram_block1a65~portadataout ),
	.ram_block1a81(\ux0120|altsyncram_component0|auto_generated|ram_block1a81~portadataout ),
	.ram_block1a97(\ux0120|altsyncram_component0|auto_generated|ram_block1a97~portadataout ),
	.ram_block1a113(\ux0120|altsyncram_component0|auto_generated|ram_block1a113~portadataout ),
	.ram_block1a33(\ux0120|altsyncram_component0|auto_generated|ram_block1a33~portadataout ),
	.ram_block1a49(\ux0120|altsyncram_component0|auto_generated|ram_block1a49~portadataout ),
	.ram_block1a1(\ux0120|altsyncram_component0|auto_generated|ram_block1a1~portadataout ),
	.ram_block1a17(\ux0120|altsyncram_component0|auto_generated|ram_block1a17~portadataout ),
	.ram_block1a66(\ux0120|altsyncram_component0|auto_generated|ram_block1a66~portadataout ),
	.ram_block1a82(\ux0120|altsyncram_component0|auto_generated|ram_block1a82~portadataout ),
	.ram_block1a98(\ux0120|altsyncram_component0|auto_generated|ram_block1a98~portadataout ),
	.ram_block1a114(\ux0120|altsyncram_component0|auto_generated|ram_block1a114~portadataout ),
	.ram_block1a34(\ux0120|altsyncram_component0|auto_generated|ram_block1a34~portadataout ),
	.ram_block1a50(\ux0120|altsyncram_component0|auto_generated|ram_block1a50~portadataout ),
	.ram_block1a2(\ux0120|altsyncram_component0|auto_generated|ram_block1a2~portadataout ),
	.ram_block1a18(\ux0120|altsyncram_component0|auto_generated|ram_block1a18~portadataout ),
	.ram_block1a67(\ux0120|altsyncram_component0|auto_generated|ram_block1a67~portadataout ),
	.ram_block1a83(\ux0120|altsyncram_component0|auto_generated|ram_block1a83~portadataout ),
	.ram_block1a99(\ux0120|altsyncram_component0|auto_generated|ram_block1a99~portadataout ),
	.ram_block1a115(\ux0120|altsyncram_component0|auto_generated|ram_block1a115~portadataout ),
	.ram_block1a35(\ux0120|altsyncram_component0|auto_generated|ram_block1a35~portadataout ),
	.ram_block1a51(\ux0120|altsyncram_component0|auto_generated|ram_block1a51~portadataout ),
	.ram_block1a3(\ux0120|altsyncram_component0|auto_generated|ram_block1a3~portadataout ),
	.ram_block1a19(\ux0120|altsyncram_component0|auto_generated|ram_block1a19~portadataout ),
	.ram_block1a68(\ux0120|altsyncram_component0|auto_generated|ram_block1a68~portadataout ),
	.ram_block1a84(\ux0120|altsyncram_component0|auto_generated|ram_block1a84~portadataout ),
	.ram_block1a100(\ux0120|altsyncram_component0|auto_generated|ram_block1a100~portadataout ),
	.ram_block1a116(\ux0120|altsyncram_component0|auto_generated|ram_block1a116~portadataout ),
	.ram_block1a36(\ux0120|altsyncram_component0|auto_generated|ram_block1a36~portadataout ),
	.ram_block1a52(\ux0120|altsyncram_component0|auto_generated|ram_block1a52~portadataout ),
	.ram_block1a4(\ux0120|altsyncram_component0|auto_generated|ram_block1a4~portadataout ),
	.ram_block1a20(\ux0120|altsyncram_component0|auto_generated|ram_block1a20~portadataout ),
	.ram_block1a69(\ux0120|altsyncram_component0|auto_generated|ram_block1a69~portadataout ),
	.ram_block1a85(\ux0120|altsyncram_component0|auto_generated|ram_block1a85~portadataout ),
	.ram_block1a101(\ux0120|altsyncram_component0|auto_generated|ram_block1a101~portadataout ),
	.ram_block1a117(\ux0120|altsyncram_component0|auto_generated|ram_block1a117~portadataout ),
	.ram_block1a37(\ux0120|altsyncram_component0|auto_generated|ram_block1a37~portadataout ),
	.ram_block1a53(\ux0120|altsyncram_component0|auto_generated|ram_block1a53~portadataout ),
	.ram_block1a5(\ux0120|altsyncram_component0|auto_generated|ram_block1a5~portadataout ),
	.ram_block1a21(\ux0120|altsyncram_component0|auto_generated|ram_block1a21~portadataout ),
	.ram_block1a70(\ux0120|altsyncram_component0|auto_generated|ram_block1a70~portadataout ),
	.ram_block1a86(\ux0120|altsyncram_component0|auto_generated|ram_block1a86~portadataout ),
	.ram_block1a102(\ux0120|altsyncram_component0|auto_generated|ram_block1a102~portadataout ),
	.ram_block1a118(\ux0120|altsyncram_component0|auto_generated|ram_block1a118~portadataout ),
	.ram_block1a38(\ux0120|altsyncram_component0|auto_generated|ram_block1a38~portadataout ),
	.ram_block1a54(\ux0120|altsyncram_component0|auto_generated|ram_block1a54~portadataout ),
	.ram_block1a6(\ux0120|altsyncram_component0|auto_generated|ram_block1a6~portadataout ),
	.ram_block1a22(\ux0120|altsyncram_component0|auto_generated|ram_block1a22~portadataout ),
	.ram_block1a71(\ux0120|altsyncram_component0|auto_generated|ram_block1a71~portadataout ),
	.ram_block1a87(\ux0120|altsyncram_component0|auto_generated|ram_block1a87~portadataout ),
	.ram_block1a103(\ux0120|altsyncram_component0|auto_generated|ram_block1a103~portadataout ),
	.ram_block1a119(\ux0120|altsyncram_component0|auto_generated|ram_block1a119~portadataout ),
	.ram_block1a39(\ux0120|altsyncram_component0|auto_generated|ram_block1a39~portadataout ),
	.ram_block1a55(\ux0120|altsyncram_component0|auto_generated|ram_block1a55~portadataout ),
	.ram_block1a7(\ux0120|altsyncram_component0|auto_generated|ram_block1a7~portadataout ),
	.ram_block1a23(\ux0120|altsyncram_component0|auto_generated|ram_block1a23~portadataout ),
	.ram_block1a72(\ux0120|altsyncram_component0|auto_generated|ram_block1a72~portadataout ),
	.ram_block1a88(\ux0120|altsyncram_component0|auto_generated|ram_block1a88~portadataout ),
	.ram_block1a104(\ux0120|altsyncram_component0|auto_generated|ram_block1a104~portadataout ),
	.ram_block1a120(\ux0120|altsyncram_component0|auto_generated|ram_block1a120~portadataout ),
	.ram_block1a40(\ux0120|altsyncram_component0|auto_generated|ram_block1a40~portadataout ),
	.ram_block1a56(\ux0120|altsyncram_component0|auto_generated|ram_block1a56~portadataout ),
	.ram_block1a8(\ux0120|altsyncram_component0|auto_generated|ram_block1a8~portadataout ),
	.ram_block1a24(\ux0120|altsyncram_component0|auto_generated|ram_block1a24~portadataout ),
	.ram_block1a73(\ux0120|altsyncram_component0|auto_generated|ram_block1a73~portadataout ),
	.ram_block1a89(\ux0120|altsyncram_component0|auto_generated|ram_block1a89~portadataout ),
	.ram_block1a105(\ux0120|altsyncram_component0|auto_generated|ram_block1a105~portadataout ),
	.ram_block1a121(\ux0120|altsyncram_component0|auto_generated|ram_block1a121~portadataout ),
	.ram_block1a41(\ux0120|altsyncram_component0|auto_generated|ram_block1a41~portadataout ),
	.ram_block1a57(\ux0120|altsyncram_component0|auto_generated|ram_block1a57~portadataout ),
	.ram_block1a9(\ux0120|altsyncram_component0|auto_generated|ram_block1a9~portadataout ),
	.ram_block1a25(\ux0120|altsyncram_component0|auto_generated|ram_block1a25~portadataout ),
	.ram_block1a74(\ux0120|altsyncram_component0|auto_generated|ram_block1a74~portadataout ),
	.ram_block1a90(\ux0120|altsyncram_component0|auto_generated|ram_block1a90~portadataout ),
	.ram_block1a106(\ux0120|altsyncram_component0|auto_generated|ram_block1a106~portadataout ),
	.ram_block1a122(\ux0120|altsyncram_component0|auto_generated|ram_block1a122~portadataout ),
	.ram_block1a42(\ux0120|altsyncram_component0|auto_generated|ram_block1a42~portadataout ),
	.ram_block1a58(\ux0120|altsyncram_component0|auto_generated|ram_block1a58~portadataout ),
	.ram_block1a10(\ux0120|altsyncram_component0|auto_generated|ram_block1a10~portadataout ),
	.ram_block1a26(\ux0120|altsyncram_component0|auto_generated|ram_block1a26~portadataout ),
	.ram_block1a75(\ux0120|altsyncram_component0|auto_generated|ram_block1a75~portadataout ),
	.ram_block1a91(\ux0120|altsyncram_component0|auto_generated|ram_block1a91~portadataout ),
	.ram_block1a107(\ux0120|altsyncram_component0|auto_generated|ram_block1a107~portadataout ),
	.ram_block1a123(\ux0120|altsyncram_component0|auto_generated|ram_block1a123~portadataout ),
	.ram_block1a43(\ux0120|altsyncram_component0|auto_generated|ram_block1a43~portadataout ),
	.ram_block1a59(\ux0120|altsyncram_component0|auto_generated|ram_block1a59~portadataout ),
	.ram_block1a11(\ux0120|altsyncram_component0|auto_generated|ram_block1a11~portadataout ),
	.ram_block1a27(\ux0120|altsyncram_component0|auto_generated|ram_block1a27~portadataout ),
	.ram_block1a76(\ux0120|altsyncram_component0|auto_generated|ram_block1a76~portadataout ),
	.ram_block1a92(\ux0120|altsyncram_component0|auto_generated|ram_block1a92~portadataout ),
	.ram_block1a108(\ux0120|altsyncram_component0|auto_generated|ram_block1a108~portadataout ),
	.ram_block1a124(\ux0120|altsyncram_component0|auto_generated|ram_block1a124~portadataout ),
	.ram_block1a44(\ux0120|altsyncram_component0|auto_generated|ram_block1a44~portadataout ),
	.ram_block1a60(\ux0120|altsyncram_component0|auto_generated|ram_block1a60~portadataout ),
	.ram_block1a12(\ux0120|altsyncram_component0|auto_generated|ram_block1a12~portadataout ),
	.ram_block1a28(\ux0120|altsyncram_component0|auto_generated|ram_block1a28~portadataout ),
	.ram_block1a77(\ux0120|altsyncram_component0|auto_generated|ram_block1a77~portadataout ),
	.ram_block1a93(\ux0120|altsyncram_component0|auto_generated|ram_block1a93~portadataout ),
	.ram_block1a109(\ux0120|altsyncram_component0|auto_generated|ram_block1a109~portadataout ),
	.ram_block1a125(\ux0120|altsyncram_component0|auto_generated|ram_block1a125~portadataout ),
	.ram_block1a45(\ux0120|altsyncram_component0|auto_generated|ram_block1a45~portadataout ),
	.ram_block1a61(\ux0120|altsyncram_component0|auto_generated|ram_block1a61~portadataout ),
	.ram_block1a13(\ux0120|altsyncram_component0|auto_generated|ram_block1a13~portadataout ),
	.ram_block1a29(\ux0120|altsyncram_component0|auto_generated|ram_block1a29~portadataout ),
	.ram_block1a78(\ux0120|altsyncram_component0|auto_generated|ram_block1a78~portadataout ),
	.ram_block1a94(\ux0120|altsyncram_component0|auto_generated|ram_block1a94~portadataout ),
	.ram_block1a110(\ux0120|altsyncram_component0|auto_generated|ram_block1a110~portadataout ),
	.ram_block1a126(\ux0120|altsyncram_component0|auto_generated|ram_block1a126~portadataout ),
	.ram_block1a46(\ux0120|altsyncram_component0|auto_generated|ram_block1a46~portadataout ),
	.ram_block1a62(\ux0120|altsyncram_component0|auto_generated|ram_block1a62~portadataout ),
	.ram_block1a14(\ux0120|altsyncram_component0|auto_generated|ram_block1a14~portadataout ),
	.ram_block1a30(\ux0120|altsyncram_component0|auto_generated|ram_block1a30~portadataout ),
	.ram_block1a79(\ux0120|altsyncram_component0|auto_generated|ram_block1a79~portadataout ),
	.ram_block1a95(\ux0120|altsyncram_component0|auto_generated|ram_block1a95~portadataout ),
	.ram_block1a111(\ux0120|altsyncram_component0|auto_generated|ram_block1a111~portadataout ),
	.ram_block1a127(\ux0120|altsyncram_component0|auto_generated|ram_block1a127~portadataout ),
	.ram_block1a47(\ux0120|altsyncram_component0|auto_generated|ram_block1a47~portadataout ),
	.ram_block1a63(\ux0120|altsyncram_component0|auto_generated|ram_block1a63~portadataout ),
	.ram_block1a15(\ux0120|altsyncram_component0|auto_generated|ram_block1a15~portadataout ),
	.ram_block1a31(\ux0120|altsyncram_component0|auto_generated|ram_block1a31~portadataout ),
	.rom_add_0(\ux009|rom_add[0]~q ),
	.rom_add_1(\ux009|rom_add[1]~q ),
	.rom_add_2(\ux009|rom_add[2]~q ),
	.rom_add_3(\ux009|rom_add[3]~q ),
	.rom_add_4(\ux009|rom_add[4]~q ),
	.rom_add_5(\ux009|rom_add[5]~q ),
	.rom_add_6(\ux009|rom_add[6]~q ),
	.rom_add_7(\ux009|rom_add[7]~q ),
	.rom_add_8(\ux009|rom_add[8]~q ),
	.rom_add_9(\ux009|rom_add[9]~q ),
	.rom_add_10(\ux009|rom_add[10]~q ),
	.rom_add_11(\ux009|rom_add[11]~q ),
	.rom_add_12(\ux009|rom_add[12]~q ),
	.rom_add_15(\ux009|rom_add[15]~q ),
	.rom_add_13(\ux009|rom_add[13]~q ),
	.rom_add_14(\ux009|rom_add[14]~q ),
	.out_address_reg_a_2(\ux0120|altsyncram_component0|auto_generated|out_address_reg_a[2]~q ),
	.out_address_reg_a_0(\ux0120|altsyncram_component0|auto_generated|out_address_reg_a[0]~q ),
	.out_address_reg_a_1(\ux0120|altsyncram_component0|auto_generated|out_address_reg_a[1]~q ),
	.clk(clk),
	.clken(clken));

endmodule

module DDS_48_v1_asj_altqmcpipe (
	data_out_12,
	pipeline_dffe_32,
	pipeline_dffe_33,
	pipeline_dffe_34,
	pipeline_dffe_35,
	pipeline_dffe_36,
	pipeline_dffe_37,
	pipeline_dffe_38,
	pipeline_dffe_39,
	pipeline_dffe_40,
	pipeline_dffe_41,
	pipeline_dffe_42,
	pipeline_dffe_43,
	pipeline_dffe_44,
	pipeline_dffe_47,
	pipeline_dffe_31,
	pipeline_dffe_45,
	pipeline_dffe_46,
	pipeline_dffe_30,
	pipeline_dffe_321,
	pipeline_dffe_29,
	pipeline_dffe_331,
	pipeline_dffe_341,
	pipeline_dffe_351,
	pipeline_dffe_361,
	pipeline_dffe_371,
	pipeline_dffe_381,
	pipeline_dffe_391,
	pipeline_dffe_401,
	pipeline_dffe_411,
	pipeline_dffe_421,
	pipeline_dffe_431,
	pipeline_dffe_441,
	pipeline_dffe_471,
	pipeline_dffe_311,
	pipeline_dffe_28,
	pipeline_dffe_451,
	pipeline_dffe_461,
	pipeline_dffe_301,
	pipeline_dffe_27,
	pipeline_dffe_291,
	pipeline_dffe_281,
	pipeline_dffe_271,
	pipeline_dffe_26,
	pipeline_dffe_25,
	pipeline_dffe_24,
	pipeline_dffe_23,
	pipeline_dffe_22,
	pipeline_dffe_21,
	pipeline_dffe_20,
	pipeline_dffe_19,
	pipeline_dffe_18,
	pipeline_dffe_17,
	pipeline_dffe_16,
	pipeline_dffe_15,
	pipeline_dffe_14,
	pipeline_dffe_13,
	pipeline_dffe_12,
	pipeline_dffe_11,
	pipeline_dffe_10,
	pipeline_dffe_9,
	pipeline_dffe_8,
	pipeline_dffe_7,
	pipeline_dffe_6,
	pipeline_dffe_5,
	pipeline_dffe_4,
	pipeline_dffe_3,
	pipeline_dffe_2,
	pipeline_dffe_1,
	pipeline_dffe_0,
	clk,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	data_out_12;
output 	pipeline_dffe_32;
output 	pipeline_dffe_33;
output 	pipeline_dffe_34;
output 	pipeline_dffe_35;
output 	pipeline_dffe_36;
output 	pipeline_dffe_37;
output 	pipeline_dffe_38;
output 	pipeline_dffe_39;
output 	pipeline_dffe_40;
output 	pipeline_dffe_41;
output 	pipeline_dffe_42;
output 	pipeline_dffe_43;
output 	pipeline_dffe_44;
output 	pipeline_dffe_47;
output 	pipeline_dffe_31;
output 	pipeline_dffe_45;
output 	pipeline_dffe_46;
output 	pipeline_dffe_30;
input 	pipeline_dffe_321;
output 	pipeline_dffe_29;
input 	pipeline_dffe_331;
input 	pipeline_dffe_341;
input 	pipeline_dffe_351;
input 	pipeline_dffe_361;
input 	pipeline_dffe_371;
input 	pipeline_dffe_381;
input 	pipeline_dffe_391;
input 	pipeline_dffe_401;
input 	pipeline_dffe_411;
input 	pipeline_dffe_421;
input 	pipeline_dffe_431;
input 	pipeline_dffe_441;
input 	pipeline_dffe_471;
input 	pipeline_dffe_311;
output 	pipeline_dffe_28;
input 	pipeline_dffe_451;
input 	pipeline_dffe_461;
input 	pipeline_dffe_301;
output 	pipeline_dffe_27;
input 	pipeline_dffe_291;
input 	pipeline_dffe_281;
input 	pipeline_dffe_271;
input 	pipeline_dffe_26;
input 	pipeline_dffe_25;
input 	pipeline_dffe_24;
input 	pipeline_dffe_23;
input 	pipeline_dffe_22;
input 	pipeline_dffe_21;
input 	pipeline_dffe_20;
input 	pipeline_dffe_19;
input 	pipeline_dffe_18;
input 	pipeline_dffe_17;
input 	pipeline_dffe_16;
input 	pipeline_dffe_15;
input 	pipeline_dffe_14;
input 	pipeline_dffe_13;
input 	pipeline_dffe_12;
input 	pipeline_dffe_11;
input 	pipeline_dffe_10;
input 	pipeline_dffe_9;
input 	pipeline_dffe_8;
input 	pipeline_dffe_7;
input 	pipeline_dffe_6;
input 	pipeline_dffe_5;
input 	pipeline_dffe_4;
input 	pipeline_dffe_3;
input 	pipeline_dffe_2;
input 	pipeline_dffe_1;
input 	pipeline_dffe_0;
input 	clk;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \phi_int_arr_reg[32]~q ;
wire \phi_int_arr_reg[33]~q ;
wire \phi_int_arr_reg[34]~q ;
wire \phi_int_arr_reg[35]~q ;
wire \phi_int_arr_reg[36]~q ;
wire \phi_int_arr_reg[37]~q ;
wire \phi_int_arr_reg[38]~q ;
wire \phi_int_arr_reg[39]~q ;
wire \phi_int_arr_reg[40]~q ;
wire \phi_int_arr_reg[41]~q ;
wire \phi_int_arr_reg[42]~q ;
wire \phi_int_arr_reg[43]~q ;
wire \phi_int_arr_reg[44]~q ;
wire \phi_int_arr_reg[47]~q ;
wire \phi_int_arr_reg[31]~q ;
wire \phi_int_arr_reg[45]~q ;
wire \phi_int_arr_reg[46]~q ;
wire \phi_int_arr_reg[30]~q ;
wire \phi_int_arr_reg[29]~q ;
wire \phi_int_arr_reg[28]~q ;
wire \phi_int_arr_reg[27]~q ;
wire \phi_int_arr_reg[26]~q ;
wire \phi_int_arr_reg[25]~q ;
wire \phi_int_arr_reg[24]~q ;
wire \phi_int_arr_reg[23]~q ;
wire \phi_int_arr_reg[22]~q ;
wire \phi_int_arr_reg[21]~q ;
wire \phi_int_arr_reg[20]~q ;
wire \phi_int_arr_reg[19]~q ;
wire \phi_int_arr_reg[18]~q ;
wire \phi_int_arr_reg[17]~q ;
wire \phi_int_arr_reg[16]~q ;
wire \phi_int_arr_reg[15]~q ;
wire \phi_int_arr_reg[14]~q ;
wire \phi_int_arr_reg[13]~q ;
wire \phi_int_arr_reg[12]~q ;
wire \phi_int_arr_reg[11]~q ;
wire \phi_int_arr_reg[10]~q ;
wire \phi_int_arr_reg[9]~q ;
wire \phi_int_arr_reg[8]~q ;
wire \phi_int_arr_reg[7]~q ;
wire \phi_int_arr_reg[6]~q ;
wire \phi_int_arr_reg[5]~q ;
wire \phi_int_arr_reg[4]~q ;
wire \phi_int_arr_reg[3]~q ;
wire \phi_int_arr_reg[2]~q ;
wire \phi_int_arr_reg[1]~q ;
wire \phi_int_arr_reg[0]~q ;


DDS_48_v1_lpm_add_sub_1 acc(
	.phi_int_arr_reg_32(\phi_int_arr_reg[32]~q ),
	.phi_int_arr_reg_33(\phi_int_arr_reg[33]~q ),
	.phi_int_arr_reg_34(\phi_int_arr_reg[34]~q ),
	.phi_int_arr_reg_35(\phi_int_arr_reg[35]~q ),
	.phi_int_arr_reg_36(\phi_int_arr_reg[36]~q ),
	.phi_int_arr_reg_37(\phi_int_arr_reg[37]~q ),
	.phi_int_arr_reg_38(\phi_int_arr_reg[38]~q ),
	.phi_int_arr_reg_39(\phi_int_arr_reg[39]~q ),
	.phi_int_arr_reg_40(\phi_int_arr_reg[40]~q ),
	.phi_int_arr_reg_41(\phi_int_arr_reg[41]~q ),
	.phi_int_arr_reg_42(\phi_int_arr_reg[42]~q ),
	.phi_int_arr_reg_43(\phi_int_arr_reg[43]~q ),
	.phi_int_arr_reg_44(\phi_int_arr_reg[44]~q ),
	.phi_int_arr_reg_47(\phi_int_arr_reg[47]~q ),
	.phi_int_arr_reg_31(\phi_int_arr_reg[31]~q ),
	.phi_int_arr_reg_45(\phi_int_arr_reg[45]~q ),
	.phi_int_arr_reg_46(\phi_int_arr_reg[46]~q ),
	.phi_int_arr_reg_30(\phi_int_arr_reg[30]~q ),
	.phi_int_arr_reg_29(\phi_int_arr_reg[29]~q ),
	.phi_int_arr_reg_28(\phi_int_arr_reg[28]~q ),
	.phi_int_arr_reg_27(\phi_int_arr_reg[27]~q ),
	.phi_int_arr_reg_26(\phi_int_arr_reg[26]~q ),
	.phi_int_arr_reg_25(\phi_int_arr_reg[25]~q ),
	.phi_int_arr_reg_24(\phi_int_arr_reg[24]~q ),
	.phi_int_arr_reg_23(\phi_int_arr_reg[23]~q ),
	.phi_int_arr_reg_22(\phi_int_arr_reg[22]~q ),
	.phi_int_arr_reg_21(\phi_int_arr_reg[21]~q ),
	.phi_int_arr_reg_20(\phi_int_arr_reg[20]~q ),
	.phi_int_arr_reg_19(\phi_int_arr_reg[19]~q ),
	.phi_int_arr_reg_18(\phi_int_arr_reg[18]~q ),
	.phi_int_arr_reg_17(\phi_int_arr_reg[17]~q ),
	.phi_int_arr_reg_16(\phi_int_arr_reg[16]~q ),
	.phi_int_arr_reg_15(\phi_int_arr_reg[15]~q ),
	.phi_int_arr_reg_14(\phi_int_arr_reg[14]~q ),
	.phi_int_arr_reg_13(\phi_int_arr_reg[13]~q ),
	.phi_int_arr_reg_12(\phi_int_arr_reg[12]~q ),
	.phi_int_arr_reg_11(\phi_int_arr_reg[11]~q ),
	.phi_int_arr_reg_10(\phi_int_arr_reg[10]~q ),
	.phi_int_arr_reg_9(\phi_int_arr_reg[9]~q ),
	.phi_int_arr_reg_8(\phi_int_arr_reg[8]~q ),
	.phi_int_arr_reg_7(\phi_int_arr_reg[7]~q ),
	.phi_int_arr_reg_6(\phi_int_arr_reg[6]~q ),
	.phi_int_arr_reg_5(\phi_int_arr_reg[5]~q ),
	.phi_int_arr_reg_4(\phi_int_arr_reg[4]~q ),
	.phi_int_arr_reg_3(\phi_int_arr_reg[3]~q ),
	.phi_int_arr_reg_2(\phi_int_arr_reg[2]~q ),
	.phi_int_arr_reg_1(\phi_int_arr_reg[1]~q ),
	.phi_int_arr_reg_0(\phi_int_arr_reg[0]~q ),
	.pipeline_dffe_32(pipeline_dffe_32),
	.pipeline_dffe_33(pipeline_dffe_33),
	.pipeline_dffe_34(pipeline_dffe_34),
	.pipeline_dffe_35(pipeline_dffe_35),
	.pipeline_dffe_36(pipeline_dffe_36),
	.pipeline_dffe_37(pipeline_dffe_37),
	.pipeline_dffe_38(pipeline_dffe_38),
	.pipeline_dffe_39(pipeline_dffe_39),
	.pipeline_dffe_40(pipeline_dffe_40),
	.pipeline_dffe_41(pipeline_dffe_41),
	.pipeline_dffe_42(pipeline_dffe_42),
	.pipeline_dffe_43(pipeline_dffe_43),
	.pipeline_dffe_44(pipeline_dffe_44),
	.pipeline_dffe_47(pipeline_dffe_47),
	.pipeline_dffe_31(pipeline_dffe_31),
	.pipeline_dffe_45(pipeline_dffe_45),
	.pipeline_dffe_46(pipeline_dffe_46),
	.pipeline_dffe_30(pipeline_dffe_30),
	.pipeline_dffe_29(pipeline_dffe_29),
	.pipeline_dffe_28(pipeline_dffe_28),
	.pipeline_dffe_27(pipeline_dffe_27),
	.clock(clk),
	.reset_n(reset_n),
	.clken(clken));

dffeas \phi_int_arr_reg[32] (
	.clk(clk),
	.d(pipeline_dffe_321),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_int_arr_reg[32]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[32] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[32] .power_up = "low";

dffeas \phi_int_arr_reg[33] (
	.clk(clk),
	.d(pipeline_dffe_331),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_int_arr_reg[33]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[33] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[33] .power_up = "low";

dffeas \phi_int_arr_reg[34] (
	.clk(clk),
	.d(pipeline_dffe_341),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_int_arr_reg[34]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[34] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[34] .power_up = "low";

dffeas \phi_int_arr_reg[35] (
	.clk(clk),
	.d(pipeline_dffe_351),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_int_arr_reg[35]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[35] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[35] .power_up = "low";

dffeas \phi_int_arr_reg[36] (
	.clk(clk),
	.d(pipeline_dffe_361),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_int_arr_reg[36]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[36] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[36] .power_up = "low";

dffeas \phi_int_arr_reg[37] (
	.clk(clk),
	.d(pipeline_dffe_371),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_int_arr_reg[37]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[37] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[37] .power_up = "low";

dffeas \phi_int_arr_reg[38] (
	.clk(clk),
	.d(pipeline_dffe_381),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_int_arr_reg[38]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[38] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[38] .power_up = "low";

dffeas \phi_int_arr_reg[39] (
	.clk(clk),
	.d(pipeline_dffe_391),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_int_arr_reg[39]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[39] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[39] .power_up = "low";

dffeas \phi_int_arr_reg[40] (
	.clk(clk),
	.d(pipeline_dffe_401),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_int_arr_reg[40]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[40] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[40] .power_up = "low";

dffeas \phi_int_arr_reg[41] (
	.clk(clk),
	.d(pipeline_dffe_411),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_int_arr_reg[41]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[41] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[41] .power_up = "low";

dffeas \phi_int_arr_reg[42] (
	.clk(clk),
	.d(pipeline_dffe_421),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_int_arr_reg[42]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[42] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[42] .power_up = "low";

dffeas \phi_int_arr_reg[43] (
	.clk(clk),
	.d(pipeline_dffe_431),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_int_arr_reg[43]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[43] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[43] .power_up = "low";

dffeas \phi_int_arr_reg[44] (
	.clk(clk),
	.d(pipeline_dffe_441),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_int_arr_reg[44]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[44] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[44] .power_up = "low";

dffeas \phi_int_arr_reg[47] (
	.clk(clk),
	.d(pipeline_dffe_471),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_int_arr_reg[47]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[47] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[47] .power_up = "low";

dffeas \phi_int_arr_reg[31] (
	.clk(clk),
	.d(pipeline_dffe_311),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_int_arr_reg[31]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[31] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[31] .power_up = "low";

dffeas \phi_int_arr_reg[45] (
	.clk(clk),
	.d(pipeline_dffe_451),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_int_arr_reg[45]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[45] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[45] .power_up = "low";

dffeas \phi_int_arr_reg[46] (
	.clk(clk),
	.d(pipeline_dffe_461),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_int_arr_reg[46]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[46] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[46] .power_up = "low";

dffeas \phi_int_arr_reg[30] (
	.clk(clk),
	.d(pipeline_dffe_301),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_int_arr_reg[30]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[30] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[30] .power_up = "low";

dffeas \phi_int_arr_reg[29] (
	.clk(clk),
	.d(pipeline_dffe_291),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_int_arr_reg[29]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[29] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[29] .power_up = "low";

dffeas \phi_int_arr_reg[28] (
	.clk(clk),
	.d(pipeline_dffe_281),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_int_arr_reg[28]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[28] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[28] .power_up = "low";

dffeas \phi_int_arr_reg[27] (
	.clk(clk),
	.d(pipeline_dffe_271),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_int_arr_reg[27]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[27] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[27] .power_up = "low";

dffeas \phi_int_arr_reg[26] (
	.clk(clk),
	.d(pipeline_dffe_26),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_int_arr_reg[26]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[26] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[26] .power_up = "low";

dffeas \phi_int_arr_reg[25] (
	.clk(clk),
	.d(pipeline_dffe_25),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_int_arr_reg[25]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[25] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[25] .power_up = "low";

dffeas \phi_int_arr_reg[24] (
	.clk(clk),
	.d(pipeline_dffe_24),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_int_arr_reg[24]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[24] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[24] .power_up = "low";

dffeas \phi_int_arr_reg[23] (
	.clk(clk),
	.d(pipeline_dffe_23),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_int_arr_reg[23]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[23] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[23] .power_up = "low";

dffeas \phi_int_arr_reg[22] (
	.clk(clk),
	.d(pipeline_dffe_22),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_int_arr_reg[22]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[22] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[22] .power_up = "low";

dffeas \phi_int_arr_reg[21] (
	.clk(clk),
	.d(pipeline_dffe_21),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_int_arr_reg[21]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[21] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[21] .power_up = "low";

dffeas \phi_int_arr_reg[20] (
	.clk(clk),
	.d(pipeline_dffe_20),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_int_arr_reg[20]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[20] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[20] .power_up = "low";

dffeas \phi_int_arr_reg[19] (
	.clk(clk),
	.d(pipeline_dffe_19),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_int_arr_reg[19]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[19] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[19] .power_up = "low";

dffeas \phi_int_arr_reg[18] (
	.clk(clk),
	.d(pipeline_dffe_18),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_int_arr_reg[18]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[18] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[18] .power_up = "low";

dffeas \phi_int_arr_reg[17] (
	.clk(clk),
	.d(pipeline_dffe_17),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_int_arr_reg[17]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[17] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[17] .power_up = "low";

dffeas \phi_int_arr_reg[16] (
	.clk(clk),
	.d(pipeline_dffe_16),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_int_arr_reg[16]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[16] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[16] .power_up = "low";

dffeas \phi_int_arr_reg[15] (
	.clk(clk),
	.d(pipeline_dffe_15),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_int_arr_reg[15]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[15] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[15] .power_up = "low";

dffeas \phi_int_arr_reg[14] (
	.clk(clk),
	.d(pipeline_dffe_14),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_int_arr_reg[14]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[14] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[14] .power_up = "low";

dffeas \phi_int_arr_reg[13] (
	.clk(clk),
	.d(pipeline_dffe_13),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_int_arr_reg[13]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[13] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[13] .power_up = "low";

dffeas \phi_int_arr_reg[12] (
	.clk(clk),
	.d(pipeline_dffe_12),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_int_arr_reg[12]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[12] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[12] .power_up = "low";

dffeas \phi_int_arr_reg[11] (
	.clk(clk),
	.d(pipeline_dffe_11),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_int_arr_reg[11]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[11] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[11] .power_up = "low";

dffeas \phi_int_arr_reg[10] (
	.clk(clk),
	.d(pipeline_dffe_10),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_int_arr_reg[10]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[10] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[10] .power_up = "low";

dffeas \phi_int_arr_reg[9] (
	.clk(clk),
	.d(pipeline_dffe_9),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_int_arr_reg[9]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[9] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[9] .power_up = "low";

dffeas \phi_int_arr_reg[8] (
	.clk(clk),
	.d(pipeline_dffe_8),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_int_arr_reg[8]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[8] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[8] .power_up = "low";

dffeas \phi_int_arr_reg[7] (
	.clk(clk),
	.d(pipeline_dffe_7),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_int_arr_reg[7]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[7] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[7] .power_up = "low";

dffeas \phi_int_arr_reg[6] (
	.clk(clk),
	.d(pipeline_dffe_6),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_int_arr_reg[6]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[6] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[6] .power_up = "low";

dffeas \phi_int_arr_reg[5] (
	.clk(clk),
	.d(pipeline_dffe_5),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_int_arr_reg[5]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[5] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[5] .power_up = "low";

dffeas \phi_int_arr_reg[4] (
	.clk(clk),
	.d(pipeline_dffe_4),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_int_arr_reg[4]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[4] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[4] .power_up = "low";

dffeas \phi_int_arr_reg[3] (
	.clk(clk),
	.d(pipeline_dffe_3),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_int_arr_reg[3]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[3] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[3] .power_up = "low";

dffeas \phi_int_arr_reg[2] (
	.clk(clk),
	.d(pipeline_dffe_2),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_int_arr_reg[2]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[2] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[2] .power_up = "low";

dffeas \phi_int_arr_reg[1] (
	.clk(clk),
	.d(pipeline_dffe_1),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_int_arr_reg[1]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[1] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[1] .power_up = "low";

dffeas \phi_int_arr_reg[0] (
	.clk(clk),
	.d(pipeline_dffe_0),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_int_arr_reg[0]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[0] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[0] .power_up = "low";

endmodule

module DDS_48_v1_lpm_add_sub_1 (
	phi_int_arr_reg_32,
	phi_int_arr_reg_33,
	phi_int_arr_reg_34,
	phi_int_arr_reg_35,
	phi_int_arr_reg_36,
	phi_int_arr_reg_37,
	phi_int_arr_reg_38,
	phi_int_arr_reg_39,
	phi_int_arr_reg_40,
	phi_int_arr_reg_41,
	phi_int_arr_reg_42,
	phi_int_arr_reg_43,
	phi_int_arr_reg_44,
	phi_int_arr_reg_47,
	phi_int_arr_reg_31,
	phi_int_arr_reg_45,
	phi_int_arr_reg_46,
	phi_int_arr_reg_30,
	phi_int_arr_reg_29,
	phi_int_arr_reg_28,
	phi_int_arr_reg_27,
	phi_int_arr_reg_26,
	phi_int_arr_reg_25,
	phi_int_arr_reg_24,
	phi_int_arr_reg_23,
	phi_int_arr_reg_22,
	phi_int_arr_reg_21,
	phi_int_arr_reg_20,
	phi_int_arr_reg_19,
	phi_int_arr_reg_18,
	phi_int_arr_reg_17,
	phi_int_arr_reg_16,
	phi_int_arr_reg_15,
	phi_int_arr_reg_14,
	phi_int_arr_reg_13,
	phi_int_arr_reg_12,
	phi_int_arr_reg_11,
	phi_int_arr_reg_10,
	phi_int_arr_reg_9,
	phi_int_arr_reg_8,
	phi_int_arr_reg_7,
	phi_int_arr_reg_6,
	phi_int_arr_reg_5,
	phi_int_arr_reg_4,
	phi_int_arr_reg_3,
	phi_int_arr_reg_2,
	phi_int_arr_reg_1,
	phi_int_arr_reg_0,
	pipeline_dffe_32,
	pipeline_dffe_33,
	pipeline_dffe_34,
	pipeline_dffe_35,
	pipeline_dffe_36,
	pipeline_dffe_37,
	pipeline_dffe_38,
	pipeline_dffe_39,
	pipeline_dffe_40,
	pipeline_dffe_41,
	pipeline_dffe_42,
	pipeline_dffe_43,
	pipeline_dffe_44,
	pipeline_dffe_47,
	pipeline_dffe_31,
	pipeline_dffe_45,
	pipeline_dffe_46,
	pipeline_dffe_30,
	pipeline_dffe_29,
	pipeline_dffe_28,
	pipeline_dffe_27,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	phi_int_arr_reg_32;
input 	phi_int_arr_reg_33;
input 	phi_int_arr_reg_34;
input 	phi_int_arr_reg_35;
input 	phi_int_arr_reg_36;
input 	phi_int_arr_reg_37;
input 	phi_int_arr_reg_38;
input 	phi_int_arr_reg_39;
input 	phi_int_arr_reg_40;
input 	phi_int_arr_reg_41;
input 	phi_int_arr_reg_42;
input 	phi_int_arr_reg_43;
input 	phi_int_arr_reg_44;
input 	phi_int_arr_reg_47;
input 	phi_int_arr_reg_31;
input 	phi_int_arr_reg_45;
input 	phi_int_arr_reg_46;
input 	phi_int_arr_reg_30;
input 	phi_int_arr_reg_29;
input 	phi_int_arr_reg_28;
input 	phi_int_arr_reg_27;
input 	phi_int_arr_reg_26;
input 	phi_int_arr_reg_25;
input 	phi_int_arr_reg_24;
input 	phi_int_arr_reg_23;
input 	phi_int_arr_reg_22;
input 	phi_int_arr_reg_21;
input 	phi_int_arr_reg_20;
input 	phi_int_arr_reg_19;
input 	phi_int_arr_reg_18;
input 	phi_int_arr_reg_17;
input 	phi_int_arr_reg_16;
input 	phi_int_arr_reg_15;
input 	phi_int_arr_reg_14;
input 	phi_int_arr_reg_13;
input 	phi_int_arr_reg_12;
input 	phi_int_arr_reg_11;
input 	phi_int_arr_reg_10;
input 	phi_int_arr_reg_9;
input 	phi_int_arr_reg_8;
input 	phi_int_arr_reg_7;
input 	phi_int_arr_reg_6;
input 	phi_int_arr_reg_5;
input 	phi_int_arr_reg_4;
input 	phi_int_arr_reg_3;
input 	phi_int_arr_reg_2;
input 	phi_int_arr_reg_1;
input 	phi_int_arr_reg_0;
output 	pipeline_dffe_32;
output 	pipeline_dffe_33;
output 	pipeline_dffe_34;
output 	pipeline_dffe_35;
output 	pipeline_dffe_36;
output 	pipeline_dffe_37;
output 	pipeline_dffe_38;
output 	pipeline_dffe_39;
output 	pipeline_dffe_40;
output 	pipeline_dffe_41;
output 	pipeline_dffe_42;
output 	pipeline_dffe_43;
output 	pipeline_dffe_44;
output 	pipeline_dffe_47;
output 	pipeline_dffe_31;
output 	pipeline_dffe_45;
output 	pipeline_dffe_46;
output 	pipeline_dffe_30;
output 	pipeline_dffe_29;
output 	pipeline_dffe_28;
output 	pipeline_dffe_27;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



DDS_48_v1_add_sub_qmh auto_generated(
	.phi_int_arr_reg_32(phi_int_arr_reg_32),
	.phi_int_arr_reg_33(phi_int_arr_reg_33),
	.phi_int_arr_reg_34(phi_int_arr_reg_34),
	.phi_int_arr_reg_35(phi_int_arr_reg_35),
	.phi_int_arr_reg_36(phi_int_arr_reg_36),
	.phi_int_arr_reg_37(phi_int_arr_reg_37),
	.phi_int_arr_reg_38(phi_int_arr_reg_38),
	.phi_int_arr_reg_39(phi_int_arr_reg_39),
	.phi_int_arr_reg_40(phi_int_arr_reg_40),
	.phi_int_arr_reg_41(phi_int_arr_reg_41),
	.phi_int_arr_reg_42(phi_int_arr_reg_42),
	.phi_int_arr_reg_43(phi_int_arr_reg_43),
	.phi_int_arr_reg_44(phi_int_arr_reg_44),
	.phi_int_arr_reg_47(phi_int_arr_reg_47),
	.phi_int_arr_reg_31(phi_int_arr_reg_31),
	.phi_int_arr_reg_45(phi_int_arr_reg_45),
	.phi_int_arr_reg_46(phi_int_arr_reg_46),
	.phi_int_arr_reg_30(phi_int_arr_reg_30),
	.phi_int_arr_reg_29(phi_int_arr_reg_29),
	.phi_int_arr_reg_28(phi_int_arr_reg_28),
	.phi_int_arr_reg_27(phi_int_arr_reg_27),
	.phi_int_arr_reg_26(phi_int_arr_reg_26),
	.phi_int_arr_reg_25(phi_int_arr_reg_25),
	.phi_int_arr_reg_24(phi_int_arr_reg_24),
	.phi_int_arr_reg_23(phi_int_arr_reg_23),
	.phi_int_arr_reg_22(phi_int_arr_reg_22),
	.phi_int_arr_reg_21(phi_int_arr_reg_21),
	.phi_int_arr_reg_20(phi_int_arr_reg_20),
	.phi_int_arr_reg_19(phi_int_arr_reg_19),
	.phi_int_arr_reg_18(phi_int_arr_reg_18),
	.phi_int_arr_reg_17(phi_int_arr_reg_17),
	.phi_int_arr_reg_16(phi_int_arr_reg_16),
	.phi_int_arr_reg_15(phi_int_arr_reg_15),
	.phi_int_arr_reg_14(phi_int_arr_reg_14),
	.phi_int_arr_reg_13(phi_int_arr_reg_13),
	.phi_int_arr_reg_12(phi_int_arr_reg_12),
	.phi_int_arr_reg_11(phi_int_arr_reg_11),
	.phi_int_arr_reg_10(phi_int_arr_reg_10),
	.phi_int_arr_reg_9(phi_int_arr_reg_9),
	.phi_int_arr_reg_8(phi_int_arr_reg_8),
	.phi_int_arr_reg_7(phi_int_arr_reg_7),
	.phi_int_arr_reg_6(phi_int_arr_reg_6),
	.phi_int_arr_reg_5(phi_int_arr_reg_5),
	.phi_int_arr_reg_4(phi_int_arr_reg_4),
	.phi_int_arr_reg_3(phi_int_arr_reg_3),
	.phi_int_arr_reg_2(phi_int_arr_reg_2),
	.phi_int_arr_reg_1(phi_int_arr_reg_1),
	.phi_int_arr_reg_0(phi_int_arr_reg_0),
	.pipeline_dffe_32(pipeline_dffe_32),
	.pipeline_dffe_33(pipeline_dffe_33),
	.pipeline_dffe_34(pipeline_dffe_34),
	.pipeline_dffe_35(pipeline_dffe_35),
	.pipeline_dffe_36(pipeline_dffe_36),
	.pipeline_dffe_37(pipeline_dffe_37),
	.pipeline_dffe_38(pipeline_dffe_38),
	.pipeline_dffe_39(pipeline_dffe_39),
	.pipeline_dffe_40(pipeline_dffe_40),
	.pipeline_dffe_41(pipeline_dffe_41),
	.pipeline_dffe_42(pipeline_dffe_42),
	.pipeline_dffe_43(pipeline_dffe_43),
	.pipeline_dffe_44(pipeline_dffe_44),
	.pipeline_dffe_47(pipeline_dffe_47),
	.pipeline_dffe_31(pipeline_dffe_31),
	.pipeline_dffe_45(pipeline_dffe_45),
	.pipeline_dffe_46(pipeline_dffe_46),
	.pipeline_dffe_30(pipeline_dffe_30),
	.pipeline_dffe_29(pipeline_dffe_29),
	.pipeline_dffe_28(pipeline_dffe_28),
	.pipeline_dffe_27(pipeline_dffe_27),
	.clock(clock),
	.reset_n(reset_n),
	.clken(clken));

endmodule

module DDS_48_v1_add_sub_qmh (
	phi_int_arr_reg_32,
	phi_int_arr_reg_33,
	phi_int_arr_reg_34,
	phi_int_arr_reg_35,
	phi_int_arr_reg_36,
	phi_int_arr_reg_37,
	phi_int_arr_reg_38,
	phi_int_arr_reg_39,
	phi_int_arr_reg_40,
	phi_int_arr_reg_41,
	phi_int_arr_reg_42,
	phi_int_arr_reg_43,
	phi_int_arr_reg_44,
	phi_int_arr_reg_47,
	phi_int_arr_reg_31,
	phi_int_arr_reg_45,
	phi_int_arr_reg_46,
	phi_int_arr_reg_30,
	phi_int_arr_reg_29,
	phi_int_arr_reg_28,
	phi_int_arr_reg_27,
	phi_int_arr_reg_26,
	phi_int_arr_reg_25,
	phi_int_arr_reg_24,
	phi_int_arr_reg_23,
	phi_int_arr_reg_22,
	phi_int_arr_reg_21,
	phi_int_arr_reg_20,
	phi_int_arr_reg_19,
	phi_int_arr_reg_18,
	phi_int_arr_reg_17,
	phi_int_arr_reg_16,
	phi_int_arr_reg_15,
	phi_int_arr_reg_14,
	phi_int_arr_reg_13,
	phi_int_arr_reg_12,
	phi_int_arr_reg_11,
	phi_int_arr_reg_10,
	phi_int_arr_reg_9,
	phi_int_arr_reg_8,
	phi_int_arr_reg_7,
	phi_int_arr_reg_6,
	phi_int_arr_reg_5,
	phi_int_arr_reg_4,
	phi_int_arr_reg_3,
	phi_int_arr_reg_2,
	phi_int_arr_reg_1,
	phi_int_arr_reg_0,
	pipeline_dffe_32,
	pipeline_dffe_33,
	pipeline_dffe_34,
	pipeline_dffe_35,
	pipeline_dffe_36,
	pipeline_dffe_37,
	pipeline_dffe_38,
	pipeline_dffe_39,
	pipeline_dffe_40,
	pipeline_dffe_41,
	pipeline_dffe_42,
	pipeline_dffe_43,
	pipeline_dffe_44,
	pipeline_dffe_47,
	pipeline_dffe_31,
	pipeline_dffe_45,
	pipeline_dffe_46,
	pipeline_dffe_30,
	pipeline_dffe_29,
	pipeline_dffe_28,
	pipeline_dffe_27,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	phi_int_arr_reg_32;
input 	phi_int_arr_reg_33;
input 	phi_int_arr_reg_34;
input 	phi_int_arr_reg_35;
input 	phi_int_arr_reg_36;
input 	phi_int_arr_reg_37;
input 	phi_int_arr_reg_38;
input 	phi_int_arr_reg_39;
input 	phi_int_arr_reg_40;
input 	phi_int_arr_reg_41;
input 	phi_int_arr_reg_42;
input 	phi_int_arr_reg_43;
input 	phi_int_arr_reg_44;
input 	phi_int_arr_reg_47;
input 	phi_int_arr_reg_31;
input 	phi_int_arr_reg_45;
input 	phi_int_arr_reg_46;
input 	phi_int_arr_reg_30;
input 	phi_int_arr_reg_29;
input 	phi_int_arr_reg_28;
input 	phi_int_arr_reg_27;
input 	phi_int_arr_reg_26;
input 	phi_int_arr_reg_25;
input 	phi_int_arr_reg_24;
input 	phi_int_arr_reg_23;
input 	phi_int_arr_reg_22;
input 	phi_int_arr_reg_21;
input 	phi_int_arr_reg_20;
input 	phi_int_arr_reg_19;
input 	phi_int_arr_reg_18;
input 	phi_int_arr_reg_17;
input 	phi_int_arr_reg_16;
input 	phi_int_arr_reg_15;
input 	phi_int_arr_reg_14;
input 	phi_int_arr_reg_13;
input 	phi_int_arr_reg_12;
input 	phi_int_arr_reg_11;
input 	phi_int_arr_reg_10;
input 	phi_int_arr_reg_9;
input 	phi_int_arr_reg_8;
input 	phi_int_arr_reg_7;
input 	phi_int_arr_reg_6;
input 	phi_int_arr_reg_5;
input 	phi_int_arr_reg_4;
input 	phi_int_arr_reg_3;
input 	phi_int_arr_reg_2;
input 	phi_int_arr_reg_1;
input 	phi_int_arr_reg_0;
output 	pipeline_dffe_32;
output 	pipeline_dffe_33;
output 	pipeline_dffe_34;
output 	pipeline_dffe_35;
output 	pipeline_dffe_36;
output 	pipeline_dffe_37;
output 	pipeline_dffe_38;
output 	pipeline_dffe_39;
output 	pipeline_dffe_40;
output 	pipeline_dffe_41;
output 	pipeline_dffe_42;
output 	pipeline_dffe_43;
output 	pipeline_dffe_44;
output 	pipeline_dffe_47;
output 	pipeline_dffe_31;
output 	pipeline_dffe_45;
output 	pipeline_dffe_46;
output 	pipeline_dffe_30;
output 	pipeline_dffe_29;
output 	pipeline_dffe_28;
output 	pipeline_dffe_27;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \op_1~189_sumout ;
wire \pipeline_dffe[0]~q ;
wire \op_1~190 ;
wire \op_1~185_sumout ;
wire \pipeline_dffe[1]~q ;
wire \op_1~186 ;
wire \op_1~181_sumout ;
wire \pipeline_dffe[2]~q ;
wire \op_1~182 ;
wire \op_1~177_sumout ;
wire \pipeline_dffe[3]~q ;
wire \op_1~178 ;
wire \op_1~173_sumout ;
wire \pipeline_dffe[4]~q ;
wire \op_1~174 ;
wire \op_1~169_sumout ;
wire \pipeline_dffe[5]~q ;
wire \op_1~170 ;
wire \op_1~165_sumout ;
wire \pipeline_dffe[6]~q ;
wire \op_1~166 ;
wire \op_1~161_sumout ;
wire \pipeline_dffe[7]~q ;
wire \op_1~162 ;
wire \op_1~157_sumout ;
wire \pipeline_dffe[8]~q ;
wire \op_1~158 ;
wire \op_1~153_sumout ;
wire \pipeline_dffe[9]~q ;
wire \op_1~154 ;
wire \op_1~149_sumout ;
wire \pipeline_dffe[10]~q ;
wire \op_1~150 ;
wire \op_1~145_sumout ;
wire \pipeline_dffe[11]~q ;
wire \op_1~146 ;
wire \op_1~141_sumout ;
wire \pipeline_dffe[12]~q ;
wire \op_1~142 ;
wire \op_1~137_sumout ;
wire \pipeline_dffe[13]~q ;
wire \op_1~138 ;
wire \op_1~133_sumout ;
wire \pipeline_dffe[14]~q ;
wire \op_1~134 ;
wire \op_1~129_sumout ;
wire \pipeline_dffe[15]~q ;
wire \op_1~130 ;
wire \op_1~125_sumout ;
wire \pipeline_dffe[16]~q ;
wire \op_1~126 ;
wire \op_1~121_sumout ;
wire \pipeline_dffe[17]~q ;
wire \op_1~122 ;
wire \op_1~117_sumout ;
wire \pipeline_dffe[18]~q ;
wire \op_1~118 ;
wire \op_1~113_sumout ;
wire \pipeline_dffe[19]~q ;
wire \op_1~114 ;
wire \op_1~109_sumout ;
wire \pipeline_dffe[20]~q ;
wire \op_1~110 ;
wire \op_1~105_sumout ;
wire \pipeline_dffe[21]~q ;
wire \op_1~106 ;
wire \op_1~101_sumout ;
wire \pipeline_dffe[22]~q ;
wire \op_1~102 ;
wire \op_1~97_sumout ;
wire \pipeline_dffe[23]~q ;
wire \op_1~98 ;
wire \op_1~93_sumout ;
wire \pipeline_dffe[24]~q ;
wire \op_1~94 ;
wire \op_1~89_sumout ;
wire \pipeline_dffe[25]~q ;
wire \op_1~90 ;
wire \op_1~85_sumout ;
wire \pipeline_dffe[26]~q ;
wire \op_1~86 ;
wire \op_1~82 ;
wire \op_1~78 ;
wire \op_1~74 ;
wire \op_1~70 ;
wire \op_1~58 ;
wire \op_1~1_sumout ;
wire \op_1~2 ;
wire \op_1~5_sumout ;
wire \op_1~6 ;
wire \op_1~9_sumout ;
wire \op_1~10 ;
wire \op_1~13_sumout ;
wire \op_1~14 ;
wire \op_1~17_sumout ;
wire \op_1~18 ;
wire \op_1~21_sumout ;
wire \op_1~22 ;
wire \op_1~25_sumout ;
wire \op_1~26 ;
wire \op_1~29_sumout ;
wire \op_1~30 ;
wire \op_1~33_sumout ;
wire \op_1~34 ;
wire \op_1~37_sumout ;
wire \op_1~38 ;
wire \op_1~41_sumout ;
wire \op_1~42 ;
wire \op_1~45_sumout ;
wire \op_1~46 ;
wire \op_1~49_sumout ;
wire \op_1~50 ;
wire \op_1~62 ;
wire \op_1~66 ;
wire \op_1~53_sumout ;
wire \op_1~57_sumout ;
wire \op_1~61_sumout ;
wire \op_1~65_sumout ;
wire \op_1~69_sumout ;
wire \op_1~73_sumout ;
wire \op_1~77_sumout ;
wire \op_1~81_sumout ;


dffeas \pipeline_dffe[32] (
	.clk(clock),
	.d(\op_1~1_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_32),
	.prn(vcc));
defparam \pipeline_dffe[32] .is_wysiwyg = "true";
defparam \pipeline_dffe[32] .power_up = "low";

dffeas \pipeline_dffe[33] (
	.clk(clock),
	.d(\op_1~5_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_33),
	.prn(vcc));
defparam \pipeline_dffe[33] .is_wysiwyg = "true";
defparam \pipeline_dffe[33] .power_up = "low";

dffeas \pipeline_dffe[34] (
	.clk(clock),
	.d(\op_1~9_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_34),
	.prn(vcc));
defparam \pipeline_dffe[34] .is_wysiwyg = "true";
defparam \pipeline_dffe[34] .power_up = "low";

dffeas \pipeline_dffe[35] (
	.clk(clock),
	.d(\op_1~13_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_35),
	.prn(vcc));
defparam \pipeline_dffe[35] .is_wysiwyg = "true";
defparam \pipeline_dffe[35] .power_up = "low";

dffeas \pipeline_dffe[36] (
	.clk(clock),
	.d(\op_1~17_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_36),
	.prn(vcc));
defparam \pipeline_dffe[36] .is_wysiwyg = "true";
defparam \pipeline_dffe[36] .power_up = "low";

dffeas \pipeline_dffe[37] (
	.clk(clock),
	.d(\op_1~21_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_37),
	.prn(vcc));
defparam \pipeline_dffe[37] .is_wysiwyg = "true";
defparam \pipeline_dffe[37] .power_up = "low";

dffeas \pipeline_dffe[38] (
	.clk(clock),
	.d(\op_1~25_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_38),
	.prn(vcc));
defparam \pipeline_dffe[38] .is_wysiwyg = "true";
defparam \pipeline_dffe[38] .power_up = "low";

dffeas \pipeline_dffe[39] (
	.clk(clock),
	.d(\op_1~29_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_39),
	.prn(vcc));
defparam \pipeline_dffe[39] .is_wysiwyg = "true";
defparam \pipeline_dffe[39] .power_up = "low";

dffeas \pipeline_dffe[40] (
	.clk(clock),
	.d(\op_1~33_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_40),
	.prn(vcc));
defparam \pipeline_dffe[40] .is_wysiwyg = "true";
defparam \pipeline_dffe[40] .power_up = "low";

dffeas \pipeline_dffe[41] (
	.clk(clock),
	.d(\op_1~37_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_41),
	.prn(vcc));
defparam \pipeline_dffe[41] .is_wysiwyg = "true";
defparam \pipeline_dffe[41] .power_up = "low";

dffeas \pipeline_dffe[42] (
	.clk(clock),
	.d(\op_1~41_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_42),
	.prn(vcc));
defparam \pipeline_dffe[42] .is_wysiwyg = "true";
defparam \pipeline_dffe[42] .power_up = "low";

dffeas \pipeline_dffe[43] (
	.clk(clock),
	.d(\op_1~45_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_43),
	.prn(vcc));
defparam \pipeline_dffe[43] .is_wysiwyg = "true";
defparam \pipeline_dffe[43] .power_up = "low";

dffeas \pipeline_dffe[44] (
	.clk(clock),
	.d(\op_1~49_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_44),
	.prn(vcc));
defparam \pipeline_dffe[44] .is_wysiwyg = "true";
defparam \pipeline_dffe[44] .power_up = "low";

dffeas \pipeline_dffe[47] (
	.clk(clock),
	.d(\op_1~53_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_47),
	.prn(vcc));
defparam \pipeline_dffe[47] .is_wysiwyg = "true";
defparam \pipeline_dffe[47] .power_up = "low";

dffeas \pipeline_dffe[31] (
	.clk(clock),
	.d(\op_1~57_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_31),
	.prn(vcc));
defparam \pipeline_dffe[31] .is_wysiwyg = "true";
defparam \pipeline_dffe[31] .power_up = "low";

dffeas \pipeline_dffe[45] (
	.clk(clock),
	.d(\op_1~61_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_45),
	.prn(vcc));
defparam \pipeline_dffe[45] .is_wysiwyg = "true";
defparam \pipeline_dffe[45] .power_up = "low";

dffeas \pipeline_dffe[46] (
	.clk(clock),
	.d(\op_1~65_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_46),
	.prn(vcc));
defparam \pipeline_dffe[46] .is_wysiwyg = "true";
defparam \pipeline_dffe[46] .power_up = "low";

dffeas \pipeline_dffe[30] (
	.clk(clock),
	.d(\op_1~69_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_30),
	.prn(vcc));
defparam \pipeline_dffe[30] .is_wysiwyg = "true";
defparam \pipeline_dffe[30] .power_up = "low";

dffeas \pipeline_dffe[29] (
	.clk(clock),
	.d(\op_1~73_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_29),
	.prn(vcc));
defparam \pipeline_dffe[29] .is_wysiwyg = "true";
defparam \pipeline_dffe[29] .power_up = "low";

dffeas \pipeline_dffe[28] (
	.clk(clock),
	.d(\op_1~77_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_28),
	.prn(vcc));
defparam \pipeline_dffe[28] .is_wysiwyg = "true";
defparam \pipeline_dffe[28] .power_up = "low";

dffeas \pipeline_dffe[27] (
	.clk(clock),
	.d(\op_1~81_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_27),
	.prn(vcc));
defparam \pipeline_dffe[27] .is_wysiwyg = "true";
defparam \pipeline_dffe[27] .power_up = "low";

arriav_lcell_comb \op_1~189 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_0),
	.datae(gnd),
	.dataf(!\pipeline_dffe[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~189_sumout ),
	.cout(\op_1~190 ),
	.shareout());
defparam \op_1~189 .extended_lut = "off";
defparam \op_1~189 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~189 .shared_arith = "off";

dffeas \pipeline_dffe[0] (
	.clk(clock),
	.d(\op_1~189_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\pipeline_dffe[0]~q ),
	.prn(vcc));
defparam \pipeline_dffe[0] .is_wysiwyg = "true";
defparam \pipeline_dffe[0] .power_up = "low";

arriav_lcell_comb \op_1~185 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_1),
	.datae(gnd),
	.dataf(!\pipeline_dffe[1]~q ),
	.datag(gnd),
	.cin(\op_1~190 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~185_sumout ),
	.cout(\op_1~186 ),
	.shareout());
defparam \op_1~185 .extended_lut = "off";
defparam \op_1~185 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~185 .shared_arith = "off";

dffeas \pipeline_dffe[1] (
	.clk(clock),
	.d(\op_1~185_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\pipeline_dffe[1]~q ),
	.prn(vcc));
defparam \pipeline_dffe[1] .is_wysiwyg = "true";
defparam \pipeline_dffe[1] .power_up = "low";

arriav_lcell_comb \op_1~181 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_2),
	.datae(gnd),
	.dataf(!\pipeline_dffe[2]~q ),
	.datag(gnd),
	.cin(\op_1~186 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~181_sumout ),
	.cout(\op_1~182 ),
	.shareout());
defparam \op_1~181 .extended_lut = "off";
defparam \op_1~181 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~181 .shared_arith = "off";

dffeas \pipeline_dffe[2] (
	.clk(clock),
	.d(\op_1~181_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\pipeline_dffe[2]~q ),
	.prn(vcc));
defparam \pipeline_dffe[2] .is_wysiwyg = "true";
defparam \pipeline_dffe[2] .power_up = "low";

arriav_lcell_comb \op_1~177 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_3),
	.datae(gnd),
	.dataf(!\pipeline_dffe[3]~q ),
	.datag(gnd),
	.cin(\op_1~182 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~177_sumout ),
	.cout(\op_1~178 ),
	.shareout());
defparam \op_1~177 .extended_lut = "off";
defparam \op_1~177 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~177 .shared_arith = "off";

dffeas \pipeline_dffe[3] (
	.clk(clock),
	.d(\op_1~177_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\pipeline_dffe[3]~q ),
	.prn(vcc));
defparam \pipeline_dffe[3] .is_wysiwyg = "true";
defparam \pipeline_dffe[3] .power_up = "low";

arriav_lcell_comb \op_1~173 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_4),
	.datae(gnd),
	.dataf(!\pipeline_dffe[4]~q ),
	.datag(gnd),
	.cin(\op_1~178 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~173_sumout ),
	.cout(\op_1~174 ),
	.shareout());
defparam \op_1~173 .extended_lut = "off";
defparam \op_1~173 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~173 .shared_arith = "off";

dffeas \pipeline_dffe[4] (
	.clk(clock),
	.d(\op_1~173_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\pipeline_dffe[4]~q ),
	.prn(vcc));
defparam \pipeline_dffe[4] .is_wysiwyg = "true";
defparam \pipeline_dffe[4] .power_up = "low";

arriav_lcell_comb \op_1~169 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_5),
	.datae(gnd),
	.dataf(!\pipeline_dffe[5]~q ),
	.datag(gnd),
	.cin(\op_1~174 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~169_sumout ),
	.cout(\op_1~170 ),
	.shareout());
defparam \op_1~169 .extended_lut = "off";
defparam \op_1~169 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~169 .shared_arith = "off";

dffeas \pipeline_dffe[5] (
	.clk(clock),
	.d(\op_1~169_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\pipeline_dffe[5]~q ),
	.prn(vcc));
defparam \pipeline_dffe[5] .is_wysiwyg = "true";
defparam \pipeline_dffe[5] .power_up = "low";

arriav_lcell_comb \op_1~165 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_6),
	.datae(gnd),
	.dataf(!\pipeline_dffe[6]~q ),
	.datag(gnd),
	.cin(\op_1~170 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~165_sumout ),
	.cout(\op_1~166 ),
	.shareout());
defparam \op_1~165 .extended_lut = "off";
defparam \op_1~165 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~165 .shared_arith = "off";

dffeas \pipeline_dffe[6] (
	.clk(clock),
	.d(\op_1~165_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\pipeline_dffe[6]~q ),
	.prn(vcc));
defparam \pipeline_dffe[6] .is_wysiwyg = "true";
defparam \pipeline_dffe[6] .power_up = "low";

arriav_lcell_comb \op_1~161 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_7),
	.datae(gnd),
	.dataf(!\pipeline_dffe[7]~q ),
	.datag(gnd),
	.cin(\op_1~166 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~161_sumout ),
	.cout(\op_1~162 ),
	.shareout());
defparam \op_1~161 .extended_lut = "off";
defparam \op_1~161 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~161 .shared_arith = "off";

dffeas \pipeline_dffe[7] (
	.clk(clock),
	.d(\op_1~161_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\pipeline_dffe[7]~q ),
	.prn(vcc));
defparam \pipeline_dffe[7] .is_wysiwyg = "true";
defparam \pipeline_dffe[7] .power_up = "low";

arriav_lcell_comb \op_1~157 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_8),
	.datae(gnd),
	.dataf(!\pipeline_dffe[8]~q ),
	.datag(gnd),
	.cin(\op_1~162 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~157_sumout ),
	.cout(\op_1~158 ),
	.shareout());
defparam \op_1~157 .extended_lut = "off";
defparam \op_1~157 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~157 .shared_arith = "off";

dffeas \pipeline_dffe[8] (
	.clk(clock),
	.d(\op_1~157_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\pipeline_dffe[8]~q ),
	.prn(vcc));
defparam \pipeline_dffe[8] .is_wysiwyg = "true";
defparam \pipeline_dffe[8] .power_up = "low";

arriav_lcell_comb \op_1~153 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_9),
	.datae(gnd),
	.dataf(!\pipeline_dffe[9]~q ),
	.datag(gnd),
	.cin(\op_1~158 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~153_sumout ),
	.cout(\op_1~154 ),
	.shareout());
defparam \op_1~153 .extended_lut = "off";
defparam \op_1~153 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~153 .shared_arith = "off";

dffeas \pipeline_dffe[9] (
	.clk(clock),
	.d(\op_1~153_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\pipeline_dffe[9]~q ),
	.prn(vcc));
defparam \pipeline_dffe[9] .is_wysiwyg = "true";
defparam \pipeline_dffe[9] .power_up = "low";

arriav_lcell_comb \op_1~149 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_10),
	.datae(gnd),
	.dataf(!\pipeline_dffe[10]~q ),
	.datag(gnd),
	.cin(\op_1~154 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~149_sumout ),
	.cout(\op_1~150 ),
	.shareout());
defparam \op_1~149 .extended_lut = "off";
defparam \op_1~149 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~149 .shared_arith = "off";

dffeas \pipeline_dffe[10] (
	.clk(clock),
	.d(\op_1~149_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\pipeline_dffe[10]~q ),
	.prn(vcc));
defparam \pipeline_dffe[10] .is_wysiwyg = "true";
defparam \pipeline_dffe[10] .power_up = "low";

arriav_lcell_comb \op_1~145 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_11),
	.datae(gnd),
	.dataf(!\pipeline_dffe[11]~q ),
	.datag(gnd),
	.cin(\op_1~150 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~145_sumout ),
	.cout(\op_1~146 ),
	.shareout());
defparam \op_1~145 .extended_lut = "off";
defparam \op_1~145 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~145 .shared_arith = "off";

dffeas \pipeline_dffe[11] (
	.clk(clock),
	.d(\op_1~145_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\pipeline_dffe[11]~q ),
	.prn(vcc));
defparam \pipeline_dffe[11] .is_wysiwyg = "true";
defparam \pipeline_dffe[11] .power_up = "low";

arriav_lcell_comb \op_1~141 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_12),
	.datae(gnd),
	.dataf(!\pipeline_dffe[12]~q ),
	.datag(gnd),
	.cin(\op_1~146 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~141_sumout ),
	.cout(\op_1~142 ),
	.shareout());
defparam \op_1~141 .extended_lut = "off";
defparam \op_1~141 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~141 .shared_arith = "off";

dffeas \pipeline_dffe[12] (
	.clk(clock),
	.d(\op_1~141_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\pipeline_dffe[12]~q ),
	.prn(vcc));
defparam \pipeline_dffe[12] .is_wysiwyg = "true";
defparam \pipeline_dffe[12] .power_up = "low";

arriav_lcell_comb \op_1~137 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_13),
	.datae(gnd),
	.dataf(!\pipeline_dffe[13]~q ),
	.datag(gnd),
	.cin(\op_1~142 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~137_sumout ),
	.cout(\op_1~138 ),
	.shareout());
defparam \op_1~137 .extended_lut = "off";
defparam \op_1~137 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~137 .shared_arith = "off";

dffeas \pipeline_dffe[13] (
	.clk(clock),
	.d(\op_1~137_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\pipeline_dffe[13]~q ),
	.prn(vcc));
defparam \pipeline_dffe[13] .is_wysiwyg = "true";
defparam \pipeline_dffe[13] .power_up = "low";

arriav_lcell_comb \op_1~133 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_14),
	.datae(gnd),
	.dataf(!\pipeline_dffe[14]~q ),
	.datag(gnd),
	.cin(\op_1~138 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~133_sumout ),
	.cout(\op_1~134 ),
	.shareout());
defparam \op_1~133 .extended_lut = "off";
defparam \op_1~133 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~133 .shared_arith = "off";

dffeas \pipeline_dffe[14] (
	.clk(clock),
	.d(\op_1~133_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\pipeline_dffe[14]~q ),
	.prn(vcc));
defparam \pipeline_dffe[14] .is_wysiwyg = "true";
defparam \pipeline_dffe[14] .power_up = "low";

arriav_lcell_comb \op_1~129 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_15),
	.datae(gnd),
	.dataf(!\pipeline_dffe[15]~q ),
	.datag(gnd),
	.cin(\op_1~134 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~129_sumout ),
	.cout(\op_1~130 ),
	.shareout());
defparam \op_1~129 .extended_lut = "off";
defparam \op_1~129 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~129 .shared_arith = "off";

dffeas \pipeline_dffe[15] (
	.clk(clock),
	.d(\op_1~129_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\pipeline_dffe[15]~q ),
	.prn(vcc));
defparam \pipeline_dffe[15] .is_wysiwyg = "true";
defparam \pipeline_dffe[15] .power_up = "low";

arriav_lcell_comb \op_1~125 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_16),
	.datae(gnd),
	.dataf(!\pipeline_dffe[16]~q ),
	.datag(gnd),
	.cin(\op_1~130 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~125_sumout ),
	.cout(\op_1~126 ),
	.shareout());
defparam \op_1~125 .extended_lut = "off";
defparam \op_1~125 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~125 .shared_arith = "off";

dffeas \pipeline_dffe[16] (
	.clk(clock),
	.d(\op_1~125_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\pipeline_dffe[16]~q ),
	.prn(vcc));
defparam \pipeline_dffe[16] .is_wysiwyg = "true";
defparam \pipeline_dffe[16] .power_up = "low";

arriav_lcell_comb \op_1~121 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_17),
	.datae(gnd),
	.dataf(!\pipeline_dffe[17]~q ),
	.datag(gnd),
	.cin(\op_1~126 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~121_sumout ),
	.cout(\op_1~122 ),
	.shareout());
defparam \op_1~121 .extended_lut = "off";
defparam \op_1~121 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~121 .shared_arith = "off";

dffeas \pipeline_dffe[17] (
	.clk(clock),
	.d(\op_1~121_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\pipeline_dffe[17]~q ),
	.prn(vcc));
defparam \pipeline_dffe[17] .is_wysiwyg = "true";
defparam \pipeline_dffe[17] .power_up = "low";

arriav_lcell_comb \op_1~117 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_18),
	.datae(gnd),
	.dataf(!\pipeline_dffe[18]~q ),
	.datag(gnd),
	.cin(\op_1~122 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~117_sumout ),
	.cout(\op_1~118 ),
	.shareout());
defparam \op_1~117 .extended_lut = "off";
defparam \op_1~117 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~117 .shared_arith = "off";

dffeas \pipeline_dffe[18] (
	.clk(clock),
	.d(\op_1~117_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\pipeline_dffe[18]~q ),
	.prn(vcc));
defparam \pipeline_dffe[18] .is_wysiwyg = "true";
defparam \pipeline_dffe[18] .power_up = "low";

arriav_lcell_comb \op_1~113 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_19),
	.datae(gnd),
	.dataf(!\pipeline_dffe[19]~q ),
	.datag(gnd),
	.cin(\op_1~118 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~113_sumout ),
	.cout(\op_1~114 ),
	.shareout());
defparam \op_1~113 .extended_lut = "off";
defparam \op_1~113 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~113 .shared_arith = "off";

dffeas \pipeline_dffe[19] (
	.clk(clock),
	.d(\op_1~113_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\pipeline_dffe[19]~q ),
	.prn(vcc));
defparam \pipeline_dffe[19] .is_wysiwyg = "true";
defparam \pipeline_dffe[19] .power_up = "low";

arriav_lcell_comb \op_1~109 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_20),
	.datae(gnd),
	.dataf(!\pipeline_dffe[20]~q ),
	.datag(gnd),
	.cin(\op_1~114 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~109_sumout ),
	.cout(\op_1~110 ),
	.shareout());
defparam \op_1~109 .extended_lut = "off";
defparam \op_1~109 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~109 .shared_arith = "off";

dffeas \pipeline_dffe[20] (
	.clk(clock),
	.d(\op_1~109_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\pipeline_dffe[20]~q ),
	.prn(vcc));
defparam \pipeline_dffe[20] .is_wysiwyg = "true";
defparam \pipeline_dffe[20] .power_up = "low";

arriav_lcell_comb \op_1~105 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_21),
	.datae(gnd),
	.dataf(!\pipeline_dffe[21]~q ),
	.datag(gnd),
	.cin(\op_1~110 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~105_sumout ),
	.cout(\op_1~106 ),
	.shareout());
defparam \op_1~105 .extended_lut = "off";
defparam \op_1~105 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~105 .shared_arith = "off";

dffeas \pipeline_dffe[21] (
	.clk(clock),
	.d(\op_1~105_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\pipeline_dffe[21]~q ),
	.prn(vcc));
defparam \pipeline_dffe[21] .is_wysiwyg = "true";
defparam \pipeline_dffe[21] .power_up = "low";

arriav_lcell_comb \op_1~101 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_22),
	.datae(gnd),
	.dataf(!\pipeline_dffe[22]~q ),
	.datag(gnd),
	.cin(\op_1~106 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~101_sumout ),
	.cout(\op_1~102 ),
	.shareout());
defparam \op_1~101 .extended_lut = "off";
defparam \op_1~101 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~101 .shared_arith = "off";

dffeas \pipeline_dffe[22] (
	.clk(clock),
	.d(\op_1~101_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\pipeline_dffe[22]~q ),
	.prn(vcc));
defparam \pipeline_dffe[22] .is_wysiwyg = "true";
defparam \pipeline_dffe[22] .power_up = "low";

arriav_lcell_comb \op_1~97 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_23),
	.datae(gnd),
	.dataf(!\pipeline_dffe[23]~q ),
	.datag(gnd),
	.cin(\op_1~102 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~97_sumout ),
	.cout(\op_1~98 ),
	.shareout());
defparam \op_1~97 .extended_lut = "off";
defparam \op_1~97 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~97 .shared_arith = "off";

dffeas \pipeline_dffe[23] (
	.clk(clock),
	.d(\op_1~97_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\pipeline_dffe[23]~q ),
	.prn(vcc));
defparam \pipeline_dffe[23] .is_wysiwyg = "true";
defparam \pipeline_dffe[23] .power_up = "low";

arriav_lcell_comb \op_1~93 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_24),
	.datae(gnd),
	.dataf(!\pipeline_dffe[24]~q ),
	.datag(gnd),
	.cin(\op_1~98 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~93_sumout ),
	.cout(\op_1~94 ),
	.shareout());
defparam \op_1~93 .extended_lut = "off";
defparam \op_1~93 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~93 .shared_arith = "off";

dffeas \pipeline_dffe[24] (
	.clk(clock),
	.d(\op_1~93_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\pipeline_dffe[24]~q ),
	.prn(vcc));
defparam \pipeline_dffe[24] .is_wysiwyg = "true";
defparam \pipeline_dffe[24] .power_up = "low";

arriav_lcell_comb \op_1~89 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_25),
	.datae(gnd),
	.dataf(!\pipeline_dffe[25]~q ),
	.datag(gnd),
	.cin(\op_1~94 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~89_sumout ),
	.cout(\op_1~90 ),
	.shareout());
defparam \op_1~89 .extended_lut = "off";
defparam \op_1~89 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~89 .shared_arith = "off";

dffeas \pipeline_dffe[25] (
	.clk(clock),
	.d(\op_1~89_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\pipeline_dffe[25]~q ),
	.prn(vcc));
defparam \pipeline_dffe[25] .is_wysiwyg = "true";
defparam \pipeline_dffe[25] .power_up = "low";

arriav_lcell_comb \op_1~85 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_26),
	.datae(gnd),
	.dataf(!\pipeline_dffe[26]~q ),
	.datag(gnd),
	.cin(\op_1~90 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~85_sumout ),
	.cout(\op_1~86 ),
	.shareout());
defparam \op_1~85 .extended_lut = "off";
defparam \op_1~85 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~85 .shared_arith = "off";

dffeas \pipeline_dffe[26] (
	.clk(clock),
	.d(\op_1~85_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\pipeline_dffe[26]~q ),
	.prn(vcc));
defparam \pipeline_dffe[26] .is_wysiwyg = "true";
defparam \pipeline_dffe[26] .power_up = "low";

arriav_lcell_comb \op_1~81 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_27),
	.datae(gnd),
	.dataf(!pipeline_dffe_27),
	.datag(gnd),
	.cin(\op_1~86 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~81_sumout ),
	.cout(\op_1~82 ),
	.shareout());
defparam \op_1~81 .extended_lut = "off";
defparam \op_1~81 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~81 .shared_arith = "off";

arriav_lcell_comb \op_1~77 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_28),
	.datae(gnd),
	.dataf(!pipeline_dffe_28),
	.datag(gnd),
	.cin(\op_1~82 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~77_sumout ),
	.cout(\op_1~78 ),
	.shareout());
defparam \op_1~77 .extended_lut = "off";
defparam \op_1~77 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~77 .shared_arith = "off";

arriav_lcell_comb \op_1~73 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_29),
	.datae(gnd),
	.dataf(!pipeline_dffe_29),
	.datag(gnd),
	.cin(\op_1~78 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~73_sumout ),
	.cout(\op_1~74 ),
	.shareout());
defparam \op_1~73 .extended_lut = "off";
defparam \op_1~73 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~73 .shared_arith = "off";

arriav_lcell_comb \op_1~69 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_30),
	.datae(gnd),
	.dataf(!pipeline_dffe_30),
	.datag(gnd),
	.cin(\op_1~74 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~69_sumout ),
	.cout(\op_1~70 ),
	.shareout());
defparam \op_1~69 .extended_lut = "off";
defparam \op_1~69 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~69 .shared_arith = "off";

arriav_lcell_comb \op_1~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_31),
	.datae(gnd),
	.dataf(!pipeline_dffe_31),
	.datag(gnd),
	.cin(\op_1~70 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~57_sumout ),
	.cout(\op_1~58 ),
	.shareout());
defparam \op_1~57 .extended_lut = "off";
defparam \op_1~57 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~57 .shared_arith = "off";

arriav_lcell_comb \op_1~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_32),
	.datae(gnd),
	.dataf(!pipeline_dffe_32),
	.datag(gnd),
	.cin(\op_1~58 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~1_sumout ),
	.cout(\op_1~2 ),
	.shareout());
defparam \op_1~1 .extended_lut = "off";
defparam \op_1~1 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~1 .shared_arith = "off";

arriav_lcell_comb \op_1~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_33),
	.datae(gnd),
	.dataf(!pipeline_dffe_33),
	.datag(gnd),
	.cin(\op_1~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~5_sumout ),
	.cout(\op_1~6 ),
	.shareout());
defparam \op_1~5 .extended_lut = "off";
defparam \op_1~5 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~5 .shared_arith = "off";

arriav_lcell_comb \op_1~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_34),
	.datae(gnd),
	.dataf(!pipeline_dffe_34),
	.datag(gnd),
	.cin(\op_1~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~9_sumout ),
	.cout(\op_1~10 ),
	.shareout());
defparam \op_1~9 .extended_lut = "off";
defparam \op_1~9 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~9 .shared_arith = "off";

arriav_lcell_comb \op_1~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_35),
	.datae(gnd),
	.dataf(!pipeline_dffe_35),
	.datag(gnd),
	.cin(\op_1~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~13_sumout ),
	.cout(\op_1~14 ),
	.shareout());
defparam \op_1~13 .extended_lut = "off";
defparam \op_1~13 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~13 .shared_arith = "off";

arriav_lcell_comb \op_1~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_36),
	.datae(gnd),
	.dataf(!pipeline_dffe_36),
	.datag(gnd),
	.cin(\op_1~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~17_sumout ),
	.cout(\op_1~18 ),
	.shareout());
defparam \op_1~17 .extended_lut = "off";
defparam \op_1~17 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~17 .shared_arith = "off";

arriav_lcell_comb \op_1~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_37),
	.datae(gnd),
	.dataf(!pipeline_dffe_37),
	.datag(gnd),
	.cin(\op_1~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~21_sumout ),
	.cout(\op_1~22 ),
	.shareout());
defparam \op_1~21 .extended_lut = "off";
defparam \op_1~21 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~21 .shared_arith = "off";

arriav_lcell_comb \op_1~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_38),
	.datae(gnd),
	.dataf(!pipeline_dffe_38),
	.datag(gnd),
	.cin(\op_1~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~25_sumout ),
	.cout(\op_1~26 ),
	.shareout());
defparam \op_1~25 .extended_lut = "off";
defparam \op_1~25 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~25 .shared_arith = "off";

arriav_lcell_comb \op_1~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_39),
	.datae(gnd),
	.dataf(!pipeline_dffe_39),
	.datag(gnd),
	.cin(\op_1~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~29_sumout ),
	.cout(\op_1~30 ),
	.shareout());
defparam \op_1~29 .extended_lut = "off";
defparam \op_1~29 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~29 .shared_arith = "off";

arriav_lcell_comb \op_1~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_40),
	.datae(gnd),
	.dataf(!pipeline_dffe_40),
	.datag(gnd),
	.cin(\op_1~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~33_sumout ),
	.cout(\op_1~34 ),
	.shareout());
defparam \op_1~33 .extended_lut = "off";
defparam \op_1~33 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~33 .shared_arith = "off";

arriav_lcell_comb \op_1~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_41),
	.datae(gnd),
	.dataf(!pipeline_dffe_41),
	.datag(gnd),
	.cin(\op_1~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~37_sumout ),
	.cout(\op_1~38 ),
	.shareout());
defparam \op_1~37 .extended_lut = "off";
defparam \op_1~37 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~37 .shared_arith = "off";

arriav_lcell_comb \op_1~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_42),
	.datae(gnd),
	.dataf(!pipeline_dffe_42),
	.datag(gnd),
	.cin(\op_1~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~41_sumout ),
	.cout(\op_1~42 ),
	.shareout());
defparam \op_1~41 .extended_lut = "off";
defparam \op_1~41 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~41 .shared_arith = "off";

arriav_lcell_comb \op_1~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_43),
	.datae(gnd),
	.dataf(!pipeline_dffe_43),
	.datag(gnd),
	.cin(\op_1~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~45_sumout ),
	.cout(\op_1~46 ),
	.shareout());
defparam \op_1~45 .extended_lut = "off";
defparam \op_1~45 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~45 .shared_arith = "off";

arriav_lcell_comb \op_1~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_44),
	.datae(gnd),
	.dataf(!pipeline_dffe_44),
	.datag(gnd),
	.cin(\op_1~46 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~49_sumout ),
	.cout(\op_1~50 ),
	.shareout());
defparam \op_1~49 .extended_lut = "off";
defparam \op_1~49 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~49 .shared_arith = "off";

arriav_lcell_comb \op_1~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_45),
	.datae(gnd),
	.dataf(!pipeline_dffe_45),
	.datag(gnd),
	.cin(\op_1~50 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~61_sumout ),
	.cout(\op_1~62 ),
	.shareout());
defparam \op_1~61 .extended_lut = "off";
defparam \op_1~61 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~61 .shared_arith = "off";

arriav_lcell_comb \op_1~65 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_46),
	.datae(gnd),
	.dataf(!pipeline_dffe_46),
	.datag(gnd),
	.cin(\op_1~62 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~65_sumout ),
	.cout(\op_1~66 ),
	.shareout());
defparam \op_1~65 .extended_lut = "off";
defparam \op_1~65 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~65 .shared_arith = "off";

arriav_lcell_comb \op_1~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_47),
	.datae(gnd),
	.dataf(!pipeline_dffe_47),
	.datag(gnd),
	.cin(\op_1~66 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~53_sumout ),
	.cout(),
	.shareout());
defparam \op_1~53 .extended_lut = "off";
defparam \op_1~53 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~53 .shared_arith = "off";

endmodule

module DDS_48_v1_asj_dxx (
	dxxpdo_5,
	dxxpdo_6,
	dxxpdo_7,
	dxxpdo_8,
	dxxpdo_9,
	dxxpdo_10,
	dxxpdo_11,
	dxxpdo_12,
	dxxpdo_13,
	dxxpdo_14,
	dxxpdo_15,
	dxxpdo_16,
	dxxpdo_17,
	dxxpdo_20,
	dxxpdo_18,
	dxxpdo_19,
	dxxrv_5,
	dxxrv_6,
	dxxrv_7,
	dxxrv_8,
	dxxrv_9,
	dxxrv_4,
	dxxrv_3,
	dxxrv_2,
	dxxrv_1,
	dxxrv_0,
	data_out_12,
	pipeline_dffe_32,
	pipeline_dffe_33,
	pipeline_dffe_34,
	pipeline_dffe_35,
	pipeline_dffe_36,
	pipeline_dffe_37,
	pipeline_dffe_38,
	pipeline_dffe_39,
	pipeline_dffe_40,
	pipeline_dffe_41,
	pipeline_dffe_42,
	pipeline_dffe_43,
	pipeline_dffe_44,
	pipeline_dffe_47,
	pipeline_dffe_31,
	pipeline_dffe_45,
	pipeline_dffe_46,
	pipeline_dffe_30,
	pipeline_dffe_29,
	pipeline_dffe_28,
	pipeline_dffe_27,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	dxxpdo_5;
output 	dxxpdo_6;
output 	dxxpdo_7;
output 	dxxpdo_8;
output 	dxxpdo_9;
output 	dxxpdo_10;
output 	dxxpdo_11;
output 	dxxpdo_12;
output 	dxxpdo_13;
output 	dxxpdo_14;
output 	dxxpdo_15;
output 	dxxpdo_16;
output 	dxxpdo_17;
output 	dxxpdo_20;
output 	dxxpdo_18;
output 	dxxpdo_19;
input 	dxxrv_5;
input 	dxxrv_6;
input 	dxxrv_7;
input 	dxxrv_8;
input 	dxxrv_9;
input 	dxxrv_4;
input 	dxxrv_3;
input 	dxxrv_2;
input 	dxxrv_1;
input 	dxxrv_0;
input 	data_out_12;
input 	pipeline_dffe_32;
input 	pipeline_dffe_33;
input 	pipeline_dffe_34;
input 	pipeline_dffe_35;
input 	pipeline_dffe_36;
input 	pipeline_dffe_37;
input 	pipeline_dffe_38;
input 	pipeline_dffe_39;
input 	pipeline_dffe_40;
input 	pipeline_dffe_41;
input 	pipeline_dffe_42;
input 	pipeline_dffe_43;
input 	pipeline_dffe_44;
input 	pipeline_dffe_47;
input 	pipeline_dffe_31;
input 	pipeline_dffe_45;
input 	pipeline_dffe_46;
input 	pipeline_dffe_30;
input 	pipeline_dffe_29;
input 	pipeline_dffe_28;
input 	pipeline_dffe_27;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Add0~82_cout ;
wire \Add0~78_cout ;
wire \Add0~74_cout ;
wire \Add0~70_cout ;
wire \Add0~58_cout ;
wire \Add0~1_sumout ;
wire \phi_dither_out_w[5]~q ;
wire \Add0~2 ;
wire \Add0~5_sumout ;
wire \phi_dither_out_w[6]~q ;
wire \Add0~6 ;
wire \Add0~9_sumout ;
wire \phi_dither_out_w[7]~q ;
wire \Add0~10 ;
wire \Add0~13_sumout ;
wire \phi_dither_out_w[8]~q ;
wire \Add0~14 ;
wire \Add0~17_sumout ;
wire \phi_dither_out_w[9]~q ;
wire \Add0~18 ;
wire \Add0~21_sumout ;
wire \phi_dither_out_w[10]~q ;
wire \Add0~22 ;
wire \Add0~25_sumout ;
wire \phi_dither_out_w[11]~q ;
wire \Add0~26 ;
wire \Add0~29_sumout ;
wire \phi_dither_out_w[12]~q ;
wire \Add0~30 ;
wire \Add0~33_sumout ;
wire \phi_dither_out_w[13]~q ;
wire \Add0~34 ;
wire \Add0~37_sumout ;
wire \phi_dither_out_w[14]~q ;
wire \Add0~38 ;
wire \Add0~41_sumout ;
wire \phi_dither_out_w[15]~q ;
wire \Add0~42 ;
wire \Add0~45_sumout ;
wire \phi_dither_out_w[16]~q ;
wire \Add0~46 ;
wire \Add0~49_sumout ;
wire \phi_dither_out_w[17]~q ;
wire \Add0~50 ;
wire \Add0~62 ;
wire \Add0~66 ;
wire \Add0~53_sumout ;
wire \phi_dither_out_w[20]~q ;
wire \Add0~61_sumout ;
wire \phi_dither_out_w[18]~q ;
wire \Add0~65_sumout ;
wire \phi_dither_out_w[19]~q ;


dffeas \dxxpdo[5] (
	.clk(clk),
	.d(\phi_dither_out_w[5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(dxxpdo_5),
	.prn(vcc));
defparam \dxxpdo[5] .is_wysiwyg = "true";
defparam \dxxpdo[5] .power_up = "low";

dffeas \dxxpdo[6] (
	.clk(clk),
	.d(\phi_dither_out_w[6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(dxxpdo_6),
	.prn(vcc));
defparam \dxxpdo[6] .is_wysiwyg = "true";
defparam \dxxpdo[6] .power_up = "low";

dffeas \dxxpdo[7] (
	.clk(clk),
	.d(\phi_dither_out_w[7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(dxxpdo_7),
	.prn(vcc));
defparam \dxxpdo[7] .is_wysiwyg = "true";
defparam \dxxpdo[7] .power_up = "low";

dffeas \dxxpdo[8] (
	.clk(clk),
	.d(\phi_dither_out_w[8]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(dxxpdo_8),
	.prn(vcc));
defparam \dxxpdo[8] .is_wysiwyg = "true";
defparam \dxxpdo[8] .power_up = "low";

dffeas \dxxpdo[9] (
	.clk(clk),
	.d(\phi_dither_out_w[9]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(dxxpdo_9),
	.prn(vcc));
defparam \dxxpdo[9] .is_wysiwyg = "true";
defparam \dxxpdo[9] .power_up = "low";

dffeas \dxxpdo[10] (
	.clk(clk),
	.d(\phi_dither_out_w[10]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(dxxpdo_10),
	.prn(vcc));
defparam \dxxpdo[10] .is_wysiwyg = "true";
defparam \dxxpdo[10] .power_up = "low";

dffeas \dxxpdo[11] (
	.clk(clk),
	.d(\phi_dither_out_w[11]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(dxxpdo_11),
	.prn(vcc));
defparam \dxxpdo[11] .is_wysiwyg = "true";
defparam \dxxpdo[11] .power_up = "low";

dffeas \dxxpdo[12] (
	.clk(clk),
	.d(\phi_dither_out_w[12]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(dxxpdo_12),
	.prn(vcc));
defparam \dxxpdo[12] .is_wysiwyg = "true";
defparam \dxxpdo[12] .power_up = "low";

dffeas \dxxpdo[13] (
	.clk(clk),
	.d(\phi_dither_out_w[13]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(dxxpdo_13),
	.prn(vcc));
defparam \dxxpdo[13] .is_wysiwyg = "true";
defparam \dxxpdo[13] .power_up = "low";

dffeas \dxxpdo[14] (
	.clk(clk),
	.d(\phi_dither_out_w[14]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(dxxpdo_14),
	.prn(vcc));
defparam \dxxpdo[14] .is_wysiwyg = "true";
defparam \dxxpdo[14] .power_up = "low";

dffeas \dxxpdo[15] (
	.clk(clk),
	.d(\phi_dither_out_w[15]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(dxxpdo_15),
	.prn(vcc));
defparam \dxxpdo[15] .is_wysiwyg = "true";
defparam \dxxpdo[15] .power_up = "low";

dffeas \dxxpdo[16] (
	.clk(clk),
	.d(\phi_dither_out_w[16]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(dxxpdo_16),
	.prn(vcc));
defparam \dxxpdo[16] .is_wysiwyg = "true";
defparam \dxxpdo[16] .power_up = "low";

dffeas \dxxpdo[17] (
	.clk(clk),
	.d(\phi_dither_out_w[17]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(dxxpdo_17),
	.prn(vcc));
defparam \dxxpdo[17] .is_wysiwyg = "true";
defparam \dxxpdo[17] .power_up = "low";

dffeas \dxxpdo[20] (
	.clk(clk),
	.d(\phi_dither_out_w[20]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(dxxpdo_20),
	.prn(vcc));
defparam \dxxpdo[20] .is_wysiwyg = "true";
defparam \dxxpdo[20] .power_up = "low";

dffeas \dxxpdo[18] (
	.clk(clk),
	.d(\phi_dither_out_w[18]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(dxxpdo_18),
	.prn(vcc));
defparam \dxxpdo[18] .is_wysiwyg = "true";
defparam \dxxpdo[18] .power_up = "low";

dffeas \dxxpdo[19] (
	.clk(clk),
	.d(\phi_dither_out_w[19]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(dxxpdo_19),
	.prn(vcc));
defparam \dxxpdo[19] .is_wysiwyg = "true";
defparam \dxxpdo[19] .power_up = "low";

arriav_lcell_comb \Add0~82 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxrv_0),
	.datae(gnd),
	.dataf(!pipeline_dffe_27),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\Add0~82_cout ),
	.shareout());
defparam \Add0~82 .extended_lut = "off";
defparam \Add0~82 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~82 .shared_arith = "off";

arriav_lcell_comb \Add0~78 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxrv_1),
	.datae(gnd),
	.dataf(!pipeline_dffe_28),
	.datag(gnd),
	.cin(\Add0~82_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\Add0~78_cout ),
	.shareout());
defparam \Add0~78 .extended_lut = "off";
defparam \Add0~78 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~78 .shared_arith = "off";

arriav_lcell_comb \Add0~74 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxrv_2),
	.datae(gnd),
	.dataf(!pipeline_dffe_29),
	.datag(gnd),
	.cin(\Add0~78_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\Add0~74_cout ),
	.shareout());
defparam \Add0~74 .extended_lut = "off";
defparam \Add0~74 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~74 .shared_arith = "off";

arriav_lcell_comb \Add0~70 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxrv_3),
	.datae(gnd),
	.dataf(!pipeline_dffe_30),
	.datag(gnd),
	.cin(\Add0~74_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\Add0~70_cout ),
	.shareout());
defparam \Add0~70 .extended_lut = "off";
defparam \Add0~70 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~70 .shared_arith = "off";

arriav_lcell_comb \Add0~58 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxrv_4),
	.datae(gnd),
	.dataf(!pipeline_dffe_31),
	.datag(gnd),
	.cin(\Add0~70_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\Add0~58_cout ),
	.shareout());
defparam \Add0~58 .extended_lut = "off";
defparam \Add0~58 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~58 .shared_arith = "off";

arriav_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxrv_5),
	.datae(gnd),
	.dataf(!pipeline_dffe_32),
	.datag(gnd),
	.cin(\Add0~58_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(\Add0~2 ),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~1 .shared_arith = "off";

dffeas \phi_dither_out_w[5] (
	.clk(clk),
	.d(\Add0~1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_dither_out_w[5]~q ),
	.prn(vcc));
defparam \phi_dither_out_w[5] .is_wysiwyg = "true";
defparam \phi_dither_out_w[5] .power_up = "low";

arriav_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxrv_6),
	.datae(gnd),
	.dataf(!pipeline_dffe_33),
	.datag(gnd),
	.cin(\Add0~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~5 .shared_arith = "off";

dffeas \phi_dither_out_w[6] (
	.clk(clk),
	.d(\Add0~5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_dither_out_w[6]~q ),
	.prn(vcc));
defparam \phi_dither_out_w[6] .is_wysiwyg = "true";
defparam \phi_dither_out_w[6] .power_up = "low";

arriav_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxrv_7),
	.datae(gnd),
	.dataf(!pipeline_dffe_34),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~9 .shared_arith = "off";

dffeas \phi_dither_out_w[7] (
	.clk(clk),
	.d(\Add0~9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_dither_out_w[7]~q ),
	.prn(vcc));
defparam \phi_dither_out_w[7] .is_wysiwyg = "true";
defparam \phi_dither_out_w[7] .power_up = "low";

arriav_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxrv_8),
	.datae(gnd),
	.dataf(!pipeline_dffe_35),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~13 .shared_arith = "off";

dffeas \phi_dither_out_w[8] (
	.clk(clk),
	.d(\Add0~13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_dither_out_w[8]~q ),
	.prn(vcc));
defparam \phi_dither_out_w[8] .is_wysiwyg = "true";
defparam \phi_dither_out_w[8] .power_up = "low";

arriav_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxrv_9),
	.datae(gnd),
	.dataf(!pipeline_dffe_36),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout());
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~17 .shared_arith = "off";

dffeas \phi_dither_out_w[9] (
	.clk(clk),
	.d(\Add0~17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_dither_out_w[9]~q ),
	.prn(vcc));
defparam \phi_dither_out_w[9] .is_wysiwyg = "true";
defparam \phi_dither_out_w[9] .power_up = "low";

arriav_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxrv_9),
	.datae(gnd),
	.dataf(!pipeline_dffe_37),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout());
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~21 .shared_arith = "off";

dffeas \phi_dither_out_w[10] (
	.clk(clk),
	.d(\Add0~21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_dither_out_w[10]~q ),
	.prn(vcc));
defparam \phi_dither_out_w[10] .is_wysiwyg = "true";
defparam \phi_dither_out_w[10] .power_up = "low";

arriav_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxrv_9),
	.datae(gnd),
	.dataf(!pipeline_dffe_38),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout());
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~25 .shared_arith = "off";

dffeas \phi_dither_out_w[11] (
	.clk(clk),
	.d(\Add0~25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_dither_out_w[11]~q ),
	.prn(vcc));
defparam \phi_dither_out_w[11] .is_wysiwyg = "true";
defparam \phi_dither_out_w[11] .power_up = "low";

arriav_lcell_comb \Add0~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxrv_9),
	.datae(gnd),
	.dataf(!pipeline_dffe_39),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout());
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~29 .shared_arith = "off";

dffeas \phi_dither_out_w[12] (
	.clk(clk),
	.d(\Add0~29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_dither_out_w[12]~q ),
	.prn(vcc));
defparam \phi_dither_out_w[12] .is_wysiwyg = "true";
defparam \phi_dither_out_w[12] .power_up = "low";

arriav_lcell_comb \Add0~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxrv_9),
	.datae(gnd),
	.dataf(!pipeline_dffe_40),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~33_sumout ),
	.cout(\Add0~34 ),
	.shareout());
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~33 .shared_arith = "off";

dffeas \phi_dither_out_w[13] (
	.clk(clk),
	.d(\Add0~33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_dither_out_w[13]~q ),
	.prn(vcc));
defparam \phi_dither_out_w[13] .is_wysiwyg = "true";
defparam \phi_dither_out_w[13] .power_up = "low";

arriav_lcell_comb \Add0~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxrv_9),
	.datae(gnd),
	.dataf(!pipeline_dffe_41),
	.datag(gnd),
	.cin(\Add0~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~37_sumout ),
	.cout(\Add0~38 ),
	.shareout());
defparam \Add0~37 .extended_lut = "off";
defparam \Add0~37 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~37 .shared_arith = "off";

dffeas \phi_dither_out_w[14] (
	.clk(clk),
	.d(\Add0~37_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_dither_out_w[14]~q ),
	.prn(vcc));
defparam \phi_dither_out_w[14] .is_wysiwyg = "true";
defparam \phi_dither_out_w[14] .power_up = "low";

arriav_lcell_comb \Add0~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxrv_9),
	.datae(gnd),
	.dataf(!pipeline_dffe_42),
	.datag(gnd),
	.cin(\Add0~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~41_sumout ),
	.cout(\Add0~42 ),
	.shareout());
defparam \Add0~41 .extended_lut = "off";
defparam \Add0~41 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~41 .shared_arith = "off";

dffeas \phi_dither_out_w[15] (
	.clk(clk),
	.d(\Add0~41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_dither_out_w[15]~q ),
	.prn(vcc));
defparam \phi_dither_out_w[15] .is_wysiwyg = "true";
defparam \phi_dither_out_w[15] .power_up = "low";

arriav_lcell_comb \Add0~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxrv_9),
	.datae(gnd),
	.dataf(!pipeline_dffe_43),
	.datag(gnd),
	.cin(\Add0~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~45_sumout ),
	.cout(\Add0~46 ),
	.shareout());
defparam \Add0~45 .extended_lut = "off";
defparam \Add0~45 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~45 .shared_arith = "off";

dffeas \phi_dither_out_w[16] (
	.clk(clk),
	.d(\Add0~45_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_dither_out_w[16]~q ),
	.prn(vcc));
defparam \phi_dither_out_w[16] .is_wysiwyg = "true";
defparam \phi_dither_out_w[16] .power_up = "low";

arriav_lcell_comb \Add0~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxrv_9),
	.datae(gnd),
	.dataf(!pipeline_dffe_44),
	.datag(gnd),
	.cin(\Add0~46 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~49_sumout ),
	.cout(\Add0~50 ),
	.shareout());
defparam \Add0~49 .extended_lut = "off";
defparam \Add0~49 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~49 .shared_arith = "off";

dffeas \phi_dither_out_w[17] (
	.clk(clk),
	.d(\Add0~49_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_dither_out_w[17]~q ),
	.prn(vcc));
defparam \phi_dither_out_w[17] .is_wysiwyg = "true";
defparam \phi_dither_out_w[17] .power_up = "low";

arriav_lcell_comb \Add0~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxrv_9),
	.datae(gnd),
	.dataf(!pipeline_dffe_45),
	.datag(gnd),
	.cin(\Add0~50 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~61_sumout ),
	.cout(\Add0~62 ),
	.shareout());
defparam \Add0~61 .extended_lut = "off";
defparam \Add0~61 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~61 .shared_arith = "off";

arriav_lcell_comb \Add0~65 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxrv_9),
	.datae(gnd),
	.dataf(!pipeline_dffe_46),
	.datag(gnd),
	.cin(\Add0~62 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~65_sumout ),
	.cout(\Add0~66 ),
	.shareout());
defparam \Add0~65 .extended_lut = "off";
defparam \Add0~65 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~65 .shared_arith = "off";

arriav_lcell_comb \Add0~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxrv_9),
	.datae(gnd),
	.dataf(!pipeline_dffe_47),
	.datag(gnd),
	.cin(\Add0~66 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~53_sumout ),
	.cout(),
	.shareout());
defparam \Add0~53 .extended_lut = "off";
defparam \Add0~53 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~53 .shared_arith = "off";

dffeas \phi_dither_out_w[20] (
	.clk(clk),
	.d(\Add0~53_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_dither_out_w[20]~q ),
	.prn(vcc));
defparam \phi_dither_out_w[20] .is_wysiwyg = "true";
defparam \phi_dither_out_w[20] .power_up = "low";

dffeas \phi_dither_out_w[18] (
	.clk(clk),
	.d(\Add0~61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_dither_out_w[18]~q ),
	.prn(vcc));
defparam \phi_dither_out_w[18] .is_wysiwyg = "true";
defparam \phi_dither_out_w[18] .power_up = "low";

dffeas \phi_dither_out_w[19] (
	.clk(clk),
	.d(\Add0~65_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_dither_out_w[19]~q ),
	.prn(vcc));
defparam \phi_dither_out_w[19] .is_wysiwyg = "true";
defparam \phi_dither_out_w[19] .power_up = "low";

endmodule

module DDS_48_v1_asj_dxx_g (
	dxxrv_5,
	dxxrv_6,
	dxxrv_7,
	dxxrv_8,
	dxxrv_9,
	dxxrv_4,
	dxxrv_3,
	dxxrv_2,
	dxxrv_1,
	dxxrv_0,
	data_out_12,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	dxxrv_5;
output 	dxxrv_6;
output 	dxxrv_7;
output 	dxxrv_8;
output 	dxxrv_9;
output 	dxxrv_4;
output 	dxxrv_3;
output 	dxxrv_2;
output 	dxxrv_1;
output 	dxxrv_0;
input 	data_out_12;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \lsfr_reg~1_combout ;
wire \lsfr_reg[12]~q ;
wire \lsfr_reg[13]~q ;
wire \lsfr_reg[14]~q ;
wire \lsfr_reg~2_combout ;
wire \lsfr_reg[15]~q ;
wire \lsfr_reg~9_combout ;
wire \lsfr_reg[0]~q ;
wire \lsfr_reg[1]~q ;
wire \lsfr_reg~8_combout ;
wire \lsfr_reg[2]~q ;
wire \lsfr_reg~7_combout ;
wire \lsfr_reg[3]~q ;
wire \lsfr_reg~6_combout ;
wire \lsfr_reg[4]~q ;
wire \lsfr_reg[5]~q ;
wire \lsfr_reg~5_combout ;
wire \lsfr_reg[6]~q ;
wire \lsfr_reg~4_combout ;
wire \lsfr_reg[7]~q ;
wire \lsfr_reg[8]~q ;
wire \lsfr_reg~3_combout ;
wire \lsfr_reg[9]~q ;
wire \lsfr_reg[10]~q ;
wire \lsfr_reg~0_combout ;
wire \lsfr_reg[11]~q ;
wire \Add0~38 ;
wire \Add0~34 ;
wire \Add0~30 ;
wire \Add0~26 ;
wire \Add0~22 ;
wire \Add0~1_sumout ;
wire \Add0~2 ;
wire \Add0~5_sumout ;
wire \Add0~6 ;
wire \Add0~9_sumout ;
wire \Add0~10 ;
wire \Add0~13_sumout ;
wire \Add0~14 ;
wire \Add0~17_sumout ;
wire \Add0~21_sumout ;
wire \Add0~25_sumout ;
wire \Add0~29_sumout ;
wire \Add0~33_sumout ;
wire \Add0~37_sumout ;


dffeas \dxxrv[5] (
	.clk(clk),
	.d(\Add0~1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(dxxrv_5),
	.prn(vcc));
defparam \dxxrv[5] .is_wysiwyg = "true";
defparam \dxxrv[5] .power_up = "low";

dffeas \dxxrv[6] (
	.clk(clk),
	.d(\Add0~5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(dxxrv_6),
	.prn(vcc));
defparam \dxxrv[6] .is_wysiwyg = "true";
defparam \dxxrv[6] .power_up = "low";

dffeas \dxxrv[7] (
	.clk(clk),
	.d(\Add0~9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(dxxrv_7),
	.prn(vcc));
defparam \dxxrv[7] .is_wysiwyg = "true";
defparam \dxxrv[7] .power_up = "low";

dffeas \dxxrv[8] (
	.clk(clk),
	.d(\Add0~13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(dxxrv_8),
	.prn(vcc));
defparam \dxxrv[8] .is_wysiwyg = "true";
defparam \dxxrv[8] .power_up = "low";

dffeas \dxxrv[9] (
	.clk(clk),
	.d(\Add0~17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(dxxrv_9),
	.prn(vcc));
defparam \dxxrv[9] .is_wysiwyg = "true";
defparam \dxxrv[9] .power_up = "low";

dffeas \dxxrv[4] (
	.clk(clk),
	.d(\Add0~21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(dxxrv_4),
	.prn(vcc));
defparam \dxxrv[4] .is_wysiwyg = "true";
defparam \dxxrv[4] .power_up = "low";

dffeas \dxxrv[3] (
	.clk(clk),
	.d(\Add0~25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(dxxrv_3),
	.prn(vcc));
defparam \dxxrv[3] .is_wysiwyg = "true";
defparam \dxxrv[3] .power_up = "low";

dffeas \dxxrv[2] (
	.clk(clk),
	.d(\Add0~29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(dxxrv_2),
	.prn(vcc));
defparam \dxxrv[2] .is_wysiwyg = "true";
defparam \dxxrv[2] .power_up = "low";

dffeas \dxxrv[1] (
	.clk(clk),
	.d(\Add0~33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(dxxrv_1),
	.prn(vcc));
defparam \dxxrv[1] .is_wysiwyg = "true";
defparam \dxxrv[1] .power_up = "low";

dffeas \dxxrv[0] (
	.clk(clk),
	.d(\Add0~37_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(dxxrv_0),
	.prn(vcc));
defparam \dxxrv[0] .is_wysiwyg = "true";
defparam \dxxrv[0] .power_up = "low";

arriav_lcell_comb \lsfr_reg~1 (
	.dataa(!reset_n),
	.datab(!\lsfr_reg[11]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lsfr_reg~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lsfr_reg~1 .extended_lut = "off";
defparam \lsfr_reg~1 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \lsfr_reg~1 .shared_arith = "off";

dffeas \lsfr_reg[12] (
	.clk(clk),
	.d(\lsfr_reg~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(data_out_12),
	.q(\lsfr_reg[12]~q ),
	.prn(vcc));
defparam \lsfr_reg[12] .is_wysiwyg = "true";
defparam \lsfr_reg[12] .power_up = "low";

dffeas \lsfr_reg[13] (
	.clk(clk),
	.d(\lsfr_reg[12]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\lsfr_reg[13]~q ),
	.prn(vcc));
defparam \lsfr_reg[13] .is_wysiwyg = "true";
defparam \lsfr_reg[13] .power_up = "low";

dffeas \lsfr_reg[14] (
	.clk(clk),
	.d(\lsfr_reg[13]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\lsfr_reg[14]~q ),
	.prn(vcc));
defparam \lsfr_reg[14] .is_wysiwyg = "true";
defparam \lsfr_reg[14] .power_up = "low";

arriav_lcell_comb \lsfr_reg~2 (
	.dataa(!reset_n),
	.datab(!\lsfr_reg[14]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lsfr_reg~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lsfr_reg~2 .extended_lut = "off";
defparam \lsfr_reg~2 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \lsfr_reg~2 .shared_arith = "off";

dffeas \lsfr_reg[15] (
	.clk(clk),
	.d(\lsfr_reg~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(data_out_12),
	.q(\lsfr_reg[15]~q ),
	.prn(vcc));
defparam \lsfr_reg[15] .is_wysiwyg = "true";
defparam \lsfr_reg[15] .power_up = "low";

arriav_lcell_comb \lsfr_reg~9 (
	.dataa(!\lsfr_reg[15]~q ),
	.datab(!\lsfr_reg[12]~q ),
	.datac(!\lsfr_reg[14]~q ),
	.datad(!\lsfr_reg[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lsfr_reg~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lsfr_reg~9 .extended_lut = "off";
defparam \lsfr_reg~9 .lut_mask = 64'h6996699669966996;
defparam \lsfr_reg~9 .shared_arith = "off";

dffeas \lsfr_reg[0] (
	.clk(clk),
	.d(\lsfr_reg~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(data_out_12),
	.q(\lsfr_reg[0]~q ),
	.prn(vcc));
defparam \lsfr_reg[0] .is_wysiwyg = "true";
defparam \lsfr_reg[0] .power_up = "low";

dffeas \lsfr_reg[1] (
	.clk(clk),
	.d(\lsfr_reg[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\lsfr_reg[1]~q ),
	.prn(vcc));
defparam \lsfr_reg[1] .is_wysiwyg = "true";
defparam \lsfr_reg[1] .power_up = "low";

arriav_lcell_comb \lsfr_reg~8 (
	.dataa(!reset_n),
	.datab(!\lsfr_reg[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lsfr_reg~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lsfr_reg~8 .extended_lut = "off";
defparam \lsfr_reg~8 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \lsfr_reg~8 .shared_arith = "off";

dffeas \lsfr_reg[2] (
	.clk(clk),
	.d(\lsfr_reg~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(data_out_12),
	.q(\lsfr_reg[2]~q ),
	.prn(vcc));
defparam \lsfr_reg[2] .is_wysiwyg = "true";
defparam \lsfr_reg[2] .power_up = "low";

arriav_lcell_comb \lsfr_reg~7 (
	.dataa(!reset_n),
	.datab(!\lsfr_reg[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lsfr_reg~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lsfr_reg~7 .extended_lut = "off";
defparam \lsfr_reg~7 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \lsfr_reg~7 .shared_arith = "off";

dffeas \lsfr_reg[3] (
	.clk(clk),
	.d(\lsfr_reg~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(data_out_12),
	.q(\lsfr_reg[3]~q ),
	.prn(vcc));
defparam \lsfr_reg[3] .is_wysiwyg = "true";
defparam \lsfr_reg[3] .power_up = "low";

arriav_lcell_comb \lsfr_reg~6 (
	.dataa(!reset_n),
	.datab(!\lsfr_reg[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lsfr_reg~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lsfr_reg~6 .extended_lut = "off";
defparam \lsfr_reg~6 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \lsfr_reg~6 .shared_arith = "off";

dffeas \lsfr_reg[4] (
	.clk(clk),
	.d(\lsfr_reg~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(data_out_12),
	.q(\lsfr_reg[4]~q ),
	.prn(vcc));
defparam \lsfr_reg[4] .is_wysiwyg = "true";
defparam \lsfr_reg[4] .power_up = "low";

dffeas \lsfr_reg[5] (
	.clk(clk),
	.d(\lsfr_reg[4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\lsfr_reg[5]~q ),
	.prn(vcc));
defparam \lsfr_reg[5] .is_wysiwyg = "true";
defparam \lsfr_reg[5] .power_up = "low";

arriav_lcell_comb \lsfr_reg~5 (
	.dataa(!reset_n),
	.datab(!\lsfr_reg[5]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lsfr_reg~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lsfr_reg~5 .extended_lut = "off";
defparam \lsfr_reg~5 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \lsfr_reg~5 .shared_arith = "off";

dffeas \lsfr_reg[6] (
	.clk(clk),
	.d(\lsfr_reg~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(data_out_12),
	.q(\lsfr_reg[6]~q ),
	.prn(vcc));
defparam \lsfr_reg[6] .is_wysiwyg = "true";
defparam \lsfr_reg[6] .power_up = "low";

arriav_lcell_comb \lsfr_reg~4 (
	.dataa(!reset_n),
	.datab(!\lsfr_reg[6]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lsfr_reg~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lsfr_reg~4 .extended_lut = "off";
defparam \lsfr_reg~4 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \lsfr_reg~4 .shared_arith = "off";

dffeas \lsfr_reg[7] (
	.clk(clk),
	.d(\lsfr_reg~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(data_out_12),
	.q(\lsfr_reg[7]~q ),
	.prn(vcc));
defparam \lsfr_reg[7] .is_wysiwyg = "true";
defparam \lsfr_reg[7] .power_up = "low";

dffeas \lsfr_reg[8] (
	.clk(clk),
	.d(\lsfr_reg[7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\lsfr_reg[8]~q ),
	.prn(vcc));
defparam \lsfr_reg[8] .is_wysiwyg = "true";
defparam \lsfr_reg[8] .power_up = "low";

arriav_lcell_comb \lsfr_reg~3 (
	.dataa(!reset_n),
	.datab(!\lsfr_reg[8]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lsfr_reg~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lsfr_reg~3 .extended_lut = "off";
defparam \lsfr_reg~3 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \lsfr_reg~3 .shared_arith = "off";

dffeas \lsfr_reg[9] (
	.clk(clk),
	.d(\lsfr_reg~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(data_out_12),
	.q(\lsfr_reg[9]~q ),
	.prn(vcc));
defparam \lsfr_reg[9] .is_wysiwyg = "true";
defparam \lsfr_reg[9] .power_up = "low";

dffeas \lsfr_reg[10] (
	.clk(clk),
	.d(\lsfr_reg[9]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\lsfr_reg[10]~q ),
	.prn(vcc));
defparam \lsfr_reg[10] .is_wysiwyg = "true";
defparam \lsfr_reg[10] .power_up = "low";

arriav_lcell_comb \lsfr_reg~0 (
	.dataa(!reset_n),
	.datab(!\lsfr_reg[10]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lsfr_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lsfr_reg~0 .extended_lut = "off";
defparam \lsfr_reg~0 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \lsfr_reg~0 .shared_arith = "off";

dffeas \lsfr_reg[11] (
	.clk(clk),
	.d(\lsfr_reg~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(data_out_12),
	.q(\lsfr_reg[11]~q ),
	.prn(vcc));
defparam \lsfr_reg[11] .is_wysiwyg = "true";
defparam \lsfr_reg[11] .power_up = "low";

arriav_lcell_comb \Add0~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\lsfr_reg[15]~q ),
	.datae(gnd),
	.dataf(!\lsfr_reg[6]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~37_sumout ),
	.cout(\Add0~38 ),
	.shareout());
defparam \Add0~37 .extended_lut = "off";
defparam \Add0~37 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~37 .shared_arith = "off";

arriav_lcell_comb \Add0~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\lsfr_reg[7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~33_sumout ),
	.cout(\Add0~34 ),
	.shareout());
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h00000000000000FF;
defparam \Add0~33 .shared_arith = "off";

arriav_lcell_comb \Add0~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\lsfr_reg[8]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout());
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h00000000000000FF;
defparam \Add0~29 .shared_arith = "off";

arriav_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\lsfr_reg[9]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout());
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h00000000000000FF;
defparam \Add0~25 .shared_arith = "off";

arriav_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\lsfr_reg[10]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout());
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h00000000000000FF;
defparam \Add0~21 .shared_arith = "off";

arriav_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\lsfr_reg[11]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(\Add0~2 ),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h00000000000000FF;
defparam \Add0~1 .shared_arith = "off";

arriav_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\lsfr_reg[12]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h00000000000000FF;
defparam \Add0~5 .shared_arith = "off";

arriav_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\lsfr_reg[13]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h00000000000000FF;
defparam \Add0~9 .shared_arith = "off";

arriav_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\lsfr_reg[14]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h00000000000000FF;
defparam \Add0~13 .shared_arith = "off";

arriav_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\lsfr_reg[15]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(),
	.shareout());
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h00000000000000FF;
defparam \Add0~17 .shared_arith = "off";

endmodule

module DDS_48_v1_asj_gal (
	rom_add_0,
	rom_add_1,
	rom_add_2,
	rom_add_3,
	rom_add_4,
	rom_add_5,
	rom_add_6,
	rom_add_7,
	rom_add_8,
	rom_add_9,
	rom_add_10,
	rom_add_11,
	rom_add_12,
	rom_add_15,
	rom_add_13,
	rom_add_14,
	data_out_12,
	pipeline_dffe_0,
	pipeline_dffe_1,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	pipeline_dffe_10,
	pipeline_dffe_11,
	pipeline_dffe_12,
	pipeline_dffe_15,
	pipeline_dffe_13,
	pipeline_dffe_14,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	rom_add_0;
output 	rom_add_1;
output 	rom_add_2;
output 	rom_add_3;
output 	rom_add_4;
output 	rom_add_5;
output 	rom_add_6;
output 	rom_add_7;
output 	rom_add_8;
output 	rom_add_9;
output 	rom_add_10;
output 	rom_add_11;
output 	rom_add_12;
output 	rom_add_15;
output 	rom_add_13;
output 	rom_add_14;
input 	data_out_12;
input 	pipeline_dffe_0;
input 	pipeline_dffe_1;
input 	pipeline_dffe_2;
input 	pipeline_dffe_3;
input 	pipeline_dffe_4;
input 	pipeline_dffe_5;
input 	pipeline_dffe_6;
input 	pipeline_dffe_7;
input 	pipeline_dffe_8;
input 	pipeline_dffe_9;
input 	pipeline_dffe_10;
input 	pipeline_dffe_11;
input 	pipeline_dffe_12;
input 	pipeline_dffe_15;
input 	pipeline_dffe_13;
input 	pipeline_dffe_14;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \rom_add[0] (
	.clk(clk),
	.d(pipeline_dffe_0),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(rom_add_0),
	.prn(vcc));
defparam \rom_add[0] .is_wysiwyg = "true";
defparam \rom_add[0] .power_up = "low";

dffeas \rom_add[1] (
	.clk(clk),
	.d(pipeline_dffe_1),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(rom_add_1),
	.prn(vcc));
defparam \rom_add[1] .is_wysiwyg = "true";
defparam \rom_add[1] .power_up = "low";

dffeas \rom_add[2] (
	.clk(clk),
	.d(pipeline_dffe_2),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(rom_add_2),
	.prn(vcc));
defparam \rom_add[2] .is_wysiwyg = "true";
defparam \rom_add[2] .power_up = "low";

dffeas \rom_add[3] (
	.clk(clk),
	.d(pipeline_dffe_3),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(rom_add_3),
	.prn(vcc));
defparam \rom_add[3] .is_wysiwyg = "true";
defparam \rom_add[3] .power_up = "low";

dffeas \rom_add[4] (
	.clk(clk),
	.d(pipeline_dffe_4),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(rom_add_4),
	.prn(vcc));
defparam \rom_add[4] .is_wysiwyg = "true";
defparam \rom_add[4] .power_up = "low";

dffeas \rom_add[5] (
	.clk(clk),
	.d(pipeline_dffe_5),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(rom_add_5),
	.prn(vcc));
defparam \rom_add[5] .is_wysiwyg = "true";
defparam \rom_add[5] .power_up = "low";

dffeas \rom_add[6] (
	.clk(clk),
	.d(pipeline_dffe_6),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(rom_add_6),
	.prn(vcc));
defparam \rom_add[6] .is_wysiwyg = "true";
defparam \rom_add[6] .power_up = "low";

dffeas \rom_add[7] (
	.clk(clk),
	.d(pipeline_dffe_7),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(rom_add_7),
	.prn(vcc));
defparam \rom_add[7] .is_wysiwyg = "true";
defparam \rom_add[7] .power_up = "low";

dffeas \rom_add[8] (
	.clk(clk),
	.d(pipeline_dffe_8),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(rom_add_8),
	.prn(vcc));
defparam \rom_add[8] .is_wysiwyg = "true";
defparam \rom_add[8] .power_up = "low";

dffeas \rom_add[9] (
	.clk(clk),
	.d(pipeline_dffe_9),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(rom_add_9),
	.prn(vcc));
defparam \rom_add[9] .is_wysiwyg = "true";
defparam \rom_add[9] .power_up = "low";

dffeas \rom_add[10] (
	.clk(clk),
	.d(pipeline_dffe_10),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(rom_add_10),
	.prn(vcc));
defparam \rom_add[10] .is_wysiwyg = "true";
defparam \rom_add[10] .power_up = "low";

dffeas \rom_add[11] (
	.clk(clk),
	.d(pipeline_dffe_11),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(rom_add_11),
	.prn(vcc));
defparam \rom_add[11] .is_wysiwyg = "true";
defparam \rom_add[11] .power_up = "low";

dffeas \rom_add[12] (
	.clk(clk),
	.d(pipeline_dffe_12),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(rom_add_12),
	.prn(vcc));
defparam \rom_add[12] .is_wysiwyg = "true";
defparam \rom_add[12] .power_up = "low";

dffeas \rom_add[15] (
	.clk(clk),
	.d(pipeline_dffe_15),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(rom_add_15),
	.prn(vcc));
defparam \rom_add[15] .is_wysiwyg = "true";
defparam \rom_add[15] .power_up = "low";

dffeas \rom_add[13] (
	.clk(clk),
	.d(pipeline_dffe_13),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(rom_add_13),
	.prn(vcc));
defparam \rom_add[13] .is_wysiwyg = "true";
defparam \rom_add[13] .power_up = "low";

dffeas \rom_add[14] (
	.clk(clk),
	.d(pipeline_dffe_14),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(rom_add_14),
	.prn(vcc));
defparam \rom_add[14] .is_wysiwyg = "true";
defparam \rom_add[14] .power_up = "low";

endmodule

module DDS_48_v1_asj_nco_as_m_cen (
	ram_block1a64,
	ram_block1a80,
	ram_block1a96,
	ram_block1a112,
	ram_block1a32,
	ram_block1a48,
	ram_block1a0,
	ram_block1a16,
	ram_block1a65,
	ram_block1a81,
	ram_block1a97,
	ram_block1a113,
	ram_block1a33,
	ram_block1a49,
	ram_block1a1,
	ram_block1a17,
	ram_block1a66,
	ram_block1a82,
	ram_block1a98,
	ram_block1a114,
	ram_block1a34,
	ram_block1a50,
	ram_block1a2,
	ram_block1a18,
	ram_block1a67,
	ram_block1a83,
	ram_block1a99,
	ram_block1a115,
	ram_block1a35,
	ram_block1a51,
	ram_block1a3,
	ram_block1a19,
	ram_block1a68,
	ram_block1a84,
	ram_block1a100,
	ram_block1a116,
	ram_block1a36,
	ram_block1a52,
	ram_block1a4,
	ram_block1a20,
	ram_block1a69,
	ram_block1a85,
	ram_block1a101,
	ram_block1a117,
	ram_block1a37,
	ram_block1a53,
	ram_block1a5,
	ram_block1a21,
	ram_block1a70,
	ram_block1a86,
	ram_block1a102,
	ram_block1a118,
	ram_block1a38,
	ram_block1a54,
	ram_block1a6,
	ram_block1a22,
	ram_block1a71,
	ram_block1a87,
	ram_block1a103,
	ram_block1a119,
	ram_block1a39,
	ram_block1a55,
	ram_block1a7,
	ram_block1a23,
	ram_block1a72,
	ram_block1a88,
	ram_block1a104,
	ram_block1a120,
	ram_block1a40,
	ram_block1a56,
	ram_block1a8,
	ram_block1a24,
	ram_block1a73,
	ram_block1a89,
	ram_block1a105,
	ram_block1a121,
	ram_block1a41,
	ram_block1a57,
	ram_block1a9,
	ram_block1a25,
	ram_block1a74,
	ram_block1a90,
	ram_block1a106,
	ram_block1a122,
	ram_block1a42,
	ram_block1a58,
	ram_block1a10,
	ram_block1a26,
	ram_block1a75,
	ram_block1a91,
	ram_block1a107,
	ram_block1a123,
	ram_block1a43,
	ram_block1a59,
	ram_block1a11,
	ram_block1a27,
	ram_block1a76,
	ram_block1a92,
	ram_block1a108,
	ram_block1a124,
	ram_block1a44,
	ram_block1a60,
	ram_block1a12,
	ram_block1a28,
	ram_block1a77,
	ram_block1a93,
	ram_block1a109,
	ram_block1a125,
	ram_block1a45,
	ram_block1a61,
	ram_block1a13,
	ram_block1a29,
	ram_block1a78,
	ram_block1a94,
	ram_block1a110,
	ram_block1a126,
	ram_block1a46,
	ram_block1a62,
	ram_block1a14,
	ram_block1a30,
	ram_block1a79,
	ram_block1a95,
	ram_block1a111,
	ram_block1a127,
	ram_block1a47,
	ram_block1a63,
	ram_block1a15,
	ram_block1a31,
	rom_add_0,
	rom_add_1,
	rom_add_2,
	rom_add_3,
	rom_add_4,
	rom_add_5,
	rom_add_6,
	rom_add_7,
	rom_add_8,
	rom_add_9,
	rom_add_10,
	rom_add_11,
	rom_add_12,
	rom_add_15,
	rom_add_13,
	rom_add_14,
	out_address_reg_a_2,
	out_address_reg_a_0,
	out_address_reg_a_1,
	clk,
	clken)/* synthesis synthesis_greybox=1 */;
output 	ram_block1a64;
output 	ram_block1a80;
output 	ram_block1a96;
output 	ram_block1a112;
output 	ram_block1a32;
output 	ram_block1a48;
output 	ram_block1a0;
output 	ram_block1a16;
output 	ram_block1a65;
output 	ram_block1a81;
output 	ram_block1a97;
output 	ram_block1a113;
output 	ram_block1a33;
output 	ram_block1a49;
output 	ram_block1a1;
output 	ram_block1a17;
output 	ram_block1a66;
output 	ram_block1a82;
output 	ram_block1a98;
output 	ram_block1a114;
output 	ram_block1a34;
output 	ram_block1a50;
output 	ram_block1a2;
output 	ram_block1a18;
output 	ram_block1a67;
output 	ram_block1a83;
output 	ram_block1a99;
output 	ram_block1a115;
output 	ram_block1a35;
output 	ram_block1a51;
output 	ram_block1a3;
output 	ram_block1a19;
output 	ram_block1a68;
output 	ram_block1a84;
output 	ram_block1a100;
output 	ram_block1a116;
output 	ram_block1a36;
output 	ram_block1a52;
output 	ram_block1a4;
output 	ram_block1a20;
output 	ram_block1a69;
output 	ram_block1a85;
output 	ram_block1a101;
output 	ram_block1a117;
output 	ram_block1a37;
output 	ram_block1a53;
output 	ram_block1a5;
output 	ram_block1a21;
output 	ram_block1a70;
output 	ram_block1a86;
output 	ram_block1a102;
output 	ram_block1a118;
output 	ram_block1a38;
output 	ram_block1a54;
output 	ram_block1a6;
output 	ram_block1a22;
output 	ram_block1a71;
output 	ram_block1a87;
output 	ram_block1a103;
output 	ram_block1a119;
output 	ram_block1a39;
output 	ram_block1a55;
output 	ram_block1a7;
output 	ram_block1a23;
output 	ram_block1a72;
output 	ram_block1a88;
output 	ram_block1a104;
output 	ram_block1a120;
output 	ram_block1a40;
output 	ram_block1a56;
output 	ram_block1a8;
output 	ram_block1a24;
output 	ram_block1a73;
output 	ram_block1a89;
output 	ram_block1a105;
output 	ram_block1a121;
output 	ram_block1a41;
output 	ram_block1a57;
output 	ram_block1a9;
output 	ram_block1a25;
output 	ram_block1a74;
output 	ram_block1a90;
output 	ram_block1a106;
output 	ram_block1a122;
output 	ram_block1a42;
output 	ram_block1a58;
output 	ram_block1a10;
output 	ram_block1a26;
output 	ram_block1a75;
output 	ram_block1a91;
output 	ram_block1a107;
output 	ram_block1a123;
output 	ram_block1a43;
output 	ram_block1a59;
output 	ram_block1a11;
output 	ram_block1a27;
output 	ram_block1a76;
output 	ram_block1a92;
output 	ram_block1a108;
output 	ram_block1a124;
output 	ram_block1a44;
output 	ram_block1a60;
output 	ram_block1a12;
output 	ram_block1a28;
output 	ram_block1a77;
output 	ram_block1a93;
output 	ram_block1a109;
output 	ram_block1a125;
output 	ram_block1a45;
output 	ram_block1a61;
output 	ram_block1a13;
output 	ram_block1a29;
output 	ram_block1a78;
output 	ram_block1a94;
output 	ram_block1a110;
output 	ram_block1a126;
output 	ram_block1a46;
output 	ram_block1a62;
output 	ram_block1a14;
output 	ram_block1a30;
output 	ram_block1a79;
output 	ram_block1a95;
output 	ram_block1a111;
output 	ram_block1a127;
output 	ram_block1a47;
output 	ram_block1a63;
output 	ram_block1a15;
output 	ram_block1a31;
input 	rom_add_0;
input 	rom_add_1;
input 	rom_add_2;
input 	rom_add_3;
input 	rom_add_4;
input 	rom_add_5;
input 	rom_add_6;
input 	rom_add_7;
input 	rom_add_8;
input 	rom_add_9;
input 	rom_add_10;
input 	rom_add_11;
input 	rom_add_12;
input 	rom_add_15;
input 	rom_add_13;
input 	rom_add_14;
output 	out_address_reg_a_2;
output 	out_address_reg_a_0;
output 	out_address_reg_a_1;
input 	clk;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



DDS_48_v1_altsyncram_1 altsyncram_component0(
	.ram_block1a64(ram_block1a64),
	.ram_block1a80(ram_block1a80),
	.ram_block1a96(ram_block1a96),
	.ram_block1a112(ram_block1a112),
	.ram_block1a32(ram_block1a32),
	.ram_block1a48(ram_block1a48),
	.ram_block1a0(ram_block1a0),
	.ram_block1a16(ram_block1a16),
	.ram_block1a65(ram_block1a65),
	.ram_block1a81(ram_block1a81),
	.ram_block1a97(ram_block1a97),
	.ram_block1a113(ram_block1a113),
	.ram_block1a33(ram_block1a33),
	.ram_block1a49(ram_block1a49),
	.ram_block1a1(ram_block1a1),
	.ram_block1a17(ram_block1a17),
	.ram_block1a66(ram_block1a66),
	.ram_block1a82(ram_block1a82),
	.ram_block1a98(ram_block1a98),
	.ram_block1a114(ram_block1a114),
	.ram_block1a34(ram_block1a34),
	.ram_block1a50(ram_block1a50),
	.ram_block1a2(ram_block1a2),
	.ram_block1a18(ram_block1a18),
	.ram_block1a67(ram_block1a67),
	.ram_block1a83(ram_block1a83),
	.ram_block1a99(ram_block1a99),
	.ram_block1a115(ram_block1a115),
	.ram_block1a35(ram_block1a35),
	.ram_block1a51(ram_block1a51),
	.ram_block1a3(ram_block1a3),
	.ram_block1a19(ram_block1a19),
	.ram_block1a68(ram_block1a68),
	.ram_block1a84(ram_block1a84),
	.ram_block1a100(ram_block1a100),
	.ram_block1a116(ram_block1a116),
	.ram_block1a36(ram_block1a36),
	.ram_block1a52(ram_block1a52),
	.ram_block1a4(ram_block1a4),
	.ram_block1a20(ram_block1a20),
	.ram_block1a69(ram_block1a69),
	.ram_block1a85(ram_block1a85),
	.ram_block1a101(ram_block1a101),
	.ram_block1a117(ram_block1a117),
	.ram_block1a37(ram_block1a37),
	.ram_block1a53(ram_block1a53),
	.ram_block1a5(ram_block1a5),
	.ram_block1a21(ram_block1a21),
	.ram_block1a70(ram_block1a70),
	.ram_block1a86(ram_block1a86),
	.ram_block1a102(ram_block1a102),
	.ram_block1a118(ram_block1a118),
	.ram_block1a38(ram_block1a38),
	.ram_block1a54(ram_block1a54),
	.ram_block1a6(ram_block1a6),
	.ram_block1a22(ram_block1a22),
	.ram_block1a71(ram_block1a71),
	.ram_block1a87(ram_block1a87),
	.ram_block1a103(ram_block1a103),
	.ram_block1a119(ram_block1a119),
	.ram_block1a39(ram_block1a39),
	.ram_block1a55(ram_block1a55),
	.ram_block1a7(ram_block1a7),
	.ram_block1a23(ram_block1a23),
	.ram_block1a72(ram_block1a72),
	.ram_block1a88(ram_block1a88),
	.ram_block1a104(ram_block1a104),
	.ram_block1a120(ram_block1a120),
	.ram_block1a40(ram_block1a40),
	.ram_block1a56(ram_block1a56),
	.ram_block1a8(ram_block1a8),
	.ram_block1a24(ram_block1a24),
	.ram_block1a73(ram_block1a73),
	.ram_block1a89(ram_block1a89),
	.ram_block1a105(ram_block1a105),
	.ram_block1a121(ram_block1a121),
	.ram_block1a41(ram_block1a41),
	.ram_block1a57(ram_block1a57),
	.ram_block1a9(ram_block1a9),
	.ram_block1a25(ram_block1a25),
	.ram_block1a74(ram_block1a74),
	.ram_block1a90(ram_block1a90),
	.ram_block1a106(ram_block1a106),
	.ram_block1a122(ram_block1a122),
	.ram_block1a42(ram_block1a42),
	.ram_block1a58(ram_block1a58),
	.ram_block1a10(ram_block1a10),
	.ram_block1a26(ram_block1a26),
	.ram_block1a75(ram_block1a75),
	.ram_block1a91(ram_block1a91),
	.ram_block1a107(ram_block1a107),
	.ram_block1a123(ram_block1a123),
	.ram_block1a43(ram_block1a43),
	.ram_block1a59(ram_block1a59),
	.ram_block1a11(ram_block1a11),
	.ram_block1a27(ram_block1a27),
	.ram_block1a76(ram_block1a76),
	.ram_block1a92(ram_block1a92),
	.ram_block1a108(ram_block1a108),
	.ram_block1a124(ram_block1a124),
	.ram_block1a44(ram_block1a44),
	.ram_block1a60(ram_block1a60),
	.ram_block1a12(ram_block1a12),
	.ram_block1a28(ram_block1a28),
	.ram_block1a77(ram_block1a77),
	.ram_block1a93(ram_block1a93),
	.ram_block1a109(ram_block1a109),
	.ram_block1a125(ram_block1a125),
	.ram_block1a45(ram_block1a45),
	.ram_block1a61(ram_block1a61),
	.ram_block1a13(ram_block1a13),
	.ram_block1a29(ram_block1a29),
	.ram_block1a78(ram_block1a78),
	.ram_block1a94(ram_block1a94),
	.ram_block1a110(ram_block1a110),
	.ram_block1a126(ram_block1a126),
	.ram_block1a46(ram_block1a46),
	.ram_block1a62(ram_block1a62),
	.ram_block1a14(ram_block1a14),
	.ram_block1a30(ram_block1a30),
	.ram_block1a79(ram_block1a79),
	.ram_block1a95(ram_block1a95),
	.ram_block1a111(ram_block1a111),
	.ram_block1a127(ram_block1a127),
	.ram_block1a47(ram_block1a47),
	.ram_block1a63(ram_block1a63),
	.ram_block1a15(ram_block1a15),
	.ram_block1a31(ram_block1a31),
	.address_a({rom_add_15,rom_add_14,rom_add_13,rom_add_12,rom_add_11,rom_add_10,rom_add_9,rom_add_8,rom_add_7,rom_add_6,rom_add_5,rom_add_4,rom_add_3,rom_add_2,rom_add_1,rom_add_0}),
	.out_address_reg_a_2(out_address_reg_a_2),
	.out_address_reg_a_0(out_address_reg_a_0),
	.out_address_reg_a_1(out_address_reg_a_1),
	.clock0(clk),
	.clocken0(clken));

endmodule

module DDS_48_v1_altsyncram_1 (
	ram_block1a64,
	ram_block1a80,
	ram_block1a96,
	ram_block1a112,
	ram_block1a32,
	ram_block1a48,
	ram_block1a0,
	ram_block1a16,
	ram_block1a65,
	ram_block1a81,
	ram_block1a97,
	ram_block1a113,
	ram_block1a33,
	ram_block1a49,
	ram_block1a1,
	ram_block1a17,
	ram_block1a66,
	ram_block1a82,
	ram_block1a98,
	ram_block1a114,
	ram_block1a34,
	ram_block1a50,
	ram_block1a2,
	ram_block1a18,
	ram_block1a67,
	ram_block1a83,
	ram_block1a99,
	ram_block1a115,
	ram_block1a35,
	ram_block1a51,
	ram_block1a3,
	ram_block1a19,
	ram_block1a68,
	ram_block1a84,
	ram_block1a100,
	ram_block1a116,
	ram_block1a36,
	ram_block1a52,
	ram_block1a4,
	ram_block1a20,
	ram_block1a69,
	ram_block1a85,
	ram_block1a101,
	ram_block1a117,
	ram_block1a37,
	ram_block1a53,
	ram_block1a5,
	ram_block1a21,
	ram_block1a70,
	ram_block1a86,
	ram_block1a102,
	ram_block1a118,
	ram_block1a38,
	ram_block1a54,
	ram_block1a6,
	ram_block1a22,
	ram_block1a71,
	ram_block1a87,
	ram_block1a103,
	ram_block1a119,
	ram_block1a39,
	ram_block1a55,
	ram_block1a7,
	ram_block1a23,
	ram_block1a72,
	ram_block1a88,
	ram_block1a104,
	ram_block1a120,
	ram_block1a40,
	ram_block1a56,
	ram_block1a8,
	ram_block1a24,
	ram_block1a73,
	ram_block1a89,
	ram_block1a105,
	ram_block1a121,
	ram_block1a41,
	ram_block1a57,
	ram_block1a9,
	ram_block1a25,
	ram_block1a74,
	ram_block1a90,
	ram_block1a106,
	ram_block1a122,
	ram_block1a42,
	ram_block1a58,
	ram_block1a10,
	ram_block1a26,
	ram_block1a75,
	ram_block1a91,
	ram_block1a107,
	ram_block1a123,
	ram_block1a43,
	ram_block1a59,
	ram_block1a11,
	ram_block1a27,
	ram_block1a76,
	ram_block1a92,
	ram_block1a108,
	ram_block1a124,
	ram_block1a44,
	ram_block1a60,
	ram_block1a12,
	ram_block1a28,
	ram_block1a77,
	ram_block1a93,
	ram_block1a109,
	ram_block1a125,
	ram_block1a45,
	ram_block1a61,
	ram_block1a13,
	ram_block1a29,
	ram_block1a78,
	ram_block1a94,
	ram_block1a110,
	ram_block1a126,
	ram_block1a46,
	ram_block1a62,
	ram_block1a14,
	ram_block1a30,
	ram_block1a79,
	ram_block1a95,
	ram_block1a111,
	ram_block1a127,
	ram_block1a47,
	ram_block1a63,
	ram_block1a15,
	ram_block1a31,
	address_a,
	out_address_reg_a_2,
	out_address_reg_a_0,
	out_address_reg_a_1,
	clock0,
	clocken0)/* synthesis synthesis_greybox=1 */;
output 	ram_block1a64;
output 	ram_block1a80;
output 	ram_block1a96;
output 	ram_block1a112;
output 	ram_block1a32;
output 	ram_block1a48;
output 	ram_block1a0;
output 	ram_block1a16;
output 	ram_block1a65;
output 	ram_block1a81;
output 	ram_block1a97;
output 	ram_block1a113;
output 	ram_block1a33;
output 	ram_block1a49;
output 	ram_block1a1;
output 	ram_block1a17;
output 	ram_block1a66;
output 	ram_block1a82;
output 	ram_block1a98;
output 	ram_block1a114;
output 	ram_block1a34;
output 	ram_block1a50;
output 	ram_block1a2;
output 	ram_block1a18;
output 	ram_block1a67;
output 	ram_block1a83;
output 	ram_block1a99;
output 	ram_block1a115;
output 	ram_block1a35;
output 	ram_block1a51;
output 	ram_block1a3;
output 	ram_block1a19;
output 	ram_block1a68;
output 	ram_block1a84;
output 	ram_block1a100;
output 	ram_block1a116;
output 	ram_block1a36;
output 	ram_block1a52;
output 	ram_block1a4;
output 	ram_block1a20;
output 	ram_block1a69;
output 	ram_block1a85;
output 	ram_block1a101;
output 	ram_block1a117;
output 	ram_block1a37;
output 	ram_block1a53;
output 	ram_block1a5;
output 	ram_block1a21;
output 	ram_block1a70;
output 	ram_block1a86;
output 	ram_block1a102;
output 	ram_block1a118;
output 	ram_block1a38;
output 	ram_block1a54;
output 	ram_block1a6;
output 	ram_block1a22;
output 	ram_block1a71;
output 	ram_block1a87;
output 	ram_block1a103;
output 	ram_block1a119;
output 	ram_block1a39;
output 	ram_block1a55;
output 	ram_block1a7;
output 	ram_block1a23;
output 	ram_block1a72;
output 	ram_block1a88;
output 	ram_block1a104;
output 	ram_block1a120;
output 	ram_block1a40;
output 	ram_block1a56;
output 	ram_block1a8;
output 	ram_block1a24;
output 	ram_block1a73;
output 	ram_block1a89;
output 	ram_block1a105;
output 	ram_block1a121;
output 	ram_block1a41;
output 	ram_block1a57;
output 	ram_block1a9;
output 	ram_block1a25;
output 	ram_block1a74;
output 	ram_block1a90;
output 	ram_block1a106;
output 	ram_block1a122;
output 	ram_block1a42;
output 	ram_block1a58;
output 	ram_block1a10;
output 	ram_block1a26;
output 	ram_block1a75;
output 	ram_block1a91;
output 	ram_block1a107;
output 	ram_block1a123;
output 	ram_block1a43;
output 	ram_block1a59;
output 	ram_block1a11;
output 	ram_block1a27;
output 	ram_block1a76;
output 	ram_block1a92;
output 	ram_block1a108;
output 	ram_block1a124;
output 	ram_block1a44;
output 	ram_block1a60;
output 	ram_block1a12;
output 	ram_block1a28;
output 	ram_block1a77;
output 	ram_block1a93;
output 	ram_block1a109;
output 	ram_block1a125;
output 	ram_block1a45;
output 	ram_block1a61;
output 	ram_block1a13;
output 	ram_block1a29;
output 	ram_block1a78;
output 	ram_block1a94;
output 	ram_block1a110;
output 	ram_block1a126;
output 	ram_block1a46;
output 	ram_block1a62;
output 	ram_block1a14;
output 	ram_block1a30;
output 	ram_block1a79;
output 	ram_block1a95;
output 	ram_block1a111;
output 	ram_block1a127;
output 	ram_block1a47;
output 	ram_block1a63;
output 	ram_block1a15;
output 	ram_block1a31;
input 	[15:0] address_a;
output 	out_address_reg_a_2;
output 	out_address_reg_a_0;
output 	out_address_reg_a_1;
input 	clock0;
input 	clocken0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



DDS_48_v1_altsyncram_c8g1 auto_generated(
	.ram_block1a641(ram_block1a64),
	.ram_block1a801(ram_block1a80),
	.ram_block1a961(ram_block1a96),
	.ram_block1a1121(ram_block1a112),
	.ram_block1a321(ram_block1a32),
	.ram_block1a481(ram_block1a48),
	.ram_block1a01(ram_block1a0),
	.ram_block1a161(ram_block1a16),
	.ram_block1a651(ram_block1a65),
	.ram_block1a811(ram_block1a81),
	.ram_block1a971(ram_block1a97),
	.ram_block1a1131(ram_block1a113),
	.ram_block1a331(ram_block1a33),
	.ram_block1a491(ram_block1a49),
	.ram_block1a128(ram_block1a1),
	.ram_block1a171(ram_block1a17),
	.ram_block1a661(ram_block1a66),
	.ram_block1a821(ram_block1a82),
	.ram_block1a981(ram_block1a98),
	.ram_block1a1141(ram_block1a114),
	.ram_block1a341(ram_block1a34),
	.ram_block1a501(ram_block1a50),
	.ram_block1a210(ram_block1a2),
	.ram_block1a181(ram_block1a18),
	.ram_block1a671(ram_block1a67),
	.ram_block1a831(ram_block1a83),
	.ram_block1a991(ram_block1a99),
	.ram_block1a1151(ram_block1a115),
	.ram_block1a351(ram_block1a35),
	.ram_block1a511(ram_block1a51),
	.ram_block1a310(ram_block1a3),
	.ram_block1a191(ram_block1a19),
	.ram_block1a681(ram_block1a68),
	.ram_block1a841(ram_block1a84),
	.ram_block1a1001(ram_block1a100),
	.ram_block1a1161(ram_block1a116),
	.ram_block1a361(ram_block1a36),
	.ram_block1a521(ram_block1a52),
	.ram_block1a410(ram_block1a4),
	.ram_block1a201(ram_block1a20),
	.ram_block1a691(ram_block1a69),
	.ram_block1a851(ram_block1a85),
	.ram_block1a1011(ram_block1a101),
	.ram_block1a1171(ram_block1a117),
	.ram_block1a371(ram_block1a37),
	.ram_block1a531(ram_block1a53),
	.ram_block1a510(ram_block1a5),
	.ram_block1a211(ram_block1a21),
	.ram_block1a701(ram_block1a70),
	.ram_block1a861(ram_block1a86),
	.ram_block1a1021(ram_block1a102),
	.ram_block1a1181(ram_block1a118),
	.ram_block1a381(ram_block1a38),
	.ram_block1a541(ram_block1a54),
	.ram_block1a610(ram_block1a6),
	.ram_block1a221(ram_block1a22),
	.ram_block1a711(ram_block1a71),
	.ram_block1a871(ram_block1a87),
	.ram_block1a1031(ram_block1a103),
	.ram_block1a1191(ram_block1a119),
	.ram_block1a391(ram_block1a39),
	.ram_block1a551(ram_block1a55),
	.ram_block1a710(ram_block1a7),
	.ram_block1a231(ram_block1a23),
	.ram_block1a721(ram_block1a72),
	.ram_block1a881(ram_block1a88),
	.ram_block1a1041(ram_block1a104),
	.ram_block1a1201(ram_block1a120),
	.ram_block1a401(ram_block1a40),
	.ram_block1a561(ram_block1a56),
	.ram_block1a810(ram_block1a8),
	.ram_block1a241(ram_block1a24),
	.ram_block1a731(ram_block1a73),
	.ram_block1a891(ram_block1a89),
	.ram_block1a1051(ram_block1a105),
	.ram_block1a1211(ram_block1a121),
	.ram_block1a411(ram_block1a41),
	.ram_block1a571(ram_block1a57),
	.ram_block1a910(ram_block1a9),
	.ram_block1a251(ram_block1a25),
	.ram_block1a741(ram_block1a74),
	.ram_block1a901(ram_block1a90),
	.ram_block1a1061(ram_block1a106),
	.ram_block1a1221(ram_block1a122),
	.ram_block1a421(ram_block1a42),
	.ram_block1a581(ram_block1a58),
	.ram_block1a1010(ram_block1a10),
	.ram_block1a261(ram_block1a26),
	.ram_block1a751(ram_block1a75),
	.ram_block1a911(ram_block1a91),
	.ram_block1a1071(ram_block1a107),
	.ram_block1a1231(ram_block1a123),
	.ram_block1a431(ram_block1a43),
	.ram_block1a591(ram_block1a59),
	.ram_block1a1110(ram_block1a11),
	.ram_block1a271(ram_block1a27),
	.ram_block1a761(ram_block1a76),
	.ram_block1a921(ram_block1a92),
	.ram_block1a1081(ram_block1a108),
	.ram_block1a1241(ram_block1a124),
	.ram_block1a441(ram_block1a44),
	.ram_block1a601(ram_block1a60),
	.ram_block1a129(ram_block1a12),
	.ram_block1a281(ram_block1a28),
	.ram_block1a771(ram_block1a77),
	.ram_block1a931(ram_block1a93),
	.ram_block1a1091(ram_block1a109),
	.ram_block1a1251(ram_block1a125),
	.ram_block1a451(ram_block1a45),
	.ram_block1a611(ram_block1a61),
	.ram_block1a131(ram_block1a13),
	.ram_block1a291(ram_block1a29),
	.ram_block1a781(ram_block1a78),
	.ram_block1a941(ram_block1a94),
	.ram_block1a1101(ram_block1a110),
	.ram_block1a1261(ram_block1a126),
	.ram_block1a461(ram_block1a46),
	.ram_block1a621(ram_block1a62),
	.ram_block1a141(ram_block1a14),
	.ram_block1a301(ram_block1a30),
	.ram_block1a791(ram_block1a79),
	.ram_block1a951(ram_block1a95),
	.ram_block1a1111(ram_block1a111),
	.ram_block1a1271(ram_block1a127),
	.ram_block1a471(ram_block1a47),
	.ram_block1a631(ram_block1a63),
	.ram_block1a151(ram_block1a15),
	.ram_block1a311(ram_block1a31),
	.address_a({address_a[15],address_a[14],address_a[13],address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.out_address_reg_a_2(out_address_reg_a_2),
	.out_address_reg_a_0(out_address_reg_a_0),
	.out_address_reg_a_1(out_address_reg_a_1),
	.clock0(clock0),
	.clocken0(clocken0));

endmodule

module DDS_48_v1_altsyncram_c8g1 (
	ram_block1a641,
	ram_block1a801,
	ram_block1a961,
	ram_block1a1121,
	ram_block1a321,
	ram_block1a481,
	ram_block1a01,
	ram_block1a161,
	ram_block1a651,
	ram_block1a811,
	ram_block1a971,
	ram_block1a1131,
	ram_block1a331,
	ram_block1a491,
	ram_block1a128,
	ram_block1a171,
	ram_block1a661,
	ram_block1a821,
	ram_block1a981,
	ram_block1a1141,
	ram_block1a341,
	ram_block1a501,
	ram_block1a210,
	ram_block1a181,
	ram_block1a671,
	ram_block1a831,
	ram_block1a991,
	ram_block1a1151,
	ram_block1a351,
	ram_block1a511,
	ram_block1a310,
	ram_block1a191,
	ram_block1a681,
	ram_block1a841,
	ram_block1a1001,
	ram_block1a1161,
	ram_block1a361,
	ram_block1a521,
	ram_block1a410,
	ram_block1a201,
	ram_block1a691,
	ram_block1a851,
	ram_block1a1011,
	ram_block1a1171,
	ram_block1a371,
	ram_block1a531,
	ram_block1a510,
	ram_block1a211,
	ram_block1a701,
	ram_block1a861,
	ram_block1a1021,
	ram_block1a1181,
	ram_block1a381,
	ram_block1a541,
	ram_block1a610,
	ram_block1a221,
	ram_block1a711,
	ram_block1a871,
	ram_block1a1031,
	ram_block1a1191,
	ram_block1a391,
	ram_block1a551,
	ram_block1a710,
	ram_block1a231,
	ram_block1a721,
	ram_block1a881,
	ram_block1a1041,
	ram_block1a1201,
	ram_block1a401,
	ram_block1a561,
	ram_block1a810,
	ram_block1a241,
	ram_block1a731,
	ram_block1a891,
	ram_block1a1051,
	ram_block1a1211,
	ram_block1a411,
	ram_block1a571,
	ram_block1a910,
	ram_block1a251,
	ram_block1a741,
	ram_block1a901,
	ram_block1a1061,
	ram_block1a1221,
	ram_block1a421,
	ram_block1a581,
	ram_block1a1010,
	ram_block1a261,
	ram_block1a751,
	ram_block1a911,
	ram_block1a1071,
	ram_block1a1231,
	ram_block1a431,
	ram_block1a591,
	ram_block1a1110,
	ram_block1a271,
	ram_block1a761,
	ram_block1a921,
	ram_block1a1081,
	ram_block1a1241,
	ram_block1a441,
	ram_block1a601,
	ram_block1a129,
	ram_block1a281,
	ram_block1a771,
	ram_block1a931,
	ram_block1a1091,
	ram_block1a1251,
	ram_block1a451,
	ram_block1a611,
	ram_block1a131,
	ram_block1a291,
	ram_block1a781,
	ram_block1a941,
	ram_block1a1101,
	ram_block1a1261,
	ram_block1a461,
	ram_block1a621,
	ram_block1a141,
	ram_block1a301,
	ram_block1a791,
	ram_block1a951,
	ram_block1a1111,
	ram_block1a1271,
	ram_block1a471,
	ram_block1a631,
	ram_block1a151,
	ram_block1a311,
	address_a,
	out_address_reg_a_2,
	out_address_reg_a_0,
	out_address_reg_a_1,
	clock0,
	clocken0)/* synthesis synthesis_greybox=1 */;
output 	ram_block1a641;
output 	ram_block1a801;
output 	ram_block1a961;
output 	ram_block1a1121;
output 	ram_block1a321;
output 	ram_block1a481;
output 	ram_block1a01;
output 	ram_block1a161;
output 	ram_block1a651;
output 	ram_block1a811;
output 	ram_block1a971;
output 	ram_block1a1131;
output 	ram_block1a331;
output 	ram_block1a491;
output 	ram_block1a128;
output 	ram_block1a171;
output 	ram_block1a661;
output 	ram_block1a821;
output 	ram_block1a981;
output 	ram_block1a1141;
output 	ram_block1a341;
output 	ram_block1a501;
output 	ram_block1a210;
output 	ram_block1a181;
output 	ram_block1a671;
output 	ram_block1a831;
output 	ram_block1a991;
output 	ram_block1a1151;
output 	ram_block1a351;
output 	ram_block1a511;
output 	ram_block1a310;
output 	ram_block1a191;
output 	ram_block1a681;
output 	ram_block1a841;
output 	ram_block1a1001;
output 	ram_block1a1161;
output 	ram_block1a361;
output 	ram_block1a521;
output 	ram_block1a410;
output 	ram_block1a201;
output 	ram_block1a691;
output 	ram_block1a851;
output 	ram_block1a1011;
output 	ram_block1a1171;
output 	ram_block1a371;
output 	ram_block1a531;
output 	ram_block1a510;
output 	ram_block1a211;
output 	ram_block1a701;
output 	ram_block1a861;
output 	ram_block1a1021;
output 	ram_block1a1181;
output 	ram_block1a381;
output 	ram_block1a541;
output 	ram_block1a610;
output 	ram_block1a221;
output 	ram_block1a711;
output 	ram_block1a871;
output 	ram_block1a1031;
output 	ram_block1a1191;
output 	ram_block1a391;
output 	ram_block1a551;
output 	ram_block1a710;
output 	ram_block1a231;
output 	ram_block1a721;
output 	ram_block1a881;
output 	ram_block1a1041;
output 	ram_block1a1201;
output 	ram_block1a401;
output 	ram_block1a561;
output 	ram_block1a810;
output 	ram_block1a241;
output 	ram_block1a731;
output 	ram_block1a891;
output 	ram_block1a1051;
output 	ram_block1a1211;
output 	ram_block1a411;
output 	ram_block1a571;
output 	ram_block1a910;
output 	ram_block1a251;
output 	ram_block1a741;
output 	ram_block1a901;
output 	ram_block1a1061;
output 	ram_block1a1221;
output 	ram_block1a421;
output 	ram_block1a581;
output 	ram_block1a1010;
output 	ram_block1a261;
output 	ram_block1a751;
output 	ram_block1a911;
output 	ram_block1a1071;
output 	ram_block1a1231;
output 	ram_block1a431;
output 	ram_block1a591;
output 	ram_block1a1110;
output 	ram_block1a271;
output 	ram_block1a761;
output 	ram_block1a921;
output 	ram_block1a1081;
output 	ram_block1a1241;
output 	ram_block1a441;
output 	ram_block1a601;
output 	ram_block1a129;
output 	ram_block1a281;
output 	ram_block1a771;
output 	ram_block1a931;
output 	ram_block1a1091;
output 	ram_block1a1251;
output 	ram_block1a451;
output 	ram_block1a611;
output 	ram_block1a131;
output 	ram_block1a291;
output 	ram_block1a781;
output 	ram_block1a941;
output 	ram_block1a1101;
output 	ram_block1a1261;
output 	ram_block1a461;
output 	ram_block1a621;
output 	ram_block1a141;
output 	ram_block1a301;
output 	ram_block1a791;
output 	ram_block1a951;
output 	ram_block1a1111;
output 	ram_block1a1271;
output 	ram_block1a471;
output 	ram_block1a631;
output 	ram_block1a151;
output 	ram_block1a311;
input 	[15:0] address_a;
output 	out_address_reg_a_2;
output 	out_address_reg_a_0;
output 	out_address_reg_a_1;
input 	clock0;
input 	clocken0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \address_reg_a[2]~q ;
wire \address_reg_a[0]~q ;
wire \address_reg_a[1]~q ;

wire [143:0] ram_block1a64_PORTADATAOUT_bus;
wire [143:0] ram_block1a80_PORTADATAOUT_bus;
wire [143:0] ram_block1a96_PORTADATAOUT_bus;
wire [143:0] ram_block1a112_PORTADATAOUT_bus;
wire [143:0] ram_block1a32_PORTADATAOUT_bus;
wire [143:0] ram_block1a48_PORTADATAOUT_bus;
wire [143:0] ram_block1a0_PORTADATAOUT_bus;
wire [143:0] ram_block1a16_PORTADATAOUT_bus;
wire [143:0] ram_block1a65_PORTADATAOUT_bus;
wire [143:0] ram_block1a81_PORTADATAOUT_bus;
wire [143:0] ram_block1a97_PORTADATAOUT_bus;
wire [143:0] ram_block1a113_PORTADATAOUT_bus;
wire [143:0] ram_block1a33_PORTADATAOUT_bus;
wire [143:0] ram_block1a49_PORTADATAOUT_bus;
wire [143:0] ram_block1a1_PORTADATAOUT_bus;
wire [143:0] ram_block1a17_PORTADATAOUT_bus;
wire [143:0] ram_block1a66_PORTADATAOUT_bus;
wire [143:0] ram_block1a82_PORTADATAOUT_bus;
wire [143:0] ram_block1a98_PORTADATAOUT_bus;
wire [143:0] ram_block1a114_PORTADATAOUT_bus;
wire [143:0] ram_block1a34_PORTADATAOUT_bus;
wire [143:0] ram_block1a50_PORTADATAOUT_bus;
wire [143:0] ram_block1a2_PORTADATAOUT_bus;
wire [143:0] ram_block1a18_PORTADATAOUT_bus;
wire [143:0] ram_block1a67_PORTADATAOUT_bus;
wire [143:0] ram_block1a83_PORTADATAOUT_bus;
wire [143:0] ram_block1a99_PORTADATAOUT_bus;
wire [143:0] ram_block1a115_PORTADATAOUT_bus;
wire [143:0] ram_block1a35_PORTADATAOUT_bus;
wire [143:0] ram_block1a51_PORTADATAOUT_bus;
wire [143:0] ram_block1a3_PORTADATAOUT_bus;
wire [143:0] ram_block1a19_PORTADATAOUT_bus;
wire [143:0] ram_block1a68_PORTADATAOUT_bus;
wire [143:0] ram_block1a84_PORTADATAOUT_bus;
wire [143:0] ram_block1a100_PORTADATAOUT_bus;
wire [143:0] ram_block1a116_PORTADATAOUT_bus;
wire [143:0] ram_block1a36_PORTADATAOUT_bus;
wire [143:0] ram_block1a52_PORTADATAOUT_bus;
wire [143:0] ram_block1a4_PORTADATAOUT_bus;
wire [143:0] ram_block1a20_PORTADATAOUT_bus;
wire [143:0] ram_block1a69_PORTADATAOUT_bus;
wire [143:0] ram_block1a85_PORTADATAOUT_bus;
wire [143:0] ram_block1a101_PORTADATAOUT_bus;
wire [143:0] ram_block1a117_PORTADATAOUT_bus;
wire [143:0] ram_block1a37_PORTADATAOUT_bus;
wire [143:0] ram_block1a53_PORTADATAOUT_bus;
wire [143:0] ram_block1a5_PORTADATAOUT_bus;
wire [143:0] ram_block1a21_PORTADATAOUT_bus;
wire [143:0] ram_block1a70_PORTADATAOUT_bus;
wire [143:0] ram_block1a86_PORTADATAOUT_bus;
wire [143:0] ram_block1a102_PORTADATAOUT_bus;
wire [143:0] ram_block1a118_PORTADATAOUT_bus;
wire [143:0] ram_block1a38_PORTADATAOUT_bus;
wire [143:0] ram_block1a54_PORTADATAOUT_bus;
wire [143:0] ram_block1a6_PORTADATAOUT_bus;
wire [143:0] ram_block1a22_PORTADATAOUT_bus;
wire [143:0] ram_block1a71_PORTADATAOUT_bus;
wire [143:0] ram_block1a87_PORTADATAOUT_bus;
wire [143:0] ram_block1a103_PORTADATAOUT_bus;
wire [143:0] ram_block1a119_PORTADATAOUT_bus;
wire [143:0] ram_block1a39_PORTADATAOUT_bus;
wire [143:0] ram_block1a55_PORTADATAOUT_bus;
wire [143:0] ram_block1a7_PORTADATAOUT_bus;
wire [143:0] ram_block1a23_PORTADATAOUT_bus;
wire [143:0] ram_block1a72_PORTADATAOUT_bus;
wire [143:0] ram_block1a88_PORTADATAOUT_bus;
wire [143:0] ram_block1a104_PORTADATAOUT_bus;
wire [143:0] ram_block1a120_PORTADATAOUT_bus;
wire [143:0] ram_block1a40_PORTADATAOUT_bus;
wire [143:0] ram_block1a56_PORTADATAOUT_bus;
wire [143:0] ram_block1a8_PORTADATAOUT_bus;
wire [143:0] ram_block1a24_PORTADATAOUT_bus;
wire [143:0] ram_block1a73_PORTADATAOUT_bus;
wire [143:0] ram_block1a89_PORTADATAOUT_bus;
wire [143:0] ram_block1a105_PORTADATAOUT_bus;
wire [143:0] ram_block1a121_PORTADATAOUT_bus;
wire [143:0] ram_block1a41_PORTADATAOUT_bus;
wire [143:0] ram_block1a57_PORTADATAOUT_bus;
wire [143:0] ram_block1a9_PORTADATAOUT_bus;
wire [143:0] ram_block1a25_PORTADATAOUT_bus;
wire [143:0] ram_block1a74_PORTADATAOUT_bus;
wire [143:0] ram_block1a90_PORTADATAOUT_bus;
wire [143:0] ram_block1a106_PORTADATAOUT_bus;
wire [143:0] ram_block1a122_PORTADATAOUT_bus;
wire [143:0] ram_block1a42_PORTADATAOUT_bus;
wire [143:0] ram_block1a58_PORTADATAOUT_bus;
wire [143:0] ram_block1a10_PORTADATAOUT_bus;
wire [143:0] ram_block1a26_PORTADATAOUT_bus;
wire [143:0] ram_block1a75_PORTADATAOUT_bus;
wire [143:0] ram_block1a91_PORTADATAOUT_bus;
wire [143:0] ram_block1a107_PORTADATAOUT_bus;
wire [143:0] ram_block1a123_PORTADATAOUT_bus;
wire [143:0] ram_block1a43_PORTADATAOUT_bus;
wire [143:0] ram_block1a59_PORTADATAOUT_bus;
wire [143:0] ram_block1a11_PORTADATAOUT_bus;
wire [143:0] ram_block1a27_PORTADATAOUT_bus;
wire [143:0] ram_block1a76_PORTADATAOUT_bus;
wire [143:0] ram_block1a92_PORTADATAOUT_bus;
wire [143:0] ram_block1a108_PORTADATAOUT_bus;
wire [143:0] ram_block1a124_PORTADATAOUT_bus;
wire [143:0] ram_block1a44_PORTADATAOUT_bus;
wire [143:0] ram_block1a60_PORTADATAOUT_bus;
wire [143:0] ram_block1a12_PORTADATAOUT_bus;
wire [143:0] ram_block1a28_PORTADATAOUT_bus;
wire [143:0] ram_block1a77_PORTADATAOUT_bus;
wire [143:0] ram_block1a93_PORTADATAOUT_bus;
wire [143:0] ram_block1a109_PORTADATAOUT_bus;
wire [143:0] ram_block1a125_PORTADATAOUT_bus;
wire [143:0] ram_block1a45_PORTADATAOUT_bus;
wire [143:0] ram_block1a61_PORTADATAOUT_bus;
wire [143:0] ram_block1a13_PORTADATAOUT_bus;
wire [143:0] ram_block1a29_PORTADATAOUT_bus;
wire [143:0] ram_block1a78_PORTADATAOUT_bus;
wire [143:0] ram_block1a94_PORTADATAOUT_bus;
wire [143:0] ram_block1a110_PORTADATAOUT_bus;
wire [143:0] ram_block1a126_PORTADATAOUT_bus;
wire [143:0] ram_block1a46_PORTADATAOUT_bus;
wire [143:0] ram_block1a62_PORTADATAOUT_bus;
wire [143:0] ram_block1a14_PORTADATAOUT_bus;
wire [143:0] ram_block1a30_PORTADATAOUT_bus;
wire [143:0] ram_block1a79_PORTADATAOUT_bus;
wire [143:0] ram_block1a95_PORTADATAOUT_bus;
wire [143:0] ram_block1a111_PORTADATAOUT_bus;
wire [143:0] ram_block1a127_PORTADATAOUT_bus;
wire [143:0] ram_block1a47_PORTADATAOUT_bus;
wire [143:0] ram_block1a63_PORTADATAOUT_bus;
wire [143:0] ram_block1a15_PORTADATAOUT_bus;
wire [143:0] ram_block1a31_PORTADATAOUT_bus;

assign ram_block1a641 = ram_block1a64_PORTADATAOUT_bus[0];

assign ram_block1a801 = ram_block1a80_PORTADATAOUT_bus[0];

assign ram_block1a961 = ram_block1a96_PORTADATAOUT_bus[0];

assign ram_block1a1121 = ram_block1a112_PORTADATAOUT_bus[0];

assign ram_block1a321 = ram_block1a32_PORTADATAOUT_bus[0];

assign ram_block1a481 = ram_block1a48_PORTADATAOUT_bus[0];

assign ram_block1a01 = ram_block1a0_PORTADATAOUT_bus[0];

assign ram_block1a161 = ram_block1a16_PORTADATAOUT_bus[0];

assign ram_block1a651 = ram_block1a65_PORTADATAOUT_bus[0];

assign ram_block1a811 = ram_block1a81_PORTADATAOUT_bus[0];

assign ram_block1a971 = ram_block1a97_PORTADATAOUT_bus[0];

assign ram_block1a1131 = ram_block1a113_PORTADATAOUT_bus[0];

assign ram_block1a331 = ram_block1a33_PORTADATAOUT_bus[0];

assign ram_block1a491 = ram_block1a49_PORTADATAOUT_bus[0];

assign ram_block1a128 = ram_block1a1_PORTADATAOUT_bus[0];

assign ram_block1a171 = ram_block1a17_PORTADATAOUT_bus[0];

assign ram_block1a661 = ram_block1a66_PORTADATAOUT_bus[0];

assign ram_block1a821 = ram_block1a82_PORTADATAOUT_bus[0];

assign ram_block1a981 = ram_block1a98_PORTADATAOUT_bus[0];

assign ram_block1a1141 = ram_block1a114_PORTADATAOUT_bus[0];

assign ram_block1a341 = ram_block1a34_PORTADATAOUT_bus[0];

assign ram_block1a501 = ram_block1a50_PORTADATAOUT_bus[0];

assign ram_block1a210 = ram_block1a2_PORTADATAOUT_bus[0];

assign ram_block1a181 = ram_block1a18_PORTADATAOUT_bus[0];

assign ram_block1a671 = ram_block1a67_PORTADATAOUT_bus[0];

assign ram_block1a831 = ram_block1a83_PORTADATAOUT_bus[0];

assign ram_block1a991 = ram_block1a99_PORTADATAOUT_bus[0];

assign ram_block1a1151 = ram_block1a115_PORTADATAOUT_bus[0];

assign ram_block1a351 = ram_block1a35_PORTADATAOUT_bus[0];

assign ram_block1a511 = ram_block1a51_PORTADATAOUT_bus[0];

assign ram_block1a310 = ram_block1a3_PORTADATAOUT_bus[0];

assign ram_block1a191 = ram_block1a19_PORTADATAOUT_bus[0];

assign ram_block1a681 = ram_block1a68_PORTADATAOUT_bus[0];

assign ram_block1a841 = ram_block1a84_PORTADATAOUT_bus[0];

assign ram_block1a1001 = ram_block1a100_PORTADATAOUT_bus[0];

assign ram_block1a1161 = ram_block1a116_PORTADATAOUT_bus[0];

assign ram_block1a361 = ram_block1a36_PORTADATAOUT_bus[0];

assign ram_block1a521 = ram_block1a52_PORTADATAOUT_bus[0];

assign ram_block1a410 = ram_block1a4_PORTADATAOUT_bus[0];

assign ram_block1a201 = ram_block1a20_PORTADATAOUT_bus[0];

assign ram_block1a691 = ram_block1a69_PORTADATAOUT_bus[0];

assign ram_block1a851 = ram_block1a85_PORTADATAOUT_bus[0];

assign ram_block1a1011 = ram_block1a101_PORTADATAOUT_bus[0];

assign ram_block1a1171 = ram_block1a117_PORTADATAOUT_bus[0];

assign ram_block1a371 = ram_block1a37_PORTADATAOUT_bus[0];

assign ram_block1a531 = ram_block1a53_PORTADATAOUT_bus[0];

assign ram_block1a510 = ram_block1a5_PORTADATAOUT_bus[0];

assign ram_block1a211 = ram_block1a21_PORTADATAOUT_bus[0];

assign ram_block1a701 = ram_block1a70_PORTADATAOUT_bus[0];

assign ram_block1a861 = ram_block1a86_PORTADATAOUT_bus[0];

assign ram_block1a1021 = ram_block1a102_PORTADATAOUT_bus[0];

assign ram_block1a1181 = ram_block1a118_PORTADATAOUT_bus[0];

assign ram_block1a381 = ram_block1a38_PORTADATAOUT_bus[0];

assign ram_block1a541 = ram_block1a54_PORTADATAOUT_bus[0];

assign ram_block1a610 = ram_block1a6_PORTADATAOUT_bus[0];

assign ram_block1a221 = ram_block1a22_PORTADATAOUT_bus[0];

assign ram_block1a711 = ram_block1a71_PORTADATAOUT_bus[0];

assign ram_block1a871 = ram_block1a87_PORTADATAOUT_bus[0];

assign ram_block1a1031 = ram_block1a103_PORTADATAOUT_bus[0];

assign ram_block1a1191 = ram_block1a119_PORTADATAOUT_bus[0];

assign ram_block1a391 = ram_block1a39_PORTADATAOUT_bus[0];

assign ram_block1a551 = ram_block1a55_PORTADATAOUT_bus[0];

assign ram_block1a710 = ram_block1a7_PORTADATAOUT_bus[0];

assign ram_block1a231 = ram_block1a23_PORTADATAOUT_bus[0];

assign ram_block1a721 = ram_block1a72_PORTADATAOUT_bus[0];

assign ram_block1a881 = ram_block1a88_PORTADATAOUT_bus[0];

assign ram_block1a1041 = ram_block1a104_PORTADATAOUT_bus[0];

assign ram_block1a1201 = ram_block1a120_PORTADATAOUT_bus[0];

assign ram_block1a401 = ram_block1a40_PORTADATAOUT_bus[0];

assign ram_block1a561 = ram_block1a56_PORTADATAOUT_bus[0];

assign ram_block1a810 = ram_block1a8_PORTADATAOUT_bus[0];

assign ram_block1a241 = ram_block1a24_PORTADATAOUT_bus[0];

assign ram_block1a731 = ram_block1a73_PORTADATAOUT_bus[0];

assign ram_block1a891 = ram_block1a89_PORTADATAOUT_bus[0];

assign ram_block1a1051 = ram_block1a105_PORTADATAOUT_bus[0];

assign ram_block1a1211 = ram_block1a121_PORTADATAOUT_bus[0];

assign ram_block1a411 = ram_block1a41_PORTADATAOUT_bus[0];

assign ram_block1a571 = ram_block1a57_PORTADATAOUT_bus[0];

assign ram_block1a910 = ram_block1a9_PORTADATAOUT_bus[0];

assign ram_block1a251 = ram_block1a25_PORTADATAOUT_bus[0];

assign ram_block1a741 = ram_block1a74_PORTADATAOUT_bus[0];

assign ram_block1a901 = ram_block1a90_PORTADATAOUT_bus[0];

assign ram_block1a1061 = ram_block1a106_PORTADATAOUT_bus[0];

assign ram_block1a1221 = ram_block1a122_PORTADATAOUT_bus[0];

assign ram_block1a421 = ram_block1a42_PORTADATAOUT_bus[0];

assign ram_block1a581 = ram_block1a58_PORTADATAOUT_bus[0];

assign ram_block1a1010 = ram_block1a10_PORTADATAOUT_bus[0];

assign ram_block1a261 = ram_block1a26_PORTADATAOUT_bus[0];

assign ram_block1a751 = ram_block1a75_PORTADATAOUT_bus[0];

assign ram_block1a911 = ram_block1a91_PORTADATAOUT_bus[0];

assign ram_block1a1071 = ram_block1a107_PORTADATAOUT_bus[0];

assign ram_block1a1231 = ram_block1a123_PORTADATAOUT_bus[0];

assign ram_block1a431 = ram_block1a43_PORTADATAOUT_bus[0];

assign ram_block1a591 = ram_block1a59_PORTADATAOUT_bus[0];

assign ram_block1a1110 = ram_block1a11_PORTADATAOUT_bus[0];

assign ram_block1a271 = ram_block1a27_PORTADATAOUT_bus[0];

assign ram_block1a761 = ram_block1a76_PORTADATAOUT_bus[0];

assign ram_block1a921 = ram_block1a92_PORTADATAOUT_bus[0];

assign ram_block1a1081 = ram_block1a108_PORTADATAOUT_bus[0];

assign ram_block1a1241 = ram_block1a124_PORTADATAOUT_bus[0];

assign ram_block1a441 = ram_block1a44_PORTADATAOUT_bus[0];

assign ram_block1a601 = ram_block1a60_PORTADATAOUT_bus[0];

assign ram_block1a129 = ram_block1a12_PORTADATAOUT_bus[0];

assign ram_block1a281 = ram_block1a28_PORTADATAOUT_bus[0];

assign ram_block1a771 = ram_block1a77_PORTADATAOUT_bus[0];

assign ram_block1a931 = ram_block1a93_PORTADATAOUT_bus[0];

assign ram_block1a1091 = ram_block1a109_PORTADATAOUT_bus[0];

assign ram_block1a1251 = ram_block1a125_PORTADATAOUT_bus[0];

assign ram_block1a451 = ram_block1a45_PORTADATAOUT_bus[0];

assign ram_block1a611 = ram_block1a61_PORTADATAOUT_bus[0];

assign ram_block1a131 = ram_block1a13_PORTADATAOUT_bus[0];

assign ram_block1a291 = ram_block1a29_PORTADATAOUT_bus[0];

assign ram_block1a781 = ram_block1a78_PORTADATAOUT_bus[0];

assign ram_block1a941 = ram_block1a94_PORTADATAOUT_bus[0];

assign ram_block1a1101 = ram_block1a110_PORTADATAOUT_bus[0];

assign ram_block1a1261 = ram_block1a126_PORTADATAOUT_bus[0];

assign ram_block1a461 = ram_block1a46_PORTADATAOUT_bus[0];

assign ram_block1a621 = ram_block1a62_PORTADATAOUT_bus[0];

assign ram_block1a141 = ram_block1a14_PORTADATAOUT_bus[0];

assign ram_block1a301 = ram_block1a30_PORTADATAOUT_bus[0];

assign ram_block1a791 = ram_block1a79_PORTADATAOUT_bus[0];

assign ram_block1a951 = ram_block1a95_PORTADATAOUT_bus[0];

assign ram_block1a1111 = ram_block1a111_PORTADATAOUT_bus[0];

assign ram_block1a1271 = ram_block1a127_PORTADATAOUT_bus[0];

assign ram_block1a471 = ram_block1a47_PORTADATAOUT_bus[0];

assign ram_block1a631 = ram_block1a63_PORTADATAOUT_bus[0];

assign ram_block1a151 = ram_block1a15_PORTADATAOUT_bus[0];

assign ram_block1a311 = ram_block1a31_PORTADATAOUT_bus[0];

arriav_ram_block ram_block1a64(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a64_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a64.clk0_core_clock_enable = "ena0";
defparam ram_block1a64.clk0_input_clock_enable = "ena0";
defparam ram_block1a64.clk0_output_clock_enable = "ena0";
defparam ram_block1a64.data_interleave_offset_in_bits = 1;
defparam ram_block1a64.data_interleave_width_in_bits = 1;
defparam ram_block1a64.init_file = "DDS_48_v1_nco_ii_0_sin.hex";
defparam ram_block1a64.init_file_layout = "port_a";
defparam ram_block1a64.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_c8g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a64.operation_mode = "rom";
defparam ram_block1a64.port_a_address_clear = "none";
defparam ram_block1a64.port_a_address_width = 13;
defparam ram_block1a64.port_a_data_out_clear = "none";
defparam ram_block1a64.port_a_data_out_clock = "clock0";
defparam ram_block1a64.port_a_data_width = 1;
defparam ram_block1a64.port_a_first_address = 32768;
defparam ram_block1a64.port_a_first_bit_number = 0;
defparam ram_block1a64.port_a_last_address = 40959;
defparam ram_block1a64.port_a_logical_ram_depth = 65536;
defparam ram_block1a64.port_a_logical_ram_width = 16;
defparam ram_block1a64.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a64.ram_block_type = "auto";
defparam ram_block1a64.mem_init3 = "783C1E1F0F8783C3C1E1E1F0F0F0F0F0F0F0F0F0F0F0E1E1E1C3C387870F1E1C3C78F0E1C3870E1C3871E3C78E1C78E1C78E3C71E38F1C70E38E1C71C71E38E38E38E38E38E38E38E39C71C718E38E71C738E31C738E71CE39C638C738C738C739C639CE318C739CE318C6318C6318C6318C6739CE6318CE7318CE6319CC67319CC673198CE633198CC6733198CC66733998CCC6673339998CCCE6663333399999CCCCCCC6666666673333333333333333333333333332666666666CCCCCCD99999333326664CCC99993336664CC999332664CD99B3266CC99B3664C99B366CC993264C99366CD9B264D9B264D9B26CD9364D9B26C9B26C9B26C9B24D93649B2";
defparam ram_block1a64.mem_init2 = "6D936C9B64DB24DB24DB24DB24DB249B6C936D9249B6C924DB6D924936DB6D924924936DB6DB6DB6DB6DB6DB6DB6DB6DB692492496DB6DA4924B6DB4925B6D2496DA496DB496DA496D24B6925B496D25B496D25B4B692D25B4B696D2DA5B4B49696D2D2DA5A5A5B4B4B4B4B4B4B4B4B4B4B4B4B4B4A5A5A5AD2D29696B4B5A5AD2D694B4A5AD296B4A5AD694A5AD694A5AD6B4A5294A52D6B5AD6B5AD6B5294A5294AD6B5294A56B5295AD6A56B5295A94AD4A56A56A56B52B52B52B56A56A56AD4AD4A95AB52A56AD5A952A56AD5AB56AD5AB56AD52A54A956AD52A55AA54AB54AB54AB54AB54AA55AA552AD56AB55AAD52AB55AAD56AA552AB552A955AA955";
defparam ram_block1a64.mem_init1 = "2AB552AA554AA9552AA554AAB556AA9556AA9554AAA555AAA9554AAAD554AAAD554AAA95556AAAD5556AAA95554AAAAD5554AAAA955556AAAAB55555AAAAAB555554AAAAAA5555554AAAAAAAD55555552AAAAAAAA95555555555AAAAAAAAAAAAAD5555555555555555556AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAD55555555555555555552AAAAAAAAAAAAA55555555555AAAAAAAAAB555555556AAAAAAA95555554AAAAAAB5555552AAAAA9555556AAAAAD55554AAAAA555552AAAAD55552AAAB55556AAAA55556AAAB5555AAAAD5552AAAD5552AAA5555AAAB5552AAA5556AAAD554AAAD556AAA5552AAB555AAAD556AA9554AAB555";
defparam ram_block1a64.mem_init0 = "AAA555AAA555AAA555AAA554AAB556AAD552AA554AA9552AA554AAD55AAB552AA556AAD54AAD54AA955AA955AA955AA954AAD54AAD56AA552AB55AA954AAD56AB552A954AA552A955AAD56AB55AA552A954AA552AD56AB54AA552AD56A954AA55AA552AD56A956AB54AB55AA55AA552AD52AD52AD52AD52A956A956A956AD52AD52AD52AD52AD5AA55AA54AB54AB56A956AD52AD5AA55AB54AB56A952AD5AA54AB56A952AD5AA54AB56A952A55AB54A952AD5AB54A952AD5AB54A952AD5AB56A952A54AB56AD5AA54A952A55AB56AD5AA54A952A54AB56AD5AB56AD5AA54A952A54A952AD5AB56AD5AB56AD5AB54A952A54A952A54A952A54A956AD5AB56AD5A";

arriav_ram_block ram_block1a80(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a80_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a80.clk0_core_clock_enable = "ena0";
defparam ram_block1a80.clk0_input_clock_enable = "ena0";
defparam ram_block1a80.clk0_output_clock_enable = "ena0";
defparam ram_block1a80.data_interleave_offset_in_bits = 1;
defparam ram_block1a80.data_interleave_width_in_bits = 1;
defparam ram_block1a80.init_file = "DDS_48_v1_nco_ii_0_sin.hex";
defparam ram_block1a80.init_file_layout = "port_a";
defparam ram_block1a80.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_c8g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a80.operation_mode = "rom";
defparam ram_block1a80.port_a_address_clear = "none";
defparam ram_block1a80.port_a_address_width = 13;
defparam ram_block1a80.port_a_data_out_clear = "none";
defparam ram_block1a80.port_a_data_out_clock = "clock0";
defparam ram_block1a80.port_a_data_width = 1;
defparam ram_block1a80.port_a_first_address = 40960;
defparam ram_block1a80.port_a_first_bit_number = 0;
defparam ram_block1a80.port_a_last_address = 49151;
defparam ram_block1a80.port_a_logical_ram_depth = 65536;
defparam ram_block1a80.port_a_logical_ram_width = 16;
defparam ram_block1a80.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a80.ram_block_type = "auto";
defparam ram_block1a80.mem_init3 = "FFFFFFFFFFFFFF80000000001FFFFFFF000000FFFFF00001FFFE0001FFF8001FFF000FFF001FFC00FFE00FFC01FF007FC01FE01FE01FE03FC07F01FC07F01F80FC07E07E07E07E07E0FC0F81F03E0F81F07C1F07C1F0783E0F07C3E1F0F87C3C1E1E0F0F0F07878787878F0F0F0E1E1C3C7870F1E3C78F1E3C78E1C38F1C78E1C70E38E1C71C70E38E38E38E38E39C71C718E38C71CE39C738E718E718E718C739C6318E739CE739CE6318C67398C67318CE63399CC673399CCE6733198CCC6673331999CCCCCE666667333333333333333333333333326666664CCCC99993332666CCD99B3266CC99B3264CD9B366CD9B264C9B364D9B26C9B26C9B26C9B24D";
defparam ram_block1a80.mem_init2 = "926C936C9B64936C926D9249B6D924936DB6DB2492492492492496DB6DB492496DB4925B6925B692DB496D25B49692D25B4B49696D2D2D25A5A5A5A5A52D2D2D69694B4A5AD296B4A5AD694A5294B5AD6B5294A52B5AD4A56B52B5A95A95A95A952B52A56AD5A952A54A956AD52A55AA55AA552AD56AB55AA954AAD55AA9552AA555AAAD552AAB5552AAA55552AAA955556AAAAA5555556AAAAAAAA55555555555555556AAAAAAAAAB55555555555555552AAAAAAAB5555552AAAAB55554AAAAD5552AAA5554AAA5552AA9552AAD55AAB552AB552A954AA552A956AB54AB54AB56A952A54A952A54A95AB52A56A56AD4AD4A56A56B52B5AD4A56B5AD4A5294A5";
defparam ram_block1a80.mem_init1 = "294B5AD6B4A52D694B5A52D696B4B4A5A5A52D2D2D2D2D2D2D25A5A5B4B49692D25A4B692DA4B692DA496D24B6D2496DB4924B6DB6924924924B6DB6DB64924924936DB6C9249B6C924DB249B64936C9B649B24D926C9B24D9364D9364C9B26CD9326CD93264C993264C9933664C99B33664CC999332666CCCD999B3333666666CCCCCCCCCC99999999999998CCCCCCCCCC666667333319998CCC666333199CCE6633198CC663399CC67319CC67398CE7318CE739CC6318C6318C6318E739C631CE718E738C718E718E31C638E71C638E31C71C738E38E38E38E38E38E3871C71C38E3871C78E1C70E3C70E3C78F1C3870E1C3C78F0E1C3C3878F0F0E1E1E1E3";
defparam ram_block1a80.mem_init0 = "C3C3C3C3C3E1E1E1E0F0F0787C3E1E0F0783C1F0F83C1F07C3E0F83E0F83F07C1F03E0FC1F83F03E07E07E0FC0FC07E07E03F01F80FE07F01FC07F00FE01FC03FC03FC03FC01FE00FF803FE007FE007FE007FF001FFC003FFC001FFF0003FFF0001FFFE0000FFFFC00003FFFFF0000003FFFFFFF00000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000FFFFFFFE000000FFFFFE00001FFFF80001FFFE0003FFF8001FFF0007FF8007FF800FFE007FF003FF003FE007FC01FF00FF807F803FC03F807F80FF01FC07F80FC07F01FC0FE07F03F03F81F81F81F81F03F03E07E0FC1F03E07C1F03E0F83E0F83E0F83E1F07C1E0F87C1E0F0";

arriav_ram_block ram_block1a96(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a96_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a96.clk0_core_clock_enable = "ena0";
defparam ram_block1a96.clk0_input_clock_enable = "ena0";
defparam ram_block1a96.clk0_output_clock_enable = "ena0";
defparam ram_block1a96.data_interleave_offset_in_bits = 1;
defparam ram_block1a96.data_interleave_width_in_bits = 1;
defparam ram_block1a96.init_file = "DDS_48_v1_nco_ii_0_sin.hex";
defparam ram_block1a96.init_file_layout = "port_a";
defparam ram_block1a96.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_c8g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a96.operation_mode = "rom";
defparam ram_block1a96.port_a_address_clear = "none";
defparam ram_block1a96.port_a_address_width = 13;
defparam ram_block1a96.port_a_data_out_clear = "none";
defparam ram_block1a96.port_a_data_out_clock = "clock0";
defparam ram_block1a96.port_a_data_width = 1;
defparam ram_block1a96.port_a_first_address = 49152;
defparam ram_block1a96.port_a_first_bit_number = 0;
defparam ram_block1a96.port_a_last_address = 57343;
defparam ram_block1a96.port_a_logical_ram_depth = 65536;
defparam ram_block1a96.port_a_logical_ram_width = 16;
defparam ram_block1a96.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a96.ram_block_type = "auto";
defparam ram_block1a96.mem_init3 = "1E0F07C3E0F07C1F0F83E0F83E0F83E0F81F07C0F81F07E0FC0F81F81F03F03F03F03F81F81FC0FE07F01FC07E03FC07F01FE03FC03F807F803FC03FE01FF007FC00FF801FF801FFC00FFE003FFC003FFC001FFF0003FFF8000FFFF00003FFFF00000FFFFFE000000FFFFFFFE0000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000001FFFFFFF8000001FFFFF800007FFFE0000FFFF0001FFF8001FFF0007FF8007FF001FFC00FFC00FFC00FF803FE00FF007F807F807F807F00FE01FC07F01FC0FE03F01F80FC0FC07E07E0FC0FC0F81F83F07E0F81F07C1F83E0F83E0F87C1F0783E1F0783C1E0F0F87C3C1E1E0F0F0F0F8787878787";
defparam ram_block1a96.mem_init2 = "8F0F0F0E1E1E3C387870E1E3C7870E1C3871E3C78E1C78E1C70E3C71C38E3871C71C38E38E38E38E38E38E39C71C718E38C71CE38C718E31CE31C639CE31CE718C739CE318C6318C6318C6739CE6319CE6339CC67319CC673398CC6633198CCE67331998CCC666333319999CCCCCC6666666666333333333333326666666666CCCCCD9999B3336666CCC999332664CD99B3264CD993264C993264C99366C99366C9B264D9364D93649B26C93649B24DB26D924DB249B64926DB24926DB6D924924924DB6DB6DA492492492DB6DA4925B6D2496DA496D24B692DA4B692DA4B49692D25A5B4B4B49696969696969694B4B4A5A5AD2D694B5A52D694A5AD6B5A529";
defparam ram_block1a96.mem_init1 = "4A5294A56B5AD4A56B5A95AD4AD4A56A56AD4AD4A95AB52A54A952A54A952AD5AA55AA55AAD52A954AA552A955AA955AAB556AA9552AA9554AAA5554AAA95556AAAA55555AAAAA9555555AAAAAAAA95555555555555555AAAAAAAAAAD5555555555555554AAAAAAAAD555554AAAAAD55552AAA95554AAA9555AAA9556AAB554AA9552AB556AA552AB55AAD56A954AB54AB54A956AD52A54A952B56AD4A95A952B52B52B52B5A95AD4A56B5A94A5295AD6B5A5294A52D6B4A5AD296B4A5A52D2D6969694B4B4B4B4B4969696D2D25A5B49692D25B496D25B692DB492DB4925B6D24925B6DB6D249249249249249B6DB6D924936DB24936C926D924DB26D926C93";
defparam ram_block1a96.mem_init0 = "649B26C9B26C9B26C9B364D9B264C9B366CD9B3664C99B3266CC99B33666CCC9999333266664CCCCCC99999999999999999999999999CCCCCCE666673331999CCC66633199CCE673399CC673398CE6319CC6339CC6318CE739CE739CE318C739C631CE31CE31CE39C738E71C638E31C71C738E38E38E38E38E1C71C70E38E1C70E3C71E3870E3C78F1E3C78F1E1C3C7870F0E1E1E1E3C3C3C3C3C1E1E1E0F0F0787C3E1F0F87C1E0F83C1F07C1F07C1F03E0F81F03E07E0FC0FC0FC0FC0FC07E03F01FC07F01FC07F80FF00FF00FF007FC01FF007FE00FFE007FF001FFE001FFF0003FFF0000FFFF00001FFFFE000001FFFFFFF00000000003FFFFFFFFFFFFFF";

arriav_ram_block ram_block1a112(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a112_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a112.clk0_core_clock_enable = "ena0";
defparam ram_block1a112.clk0_input_clock_enable = "ena0";
defparam ram_block1a112.clk0_output_clock_enable = "ena0";
defparam ram_block1a112.data_interleave_offset_in_bits = 1;
defparam ram_block1a112.data_interleave_width_in_bits = 1;
defparam ram_block1a112.init_file = "DDS_48_v1_nco_ii_0_sin.hex";
defparam ram_block1a112.init_file_layout = "port_a";
defparam ram_block1a112.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_c8g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a112.operation_mode = "rom";
defparam ram_block1a112.port_a_address_clear = "none";
defparam ram_block1a112.port_a_address_width = 13;
defparam ram_block1a112.port_a_data_out_clear = "none";
defparam ram_block1a112.port_a_data_out_clock = "clock0";
defparam ram_block1a112.port_a_data_width = 1;
defparam ram_block1a112.port_a_first_address = 57344;
defparam ram_block1a112.port_a_first_bit_number = 0;
defparam ram_block1a112.port_a_last_address = 65535;
defparam ram_block1a112.port_a_logical_ram_depth = 65536;
defparam ram_block1a112.port_a_logical_ram_width = 16;
defparam ram_block1a112.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a112.ram_block_type = "auto";
defparam ram_block1a112.mem_init3 = "B56AD5AB56AD52A54A952A54A952A54A952A55AB56AD5AB56AD5AB56A952A54A952A54AB56AD5AB56AD5AA54A952A54AB56AD5AB54A952A54AB56AD5AA54A952AD5AB56A952A55AB56A952A55AB56A952A55AB54A952AD5AA54AB56A952AD5AA54AB56A952AD5AA55AB54AB56A956AD52AD5AA55AA54AB54AB56A956A956A956A956AD52AD52AD52A956A956A956A956A954AB54AB55AA55AAD52AD56A954AB54AA552AD56A954AA55AAD56A954AA552A954AB55AAD56AB552A954AA552A955AAD56AA552AB55AA954AAD56AA556AA552AB552AB552AB552AA556AA556AAD54AA955AAB556AA554AA9552AA554AA9556AAD55AAA554AAB554AAB554AAB554AAB";
defparam ram_block1a112.mem_init2 = "555AAA5552AAD556AAB555AAA9554AAAD556AAA5556AAAD554AAA9555AAAB5554AAA95556AAA95556AAAB5555AAAAD5554AAAAD5555AAAA955556AAAA955554AAAAA555556AAAAAD555552AAAAA9555555AAAAAAA55555552AAAAAAAD55555555AAAAAAAAAB55555555554AAAAAAAAAAAAA955555555555555555556AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAD5555555555555555556AAAAAAAAAAAAB55555555552AAAAAAAA955555556AAAAAAA5555554AAAAAA555555AAAAAB55555AAAAAD55552AAAA55556AAAA55552AAAD5556AAAD5552AAA5556AAA5556AAA5552AAB554AAA5552AAD552AAD55AAA554AA9552AA554AA955AA9";
defparam ram_block1a112.mem_init1 = "552AB552A955AA954AAD56AB55AA956AB55AAD56A954AB54AA55AA55AA55AA55AA54AB54A956AD52A54A956AD5AB56AD5AB56AD4A952B56AD4A95AB52A56A56AD4AD4AD5A95A95A95AD4AD4AD4A56A52B5295AD4AD6B5295AD4A5295AD6A5294A5295AD6B5AD6B5AD694A5294A5AD6B4A52D6B4A52D6B4A5AD296B4A5A52D696B4B5A5AD2D29696B4B4B4A5A5A5A5A5A5A5A5A5A5A5A5A5A5B4B4B4B69696D2D25A5B4B696D2DA5B49692DA5B496D25B496D25B492DA496D24B6D25B6D24B6D2496DB4925B6DA4924B6DB6D2492492DB6DB6DB6DB6DB6DB6DB6DB6DB6D924924936DB6D924936DB64926DB24936D926DB249B649B649B649B649B64DB26D936C";
defparam ram_block1a112.mem_init0 = "9B24D93649B26C9B26C9B26C9B364D9366C9B364C9B364C9B366CD93264C993266CD9B3264CD9B3266CC99B33664CC999332664CCD99933326664CCC99999333336666666CCCCCCCCC9999999999999999999999999999CCCCCCCCC66666673333399998CCCE6663333999CCC66633399CCC6633199CC6633198CE63319CC67319CC67318CE6319CE6318CE739CC6318C6318C6318C6318E739C6318E738C739C639C639C638C738E71CE39C718E39C71CE38E31C71C738E38E38E38E38E38E38E38F1C71C70E38E1C71E38F1C78E3C70E3C70E3C78F1C3870E1C3870E1E3C7870F1E1C3C387870F0F0E1E1E1E1E1E1E1E1E1E1E1F0F0F078783C3E1F0F0783C";

arriav_ram_block ram_block1a32(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a32_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a32.clk0_core_clock_enable = "ena0";
defparam ram_block1a32.clk0_input_clock_enable = "ena0";
defparam ram_block1a32.clk0_output_clock_enable = "ena0";
defparam ram_block1a32.data_interleave_offset_in_bits = 1;
defparam ram_block1a32.data_interleave_width_in_bits = 1;
defparam ram_block1a32.init_file = "DDS_48_v1_nco_ii_0_sin.hex";
defparam ram_block1a32.init_file_layout = "port_a";
defparam ram_block1a32.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_c8g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a32.operation_mode = "rom";
defparam ram_block1a32.port_a_address_clear = "none";
defparam ram_block1a32.port_a_address_width = 13;
defparam ram_block1a32.port_a_data_out_clear = "none";
defparam ram_block1a32.port_a_data_out_clock = "clock0";
defparam ram_block1a32.port_a_data_width = 1;
defparam ram_block1a32.port_a_first_address = 16384;
defparam ram_block1a32.port_a_first_bit_number = 0;
defparam ram_block1a32.port_a_last_address = 24575;
defparam ram_block1a32.port_a_logical_ram_depth = 65536;
defparam ram_block1a32.port_a_logical_ram_width = 16;
defparam ram_block1a32.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a32.ram_block_type = "auto";
defparam ram_block1a32.mem_init3 = "1E0F07C3E0F07C1F0F83E0F83E0F83E0F81F07C0F81F07E0FC0F81F81F03F03F03F03F81F81FC0FE07F01FC07E03FC07F01FE03FC03F807F803FC03FE01FF007FC00FF801FF801FFC00FFE003FFC003FFC001FFF0003FFF8000FFFF00003FFFF00000FFFFFE000000FFFFFFFE0000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000001FFFFFFF8000001FFFFF800007FFFE0000FFFF0001FFF8001FFF0007FF8007FF001FFC00FFC00FFC00FF803FE00FF007F807F807F807F00FE01FC07F01FC0FE03F01F80FC0FC07E07E0FC0FC0F81F83F07E0F81F07C1F83E0F83E0F87C1F0783E1F0783C1E0F0F87C3C1E1E0F0F0F0F8787878787";
defparam ram_block1a32.mem_init2 = "8F0F0F0E1E1E3C387870E1E3C7870E1C3871E3C78E1C78E1C70E3C71C38E3871C71C38E38E38E38E38E38E39C71C718E38C71CE38C718E31CE31C639CE31CE718C739CE318C6318C6318C6739CE6319CE6339CC67319CC673398CC6633198CCE67331998CCC666333319999CCCCCC6666666666333333333333326666666666CCCCCD9999B3336666CCC999332664CD99B3264CD993264C993264C99366C99366C9B264D9364D93649B26C93649B24DB26D924DB249B64926DB24926DB6D924924924DB6DB6DA492492492DB6DA4925B6D2496DA496D24B692DA4B692DA4B49692D25A5B4B4B49696969696969694B4B4A5A5AD2D694B5A52D694A5AD6B5A529";
defparam ram_block1a32.mem_init1 = "4A5294A56B5AD4A56B5A95AD4AD4A56A56AD4AD4A95AB52A54A952A54A952AD5AA55AA55AAD52A954AA552A955AA955AAB556AA9552AA9554AAA5554AAA95556AAAA55555AAAAA9555555AAAAAAAA95555555555555555AAAAAAAAAAD5555555555555554AAAAAAAAD555554AAAAAD55552AAA95554AAA9555AAA9556AAB554AA9552AB556AA552AB55AAD56A954AB54AB54A956AD52A54A952B56AD4A95A952B52B52B52B5A95AD4A56B5A94A5295AD6B5A5294A52D6B4A5AD296B4A5A52D2D6969694B4B4B4B4B4969696D2D25A5B49692D25B496D25B692DB492DB4925B6D24925B6DB6D249249249249249B6DB6D924936DB24936C926D924DB26D926C93";
defparam ram_block1a32.mem_init0 = "649B26C9B26C9B26C9B364D9B264C9B366CD9B3664C99B3266CC99B33666CCC9999333266664CCCCCC99999999999999999999999999CCCCCCE666673331999CCC66633199CCE673399CC673398CE6319CC6339CC6318CE739CE739CE318C739C631CE31CE31CE39C738E71C638E31C71C738E38E38E38E38E1C71C70E38E1C70E3C71E3870E3C78F1E3C78F1E1C3C7870F0E1E1E1E3C3C3C3C3C1E1E1E0F0F0787C3E1F0F87C1E0F83C1F07C1F07C1F03E0F81F03E07E0FC0FC0FC0FC0FC07E03F01FC07F01FC07F80FF00FF00FF007FC01FF007FE00FFE007FF001FFE001FFF0003FFF0000FFFF00001FFFFE000001FFFFFFF00000000003FFFFFFFFFFFFFF";

arriav_ram_block ram_block1a48(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a48_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a48.clk0_core_clock_enable = "ena0";
defparam ram_block1a48.clk0_input_clock_enable = "ena0";
defparam ram_block1a48.clk0_output_clock_enable = "ena0";
defparam ram_block1a48.data_interleave_offset_in_bits = 1;
defparam ram_block1a48.data_interleave_width_in_bits = 1;
defparam ram_block1a48.init_file = "DDS_48_v1_nco_ii_0_sin.hex";
defparam ram_block1a48.init_file_layout = "port_a";
defparam ram_block1a48.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_c8g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a48.operation_mode = "rom";
defparam ram_block1a48.port_a_address_clear = "none";
defparam ram_block1a48.port_a_address_width = 13;
defparam ram_block1a48.port_a_data_out_clear = "none";
defparam ram_block1a48.port_a_data_out_clock = "clock0";
defparam ram_block1a48.port_a_data_width = 1;
defparam ram_block1a48.port_a_first_address = 24576;
defparam ram_block1a48.port_a_first_bit_number = 0;
defparam ram_block1a48.port_a_last_address = 32767;
defparam ram_block1a48.port_a_logical_ram_depth = 65536;
defparam ram_block1a48.port_a_logical_ram_width = 16;
defparam ram_block1a48.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a48.ram_block_type = "auto";
defparam ram_block1a48.mem_init3 = "B56AD5AB56AD52A54A952A54A952A54A952A55AB56AD5AB56AD5AB56A952A54A952A54AB56AD5AB56AD5AA54A952A54AB56AD5AB54A952A54AB56AD5AA54A952AD5AB56A952A55AB56A952A55AB56A952A55AB54A952AD5AA54AB56A952AD5AA54AB56A952AD5AA55AB54AB56A956AD52AD5AA55AA54AB54AB56A956A956A956A956AD52AD52AD52A956A956A956A956A954AB54AB55AA55AAD52AD56A954AB54AA552AD56A954AA55AAD56A954AA552A954AB55AAD56AB552A954AA552A955AAD56AA552AB55AA954AAD56AA556AA552AB552AB552AB552AA556AA556AAD54AA955AAB556AA554AA9552AA554AA9556AAD55AAA554AAB554AAB554AAB554AAB";
defparam ram_block1a48.mem_init2 = "555AAA5552AAD556AAB555AAA9554AAAD556AAA5556AAAD554AAA9555AAAB5554AAA95556AAA95556AAAB5555AAAAD5554AAAAD5555AAAA955556AAAA955554AAAAA555556AAAAAD555552AAAAA9555555AAAAAAA55555552AAAAAAAD55555555AAAAAAAAAB55555555554AAAAAAAAAAAAA955555555555555555556AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAD5555555555555555556AAAAAAAAAAAAB55555555552AAAAAAAA955555556AAAAAAA5555554AAAAAA555555AAAAAB55555AAAAAD55552AAAA55556AAAA55552AAAD5556AAAD5552AAA5556AAA5556AAA5552AAB554AAA5552AAD552AAD55AAA554AA9552AA554AA955AA9";
defparam ram_block1a48.mem_init1 = "552AB552A955AA954AAD56AB55AA956AB55AAD56A954AB54AA55AA55AA55AA55AA54AB54A956AD52A54A956AD5AB56AD5AB56AD4A952B56AD4A95AB52A56A56AD4AD4AD5A95A95A95AD4AD4AD4A56A52B5295AD4AD6B5295AD4A5295AD6A5294A5295AD6B5AD6B5AD694A5294A5AD6B4A52D6B4A52D6B4A5AD296B4A5A52D696B4B5A5AD2D29696B4B4B4A5A5A5A5A5A5A5A5A5A5A5A5A5A5B4B4B4B69696D2D25A5B4B696D2DA5B49692DA5B496D25B496D25B492DA496D24B6D25B6D24B6D2496DB4925B6DA4924B6DB6D2492492DB6DB6DB6DB6DB6DB6DB6DB6DB6D924924936DB6D924936DB64926DB24936D926DB249B649B649B649B649B64DB26D936C";
defparam ram_block1a48.mem_init0 = "9B24D93649B26C9B26C9B26C9B364D9366C9B364C9B364C9B366CD93264C993266CD9B3264CD9B3266CC99B33664CC999332664CCD99933326664CCC99999333336666666CCCCCCCCC9999999999999999999999999999CCCCCCCCC66666673333399998CCCE6663333999CCC66633399CCC6633199CC6633198CE63319CC67319CC67318CE6319CE6318CE739CC6318C6318C6318C6318E739C6318E738C739C639C639C638C738E71CE39C718E39C71CE38E31C71C738E38E38E38E38E38E38E38F1C71C70E38E1C71E38F1C78E3C70E3C70E3C78F1C3870E1C3870E1E3C7870F1E1C3C387870F0F0E1E1E1E1E1E1E1E1E1E1E1F0F0F078783C3E1F0F0783C";

arriav_ram_block ram_block1a0(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a0_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.clk0_input_clock_enable = "ena0";
defparam ram_block1a0.clk0_output_clock_enable = "ena0";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.init_file = "DDS_48_v1_nco_ii_0_sin.hex";
defparam ram_block1a0.init_file_layout = "port_a";
defparam ram_block1a0.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_c8g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.operation_mode = "rom";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 13;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "clock0";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 8191;
defparam ram_block1a0.port_a_logical_ram_depth = 65536;
defparam ram_block1a0.port_a_logical_ram_width = 16;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.ram_block_type = "auto";
defparam ram_block1a0.mem_init3 = "783C1E1F0F8783C3C1E1E1F0F0F0F0F0F0F0F0F0F0F0E1E1E1C3C387870F1E1C3C78F0E1C3870E1C3871E3C78E1C78E1C78E3C71E38F1C70E38E1C71C71E38E38E38E38E38E38E38E39C71C718E38E71C738E31C738E71CE39C638C738C738C739C639CE318C739CE318C6318C6318C6318C6739CE6318CE7318CE6319CC67319CC673198CE633198CC6733198CC66733998CCC6673339998CCCE6663333399999CCCCCCC6666666673333333333333333333333333332666666666CCCCCCD99999333326664CCC99993336664CC999332664CD99B3266CC99B3664C99B366CC993264C99366CD9B264D9B264D9B26CD9364D9B26C9B26C9B26C9B24D93649B2";
defparam ram_block1a0.mem_init2 = "6D936C9B64DB24DB24DB24DB24DB249B6C936D9249B6C924DB6D924936DB6D924924936DB6DB6DB6DB6DB6DB6DB6DB6DB692492496DB6DA4924B6DB4925B6D2496DA496DB496DA496D24B6925B496D25B496D25B4B692D25B4B696D2DA5B4B49696D2D2DA5A5A5B4B4B4B4B4B4B4B4B4B4B4B4B4B4A5A5A5AD2D29696B4B5A5AD2D694B4A5AD296B4A5AD694A5AD694A5AD6B4A5294A52D6B5AD6B5AD6B5294A5294AD6B5294A56B5295AD6A56B5295A94AD4A56A56A56B52B52B52B56A56A56AD4AD4A95AB52A56AD5A952A56AD5AB56AD5AB56AD52A54A956AD52A55AA54AB54AB54AB54AB54AA55AA552AD56AB55AAD52AB55AAD56AA552AB552A955AA955";
defparam ram_block1a0.mem_init1 = "2AB552AA554AA9552AA554AAB556AA9556AA9554AAA555AAA9554AAAD554AAAD554AAA95556AAAD5556AAA95554AAAAD5554AAAA955556AAAAB55555AAAAAB555554AAAAAA5555554AAAAAAAD55555552AAAAAAAA95555555555AAAAAAAAAAAAAD5555555555555555556AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAD55555555555555555552AAAAAAAAAAAAA55555555555AAAAAAAAAB555555556AAAAAAA95555554AAAAAAB5555552AAAAA9555556AAAAAD55554AAAAA555552AAAAD55552AAAB55556AAAA55556AAAB5555AAAAD5552AAAD5552AAA5555AAAB5552AAA5556AAAD554AAAD556AAA5552AAB555AAAD556AA9554AAB555";
defparam ram_block1a0.mem_init0 = "AAA555AAA555AAA555AAA554AAB556AAD552AA554AA9552AA554AAD55AAB552AA556AAD54AAD54AA955AA955AA955AA954AAD54AAD56AA552AB55AA954AAD56AB552A954AA552A955AAD56AB55AA552A954AA552AD56AB54AA552AD56A954AA55AA552AD56A956AB54AB55AA55AA552AD52AD52AD52AD52A956A956A956AD52AD52AD52AD52AD5AA55AA54AB54AB56A956AD52AD5AA55AB54AB56A952AD5AA54AB56A952AD5AA54AB56A952A55AB54A952AD5AB54A952AD5AB54A952AD5AB56A952A54AB56AD5AA54A952A55AB56AD5AA54A952A54AB56AD5AB56AD5AA54A952A54A952AD5AB56AD5AB56AD5AB54A952A54A952A54A952A54A956AD5AB56AD5A";

arriav_ram_block ram_block1a16(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a16_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a16.clk0_core_clock_enable = "ena0";
defparam ram_block1a16.clk0_input_clock_enable = "ena0";
defparam ram_block1a16.clk0_output_clock_enable = "ena0";
defparam ram_block1a16.data_interleave_offset_in_bits = 1;
defparam ram_block1a16.data_interleave_width_in_bits = 1;
defparam ram_block1a16.init_file = "DDS_48_v1_nco_ii_0_sin.hex";
defparam ram_block1a16.init_file_layout = "port_a";
defparam ram_block1a16.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_c8g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a16.operation_mode = "rom";
defparam ram_block1a16.port_a_address_clear = "none";
defparam ram_block1a16.port_a_address_width = 13;
defparam ram_block1a16.port_a_data_out_clear = "none";
defparam ram_block1a16.port_a_data_out_clock = "clock0";
defparam ram_block1a16.port_a_data_width = 1;
defparam ram_block1a16.port_a_first_address = 8192;
defparam ram_block1a16.port_a_first_bit_number = 0;
defparam ram_block1a16.port_a_last_address = 16383;
defparam ram_block1a16.port_a_logical_ram_depth = 65536;
defparam ram_block1a16.port_a_logical_ram_width = 16;
defparam ram_block1a16.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a16.ram_block_type = "auto";
defparam ram_block1a16.mem_init3 = "FFFFFFFFFFFFFF80000000001FFFFFFF000000FFFFF00001FFFE0001FFF8001FFF000FFF001FFC00FFE00FFC01FF007FC01FE01FE01FE03FC07F01FC07F01F80FC07E07E07E07E07E0FC0F81F03E0F81F07C1F07C1F0783E0F07C3E1F0F87C3C1E1E0F0F0F07878787878F0F0F0E1E1C3C7870F1E3C78F1E3C78E1C38F1C78E1C70E38E1C71C70E38E38E38E38E39C71C718E38C71CE39C738E718E718E718C739C6318E739CE739CE6318C67398C67318CE63399CC673399CCE6733198CCC6673331999CCCCCE666667333333333333333333333333326666664CCCC99993332666CCD99B3266CC99B3264CD9B366CD9B264C9B364D9B26C9B26C9B26C9B24D";
defparam ram_block1a16.mem_init2 = "926C936C9B64936C926D9249B6D924936DB6DB2492492492492496DB6DB492496DB4925B6925B692DB496D25B49692D25B4B49696D2D2D25A5A5A5A5A52D2D2D69694B4A5AD296B4A5AD694A5294B5AD6B5294A52B5AD4A56B52B5A95A95A95A952B52A56AD5A952A54A956AD52A55AA55AA552AD56AB55AA954AAD55AA9552AA555AAAD552AAB5552AAA55552AAA955556AAAAA5555556AAAAAAAA55555555555555556AAAAAAAAAB55555555555555552AAAAAAAB5555552AAAAB55554AAAAD5552AAA5554AAA5552AA9552AAD55AAB552AB552A954AA552A956AB54AB54AB56A952A54A952A54A95AB52A56A56AD4AD4A56A56B52B5AD4A56B5AD4A5294A5";
defparam ram_block1a16.mem_init1 = "294B5AD6B4A52D694B5A52D696B4B4A5A5A52D2D2D2D2D2D2D25A5A5B4B49692D25A4B692DA4B692DA496D24B6D2496DB4924B6DB6924924924B6DB6DB64924924936DB6C9249B6C924DB249B64936C9B649B24D926C9B24D9364D9364C9B26CD9326CD93264C993264C9933664C99B33664CC999332666CCCD999B3333666666CCCCCCCCCC99999999999998CCCCCCCCCC666667333319998CCC666333199CCE6633198CC663399CC67319CC67398CE7318CE739CC6318C6318C6318E739C631CE718E738C718E718E31C638E71C638E31C71C738E38E38E38E38E38E3871C71C38E3871C78E1C70E3C70E3C78F1C3870E1C3C78F0E1C3C3878F0F0E1E1E1E3";
defparam ram_block1a16.mem_init0 = "C3C3C3C3C3E1E1E1E0F0F0787C3E1E0F0783C1F0F83C1F07C3E0F83E0F83F07C1F03E0FC1F83F03E07E07E0FC0FC07E07E03F01F80FE07F01FC07F00FE01FC03FC03FC03FC01FE00FF803FE007FE007FE007FF001FFC003FFC001FFF0003FFF0001FFFE0000FFFFC00003FFFFF0000003FFFFFFF00000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000FFFFFFFE000000FFFFFE00001FFFF80001FFFE0003FFF8001FFF0007FF8007FF800FFE007FF003FF003FE007FC01FF00FF807F803FC03F807F80FF01FC07F80FC07F01FC0FE07F03F03F81F81F81F81F03F03E07E0FC1F03E07C1F03E0F83E0F83E0F83E1F07C1E0F87C1E0F0";

arriav_ram_block ram_block1a65(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a65_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a65.clk0_core_clock_enable = "ena0";
defparam ram_block1a65.clk0_input_clock_enable = "ena0";
defparam ram_block1a65.clk0_output_clock_enable = "ena0";
defparam ram_block1a65.data_interleave_offset_in_bits = 1;
defparam ram_block1a65.data_interleave_width_in_bits = 1;
defparam ram_block1a65.init_file = "DDS_48_v1_nco_ii_0_sin.hex";
defparam ram_block1a65.init_file_layout = "port_a";
defparam ram_block1a65.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_c8g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a65.operation_mode = "rom";
defparam ram_block1a65.port_a_address_clear = "none";
defparam ram_block1a65.port_a_address_width = 13;
defparam ram_block1a65.port_a_data_out_clear = "none";
defparam ram_block1a65.port_a_data_out_clock = "clock0";
defparam ram_block1a65.port_a_data_width = 1;
defparam ram_block1a65.port_a_first_address = 32768;
defparam ram_block1a65.port_a_first_bit_number = 1;
defparam ram_block1a65.port_a_last_address = 40959;
defparam ram_block1a65.port_a_logical_ram_depth = 65536;
defparam ram_block1a65.port_a_logical_ram_width = 16;
defparam ram_block1a65.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a65.ram_block_type = "auto";
defparam ram_block1a65.mem_init3 = "52A954AA552AD56A954AB55AA55AA55AA55AA55AA55AB54AB56A952AD5AA54A956AD5AB56AD5AB56AD5AB56AD4A952B56AD4A95AB52A56A54AD4A95A95AB52B52B52B52B52B52B52B5295A95AD4AD4A56A52B5A95AD4A56B5294AD6A5295AD6A5294AD6B5AD6A5294A5294A5294A5294A5294A5294B5AD6B5A5294B5AD694A5AD694A5AD294B5A52D694A5A52D694B5A52D29694B5A5AD2D29694B4B5A5A52D2D296969694B4B4B4B5A5A5A5A5A5A5A5A5A5A5A5A5A5A4B4B4B4B4B6969696D2D2DA5A5B4B49696D2D25A5B4B696D2DA5B4B696D2DA4B496D2DA4B692D25B496D25B496D25B496D24B692DB496D24B6925B692DB492DB492DB492DB6925B6D24";
defparam ram_block1a65.mem_init2 = "B6DA492DB692496DB692496DB692492DB6DA492492DB6DB6924924925B6DB6DB6DB6DA4924924924924924924924924924DB6DB6DB6DB6C924924926DB6DB64924936DB6D924936DB64924DB6D9249B6D9249B6D924DB64926DB249B6C926D924DB649B6C936C926D926D926D926D926D926D926D936C936C9B64DB24D926C93649B26D936C9B24D936C9B26C9364D936C9B26C9B26C9B64D9364D9364D9B26C9B26C9B264D9364D9B26C9B364D9B26CD9366C9B364C9B264D9B264D9B364C9B366C99326CD9B364C993264C9B366CD9B366CD9B3664C993264C99B366CC993266CD993266CD993366CC99B3664CD9933664CD9933664CC99B32664CD9933266";
defparam ram_block1a65.mem_init1 = "4CD99B33666CCD99B33666CCD99B332664CCD999333666CCCD9993336666CCC999933326664CCC9999B33326666CCCC999993333266664CCCCD99999333332666666CCCCCC99999993333333666666664CCCCCCCCD9999999999333333333333366666666666666666664CCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCE66666666666666666663333333333333399999999999CCCCCCCCCC666666667333333319999998CCCCCCC6666663333331999998CCCCCE666673333399999CCCCCE66663333399998CCCC6666733339999CCCCE66633331999CCCC66663333999CCCC66673331998CCCE667333999CCCC6663331998CCE667333999";
defparam ram_block1a65.mem_init0 = "CCC666333999CCC666333998CCC66733199CCC66733199CCC66733199CCC66333998CCE6733198CCE6633199CCE6633198CCE6733198CC6633399CCE6733198CC6633198CC6633199CCE673399CC6633198CC6633198CC673399CCE673198CC663399CCE673198CC673399CC663399CCE63319CCE63319CCE673198CE67319CCE63319CCE63319CC663398CC673398CE67319CCE63399CC673398CE63319CC673398CE63319CC673398CE63399CC67319CCE63398CE63319CC67319CCE63398CE63398CC67319CC67319CC663398CE63398CE63398CC67319CC67319CC67319CC67319CCE63398CE63398CE63398CE63398CE63398CE63398CE67319CC67319C";

arriav_ram_block ram_block1a81(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a81_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a81.clk0_core_clock_enable = "ena0";
defparam ram_block1a81.clk0_input_clock_enable = "ena0";
defparam ram_block1a81.clk0_output_clock_enable = "ena0";
defparam ram_block1a81.data_interleave_offset_in_bits = 1;
defparam ram_block1a81.data_interleave_width_in_bits = 1;
defparam ram_block1a81.init_file = "DDS_48_v1_nco_ii_0_sin.hex";
defparam ram_block1a81.init_file_layout = "port_a";
defparam ram_block1a81.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_c8g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a81.operation_mode = "rom";
defparam ram_block1a81.port_a_address_clear = "none";
defparam ram_block1a81.port_a_address_width = 13;
defparam ram_block1a81.port_a_data_out_clear = "none";
defparam ram_block1a81.port_a_data_out_clock = "clock0";
defparam ram_block1a81.port_a_data_width = 1;
defparam ram_block1a81.port_a_first_address = 40960;
defparam ram_block1a81.port_a_first_bit_number = 1;
defparam ram_block1a81.port_a_last_address = 49151;
defparam ram_block1a81.port_a_logical_ram_depth = 65536;
defparam ram_block1a81.port_a_logical_ram_width = 16;
defparam ram_block1a81.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a81.ram_block_type = "auto";
defparam ram_block1a81.mem_init3 = "000000000000007FFFFFFFFFFFFFFFFF00000000000FFFFFFFFE00000007FFFFFF000000FFFFFC00001FFFFC0000FFFFC0001FFFE0001FFFC000FFFC000FFF8003FFE001FFE001FFE003FF800FFE007FF003FF003FF007FE00FFC01FF007FC03FE01FF00FF007F807F807F00FF01FE03FC07F00FE03F80FE03F81FC07F03F81FC0FE07E03F03F01F81F81F81F81F83F03F07E07C0FC1F83F07E0F81F07E0F83F07C1F07E0F83E0F83E1F07C1F0783E0F07C1E0F87C3E0F0783C1E0F0F87C3C1E0F0F0787C3C3C1E1E1E0F0F0F0F0F0F0F0F0F0F0F0F0F1E1E1E1C3C3C7878F0F1E1E3C3878F1E1C3878F1E3C3870E1C3871E3C78F1C3871E3871E3871E3871C3";
defparam ram_block1a81.mem_init2 = "8E1C70E3871C70E38E1C71C78E38E38F1C71C71C71C71C71C71C71C71C738E38E38C71C718E38E71C738E31C738E71CE38C738E71CE31CE39C639C639CE31CE318E738C639CE718C639CE739CE738C6318CE739CE739CC6318CE7398C67398C67318CE6319CC67319CC67319CCE63399CC663319CCE6733998CC66333998CCE66333999CCCE6673331999CCCCE66673333199999CCCCCCE666666663333333333333333199999999993333333333333333666666666CCCCCC9999993333266664CCC99993332666CCC999B336664CC99933666CC99B3266CC99B3266CD993266CD9B366CD9B366CD9B366C99326CD9B264D9326CD9366C9B26CD9364D9364D93";
defparam ram_block1a81.mem_init1 = "64D9364D926C9B24D936C9B24D926D936C93649B649B649B64936C936D924DB64936D9249B6D9249B6DB24926DB6DB24924926DB6DB6DB6DB6D92492492DB6DB6DB6DB6DA4924925B6DB692492DB6DA492DB6924B6DA496DB492DB492DA496DA4B6925B496D25B496D25B496D2DA4B696D2DA5B4B696D2DA5A4B4B69696D2D2D25A5A5A5A5A4B4B4B4B4B4B4A5A5A5A5A5AD2D2D29696B4B4A5A52D29694B4A5AD296B4A5AD296B4A52D6B4A52D6B5A5294A5AD6B5AD6B5AD6B5AD6B5AD6B5294A52B5AD6A52B5AD4A56B5295AD4AD6A56B52B5295A95A95A95A95A95A952B52B56A56AD4AD5AB52A56AD5A952A54A952A54A952A55AB56A952A55AA54AB54A9";
defparam ram_block1a81.mem_init0 = "56A956A956AB54AB55AA552AD56AB55AAD56AB55AA954AAD56AA556AA556AAD54AA955AAB556AA9552AAD55AAA5552AAD556AAB555AAAD554AAAD555AAAB5556AAA95556AAAB5555AAAA955552AAAAD55552AAAAB555556AAAAAB5555556AAAAAAB55555555AAAAAAAAA9555555555556AAAAAAAAAAAAAAAAAD555555555555555555555555555555555555555554AAAAAAAAAAAAAAAAAB555555555554AAAAAAAAAD55555554AAAAAAAD555555AAAAAAD555552AAAAB55555AAAAA55554AAAA95555AAAAD5552AAA95552AAAD555AAA95552AA9555AAA9554AAA555AAAD552AAD552AA555AAB554AA955AAB556AA554AAD54AAD54AAD54AA556AB552A954AA5";

arriav_ram_block ram_block1a97(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a97_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a97.clk0_core_clock_enable = "ena0";
defparam ram_block1a97.clk0_input_clock_enable = "ena0";
defparam ram_block1a97.clk0_output_clock_enable = "ena0";
defparam ram_block1a97.data_interleave_offset_in_bits = 1;
defparam ram_block1a97.data_interleave_width_in_bits = 1;
defparam ram_block1a97.init_file = "DDS_48_v1_nco_ii_0_sin.hex";
defparam ram_block1a97.init_file_layout = "port_a";
defparam ram_block1a97.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_c8g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a97.operation_mode = "rom";
defparam ram_block1a97.port_a_address_clear = "none";
defparam ram_block1a97.port_a_address_width = 13;
defparam ram_block1a97.port_a_data_out_clear = "none";
defparam ram_block1a97.port_a_data_out_clock = "clock0";
defparam ram_block1a97.port_a_data_width = 1;
defparam ram_block1a97.port_a_first_address = 49152;
defparam ram_block1a97.port_a_first_bit_number = 1;
defparam ram_block1a97.port_a_last_address = 57343;
defparam ram_block1a97.port_a_logical_ram_depth = 65536;
defparam ram_block1a97.port_a_logical_ram_width = 16;
defparam ram_block1a97.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a97.ram_block_type = "auto";
defparam ram_block1a97.mem_init3 = "4AA552A955AAD54AA556AA556AA556AA554AAD55AAB552AA555AAB554AA9556AA9556AAB554AAA5552AAB5552AA95552AAB5556AAA95552AAA95556AAAB55552AAAA55554AAAAB55555AAAAA9555556AAAAAB5555556AAAAAAA555555556AAAAAAAAA555555555555AAAAAAAAAAAAAAAAAA5555555555555555555555555555555555555555556AAAAAAAAAAAAAAAAAD555555555552AAAAAAAAB55555555AAAAAAAD555555AAAAAAD55555AAAAA955556AAAA955552AAAB5555AAAAD5552AAAD555AAAB5556AAA5556AAB555AAAD556AA9554AAB556AA9552AAD55AAB552AA556AAD54AAD54AAD56AA552AB55AAD56AB55AAD56A954AB55AA55AAD52AD52AD5";
defparam ram_block1a97.mem_init2 = "2A55AA54AB54A952AD5AB54A952A54A952A54A952B56AD4A95AB56A56AD4AD5A95A952B52B52B52B52B52B5295A95AD4AD6A56B5295AD4A56B5A94AD6B5A94A5295AD6B5AD6B5AD6B5AD6B5AD6B4A5294B5AD694A5AD694A5AD296B4A5AD296B4A5A52D29694B4A5A5AD2D2969696B4B4B4B4B4A5A5A5A5A5A5A4B4B4B4B4B4969696D2D2DA5A4B4B696D2DA5B4B696D2DA4B696D25B496D25B496D25B492DA4B6D24B6925B6925B6D24B6DA492DB6924B6DB692492DB6DB4924924B6DB6DB6DB6DB6924924936DB6DB6DB6DB6C9249249B6DB6C9249B6DB24936DB24936D924DB64936D926D924DB24DB24DB24D926D936C93649B26D93649B26C9364D9364D";
defparam ram_block1a97.mem_init1 = "9364D9364D9366C9B26CD9366C99364C9B366C99326CD9B366CD9B366CD9B366CC993366CC99B3266CC99B3266CCD99332664CCD99B332666CCC999933326664CCCC99999333332666666CCCCCCCCD9999999999999999333333333319999999999999998CCCCCCCCE6666673333319999CCCCE66673331999CCCE667333998CCE66333998CC6633399CCE673198CC673398CE67319CC67319CC67318CE6319CC6339CC6339CE6318C6739CE739CE6318C639CE739CE738C631CE738C639CE318E718E738C738C738E718E71CE39C638E71CE39C718E39C71CE38E31C71C638E38E39C71C71C71C71C71C71C71C71C71E38E38E3C71C70E38E1C71C38E1C70E3";
defparam ram_block1a97.mem_init0 = "871C38F1C38F1C38F1C3871E3C78F1C3870E1C3878F1E3C3870F1E3C3878F0F1E1E3C3C787870F0F0F1E1E1E1E1E1E1E1E1E1E1E1E1E0F0F0F078787C3C1E1E0F0787C3E1E0F0783C1E0F87C3E0F07C1E0F83C1F07C1F0F83E0F83E0FC1F07C1F83E0FC1F03E0FC1F83F07E07C0FC1F81F83F03F03F03F03F01F81F80FC0FE07F03F81FC07F03F80FE03F80FE01FC07F80FF01FE01FC03FC03FC01FE01FF00FF807FC01FF007FE00FFC01FF801FF801FFC00FFE003FF800FFF000FFF000FFF8003FFE0007FFE0007FFF0000FFFF00007FFFE00007FFFF000007FFFFE000001FFFFFFC0000000FFFFFFFFE00000000001FFFFFFFFFFFFFFFFFC00000000000000";

arriav_ram_block ram_block1a113(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a113_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a113.clk0_core_clock_enable = "ena0";
defparam ram_block1a113.clk0_input_clock_enable = "ena0";
defparam ram_block1a113.clk0_output_clock_enable = "ena0";
defparam ram_block1a113.data_interleave_offset_in_bits = 1;
defparam ram_block1a113.data_interleave_width_in_bits = 1;
defparam ram_block1a113.init_file = "DDS_48_v1_nco_ii_0_sin.hex";
defparam ram_block1a113.init_file_layout = "port_a";
defparam ram_block1a113.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_c8g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a113.operation_mode = "rom";
defparam ram_block1a113.port_a_address_clear = "none";
defparam ram_block1a113.port_a_address_width = 13;
defparam ram_block1a113.port_a_data_out_clear = "none";
defparam ram_block1a113.port_a_data_out_clock = "clock0";
defparam ram_block1a113.port_a_data_width = 1;
defparam ram_block1a113.port_a_first_address = 57344;
defparam ram_block1a113.port_a_first_bit_number = 1;
defparam ram_block1a113.port_a_last_address = 65535;
defparam ram_block1a113.port_a_logical_ram_depth = 65536;
defparam ram_block1a113.port_a_logical_ram_width = 16;
defparam ram_block1a113.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a113.ram_block_type = "auto";
defparam ram_block1a113.mem_init3 = "7319CC67319CCE63398CE63398CE63398CE63398CE63398CE63398CE67319CC67319CC67319CC67319CC663398CE63398CE63398CC67319CC67319CC663398CE63398CE67319CC673198CE63398CE67319CC673398CE63399CC673198CE63399CC673198CE63399CC673398CE67319CCE63399CC663398CC673198CE673198CE67319CCE63319CCE673198CE673198CE673398CC673399CC663319CCE673398CC663319CCE673399CC6633198CC6633198CC673399CCE6733198CC6633198CC6633199CCE6733998CC6633199CCE6633198CCE6733198CCE6633199CCE66333998CC66733199CCC66733199CCC66733199CCC666333998CCC667333998CCC667";
defparam ram_block1a113.mem_init2 = "333999CCCE663331998CCC6667333999CCCE6663331999CCCC66673339998CCCC666733319998CCCE666733339999CCCCC66663333399998CCCCE666673333399999CCCCCE666663333331999998CCCCCC6666666333333319999999CCCCCCCCC66666666673333333333399999999999998CCCCCCCCCCCCCCCCCCCE6666666666666666666666666666666666666666666666666664CCCCCCCCCCCCCCCCCCD999999999999933333333336666666664CCCCCCCD99999993333332666666CCCCCC99999933333666664CCCC99999333326666CCCC9999B33326664CCC99993332666CCCD9993336666CCD9993336664CC999B33666CCD99B33666CCD99B33664";
defparam ram_block1a113.mem_init1 = "CC99933664CC99B32664CD9933664CD9933664CD9B3266CD993366CC993366CC993266CD9B3264C993264CD9B366CD9B366CD9B264C993264D9B366C99326CD9B264D9B364C9B364C9B264D9B26CD9366C9B364D9B26C9B364D9364C9B26C9B26C9B364D9364D9364DB26C9B26C9B26D9364D926C9B26D93649B26D936C9B24D926C93649B64DB26D926D936C936C936C936C936C936C936C926D926DB24DB64936C926DB249B6C924DB64936DB24936DB24936DB64924DB6D924936DB6D924924DB6DB6C924924926DB6DB6DB6DB64924924924924924924924924924B6DB6DB6DB6DB492492492DB6DB6924924B6DB692492DB6D2492DB6D2492DB6924B6DA";
defparam ram_block1a113.mem_init0 = "496DB492DB6925B6925B6925B692DB492DA496D25B692DA496D25B496D25B496D25B49692DA4B696D25A4B696D2DA5B4B696D2DA5B4B49696D2D25A5B4B4B69696D2D2D2DA5A5A5A5A4B4B4B4B4B4B4B4B4B4B4B4B4B4B5A5A5A5A52D2D2D2969694B4B5A5A52D29696B4B5A52D29694B5A52D694B4A52D694B5A5296B4A52D6B4A52D6B5A5294B5AD6B5A5294A5294A5294A5294A5294A5294AD6B5AD6A5294AD6B5294AD6A5295AD4A56B52B5A94AD4A56A56B52B5295A95A95A95A95A95A95A95AB52B52A56A54AD4A95AB52A56AD5A952A56AD5AB56AD5AB56AD5AB56AD52A54AB56A952AD5AA55AB54AB54AB54AB54AB54AB55AA552AD56A954AA552A95";

arriav_ram_block ram_block1a33(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a33_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a33.clk0_core_clock_enable = "ena0";
defparam ram_block1a33.clk0_input_clock_enable = "ena0";
defparam ram_block1a33.clk0_output_clock_enable = "ena0";
defparam ram_block1a33.data_interleave_offset_in_bits = 1;
defparam ram_block1a33.data_interleave_width_in_bits = 1;
defparam ram_block1a33.init_file = "DDS_48_v1_nco_ii_0_sin.hex";
defparam ram_block1a33.init_file_layout = "port_a";
defparam ram_block1a33.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_c8g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a33.operation_mode = "rom";
defparam ram_block1a33.port_a_address_clear = "none";
defparam ram_block1a33.port_a_address_width = 13;
defparam ram_block1a33.port_a_data_out_clear = "none";
defparam ram_block1a33.port_a_data_out_clock = "clock0";
defparam ram_block1a33.port_a_data_width = 1;
defparam ram_block1a33.port_a_first_address = 16384;
defparam ram_block1a33.port_a_first_bit_number = 1;
defparam ram_block1a33.port_a_last_address = 24575;
defparam ram_block1a33.port_a_logical_ram_depth = 65536;
defparam ram_block1a33.port_a_logical_ram_width = 16;
defparam ram_block1a33.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a33.ram_block_type = "auto";
defparam ram_block1a33.mem_init3 = "54AA556AB55AA955AAD54AAD54AAD54AAD55AA9552AA554AA9552AAD55AAA555AAA5552AAD556AAB555AAA9554AAA9555AAAB5556AAAD5552AAA95554AAAA55556AAAAD55552AAAA955554AAAAA9555556AAAAAA55555552AAAAAAA555555555AAAAAAAAAAB55555555555554AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAB55555555555554AAAAAAAAAAD55555555AAAAAAAB5555554AAAAAAD555552AAAAB55555AAAAA55555AAAA95555AAAAD5552AAAD5552AAA5554AAAD554AAA5556AAB555AAA5552AAD55AAA555AAB556AAD55AAB552AB556AA556AA552AB552A954AAD56AB55AA552A954AB55AA55AA552AD52AD52";
defparam ram_block1a33.mem_init2 = "A55AA55AB54A956AD52A54A952AD5AB56AD4A952A54AD5AB52A56AD4A95A952B52B56A56A56A56A56A56A56B52B52B5A95AD4A56A52B5A94A56B5294A56B5AD4A5294A56B5AD6B5AD6B5AD294A5294B5AD694A52D6B4A52D694A5AD296B4A5A52D694B4A5A52D29696B4B4B5A5A5AD2D2D2D2D296969696969696D2D2D2D2D25A5A5B4B4B69692D2DA5A4B49692D25B4B696D25B4B692DA4B692DA4B6D25B492DA496D24B6D24B6D2496DA492DB692496DB492496DB6D2492496DB6DB6DB49249249249249249249249249B6DB6DB6C924924DB6DB24926DB64926DB64926DB249B6C936D926DB24DB24DB24DB24D926D936C9B64DB26C9364DB26C9B26C9364";
defparam ram_block1a33.mem_init1 = "D9364D9326C9B26CD9364C9B264D9326CD9B264D9B366C993264C993264C99B366CC9933664C99B3266CC99B33664CC999332664CC999B332666CCCD999B33326666CCCCC99999B333333666666664CCCCCCCCCCCCCCCC9999999999CCCCCCCCCCCCCCCCC66666666333333399999CCCCCE666733339998CCC6667331998CCC66733198CCE6633198CC6633198CC673398CC67319CCE63398CE7319CC67398CE7318CE7318C6739CC6318C6739CE739CE739CE739CE318C639CE718C639CE31CE718E738C738C738C718E71CE31C638C718E31C738E31C718E38C71C738E38E31C71C71C71CE38E38E38E38E3871C71C71C70E38E38F1C71E38E3C71E38E1C70";
defparam ram_block1a33.mem_init0 = "E3871E3871E3871E3870E3C78E1C3870E1C3870E1C3878F1E1C3878F0E1E3C387870F0E1E1E3C3C3C387878787878787878787878787C3C3C3E1E1E0F0F0787C3C1E1F0F87C3E1F0F87C3E0F0783E1F07C3E0F83C1F07C1F07C1F07C1F07C0F83E0FC1F03E0FC1F83F07E0FC1F81F03F03F07E07E07E07E07E03F03F01F81FC0FE03F01F80FE03F80FE03F80FE03FC07F00FE01FE01FC03FC03FC01FE01FF00FF803FE00FF803FE007FC00FFC00FFC00FFE007FF001FFE003FFC003FFC003FFE000FFFC000FFFC0007FFF0000FFFF00003FFFF00001FFFFE00000FFFFFE000000FFFFFFF00000000FFFFFFFFFE0000000000000FFFFFFFFFFFFFFFFFFFFFFFFF";

arriav_ram_block ram_block1a49(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a49_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a49.clk0_core_clock_enable = "ena0";
defparam ram_block1a49.clk0_input_clock_enable = "ena0";
defparam ram_block1a49.clk0_output_clock_enable = "ena0";
defparam ram_block1a49.data_interleave_offset_in_bits = 1;
defparam ram_block1a49.data_interleave_width_in_bits = 1;
defparam ram_block1a49.init_file = "DDS_48_v1_nco_ii_0_sin.hex";
defparam ram_block1a49.init_file_layout = "port_a";
defparam ram_block1a49.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_c8g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a49.operation_mode = "rom";
defparam ram_block1a49.port_a_address_clear = "none";
defparam ram_block1a49.port_a_address_width = 13;
defparam ram_block1a49.port_a_data_out_clear = "none";
defparam ram_block1a49.port_a_data_out_clock = "clock0";
defparam ram_block1a49.port_a_data_width = 1;
defparam ram_block1a49.port_a_first_address = 24576;
defparam ram_block1a49.port_a_first_bit_number = 1;
defparam ram_block1a49.port_a_last_address = 32767;
defparam ram_block1a49.port_a_logical_ram_depth = 65536;
defparam ram_block1a49.port_a_logical_ram_width = 16;
defparam ram_block1a49.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a49.ram_block_type = "auto";
defparam ram_block1a49.mem_init3 = "C67319CC67319CC67319CC67319CC67319CC663398CE63398CE63398CE63398CE63398CC67319CC67319CC67319CC673398CE63398CE63398CC67319CC67319CCE63398CE63399CC67319CC663398CE63399CC67319CCE63398CC67319CCE63398CC67319CCE63399CC673398CE67319CCE63399CC673398CC673198CE673198CE67319CCE63319CCE673198CE673198CE673398CC663399CCE633198CE673398CC6633198CE673399CCE673198CC6633198CC6633198CC6633198CC6633199CCE673399CCC6633198CCE6733998CC6633399CCC6633399CCC66733998CCE6733199CCC66733998CCE66333998CCE66733199CCC667333998CCC667333998CCC";
defparam ram_block1a49.mem_init2 = "666333999CCCE667333999CCCE6673331998CCC66673331998CCCE66633339998CCCE666733319998CCCC6666333319998CCCCE66663333199998CCCCE6666733333999998CCCCCE666663333331999999CCCCCCC666666633333333199999999CCCCCCCCCC666666666673333333333333199999999999999999998CCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCC9999999999999999999B333333333333266666666664CCCCCCCCD9999999B33333336666666CCCCCC99999933333266666CCCCC99999B333366664CCCC9999B33366664CCC9999B3336664CCC999B3336664CCD9993336664CC999B33666CCC999332664CC99933266CCD";
defparam ram_block1a49.mem_init1 = "99B32664CD9933266CC99B3266CCD9B3266CC99B3266CD993366CC993366CC993366CD993264C99B366CD9B366CD9B366CD9B366CD9B264C99326CD9B364C9B366C99366CD9326CD9366C99366C9B364D9B26C99364D9B26C99364D9364C9B26C9B26C9B26C9B26C9B26C9B26C9364D93649B26C9B64D936C9B24D936C9B64DB26D936C9B64DB24D926D936C936C936C936C936C936C936C926D926DB24DB649B6C926DB249B6C926DB24936D9249B6D9249B6D924936DB649249B6DB649249B6DB6D924924936DB6DB6DB64924924924924924924924924924924924924924925B6DB6DB6DA4924924B6DB6DA4924B6DB6D2492DB6D2492DB6D2496DB4925B6";
defparam ram_block1a49.mem_init0 = "D2496DA492DB492DB492DB492DA496DA4B6D25B692DA496D25B496DA4B692DA4B496D25B49692DA4B496D2DA5B49692D25A4B49696D2DA5A4B4B69692D2D25A5A5B4B4B4B696969696D2D2D2D2D2D2D2D2D2D2D2D2D2D29696969694B4B4B5A5A5AD2D2D696B4B4A5A52D29694B4A5AD29694B5A52D694B5A52D6B4A5AD694A5AD694A5AD6B4A5294B5AD6B5AD694A5294A5294A5294A52B5AD6B5AD4A5295AD6B5294AD6B5295AD4A56B5295AD4AD6A56B52B5A95A95AD4AD4AD4AD4AD4AD4AD4AD5A95A95AB52B56A54AD5A952B56A54A95AB56AD5A952A54A952A54AB56AD5AA54A956AD52A55AA54AB54AB54AB54AB54AB54AA55AA552AD56AB55AA552A9";

arriav_ram_block ram_block1a1(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a1_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.clk0_input_clock_enable = "ena0";
defparam ram_block1a1.clk0_output_clock_enable = "ena0";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.init_file = "DDS_48_v1_nco_ii_0_sin.hex";
defparam ram_block1a1.init_file_layout = "port_a";
defparam ram_block1a1.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_c8g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.operation_mode = "rom";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 13;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "clock0";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 8191;
defparam ram_block1a1.port_a_logical_ram_depth = 65536;
defparam ram_block1a1.port_a_logical_ram_width = 16;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.ram_block_type = "auto";
defparam ram_block1a1.mem_init3 = "2A954AB55AAD56A954AB54AA55AA55AA55AA55AA55AA54AB54A956AD52A54AB56AD5AA54A952A54A952B56AD5AB52A54AD5A952B56A54AD5A95AB52B52B56A56A56A56A56A56A56A56B52B52B5A95AD4AD6A56B5295AD4A56B5295AD6A5295AD6B5294A56B5AD6B5A94A5294A5294A5294A52D6B5AD6B5A5294A5AD6B4A52D6B4A52D6B4A5AD694B5A52D694B5A52D296B4A5A52D29694B4A5A5AD2D69696B4B4B5A5A5A52D2D2D2D29696969696969696969696969696D2D2D2D2DA5A5A5B4B4B4969692D2DA5A4B4B696D2D25A4B49692D25B4B696D25A4B692D25B496D25A4B692DA4B6D25B496D24B692DB496DA4B6D24B6925B6925B6925B6924B6D2496";
defparam ram_block1a1.mem_init2 = "DB4925B6D2496DB692496DB692496DB6DA4924B6DB6DA4924924B6DB6DB6DB4924924924924924924924924924924924924924924DB6DB6DB6D924924936DB6DB24924DB6DB24924DB6D924936DB24936DB24936D9249B6C926DB249B6C926DB24DB649B6C936C926D926D926D926D926D926D926D936C93649B64DB26D936C9B64DB26D93649B26D9364DB26C9B24D9364D926C9B26C9B26C9B26C9B26C9B26C9B264D9364D9326C9B364D9326C9B364D9B26CD9326CD9366C99366CD9326CD9B264D9B366C993264C9B366CD9B366CD9B366CD9B366CD9B3264C993366CD993266CD993266CD993366CC99B3266CC99B3666CC99B3266CC99933664CC99B33";
defparam ram_block1a1.mem_init1 = "666CC999332664CC999332666CCD99B332664CCD9993336664CCD999B3326664CCD999B33326664CCCD999B333266664CCCD9999B3333266666CCCCC999999333332666666CCCCCCD9999999B33333336666666664CCCCCCCCCC9999999999999B33333333333333333326666666666666666666666666666666666666666666666666663333333333333333333319999999999999CCCCCCCCCCC666666666733333333199999998CCCCCCC66666673333331999998CCCCCE6666633333399999CCCCCE66663333319998CCCCE6666333319998CCCC666633331999CCCCE66633339998CCCE6663331999CCCC6663331999CCCE667333999CCCE667333998CCC";
defparam ram_block1a1.mem_init0 = "666333999CCC666333999CCC66733199CCCE66333998CCE6633399CCC66733199CCE6633399CCC66733998CC66733998CC6633399CCE6633198CC6673399CCE6733198CC6633198CC6633198CC6633198CC663319CCE673399CCE633198CC663399CCE633198CE673398CC663399CCE63319CCE63319CCE673198CE67319CCE63319CCE63319CC663399CC673398CE67319CCE63399CC673398CE67319CC663398CE67319CC663398CE67319CC673398CE63398CC67319CC673398CE63398CE67319CC67319CC663398CE63398CE63399CC67319CC67319CC67319CC663398CE63398CE63398CE63398CE63398CC67319CC67319CC67319CC67319CC67319CC6";

arriav_ram_block ram_block1a17(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a17_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a17.clk0_core_clock_enable = "ena0";
defparam ram_block1a17.clk0_input_clock_enable = "ena0";
defparam ram_block1a17.clk0_output_clock_enable = "ena0";
defparam ram_block1a17.data_interleave_offset_in_bits = 1;
defparam ram_block1a17.data_interleave_width_in_bits = 1;
defparam ram_block1a17.init_file = "DDS_48_v1_nco_ii_0_sin.hex";
defparam ram_block1a17.init_file_layout = "port_a";
defparam ram_block1a17.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_c8g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a17.operation_mode = "rom";
defparam ram_block1a17.port_a_address_clear = "none";
defparam ram_block1a17.port_a_address_width = 13;
defparam ram_block1a17.port_a_data_out_clear = "none";
defparam ram_block1a17.port_a_data_out_clock = "clock0";
defparam ram_block1a17.port_a_data_width = 1;
defparam ram_block1a17.port_a_first_address = 8192;
defparam ram_block1a17.port_a_first_bit_number = 1;
defparam ram_block1a17.port_a_last_address = 16383;
defparam ram_block1a17.port_a_logical_ram_depth = 65536;
defparam ram_block1a17.port_a_logical_ram_width = 16;
defparam ram_block1a17.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a17.ram_block_type = "auto";
defparam ram_block1a17.mem_init3 = "FFFFFFFFFFFFFFFFFFFFFFFFE0000000000000FFFFFFFFFE00000001FFFFFFE000000FFFFFE00000FFFFF00001FFFF80001FFFE0001FFFC0007FFE0007FFE000FFF8007FF8007FF800FFF001FFC00FFE007FE007FE007FC00FF803FE00FF803FE01FF00FF007F807F807F00FF00FE01FC07F80FE03F80FE03F80FE03F01F80FE07F03F01F81F80FC0FC0FC0FC0FC1F81F81F03F07E0FC1F83F07E0F81F07E0F83E07C1F07C1F07C1F07C1F0783E0F87C1F0F83C1E0F87C3E1F0F87C3E1F0F0787C3C1E1E0F0F0F878787C3C3C3C3C3C3C3C3C3C3C3C3C38787878F0F0E1E1C3C3878F0E1E3C3870F1E3C3870E1C3870E1C3870E3C78E1C38F1C38F1C38F1C38E";
defparam ram_block1a17.mem_init2 = "1C70E38F1C78E38F1C71E38E38E1C71C71C71C38E38E38E38E38E71C71C71C718E38E39C71C638E31C718E39C718E31C638C718E71CE31C639C639C639CE31CE718E738C631CE738C6318E739CE739CE739CE739CC6318C6739CC6319CE6319CE6339CC67319CE63398CE67319CC663399CC6633198CC6633198CCE6633199CCC666333199CCCC66633339999CCCCE66667333339999998CCCCCCCC66666666666666667333333333266666666666666664CCCCCCCD999999B3333266666CCCC9999B3336666CCC999B332664CC999332664CD99B3266CC99B3264CD993266CD9B3264C993264C99326CD9B364C9B366C99364C9B264D9366C9B26C99364D936";
defparam ram_block1a17.mem_init1 = "4D926C9B26C9B64D926C9B64DB26D936C93649B649B649B649B6C936D926DB249B6C924DB6C924DB6C9249B6DB64924926DB6DB6DB24924924924924924924924925B6DB6DB6D2492496DB6D24925B6D2492DB6924B6D2496DA496DA496D24B6925B496DA4B692DA4B692DA5B496D2DA5B49692D25A4B4B69692D2DA5A5B4B4B49696969696D2D2D2D2D2D2D29696969696B4B4B5A5A5AD2D29694B4A5A52D694B4A5AD296B4A52D694A5AD694A52D6B5A5294A5296B5AD6B5AD6B5AD4A5294A56B5AD4A5295AD4A52B5A94AD4A56B52B5A95A95AD4AD4AD4AD4AD4AD4AD5A95A952B52A56AD4A95AB56A54A952A56AD5AB56A952A54A956AD52A55AB54AB54A";
defparam ram_block1a17.mem_init0 = "956A956A954AB54AB55AA552A954AB55AAD56AA552A955AA954AAD54AAD55AA955AAB556AAD55AAB554AAB556AA9554AAB555AAAD554AAA5556AAA5554AAA95556AAA95556AAAB55552AAAB55554AAAAB55555AAAAA9555556AAAAAA5555555AAAAAAAB555555556AAAAAAAAAA55555555555555AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA55555555555555AAAAAAAAAAB555555554AAAAAAA95555554AAAAAAD555552AAAAA555552AAAA955556AAAAD5554AAAA55552AAA95556AAAD555AAAB5552AAA5552AAB555AAAD556AA9554AAB554AAB556AA9552AA554AA9552AB556AA556AA556AA556AB552AB55AAD54AA55";

arriav_ram_block ram_block1a66(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a66_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a66.clk0_core_clock_enable = "ena0";
defparam ram_block1a66.clk0_input_clock_enable = "ena0";
defparam ram_block1a66.clk0_output_clock_enable = "ena0";
defparam ram_block1a66.data_interleave_offset_in_bits = 1;
defparam ram_block1a66.data_interleave_width_in_bits = 1;
defparam ram_block1a66.init_file = "DDS_48_v1_nco_ii_0_sin.hex";
defparam ram_block1a66.init_file_layout = "port_a";
defparam ram_block1a66.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_c8g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a66.operation_mode = "rom";
defparam ram_block1a66.port_a_address_clear = "none";
defparam ram_block1a66.port_a_address_width = 13;
defparam ram_block1a66.port_a_data_out_clear = "none";
defparam ram_block1a66.port_a_data_out_clock = "clock0";
defparam ram_block1a66.port_a_data_width = 1;
defparam ram_block1a66.port_a_first_address = 32768;
defparam ram_block1a66.port_a_first_bit_number = 2;
defparam ram_block1a66.port_a_last_address = 40959;
defparam ram_block1a66.port_a_logical_ram_depth = 65536;
defparam ram_block1a66.port_a_logical_ram_width = 16;
defparam ram_block1a66.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a66.ram_block_type = "auto";
defparam ram_block1a66.mem_init3 = "3664CD9933664CD9B3266CC993366CC993366CC993366CD993264C99B366CD9B3264C993264C993264C993264D9B366CD9B264C99366CD93264D9B364C99366C99366C99366C99366C9B364C9B264D9326C99364C9B26CD9364D9B26C9B364D9364D9B26C9B26C9B26C9B26C9B26C9B26C9B26C9B26C9B26C9364D9364DB26C9B24D93649B26C9364DB26C9364DB26C93649B24D936C9B649B24D926C936C9B649B24DB24D926D926C936C936C936C936C936C936C936D926D926D924DB24DB649B6C936D924DB249B6C936D924DB64936D924DB64926DB249B6D9249B6C924DB6C924DB6C924DB6D9249B6DB24926DB6C9249B6DB649249B6DB64924936DB6D";
defparam ram_block1a66.mem_init2 = "9249249B6DB6DB24924924DB6DB6DB649249249249B6DB6DB6DB6DB6C924924924924924924924924924924924924924924924924924925B6DB6DB6DB6DB6D24924924924B6DB6DB6D24924924B6DB6DB4924924B6DB6D2492496DB6DA4924B6DB6D24925B6DA4924B6DB4924B6DB4924B6DB4924B6DA4925B6D2496DB4925B6D2496DB4925B6924B6DA496DA492DB4925B6925B6925B6D24B6D24B6D24B6925B6925B692DB492DB496DA496D24B6925B492DA496D25B692DB496D24B692DA496D25B496DA4B692DA4B692DA496D25B496D25B496D2DA4B692DA4B692DA5B496D25B4B692DA4B496D25A4B692D25B4B692D25B4B692D25A4B696D2DA4B49692D";
defparam ram_block1a66.mem_init1 = "25B4B696D2DA5B4B696D2DA5B4B69692D25A4B4B696D2DA5A4B4B696D2D25A5B4B49696D2D25A5B4B4969692D2DA5A5B4B4B69696D2D2DA5A5B4B4B4969696D2D2D25A5A5A4B4B4B496969692D2D2D2D25A5A5A5A4B4B4B4B4B496969696969692D2D2D2D2D2D2D2D2D2DA5A5A5A5A5A5A5A5A5A5A5A5A5A5A5A5A5A5A5A5A5A5A5A5A5A52D2D2D2D2D2D2D2D2D296969696969696B4B4B4B4B4B5A5A5A5A5AD2D2D2D2D6969696B4B4B4B5A5A5A5AD2D2D2969696B4B4B4A5A5A5AD2D2D69696B4B4B5A5A5AD2D2969694B4B5A5A52D2D29696B4B4A5A5AD2D69694B4B5A5AD2D29696B4B5A5AD2D29694B4A5A5AD2D696B4B5A5AD2D696B4B5A5AD2D696B4B";
defparam ram_block1a66.mem_init0 = "5A52D29694B4A5AD2D696B4A5A52D296B4B5A52D296B4B5A52D296B4B5A52D696B4A5A52D694B5A5AD296B4B5A52D694B5A5AD296B4A5AD29694B5A52D694B5A52D694B5A52D694B4A5AD296B4A52D694B5A52D694B5A52D694B5A52D6B4A5AD296B4A5AD294B5A52D694B5AD296B4A5AD694B5A5296B4A5AD294B5A52D6B4A5AD694B5A5296B4A52D694A5AD296B5A52D6B4A5AD694B5AD296B5A5296B4A52D694A5AD694B5AD296B5A5296B4A52D6B4A5AD694A5AD694B5AD294B5A5296B5A5296B5A52D6B4A52D6B4A52D694A5AD694A5AD694A5AD294B5AD294B5AD294B5AD294B5A5296B5A5296B5A5296B5A5296B5A5296B5A5296B5A52D6B4A52D6B4A";

arriav_ram_block ram_block1a82(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a82_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a82.clk0_core_clock_enable = "ena0";
defparam ram_block1a82.clk0_input_clock_enable = "ena0";
defparam ram_block1a82.clk0_output_clock_enable = "ena0";
defparam ram_block1a82.data_interleave_offset_in_bits = 1;
defparam ram_block1a82.data_interleave_width_in_bits = 1;
defparam ram_block1a82.init_file = "DDS_48_v1_nco_ii_0_sin.hex";
defparam ram_block1a82.init_file_layout = "port_a";
defparam ram_block1a82.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_c8g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a82.operation_mode = "rom";
defparam ram_block1a82.port_a_address_clear = "none";
defparam ram_block1a82.port_a_address_width = 13;
defparam ram_block1a82.port_a_data_out_clear = "none";
defparam ram_block1a82.port_a_data_out_clock = "clock0";
defparam ram_block1a82.port_a_data_width = 1;
defparam ram_block1a82.port_a_first_address = 40960;
defparam ram_block1a82.port_a_first_bit_number = 2;
defparam ram_block1a82.port_a_last_address = 49151;
defparam ram_block1a82.port_a_logical_ram_depth = 65536;
defparam ram_block1a82.port_a_logical_ram_width = 16;
defparam ram_block1a82.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a82.ram_block_type = "auto";
defparam ram_block1a82.mem_init3 = "00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFE00000000000000FFFFFFFFFFFC0000000003FFFFFFFFC00000001FFFFFFFC0000003FFFFFF8000001FFFFFE000001FFFFF800001FFFFF00000FFFFF00001FFFFC0000FFFFC0001FFFF0000FFFF80007FFF0000FFFE0003FFF0001FFF8001FFF8003FFF0007FFC001FFE000FFF0007FF8007FF8007FF000FFE003FFC007FF001FF800FFE007FF003FF001FF801FF801FF003FF007FE00FFC01FF803FE00FF803FE00FF803FC01FF00FF803FC03FE01FE00FF00FF00FF00FF00FF00FF00FE01FE03FC03F807F00FE01FC07F80FE03F807F01FC07F01FC07F01FC07F03F80FE07F01F80FE07F03F";
defparam ram_block1a82.mem_init2 = "81FC0FE07F03F01F81FC0FC07E07E07F03F03F03F03F03F03F03F03F03F07E07E07C0FC0F81F81F03F07E0FC0F81F03E07C0F81F03E0FC1F83E07C1F83E0FC1F07E0F83E07C1F07C1F83E0F83E0F83E0F83E0F83E0F83C1F07C1F0783E0F87C1F0F83E1F07C3E0F07C3E0F07C3E1F0783C1E0F07C3E1F0F8783C1E0F0787C3E1E0F0787C3C1E1F0F0F8783C3C1E1E0F0F0F878783C3C3C1E1E1E1E1F0F0F0F0F0F0F0F0F87878787870F0F0F0F0F0F0F0F1E1E1E1E1C3C3C38787870F0F1E1E1C3C387870F0E1E1C3C7878F0E1E3C3878F0E1E3C7870E1E3C7870E1E3C78F1E1C3870E1C3870E1C3870E1C78F1E3C78E1C38F1E3C70E1C78E1C38F1C38F1C38F";
defparam ram_block1a82.mem_init1 = "1C38F1C38E1C78E3C70E3871C38E1C70E38F1C78E3871C78E38F1C70E38E3C71C70E38E3871C71C78E38E38E1C71C71C71C71E38E38E38E38E38E38E38E38E38E38E38E39C71C71C71C718E38E38E39C71C718E38E39C71C738E38C71C638E39C718E38C71CE38C71CE38C71CE39C718E31C638C718E31C639C738E718E31CE31C639C639C638C738C738C739C639C639C631CE318E718C739C631CE718C739C6318E739C6318E739CE318C631CE739CE739C6318C6318C6318C6318C6318CE739CE739CE6318C6339CE7318C6339CE6318CE7318C67398C67398C67398CE7318CE6319CC63398CE6319CC67319CC67319CC67319CC673198CE63399CC673398";
defparam ram_block1a82.mem_init0 = "CE673198CE673398CC663319CCE673399CCE6733998CC6633199CCE6633199CCC66733998CCE66733199CCC666333199CCCE667333999CCCC66633339998CCCE666733319998CCCC66667333319999CCCCCE66667333331999998CCCCCCE6666667333333339999999998CCCCCCCCCCCE666666666666666663333333333333333333333333333333333333333332666666666666666666CCCCCCCCCCCD999999999B3333333266666664CCCCCC999999B33333666666CCCCC999993333266664CCCC9999B33366664CCC9999B3336664CCC999B3336664CCD9993336664CC999B33666CCC999332664CC99933266CCD99B32664CD99B3266CCD9933664CD993";

arriav_ram_block ram_block1a98(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a98_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a98.clk0_core_clock_enable = "ena0";
defparam ram_block1a98.clk0_input_clock_enable = "ena0";
defparam ram_block1a98.clk0_output_clock_enable = "ena0";
defparam ram_block1a98.data_interleave_offset_in_bits = 1;
defparam ram_block1a98.data_interleave_width_in_bits = 1;
defparam ram_block1a98.init_file = "DDS_48_v1_nco_ii_0_sin.hex";
defparam ram_block1a98.init_file_layout = "port_a";
defparam ram_block1a98.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_c8g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a98.operation_mode = "rom";
defparam ram_block1a98.port_a_address_clear = "none";
defparam ram_block1a98.port_a_address_width = 13;
defparam ram_block1a98.port_a_data_out_clear = "none";
defparam ram_block1a98.port_a_data_out_clock = "clock0";
defparam ram_block1a98.port_a_data_width = 1;
defparam ram_block1a98.port_a_first_address = 49152;
defparam ram_block1a98.port_a_first_bit_number = 2;
defparam ram_block1a98.port_a_last_address = 57343;
defparam ram_block1a98.port_a_logical_ram_depth = 65536;
defparam ram_block1a98.port_a_logical_ram_width = 16;
defparam ram_block1a98.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a98.ram_block_type = "auto";
defparam ram_block1a98.mem_init3 = "933664CD9933666CC99B33664CC99B33666CC999332664CC999332666CCD99B332664CCD9993336664CCD999B3326664CCD999B33326664CCCD999B333266664CCCC999993333266666CCCCCD99999B3333326666664CCCCCCC99999999B333333333666666666666CCCCCCCCCCCCCCCCCC9999999999999999999999999999999999999999998CCCCCCCCCCCCCCCCCE66666666666333333333399999999CCCCCCCE666666333333199999CCCCCE66667333319999CCCCC666633331999CCCCE66633339998CCC6667333999CCCE667331998CCC66733199CCCE6633399CCC66733198CCE6733198CC6633399CCE673399CCE673198CC663399CCE63319CCE6";
defparam ram_block1a98.mem_init2 = "3399CC673398CE63319CC67319CC67319CC67319CC67318CE63398C67318CE6319CE6339CC6339CC6339CC6319CE6318CE7398C6319CE7398C6318CE739CE739CE6318C6318C6318C6318C6318C739CE739CE718C6318E739CE318C739CE318C739C631CE718C739C631CE318E718C738C738C739C639C639C638C738C738C718E718E31CE39C738C718E31C638C718E31C738E71C638E71C638E71C638E31C738E38C71C638E39C71C738E38E31C71C738E38E38E31C71C71C71C738E38E38E38E38E38E38E38E38E38E38E38F1C71C71C71C70E38E38E3C71C71C38E38E1C71C78E38E1C71E38E3C71C38E3C71E38E1C70E3871C38E1C78E3C70E3871E3871";
defparam ram_block1a98.mem_init1 = "E3871E3871E3870E3C70E1C78F1E3870E3C78F1E3C70E1C3870E1C3870E1C3870F1E3C78F0E1C3C78F0E1C3C78F0E1E3C3878F0E1E3C3C7870F0E1E1C3C387870F0F1E1E1C3C3C38787870F0F0F0F1E1E1E1E1E1E1E1E1C3C3C3C3C3E1E1E1E1E1E1E1E1F0F0F0F0F07878783C3C3E1E1E0F0F078783C3E1E1F0F0787C3C1E0F0F87C3C1E0F0783C3E1F0F87C1E0F0783C1F0F87C1E0F87C1E0F87C1F0F83E1F07C3E0F83C1F07C1F0783E0F83E0F83E0F83E0F83E0F83F07C1F07C0F83E0FC1F07E0F83F07C0F83F07E0F81F03E07C0F81F03E07E0FC1F81F03F03E07E07C0FC0FC1F81F81F81F81F81F81F81F81F81FC0FC0FC07E07F03F01F81FC0FE07F03";
defparam ram_block1a98.mem_init0 = "F81FC0FE03F01FC0FE03F81FC07F01FC07F01FC07F01FC03F80FE03FC07F00FE01FC03F807F80FF00FE01FE01FE01FE01FE01FE01FE00FF00FF807F803FE01FF007F803FE00FF803FE00FF803FF007FE00FFC01FF801FF003FF003FF001FF801FFC00FFE003FF001FFC007FF800FFE001FFC003FFC003FFC001FFE000FFF0007FFC001FFF8003FFF0003FFF0001FFF8000FFFE0001FFFC0003FFFE0001FFFF00007FFFE00007FFFF00001FFFFE00001FFFFF000003FFFFF000000FFFFFF0000003FFFFFF80000007FFFFFFF000000007FFFFFFFF80000000007FFFFFFFFFFE00000000000000FFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000";

arriav_ram_block ram_block1a114(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a114_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a114.clk0_core_clock_enable = "ena0";
defparam ram_block1a114.clk0_input_clock_enable = "ena0";
defparam ram_block1a114.clk0_output_clock_enable = "ena0";
defparam ram_block1a114.data_interleave_offset_in_bits = 1;
defparam ram_block1a114.data_interleave_width_in_bits = 1;
defparam ram_block1a114.init_file = "DDS_48_v1_nco_ii_0_sin.hex";
defparam ram_block1a114.init_file_layout = "port_a";
defparam ram_block1a114.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_c8g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a114.operation_mode = "rom";
defparam ram_block1a114.port_a_address_clear = "none";
defparam ram_block1a114.port_a_address_width = 13;
defparam ram_block1a114.port_a_data_out_clear = "none";
defparam ram_block1a114.port_a_data_out_clock = "clock0";
defparam ram_block1a114.port_a_data_width = 1;
defparam ram_block1a114.port_a_first_address = 57344;
defparam ram_block1a114.port_a_first_bit_number = 2;
defparam ram_block1a114.port_a_last_address = 65535;
defparam ram_block1a114.port_a_logical_ram_depth = 65536;
defparam ram_block1a114.port_a_logical_ram_width = 16;
defparam ram_block1a114.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a114.ram_block_type = "auto";
defparam ram_block1a114.mem_init3 = "A5AD694A5AD694B5AD294B5AD294B5AD294B5AD294B5AD294B5AD294B5A5296B5A5296B5A5296B5A5296B4A52D6B4A52D6B4A52D694A5AD694A5AD694B5AD294B5AD294B5A5296B5A52D6B4A52D6B4A5AD694A5AD294B5AD296B5A52D6B4A52D694A5AD294B5AD296B5A52D6B4A5AD694B5AD296B4A52D694A5AD294B5A52D6B4A5AD694B5A5296B4A5AD294B5A52D6B4A5AD296B5A52D694B5A5296B4A5AD296B4A5AD694B5A52D694B5A52D694B5A52D694A5AD296B4A5A52D694B5A52D694B5A52D694B5A52D296B4A5AD296B4B5A52D694B5A5AD296B4B5A52D694B4A5AD2D694B5A5AD29694B5A5AD29694B5A5AD29694B4A5AD2D696B4A5A52D29694B5";
defparam ram_block1a114.mem_init2 = "A5AD2D696B4B5A5AD2D696B4B5A5AD2D696B4B4A5A52D29696B4B5A5AD2D29696B4B5A5A52D2D696B4B4A5A5AD2D2969694B4B5A5A52D2D29696B4B4B5A5A5AD2D2D69696B4B4B4A5A5A5AD2D2D2969696B4B4B4B5A5A5A5AD2D2D2D696969696B4B4B4B4B5A5A5A5A5A5AD2D2D2D2D2D2D296969696969696969694B4B4B4B4B4B4B4B4B4B4B4B4B4B4B4B4B4B4B4B4B4B4B4B4B4B696969696969696969692D2D2D2D2D2D25A5A5A5A5A4B4B4B4B49696969692D2D2D25A5A5A4B4B4B4969696D2D2D25A5A5B4B4B69696D2D2DA5A5B4B4B69692D2D25A5B4B49696D2D25A5B4B49696D2DA5A4B4B696D2DA5A4B49692D2DA5B4B696D2DA5B4B696D2DA5B49";
defparam ram_block1a114.mem_init1 = "692D25A4B696D2DA4B49692DA5B49692DA5B49692DA4B496D25A4B692DA5B496D25B4B692DA4B692DA4B696D25B496D25B496D24B692DA4B692DA4B6D25B496D24B692DA496D25B692DB496D24B6925B492DA496D24B6D25B6925B692DB492DB492DA496DA496DA496DB492DB492DB4925B6924B6D24B6DA492DB4925B6D2496DB4925B6D2496DB4924B6DA4925B6DA4925B6DA4925B6DA4924B6DB492496DB6DA4924B6DB6D2492496DB6DA4924925B6DB6DA492492496DB6DB6DA492492492496DB6DB6DB6DB6DB4924924924924924924924924924924924924924924924924924926DB6DB6DB6DB6DB24924924924DB6DB6DB649249249B6DB6DB2492493";
defparam ram_block1a114.mem_init0 = "6DB6D924924DB6DB24924DB6DB24926DB6C9249B6DB24936DB64926DB64926DB64926DB24936DB249B6C924DB64936D924DB64936D926DB249B64936D926DB24DB649B64936C936C936D926D926D926D926D926D926D926C936C93649B649B24DB26D926C93649B24DB26D93649B24D926C9B64D926C9B64D926C9B24D93649B26C9B64D9364D926C9B26C9B26C9B26C9B26C9B26C9B26C9B26C9B26C9B364D9364D9B26C9B364D9366C9B264D9326C99364C9B264D9B26CD9326CD9326CD9326CD93264D9B364C99366CD93264C9B366CD9B364C993264C993264C993264C99B366CD9B3264C993366CD993266CD993266CD993266CC99B3664CD9933664CD9";

arriav_ram_block ram_block1a34(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a34_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a34.clk0_core_clock_enable = "ena0";
defparam ram_block1a34.clk0_input_clock_enable = "ena0";
defparam ram_block1a34.clk0_output_clock_enable = "ena0";
defparam ram_block1a34.data_interleave_offset_in_bits = 1;
defparam ram_block1a34.data_interleave_width_in_bits = 1;
defparam ram_block1a34.init_file = "DDS_48_v1_nco_ii_0_sin.hex";
defparam ram_block1a34.init_file_layout = "port_a";
defparam ram_block1a34.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_c8g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a34.operation_mode = "rom";
defparam ram_block1a34.port_a_address_clear = "none";
defparam ram_block1a34.port_a_address_width = 13;
defparam ram_block1a34.port_a_data_out_clear = "none";
defparam ram_block1a34.port_a_data_out_clock = "clock0";
defparam ram_block1a34.port_a_data_width = 1;
defparam ram_block1a34.port_a_first_address = 16384;
defparam ram_block1a34.port_a_first_bit_number = 2;
defparam ram_block1a34.port_a_last_address = 24575;
defparam ram_block1a34.port_a_logical_ram_depth = 65536;
defparam ram_block1a34.port_a_logical_ram_width = 16;
defparam ram_block1a34.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a34.ram_block_type = "auto";
defparam ram_block1a34.mem_init3 = "CD9933266CC99B33664CD99B32664CD99B33664CC999332664CC999B33666CCC9993336664CCD9993336664CCD999B3336666CCCD999B33366664CCCD99993333266664CCCC99999B33332666664CCCCCD999999333333366666666CCCCCCCCC9999999999933333333333332666666666666666666666666666666666666666666666666666666666666667333333333333339999999999CCCCCCCCC666666673333333999999CCCCCCE666673333399999CCCCC6666733339999CCCCE66633331999CCCC6663333999CCCE667333999CCCE66333999CCC66733199CCC66733198CCE6633199CCE6733198CC6633198CC6633198CC673399CC663319CCE6331";
defparam ram_block1a34.mem_init2 = "9CC663398CC67319CCE63398CE63398CE63398CE6339CC67319CE63398C67318CE7319CE6319CE6319CE6318CE7318C6739CC6319CE7398C6318CE739CE739CC6318C6318C6318C6318C6318C6318C739CE739CE318C631CE739C6318E739C631CE738C639CE318E718C738C639C631CE31CE318E718E718E718E31CE31CE31C639C738C718E71CE39C638C718E31C738E71CE38C718E39C718E39C71CE38C71C638E31C71CE38E31C71C638E38E71C71C738E38E38E31C71C71C71C71C738E38E38E38E38E38E38E38E3871C71C71C71C71C38E38E38E1C71C71E38E38E1C71C78E38F1C71E38E3C71C38E3C71C38E1C70E3871C38E1C70E3C71E3871E38F1C";
defparam ram_block1a34.mem_init1 = "38F1C38F1E3871E3C70E3C78E1C38F1E3C78E1C3870E1C78F1E3C78F1E3C7870E1C3870F1E3C7870E1E3C7870F1E3C3878F0E1E3C387870F1E1E3C3C7878F0F1E1E1C3C3C787878F0F0F0E1E1E1E1C3C3C3C3C3C3C3C3C78787878783C3C3C3C3C3C3C3C3E1E1E1E1F0F0F0F878783C3C3E1E1F0F0F8787C3C1E1F0F0787C3C1E0F0F87C3E1E0F0783C1E0F0783C1F0F87C3E0F07C3E1F0783E0F07C3E0F87C1F0F83E0F07C1F07C3E0F83E0F83E0F83E0F83E0F83E0F83E07C1F07C1F83E0FC1F07E0F83F07C0F83F07E0FC1F03E07C0F81F03F07E0FC0F81F83F03F07E07E0FC0FC0FC0FC1F81F81F81F81F80FC0FC0FC0FE07E07F03F01F81FC0FE07E03F0";
defparam ram_block1a34.mem_init0 = "1F80FE07F01F80FE07F01FC07E03F80FE03F80FE03F807F01FC07F80FE01FC07F80FF01FE01FC03FC07F807F807F807F807F807F807FC03FC01FE01FF00FF803FC01FF007FC01FF007FC01FF007FE00FFC01FF803FF003FF003FF003FF003FF801FFC00FFE003FF800FFE003FF800FFF000FFE001FFE001FFE000FFF0007FFC001FFF0007FFE0007FFE0007FFE0003FFF0001FFFE0003FFFC0003FFFE0000FFFF80001FFFF80001FFFFC00003FFFFC00001FFFFF000001FFFFFC000003FFFFFE0000003FFFFFFC0000000FFFFFFFF000000000FFFFFFFFFE00000000001FFFFFFFFFFFFF000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

arriav_ram_block ram_block1a50(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a50_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a50.clk0_core_clock_enable = "ena0";
defparam ram_block1a50.clk0_input_clock_enable = "ena0";
defparam ram_block1a50.clk0_output_clock_enable = "ena0";
defparam ram_block1a50.data_interleave_offset_in_bits = 1;
defparam ram_block1a50.data_interleave_width_in_bits = 1;
defparam ram_block1a50.init_file = "DDS_48_v1_nco_ii_0_sin.hex";
defparam ram_block1a50.init_file_layout = "port_a";
defparam ram_block1a50.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_c8g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a50.operation_mode = "rom";
defparam ram_block1a50.port_a_address_clear = "none";
defparam ram_block1a50.port_a_address_width = 13;
defparam ram_block1a50.port_a_data_out_clear = "none";
defparam ram_block1a50.port_a_data_out_clock = "clock0";
defparam ram_block1a50.port_a_data_width = 1;
defparam ram_block1a50.port_a_first_address = 24576;
defparam ram_block1a50.port_a_first_bit_number = 2;
defparam ram_block1a50.port_a_last_address = 32767;
defparam ram_block1a50.port_a_logical_ram_depth = 65536;
defparam ram_block1a50.port_a_logical_ram_width = 16;
defparam ram_block1a50.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a50.ram_block_type = "auto";
defparam ram_block1a50.mem_init3 = "52D6B4A52D6B4A52D6B4A52D6B4A52D6B4A52D694A5AD694A5AD694A5AD694A5AD694A5AD294B5AD294B5AD294B5AD296B5A5296B5A5296B5A52D6B4A52D6B4A5AD694A5AD694B5AD294B5AD296B5A5296B4A52D6B4A5AD694A5AD294B5A5296B5A52D6B4A5AD694B5AD296B5A52D6B4A5AD694B5AD296B5A52D6B4A5AD294B5A52D6B4A5AD694B5A52D6B4A5AD294B5A52D694A5AD296B4A5AD694B5A52D694A5AD296B4A5AD296B4A5AD294B5A52D694B5A52D694B5A52D694B5A52D694B4A5AD296B4A5AD296B4A5A52D694B5A52D696B4A5AD29694B5A52D296B4A5A52D694B4A5AD2D694B5A5AD29694B5A5AD2D694B4A5AD2D696B4A5A52D29694B5A5A";
defparam ram_block1a50.mem_init2 = "D2D696B4B5A5AD2D696B4B5A5AD2D696B4B5A5AD2D29694B4A5A5AD2D69694B4A5A5AD2D29694B4B5A5A52D2D69694B4B5A5A5AD2D29696B4B4B5A5A5AD2D2D69696B4B4B5A5A5A52D2D2969696B4B4B4B5A5A5A52D2D2D296969696B4B4B4B4B5A5A5A5A5AD2D2D2D2D2D6969696969696B4B4B4B4B4B4B4B4B4B4A5A5A5A5A5A5A5A5A5A5A5A5A5A5A5A5A5A5A5A5A5A5A5A5A5A5B4B4B4B4B4B4B4B4B4B696969696969692D2D2D2D2D25A5A5A5A4B4B4B4B696969692D2D2D25A5A5A4B4B4B6969692D2D25A5A5B4B4B69696D2D2DA5A5B4B49696D2D2DA5A4B4B69692D2DA5A4B49696D2D25A4B4B696D2D25A4B49692D25A5B4B696D2DA5B4B696D25A4";
defparam ram_block1a50.mem_init1 = "B49692D25B4B696D25A4B696D25A4B696D25A4B696D25B4B692DA5B496D25A4B692DA4B496D25B496D25B496D25B496D25B496D25B496D25B496DA4B692DA496D25B492DA4B6925B492DA4B6D25B692DB496DA4B6D24B6925B492DB492DA496DA496DA496DA496DA496DA496DA492DB492DB6925B6D24B6DA496DB4925B6D2496DB4925B6D2496DB4924B6DA4925B6DA4925B6DA4925B6DA4924B6DB692492DB6DA492496DB6DA492496DB6DB4924924B6DB6DB492492492DB6DB6DB6D24924924924B6DB6DB6DB6DB6DB6D24924924924924924924924924924924924924924936DB6DB6DB6DB6DB6D924924924926DB6DB6DB649249249B6DB6DB24924936D";
defparam ram_block1a50.mem_init0 = "B6DB249249B6DB649249B6DB64924DB6D924936DB64924DB6C924DB6D9249B6D924DB6C924DB64926DB249B6C924DB64936D924DB249B6C926D924DB649B6C936C926D926DB24DB24DB649B649B649B649B649B649B649B24DB24DB26D926C936C9B649B24D926D936C9B64DB26D93649B24D936C9B24D936C9B26D9364DB26C9B24D9364D926C9B26C9B26C9B24D9364D9364D9364D9366C9B26C9B26C9B364D9364D9B26C9B364D9326C9B364D9B26CD9366C9B364C9B264D9B264D9B264D9B264C9B364C99366CD93264C9B366CD93264C993264C9B366CD9B366CD993264C993264CD9B366CC993266CD993266CD993266CD993366CC99B3266CC9933664";

arriav_ram_block ram_block1a2(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a2_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.clk0_input_clock_enable = "ena0";
defparam ram_block1a2.clk0_output_clock_enable = "ena0";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.init_file = "DDS_48_v1_nco_ii_0_sin.hex";
defparam ram_block1a2.init_file_layout = "port_a";
defparam ram_block1a2.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_c8g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.operation_mode = "rom";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 13;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "clock0";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 8191;
defparam ram_block1a2.port_a_logical_ram_depth = 65536;
defparam ram_block1a2.port_a_logical_ram_width = 16;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.ram_block_type = "auto";
defparam ram_block1a2.mem_init3 = "4CD993266CC99B3266CD993366CC993366CC993366CC993266CD9B3664C993264C993366CD9B366CD9B264C993264C99366CD9B264C99366CD93264D9B264C9B364C9B364C9B364C9B264D9B26CD9366C9B364D9B26C99364D9B26C9B364D9364D9B26C9B26C9B26CD9364D9364D9364D93649B26C9B26C9B26C9364D93649B26C9B64D936C9B26D93649B26D93649B24D936C9B64DB26D936C93649B24DB26D926C936C9B649B649B24DB24DB24DB24DB24DB24DB24DB649B649B6C936C926D926DB24DB64936C926DB249B64936D924DB64926DB249B6C924DB64926DB64936DB24936DB64926DB64924DB6D924936DB64924DB6DB24924DB6DB249249B6DB";
defparam ram_block1a2.mem_init2 = "6D9249249B6DB6DB24924924DB6DB6DB6C924924924936DB6DB6DB6DB6DB6D92492492492492492492492492492492492492492496DB6DB6DB6DB6DB6DA492492492496DB6DB6DB6924924925B6DB6DA4924925B6DB6D24924B6DB6D24924B6DB692492DB6DA4924B6DB4924B6DB4924B6DB4924B6DA4925B6D2496DB4925B6D2496DB4925B6D24B6DA496DB492DB6925B6924B6D24B6D24B6D24B6D24B6D24B6D24B6925B6925B492DA496DA4B6D25B692DB496DA4B6925B492DA4B6925B496D24B692DA4B6D25B496D25B496D25B496D25B496D25B496D25B496D25A4B692DA4B496D25B4B692DA5B496D2DA4B496D2DA4B496D2DA4B496D2DA5B49692D25A";
defparam ram_block1a2.mem_init1 = "4B496D2DA5B4B696D2DA5B4B49692D25A4B49696D2DA5A4B49696D2D25A4B4B69692D2DA5A4B4B69696D2D25A5B4B4B69696D2D2DA5A5B4B4B4969692D2D2DA5A5A4B4B4B496969692D2D2D2DA5A5A5A4B4B4B4B4969696969692D2D2D2D2D2D2DA5A5A5A5A5A5A5A5A5B4B4B4B4B4B4B4B4B4B4B4B4B4B4B4B4B4B4B4B4B4B4B4B4B4B4A5A5A5A5A5A5A5A5A5A5AD2D2D2D2D2D2D69696969696B4B4B4B4B5A5A5A5A5AD2D2D2D296969694B4B4B5A5A5A5AD2D2D2969694B4B4B5A5A5AD2D2D69696B4B4B5A5A5AD2D29696B4B4B5A5A52D2D69694B4B5A5A52D29696B4B4A5A52D2D696B4B4A5A52D29696B4B5A5AD2D696B4B5A5AD2D696B4B5A5AD2D696";
defparam ram_block1a2.mem_init0 = "B4B5A52D29694B4A5AD2D696B4A5A52D696B4B5A52D296B4B5A52D696B4A5A52D694B4A5AD29694B5A52D296B4A5AD2D694B5A52D694B4A5AD296B4A5AD296B4A5A52D694B5A52D694B5A52D694B5A52D694B5A5296B4A5AD296B4A5AD296B4A52D694B5A52D6B4A5AD296B4A52D694B5A5296B4A5AD694B5A52D6B4A5AD694B5A5296B4A5AD694B5AD296B5A52D6B4A5AD694B5AD296B5A52D6B4A5AD694B5AD294B5A5296B4A52D6B4A5AD694A5AD294B5AD296B5A5296B5A52D6B4A52D6B4A5AD694A5AD694B5AD294B5AD294B5AD296B5A5296B5A5296B5A5296B4A52D6B4A52D6B4A52D6B4A52D6B4A52D694A5AD694A5AD694A5AD694A5AD694A5AD694";

arriav_ram_block ram_block1a18(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a18_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a18.clk0_core_clock_enable = "ena0";
defparam ram_block1a18.clk0_input_clock_enable = "ena0";
defparam ram_block1a18.clk0_output_clock_enable = "ena0";
defparam ram_block1a18.data_interleave_offset_in_bits = 1;
defparam ram_block1a18.data_interleave_width_in_bits = 1;
defparam ram_block1a18.init_file = "DDS_48_v1_nco_ii_0_sin.hex";
defparam ram_block1a18.init_file_layout = "port_a";
defparam ram_block1a18.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_c8g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a18.operation_mode = "rom";
defparam ram_block1a18.port_a_address_clear = "none";
defparam ram_block1a18.port_a_address_width = 13;
defparam ram_block1a18.port_a_data_out_clear = "none";
defparam ram_block1a18.port_a_data_out_clock = "clock0";
defparam ram_block1a18.port_a_data_width = 1;
defparam ram_block1a18.port_a_first_address = 8192;
defparam ram_block1a18.port_a_first_bit_number = 2;
defparam ram_block1a18.port_a_last_address = 16383;
defparam ram_block1a18.port_a_logical_ram_depth = 65536;
defparam ram_block1a18.port_a_logical_ram_width = 16;
defparam ram_block1a18.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a18.ram_block_type = "auto";
defparam ram_block1a18.mem_init3 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000001FFFFFFFFFFFFF00000000000FFFFFFFFFE000000001FFFFFFFE00000007FFFFFF8000000FFFFFF8000007FFFFF000001FFFFF000007FFFF800007FFFF00003FFFF00003FFFE0000FFFF80007FFF8000FFFF0001FFF8000FFFC000FFFC000FFFC001FFF0007FFC001FFE000FFF000FFF000FFE001FFE003FF800FFE003FF800FFE007FF003FF801FF801FF801FF801FF803FF007FE00FFC01FF007FC01FF007FC01FF007F803FE01FF00FF007F807FC03FC03FC03FC03FC03FC03FC07F807F00FF01FE03FC07F00FE03FC07F01FC03F80FE03F80FE03F80FC07F01FC0FE03F01FC0FE03F0";
defparam ram_block1a18.mem_init2 = "1F80FC0FE07F03F01F81FC0FC0FE07E07E07E03F03F03F03F03F07E07E07E07E0FC0FC1F81F83F03E07E0FC1F81F03E07C0F81F07E0FC1F83E07C1F83E0FC1F07E0F83F07C1F07C0F83E0F83E0F83E0F83E0F83E0F83E0F87C1F07C1E0F83E1F07C3E0F87C1E0F83C1F0F87C1E0F87C3E1F0783C1E0F0783C1E0F0F87C3E1E0F0787C3C1E1F0F0787C3C3E1E1F0F0F878783C3C3E1E1E1F0F0F0F0F878787878787878783C3C3C3C3C787878787878787870F0F0F0E1E1E1E3C3C3C787870F0F1E1E3C3C7878F0F1E1C3C3878F0E1E3C3878F1E1C3C78F0E1C3C78F1E1C3870E1C3C78F1E3C78F1E3C70E1C3870E3C78F1E3870E3C78E1C78F1C38F1E3871E38";
defparam ram_block1a18.mem_init1 = "71E38F1C38F1C78E1C70E3871C38E1C70E3871C78E3871C78E38F1C71E38E3C71C70E38E38F1C71C70E38E38E3871C71C71C71C71C38E38E38E38E38E38E38E38E39C71C71C71C71C718E38E38E39C71C71CE38E38C71C718E38E71C718E38C71C638E71C738E31C738E31C638E71CE39C718E31C638C738E71CE31C639C738C718E718E718E31CE31CE31CE318E718E718C738C639C631CE318E738C639CE718C739CE318C739CE718C6318E739CE739C6318C6318C6318C6318C6318C6318C6739CE739CE6318C6339CE7318C6739CC6319CE6318CE7318CE7318CE7319CE6319CC63398CE7319CC67398CE63398CE63398CE63398CE67319CC663398CC673";
defparam ram_block1a18.mem_init0 = "198CE673198CC673399CC6633198CC6633198CC6633199CCE6733198CCE6633199CCC66733199CCC667333998CCE667333999CCCE6673339998CCC666733319998CCCE666733339999CCCCC666673333399999CCCCCE6666673333339999999CCCCCCCC666666667333333333399999999999999CCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCC9999999999999933333333332666666666CCCCCCCD99999993333336666664CCCCC99999B3333266664CCCC99999333366664CCCD999B3336666CCCD999B3336664CCD9993336664CCD999332666CCD99B332664CC999332664CD99B33664CC99B33664CD99B3266CC9993366";

arriav_ram_block ram_block1a67(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a67_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a67.clk0_core_clock_enable = "ena0";
defparam ram_block1a67.clk0_input_clock_enable = "ena0";
defparam ram_block1a67.clk0_output_clock_enable = "ena0";
defparam ram_block1a67.data_interleave_offset_in_bits = 1;
defparam ram_block1a67.data_interleave_width_in_bits = 1;
defparam ram_block1a67.init_file = "DDS_48_v1_nco_ii_0_sin.hex";
defparam ram_block1a67.init_file_layout = "port_a";
defparam ram_block1a67.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_c8g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a67.operation_mode = "rom";
defparam ram_block1a67.port_a_address_clear = "none";
defparam ram_block1a67.port_a_address_width = 13;
defparam ram_block1a67.port_a_data_out_clear = "none";
defparam ram_block1a67.port_a_data_out_clock = "clock0";
defparam ram_block1a67.port_a_data_width = 1;
defparam ram_block1a67.port_a_first_address = 32768;
defparam ram_block1a67.port_a_first_bit_number = 3;
defparam ram_block1a67.port_a_last_address = 40959;
defparam ram_block1a67.port_a_logical_ram_depth = 65536;
defparam ram_block1a67.port_a_logical_ram_width = 16;
defparam ram_block1a67.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a67.ram_block_type = "auto";
defparam ram_block1a67.mem_init3 = "0E1C3C78F0E1C3C78F1E1C3870F1E3C78F0E1C3870F1E3C78F1E3C7870E1C3870E1C3870E1C3870E1C3870E1C3870E1C3871E3C78F1E3C70E1C3870E3C78F1E3870E1C78F1E3870E1C78F1C3871E3C70E1C78F1C3871E3C70E3C78E1C78F1C38F1C3871E3871E3871E3871E3871E3871E3871E3871E3871E38F1C38F1C38E1C78E3C70E3871E38F1C38E1C70E3C71E38F1C78E3C70E3871C78E3C71E38F1C78E3871C38E3C71E38E1C70E38F1C70E38F1C70E38F1C70E38E1C71E38E3C71C38E3871C70E38E3C71C78E38F1C71C38E38F1C71C38E38E1C71C78E38E3871C71C38E38E3C71C71C38E38E3871C71C71E38E38E3871C71C71C78E38E38E38F1C71C";
defparam ram_block1a67.mem_init2 = "71C71C78E38E38E38E38E3C71C71C71C71C71C71C78E38E38E38E38E38E38E38E38E38E38E38E38E38E38E38E38E38E38E38E38E38E38E38E38E38E38E38E31C71C71C71C71C71C71CE38E38E38E38E38C71C71C71C71CE38E38E38E39C71C71C71CE38E38E39C71C71C738E38E38C71C71C738E38E39C71C71CE38E38C71C71CE38E38C71C718E38E39C71C638E38C71C718E38E71C71CE38E31C71CE38E71C718E38E71C738E38C71C638E31C718E38C71C638E31C718E38C71CE38E71C638E31C738E39C718E39C718E39C71CE38C71CE38C71CE39C718E39C718E39C738E31C738E71C638C71CE39C718E31C738E71CE38C718E31C638E71CE39C738E71C";
defparam ram_block1a67.mem_init1 = "E38C718E31C638C718E31C638C718E71CE39C738E71CE39C638C718E31CE39C738C718E31CE39C738C718E71CE39C638C738E718E31CE39C638C738C718E71CE31CE39C639C738C738E718E71CE31CE31C639C639C738C738C738E718E718E718E31CE31CE31CE31CE31C639C639C639C639C639C639C639C639C639C639C639C639C639CE31CE31CE31CE31CE318E718E718E718E738C738C738C639C639C631CE31CE318E718E738C738C639C639CE31CE718E718C738C639C639CE31CE718E738C739C639CE318E718C738C639CE31CE718E738C639C631CE718C738C639CE318E718C739C631CE718C739C639CE318E738C639CE318E738C639CE318E738";
defparam ram_block1a67.mem_init0 = "C631CE718C739C631CE718C639CE318E738C631CE718C739CE318E738C631CE718C639CE318C739C6318E738C631CE738C639CE718C639CE718C739CE318C739CE318C739CE318C739C6318E739CE318C739CE318C739CE318C739CE318C639CE718C639CE738C631CE738C6318E739C6318C739CE718C639CE738C631CE739C6318C739CE718C631CE739C6318E739CE318C639CE738C6318E739CE718C631CE739C6318C739CE718C6318E739CE318C639CE739C6318C739CE738C6318E739CE718C631CE739CE318C631CE739C6318C639CE739C6318C739CE738C6318C739CE738C6318E739CE718C6318E739CE718C6318E739CE718C631CE739CE318C6";

arriav_ram_block ram_block1a83(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a83_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a83.clk0_core_clock_enable = "ena0";
defparam ram_block1a83.clk0_input_clock_enable = "ena0";
defparam ram_block1a83.clk0_output_clock_enable = "ena0";
defparam ram_block1a83.data_interleave_offset_in_bits = 1;
defparam ram_block1a83.data_interleave_width_in_bits = 1;
defparam ram_block1a83.init_file = "DDS_48_v1_nco_ii_0_sin.hex";
defparam ram_block1a83.init_file_layout = "port_a";
defparam ram_block1a83.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_c8g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a83.operation_mode = "rom";
defparam ram_block1a83.port_a_address_clear = "none";
defparam ram_block1a83.port_a_address_width = 13;
defparam ram_block1a83.port_a_data_out_clear = "none";
defparam ram_block1a83.port_a_data_out_clock = "clock0";
defparam ram_block1a83.port_a_data_width = 1;
defparam ram_block1a83.port_a_first_address = 40960;
defparam ram_block1a83.port_a_first_bit_number = 3;
defparam ram_block1a83.port_a_last_address = 49151;
defparam ram_block1a83.port_a_logical_ram_depth = 65536;
defparam ram_block1a83.port_a_logical_ram_width = 16;
defparam ram_block1a83.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a83.ram_block_type = "auto";
defparam ram_block1a83.mem_init3 = "0000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000003FFFFFFFFFFFFFFFC00000000000007FFFFFFFFFFFE000000000007FFFFFFFFFF0000000000FFFFFFFFFC000000003FFFFFFFF000000007FFFFFFF00000001FFFFFFF00000007FFFFFF8000000FFFFFFC000001FFFFFF0000007FFFFF800000FFFFFE000003FFFFF000007FFFFE00000FFFFF000007FFFF80000FFFFF00001FFFFC00007FFFE00007FFFE00007FFFC0000FFFF80003FFFE0001FFFF0000FFFF0000FFFF0000FFFE0001FFFC0007FFF0001FFFC0007FFE0007FFF0003FFF0003FFF0003FFF0007FFE000FFF8001FFF000";
defparam ram_block1a83.mem_init2 = "7FFC001FFF000FFF8003FFC001FFE000FFF000FFF000FFF000FFF000FFF001FFE003FFC007FF800FFF001FFC007FF001FFC007FF001FFC007FE003FF801FFC00FFE007FE003FF003FF801FF801FF801FF801FF801FF803FF003FF007FE007FC00FF801FF003FE00FFC01FF003FE00FF803FE00FFC01FF007F803FE00FF803FE01FF007FC03FE00FF007F803FC01FE00FF007F807FC03FC01FE01FE00FF00FF00FF00FF007F807F807F00FF00FF00FF00FF01FE01FE03FC03F807F80FF00FE01FC03F807F00FE01FC03F807F01FE03F807F01FE03F80FE01FC07F01FE03F80FE03F80FE03F80FE03F80FE03F80FE03F81FC07F01FC0FE03F81FC07F03F80FC07F";
defparam ram_block1a83.mem_init1 = "03F80FC07E03F81FC0FE07F03F81FC0FE07F03F81F80FC07E07F03F01F81FC0FC0FE07E07F03F03F81F81F81FC0FC0FC0FC0FE07E07E07E07E07E07E07E07E07E07E07E07C0FC0FC0FC0F81F81F81F83F03F07E07E07C0FC0F81F83F03E07E07C0F81F83F03E07C0FC1F83F03E07C0F81F03E07C0F81F03E07C0F81F07E0FC1F03E07C1F83E07C0F83F07C0F83E07C1F83E0FC1F07E0F83F07C1F03E0F83F07C1F07E0F83E0F81F07C1F07C1F03E0F83E0F83E0F83E0F83E0F83E0F83E0F83E0F83E0F83E1F07C1F07C1F0F83E0F83E1F07C1F0F83E0F87C1F0783E0F87C1F0F83E1F07C3E0F87C1E0F83C1F0F83C1F0F83C1F0F83C1F0F87C1E0F87C3E0F078";
defparam ram_block1a83.mem_init0 = "3E1F0F87C1E0F0783C1E0F07C3E1F0F87C3E1F0F8783C1E0F0783C1E1F0F87C3C1E0F0787C3E1E0F0F87C3C1E1F0F0783C3E1E0F0F8783C3C1E1F0F078783C3E1E1F0F0F8787C3C3E1E1F0F0F078783C3C3E1E1E0F0F0F07878783C3C3C1E1E1E1F0F0F0F0F8787878787C3C3C3C3C3C1E1E1E1E1E1E1E1E1E0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F1E1E1E1E1E1E1E1E1E1C3C3C3C3C3C387878787870F0F0F0E1E1E1E1C3C3C3C78787870F0F0E1E1E1C3C3C787870F0F1E1E1C3C3C787870F0E1E1C3C387878F0F1E1C3C387870F0E1E3C3C7870F0E1E3C387870F1E1C3C7870F1E1C3C7870F1E1C3C7870E1E3C3878F1E1C3C78F0E1C3C78F";

arriav_ram_block ram_block1a99(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a99_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a99.clk0_core_clock_enable = "ena0";
defparam ram_block1a99.clk0_input_clock_enable = "ena0";
defparam ram_block1a99.clk0_output_clock_enable = "ena0";
defparam ram_block1a99.data_interleave_offset_in_bits = 1;
defparam ram_block1a99.data_interleave_width_in_bits = 1;
defparam ram_block1a99.init_file = "DDS_48_v1_nco_ii_0_sin.hex";
defparam ram_block1a99.init_file_layout = "port_a";
defparam ram_block1a99.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_c8g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a99.operation_mode = "rom";
defparam ram_block1a99.port_a_address_clear = "none";
defparam ram_block1a99.port_a_address_width = 13;
defparam ram_block1a99.port_a_data_out_clear = "none";
defparam ram_block1a99.port_a_data_out_clock = "clock0";
defparam ram_block1a99.port_a_data_width = 1;
defparam ram_block1a99.port_a_first_address = 49152;
defparam ram_block1a99.port_a_first_bit_number = 3;
defparam ram_block1a99.port_a_last_address = 57343;
defparam ram_block1a99.port_a_logical_ram_depth = 65536;
defparam ram_block1a99.port_a_logical_ram_width = 16;
defparam ram_block1a99.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a99.ram_block_type = "auto";
defparam ram_block1a99.mem_init3 = "E3C7870E1E3C7870F1E3C3878F0E1C3C7870F1E1C3C7870F1E1C3C7870F1E1C3C3878F0E1E1C3C7878F0E1E1C3C387870F1E1E3C3C387870F0E1E1C3C3C787870F0F1E1E1C3C3C787870F0F0E1E1E1C3C3C3C78787870F0F0F0E1E1E1E1C3C3C3C3C38787878787870F0F0F0F0F0F0F0F0F1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E0F0F0F0F0F0F0F0F0F078787878787C3C3C3C3C3E1E1E1E1F0F0F0F07878783C3C3C1E1E1E0F0F0F878783C3C1E1E1F0F0F8787C3C3E1E1F0F0F8783C3C1E1F0F078783C3E1E0F0F8783C1E1F0F0787C3E1E0F0F87C3C1E0F0787C3E1F0F0783C1E0F0783C3E1F0F87C3E1F0F87C1E0F0783C1E0F07C3E1F0F8";
defparam ram_block1a99.mem_init2 = "3C1E0F87C3E0F07C3E1F0783E1F0783E1F0783E1F0783E0F07C3E0F87C1F0F83E1F07C3E0F83C1F07C3E0F83E1F07C1F0F83E0F83E1F07C1F07C1F0F83E0F83E0F83E0F83E0F83E0F83E0F83E0F83E0F83E0F81F07C1F07C1F03E0F83E0FC1F07C1F83E0F81F07C1F83E0FC1F07E0F83F07C0F83E07C1F83E07C0F83F07C0F81F07E0FC1F03E07C0F81F03E07C0F81F03E07C0F81F83F07E07C0F81F83F03E07C0FC0F81F83F03E07E07C0FC0FC1F81F83F03F03F03E07E07E07E07C0FC0FC0FC0FC0FC0FC0FC0FC0FC0FC0FC0FE07E07E07E07F03F03F03F81F81FC0FC0FE07E07F03F01F81FC0FC07E03F03F81FC0FE07F03F81FC0FE07F03F80FC07E03F81";
defparam ram_block1a99.mem_init1 = "FC07E03F81FC07F03F80FE07F01FC07F03F80FE03F80FE03F80FE03F80FE03F80FE03F80FF01FC07F00FE03F80FF01FC03F80FF01FC03F807F00FE01FC03F807F00FE01FE03FC03F807F80FF00FF01FE01FE01FE01FE01FC03FC03FC01FE01FE01FE01FE00FF00FF007F807FC03FC01FE00FF007F803FC01FE00FF807FC01FF00FF803FE00FF803FC01FF007FE00FF803FE00FF801FF007FE00FF801FF003FE007FC00FFC01FF801FF803FF003FF003FF003FF003FF003FF801FF800FFC00FFE007FF003FF800FFC007FF001FFC007FF001FFC007FF001FFE003FFC007FF800FFF001FFE001FFE001FFE001FFE001FFE000FFF0007FF8003FFE001FFF0007FFC";
defparam ram_block1a99.mem_init0 = "001FFF0003FFE000FFFC001FFF8001FFF8001FFF8001FFFC000FFFC0007FFF0001FFFC0007FFF0000FFFE0001FFFE0001FFFE0001FFFF0000FFFF80003FFFE00007FFFC0000FFFFC0000FFFFC00007FFFF00001FFFFE00003FFFFC00001FFFFE00000FFFFFC00001FFFFF800000FFFFFE000003FFFFFC000001FFFFFF0000007FFFFFE0000003FFFFFFC0000001FFFFFFF00000001FFFFFFFC00000001FFFFFFFF8000000007FFFFFFFFE0000000001FFFFFFFFFFC00000000000FFFFFFFFFFFFC00000000000007FFFFFFFFFFFFFFF80000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000000000000000000000000000";

arriav_ram_block ram_block1a115(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a115_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a115.clk0_core_clock_enable = "ena0";
defparam ram_block1a115.clk0_input_clock_enable = "ena0";
defparam ram_block1a115.clk0_output_clock_enable = "ena0";
defparam ram_block1a115.data_interleave_offset_in_bits = 1;
defparam ram_block1a115.data_interleave_width_in_bits = 1;
defparam ram_block1a115.init_file = "DDS_48_v1_nco_ii_0_sin.hex";
defparam ram_block1a115.init_file_layout = "port_a";
defparam ram_block1a115.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_c8g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a115.operation_mode = "rom";
defparam ram_block1a115.port_a_address_clear = "none";
defparam ram_block1a115.port_a_address_width = 13;
defparam ram_block1a115.port_a_data_out_clear = "none";
defparam ram_block1a115.port_a_data_out_clock = "clock0";
defparam ram_block1a115.port_a_data_width = 1;
defparam ram_block1a115.port_a_first_address = 57344;
defparam ram_block1a115.port_a_first_bit_number = 3;
defparam ram_block1a115.port_a_last_address = 65535;
defparam ram_block1a115.port_a_logical_ram_depth = 65536;
defparam ram_block1a115.port_a_logical_ram_width = 16;
defparam ram_block1a115.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a115.ram_block_type = "auto";
defparam ram_block1a115.mem_init3 = "C6318E739CE718C631CE739CE318C631CE739CE318C631CE739CE318C639CE739C6318C639CE739C6318C739CE738C6318C739CE718C6318E739CE718C631CE739CE318C639CE739C6318C739CE738C6318E739CE318C631CE739C6318C739CE718C631CE739CE318C639CE738C6318E739CE318C739CE718C631CE739C6318C739CE718C639CE738C631CE739C6318C739CE318C639CE718C639CE738C631CE738C6318E739C6318E739C6318E739C6318E739CE318C739C6318E739C6318E739C6318E739C631CE738C631CE738C639CE718C639CE318C739C6318E738C631CE718C639CE318E739C631CE718C639CE318E738C631CE718C739C631CE718C6";
defparam ram_block1a115.mem_init2 = "39CE318E738C639CE318E738C639CE318E738C739C631CE718C739C631CE318E738C639C631CE718C738C639CE31CE718E738C639C631CE318E738C739C639CE31CE718E738C738C639C631CE31CE718E738C738C639C639CE31CE318E718E718C738C738C639C639C639CE31CE31CE31CE318E718E718E718E718E738C738C738C738C738C738C738C738C738C738C738C738C738C718E718E718E718E718E31CE31CE31CE39C639C639C738C738C718E718E71CE31CE39C639C738C738E718E71CE31C639C638C738E718E31CE39C638C738E71CE31C639C738E718E31C639C738E718E31C638C738E71CE39C738E71CE31C638C718E31C638C718E31C638E";
defparam ram_block1a115.mem_init1 = "71CE39C738E71CE38C718E31C638E71CE39C718E31C738E71C638C71CE39C718E39C738E31C738E31C738E71C638E71C638E71C738E31C738E31C738E39C718E38C71CE38E71C638E31C718E38C71C638E31C718E38C71C638E39C71CE38E31C71CE38E71C718E38E71C71CE38E31C71C638E38C71C738E38E31C71C638E38E71C71C638E38E71C71C738E38E39C71C71C638E38E39C71C71C738E38E38E71C71C71C738E38E38E38E71C71C71C71C638E38E38E38E38E71C71C71C71C71C71C718E38E38E38E38E38E38E38E38E38E38E38E38E38E38E38E38E38E38E38E38E38E38E38E38E38E38E38E3C71C71C71C71C71C71C78E38E38E38E38E3C71C71C";
defparam ram_block1a115.mem_init0 = "71C71E38E38E38E3C71C71C71C38E38E38F1C71C71C38E38E3871C71C78E38E3871C71C38E38E3C71C70E38E3871C71E38E3871C71E38E3C71C78E38E1C71C38E3871C78E38F1C70E38E1C71E38E1C71E38E1C71E38E1C70E38F1C78E3871C38E3C71E38F1C78E3C71C38E1C78E3C71E38F1C78E1C70E3871E38F1C38E1C78E3C70E3871E3871E38F1C38F1C38F1C38F1C38F1C38F1C38F1C38F1C38F1C3871E3871E3C70E3C78E1C78F1C3871E3C70E1C78F1C3871E3C70E1C38F1E3C70E1C38F1E3C78E1C3870E1C78F1E3C78F1C3870E1C3870E1C3870E1C3870E1C3870E1C3870E1C3C78F1E3C78F1E1C3870E1E3C78F1E1C3870F1E3C7870E1E3C7870E1";

arriav_ram_block ram_block1a35(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a35_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a35.clk0_core_clock_enable = "ena0";
defparam ram_block1a35.clk0_input_clock_enable = "ena0";
defparam ram_block1a35.clk0_output_clock_enable = "ena0";
defparam ram_block1a35.data_interleave_offset_in_bits = 1;
defparam ram_block1a35.data_interleave_width_in_bits = 1;
defparam ram_block1a35.init_file = "DDS_48_v1_nco_ii_0_sin.hex";
defparam ram_block1a35.init_file_layout = "port_a";
defparam ram_block1a35.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_c8g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a35.operation_mode = "rom";
defparam ram_block1a35.port_a_address_clear = "none";
defparam ram_block1a35.port_a_address_width = 13;
defparam ram_block1a35.port_a_data_out_clear = "none";
defparam ram_block1a35.port_a_data_out_clock = "clock0";
defparam ram_block1a35.port_a_data_width = 1;
defparam ram_block1a35.port_a_first_address = 16384;
defparam ram_block1a35.port_a_first_bit_number = 3;
defparam ram_block1a35.port_a_last_address = 24575;
defparam ram_block1a35.port_a_logical_ram_depth = 65536;
defparam ram_block1a35.port_a_logical_ram_width = 16;
defparam ram_block1a35.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a35.ram_block_type = "auto";
defparam ram_block1a35.mem_init3 = "3C78F0E1E3C7870F1E3C3878F1E1C3C7870F1E3C3878F0E1E3C387870F1E1C3C7870F0E1E3C3C7870F0E1E3C3C7878F0F1E1E3C3C7878F0F1E1E3C3C387870F0F1E1E1C3C3C787878F0F0E1E1E1C3C3C3C787878F0F0F0F1E1E1E1E3C3C3C3C387878787878F0F0F0F0F0F0F1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1F0F0F0F0F0F0F0F8787878787C3C3C3C3C1E1E1E1F0F0F0F07878783C3C3C1E1E1F0F0F078787C3C3C1E1E0F0F078783C3C1E1E0F0F0787C3C3E1E0F0F8783C3E1E0F0F8783C3E1E0F0787C3C1E0F0F87C3C1E0F0F87C3E1E0F0783C1E0F0F87C3E1F0F87C3E1F0F87C3E0F0783C1E0F07C3E1F0F";
defparam ram_block1a35.mem_init2 = "83C1E0F87C3E0F07C3E1F0783E1F0783E1F0783E1F07C3E0F07C1E0F87C1F0F83E0F07C1E0F83E1F07C1E0F83E0F07C1F07C3E0F83E0F87C1F07C1F07C1F07C3E0F83E0F83E0F83E0F83E0F83E0F83F07C1F07C1F07C1F03E0F83E0F81F07C1F03E0F83E07C1F07E0F83F07C1F83E0FC1F03E0F81F07E0F81F07E0FC1F03E0FC1F83F07C0F81F03E07C1F83F07E0FC0F81F03E07C0F81F83F07E07C0FC1F83F03E07E0FC0FC1F81F03F03E07E07E0FC0FC0F81F81F81F03F03F03F03F03F07E07E07E07E07E07E07E07E07F03F03F03F03F03F81F81F81FC0FC0FE07E07E03F03F81F80FC0FE07E03F03F81FC0FC07E03F01F80FC07E03F01FC0FE07F01F80FC";
defparam ram_block1a35.mem_init1 = "07F03F80FE07F01FC0FE03F81FC07F01FC07E03F80FE03F80FE03F80FE03F80FE03F80FF01FC07F01FE03F80FF01FC07F80FE01FC07F80FF01FE03FC07F80FF01FE03FC03F807F80FF00FE01FE01FC03FC03FC03FC03FC07F807F807FC03FC03FC03FC03FE01FE01FF00FF007F807FC03FE01FF00FF807FC03FE00FF007FC03FE00FF803FE01FF007FC01FF007FC00FF803FE00FFC01FF007FE00FFC01FF803FF007FE00FFC00FFC01FF801FF801FF801FF801FF801FF801FFC00FFC007FE003FF001FF800FFC007FF001FFC00FFE003FF800FFF001FFC007FF800FFF001FFE003FFC003FFC007FF8007FF8007FFC003FFC001FFE000FFF0007FFC001FFE000F";
defparam ram_block1a35.mem_init0 = "FF8001FFF0007FFE000FFFC001FFF8001FFF8001FFF8000FFFC0007FFE0003FFF8000FFFE0003FFFC0007FFF80007FFF80007FFF80003FFFC0001FFFF00007FFFC0000FFFFC0000FFFFC0000FFFFE00003FFFF80000FFFFF00000FFFFF000007FFFFC00001FFFFF800001FFFFF800000FFFFFE000001FFFFFE000000FFFFFFC000000FFFFFFE0000001FFFFFFE0000000FFFFFFFE00000003FFFFFFFE000000007FFFFFFFF8000000003FFFFFFFFFC0000000000FFFFFFFFFFFC000000000001FFFFFFFFFFFFFC000000000000000FFFFFFFFFFFFFFFFFFE000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

arriav_ram_block ram_block1a51(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a51_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a51.clk0_core_clock_enable = "ena0";
defparam ram_block1a51.clk0_input_clock_enable = "ena0";
defparam ram_block1a51.clk0_output_clock_enable = "ena0";
defparam ram_block1a51.data_interleave_offset_in_bits = 1;
defparam ram_block1a51.data_interleave_width_in_bits = 1;
defparam ram_block1a51.init_file = "DDS_48_v1_nco_ii_0_sin.hex";
defparam ram_block1a51.init_file_layout = "port_a";
defparam ram_block1a51.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_c8g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a51.operation_mode = "rom";
defparam ram_block1a51.port_a_address_clear = "none";
defparam ram_block1a51.port_a_address_width = 13;
defparam ram_block1a51.port_a_data_out_clear = "none";
defparam ram_block1a51.port_a_data_out_clock = "clock0";
defparam ram_block1a51.port_a_data_width = 1;
defparam ram_block1a51.port_a_first_address = 24576;
defparam ram_block1a51.port_a_first_bit_number = 3;
defparam ram_block1a51.port_a_last_address = 32767;
defparam ram_block1a51.port_a_logical_ram_depth = 65536;
defparam ram_block1a51.port_a_logical_ram_width = 16;
defparam ram_block1a51.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a51.ram_block_type = "auto";
defparam ram_block1a51.mem_init3 = "31CE739CE318C631CE739CE318C631CE739CE318C639CE739C6318C639CE739C6318C639CE738C6318C739CE738C6318E739CE718C6318E739CE318C631CE739C6318C639CE738C6318C739CE718C6318E739CE318C639CE739C6318C739CE718C631CE739C6318C739CE718C631CE739C6318C739CE718C631CE739C6318C739CE318C639CE738C631CE739C6318C739CE318C639CE718C639CE738C631CE739C6318E739C6318E739C6318C739CE318C739CE318C739CE318C739CE318C739C6318E739C6318E739C631CE738C631CE718C639CE718C739CE318E739C631CE738C639CE318C739C6318E738C639CE318C739C631CE718C639CE318E738C639";
defparam ram_block1a51.mem_init2 = "CE318E738C639CE318E738C639CE318E738C639CE318E738C639C631CE718C739C639CE318E738C739C631CE318E738C739C639CE318E718C738C639C631CE318E718C738C639C631CE318E718E738C738C639C631CE31CE718E718E738C738C739C639C639CE31CE31CE318E718E718E718C738C738C738C738C739C639C639C639C639C639C639C639C639C639C639C639C639C638C738C738C738C738C718E718E718E718E31CE31CE31C639C639C738C738E718E718E31CE31C639C638C738E718E71CE31C639C738C718E71CE31C639C738C718E31CE39C638C718E71CE39C638C718E31CE39C738E71CE31C638C718E31C638C718E31C638C718E31C63";
defparam ram_block1a51.mem_init1 = "8C718E31C738E71CE39C718E31C638E71CE39C718E31C738E71C638C71CE39C718E39C738E31C738E31C738E31C738E31C738E31C738E31C738E39C718E39C71CE38C71C638E71C738E39C71CE38E71C738E39C71CE38E71C738E38C71C638E39C71C638E39C71C638E39C71C638E38C71C718E38E31C71C638E38C71C71CE38E38C71C71CE38E38C71C71C638E38E39C71C71C638E38E39C71C71C718E38E38E39C71C71C71C638E38E38E38C71C71C71C71C738E38E38E38E38E38E31C71C71C71C71C71C71C71C71C71CE38E38E38E38E38E38E38E38E38E38E38E38E38E38F1C71C71C71C71C71C71C71C71C71E38E38E38E38E38E3871C71C71C71C70E3";
defparam ram_block1a51.mem_init0 = "8E38E38E3871C71C71C78E38E38E3C71C71C70E38E38E3C71C71C38E38E3871C71C38E38E3C71C71E38E3871C71C38E38F1C71C38E3871C71E38E3C71C78E38F1C71E38E1C71C38E3C71C78E3871C78E3871C78E3871C78E3C71C38E1C71E38F1C78E3871C38E1C70E3871C38E1C70E3871C38F1C78E3C70E3871E38F1C38E1C78E3C70E3C71E3871E3871E3871C38F1C38F1C38F1C38F1E3871E3871E3870E3C70E3C78E1C78F1C38F1E3870E3C78E1C38F1E3870E3C78E1C3871E3C78E1C3871E3C78F1C3870E1C38F1E3C78F1E3C70E1C3870E1C3870E1C3870E1C3870E1C3870E1C3C78F1E3C78F1E1C3870E1E3C78F1E1C3870F1E3C7870E1E3C78F0E1C";

arriav_ram_block ram_block1a3(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a3_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.clk0_input_clock_enable = "ena0";
defparam ram_block1a3.clk0_output_clock_enable = "ena0";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.init_file = "DDS_48_v1_nco_ii_0_sin.hex";
defparam ram_block1a3.init_file_layout = "port_a";
defparam ram_block1a3.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_c8g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.operation_mode = "rom";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 13;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "clock0";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 8191;
defparam ram_block1a3.port_a_logical_ram_depth = 65536;
defparam ram_block1a3.port_a_logical_ram_width = 16;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.ram_block_type = "auto";
defparam ram_block1a3.mem_init3 = "70E1E3C78F0E1C3C78F1E1C3870F1E3C78F0E1C3870F1E3C78F1E3C7870E1C3870E1C3870E1C3870E1C3870E1C3870E1C78F1E3C78F1E3870E1C3871E3C78F1C3870E3C78F1C3870E3C78E1C38F1E3870E3C78E1C38F1E3871E3C70E3C78E1C78E1C38F1C38F1C38F1E3871E3871E3871E3871C38F1C38F1C38F1C78E1C78E3C70E3871E38F1C38E1C78E3C71E3871C38E1C70E3871C38E1C70E3871C38E3C71E38F1C70E3871C78E3C71C38E3C71C38E3C71C38E3C71C78E3871C70E38F1C71E38E3C71C78E38F1C71C38E3871C71E38E3871C71C38E38F1C71C78E38E3871C71C38E38E3871C71C78E38E38E1C71C71C78E38E38E3C71C71C71C38E38E38E3";
defparam ram_block1a3.mem_init2 = "8E1C71C71C71C71C38E38E38E38E38E38F1C71C71C71C71C71C71C71C71C71E38E38E38E38E38E38E38E38E38E38E38E38E38E38E71C71C71C71C71C71C71C71C71C718E38E38E38E38E38E39C71C71C71C71C638E38E38E38C71C71C71C738E38E38E31C71C71C738E38E38C71C71C738E38E38C71C71C638E38E71C71C638E38E71C71C638E38C71C718E38E31C71C638E38C71C738E38C71C738E38C71C738E38C71C638E39C71CE38E71C738E39C71CE38E71C738E39C71CE38C71C638E71C738E31C738E39C718E39C718E39C718E39C718E39C718E39C718E39C738E31C738E71C638C71CE39C718E31C738E71CE38C718E31C738E71CE39C718E31C63";
defparam ram_block1a3.mem_init1 = "8C718E31C638C718E31C638C718E31C638C718E71CE39C738E718E31C638C738E71CE31C638C738E718E31C639C738C718E71CE31C639C738C718E71CE31CE39C638C738C718E718E31CE31CE39C639C738C738C718E718E718E31CE31CE31CE31C639C639C639C639C638C738C738C738C738C738C738C738C738C738C738C738C738C739C639C639C639C639C631CE31CE31CE318E718E718E738C738C739C639C639CE31CE31CE718E718C738C639C639CE31CE318E718C738C639C631CE318E718C738C639C631CE318E738C739C639CE318E718C739C639CE318E738C739C631CE718C738C639CE318E738C639CE318E738C639CE318E738C639CE318E7";
defparam ram_block1a3.mem_init0 = "38C639CE318E738C631CE718C739C6318E738C639CE318C739C6318E738C639CE718C739CE318E739C631CE738C631CE718C639CE718C739CE318C739CE318C739C6318E739C6318E739C6318E739C6318E739C6318C739CE318C739CE318C739CE718C639CE738C631CE738C6318E739C6318C739CE718C639CE738C6318E739C6318C739CE718C631CE739C6318C739CE718C631CE739C6318C739CE718C631CE739C6318C739CE738C6318E739CE318C631CE739C6318C639CE738C6318C739CE718C6318E739CE318C631CE739CE318C639CE739C6318C639CE738C6318C739CE738C6318C739CE738C6318E739CE718C6318E739CE718C6318E739CE718";

arriav_ram_block ram_block1a19(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a19_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a19.clk0_core_clock_enable = "ena0";
defparam ram_block1a19.clk0_input_clock_enable = "ena0";
defparam ram_block1a19.clk0_output_clock_enable = "ena0";
defparam ram_block1a19.data_interleave_offset_in_bits = 1;
defparam ram_block1a19.data_interleave_width_in_bits = 1;
defparam ram_block1a19.init_file = "DDS_48_v1_nco_ii_0_sin.hex";
defparam ram_block1a19.init_file_layout = "port_a";
defparam ram_block1a19.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_c8g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a19.operation_mode = "rom";
defparam ram_block1a19.port_a_address_clear = "none";
defparam ram_block1a19.port_a_address_width = 13;
defparam ram_block1a19.port_a_data_out_clear = "none";
defparam ram_block1a19.port_a_data_out_clock = "clock0";
defparam ram_block1a19.port_a_data_width = 1;
defparam ram_block1a19.port_a_first_address = 8192;
defparam ram_block1a19.port_a_first_bit_number = 3;
defparam ram_block1a19.port_a_last_address = 16383;
defparam ram_block1a19.port_a_logical_ram_depth = 65536;
defparam ram_block1a19.port_a_logical_ram_width = 16;
defparam ram_block1a19.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a19.ram_block_type = "auto";
defparam ram_block1a19.mem_init3 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000FFFFFFFFFFFFFFFFFFE0000000000000007FFFFFFFFFFFFF0000000000007FFFFFFFFFFE00000000007FFFFFFFFF8000000003FFFFFFFFC00000000FFFFFFFF80000000FFFFFFFE0000000FFFFFFF0000000FFFFFFE0000007FFFFFE000000FFFFFF000000FFFFFE000003FFFFF000003FFFFF000007FFFFC00001FFFFE00001FFFFE00003FFFF80000FFFFE00007FFFE00007FFFE00007FFFC0001FFFF00007FFF80003FFFC0003FFFC0003FFFC0007FFF8000FFFE0003FFF8000FFFC0007FFE0003FFF0003FFF0003FFF0007FFE000FFFC001FFF0003FF";
defparam ram_block1a19.mem_init2 = "E000FFF0007FFC001FFE000FFF0007FF8007FFC003FFC003FFC007FF8007FF800FFF001FFE003FFC007FF001FFE003FF800FFE007FF001FFC007FE003FF001FF800FFC007FE007FF003FF003FF003FF003FF003FF003FF007FE007FE00FFC01FF803FF007FE00FFC01FF007FE00FF803FE007FC01FF007FC01FF00FF803FE00FF807FC01FE00FF807FC03FE01FF00FF807FC03FC01FE01FF00FF00FF807F807F807F807FC03FC03FC07F807F807F807F807F00FF00FE01FE03FC03F807F80FF01FE03FC07F80FF01FE03FC07F00FE03FC07F01FE03F80FF01FC07F01FE03F80FE03F80FE03F80FE03F80FE03F80FC07F01FC07F03F80FE07F01FC0FE03F81FC0";
defparam ram_block1a19.mem_init1 = "7E03F01FC0FE07F01F80FC07E03F01F80FC07E07F03F81F80FC0FE07E03F03F81F80FC0FC0FE07E07F03F03F03F81F81F81F81F81FC0FC0FC0FC0FC0FC0FC0FC0FC1F81F81F81F81F81F03F03F03E07E07E0FC0FC0F81F81F03F07E07E0FC0F81F83F07E07C0FC1F83F03E07C0F81F03E07E0FC1F83F07C0F81F03E07C1F83F07E0F81F07E0FC1F03E0FC1F03E0F81F07E0F83F07C1F83E0FC1F07C0F83E0F81F07C1F03E0F83E0F81F07C1F07C1F07C1F83E0F83E0F83E0F83E0F83E0F83E0F87C1F07C1F07C1F07C3E0F83E0F87C1F07C1E0F83E0F07C1F0F83E0F07C1E0F83E1F07C3E0F07C1E0F87C1F0F83C1F0F83C1F0F83C1F0F87C1E0F87C3E0F0783";
defparam ram_block1a19.mem_init0 = "E1F0F87C1E0F0783C1E0F87C3E1F0F87C3E1F0F87C3E1E0F0783C1E0F0F87C3E1E0F0787C3E1E0F0787C3C1E0F0F8783C3E1E0F0F8783C3E1E0F0F8787C3C1E1E0F0F078783C3C1E1E0F0F078787C3C3C1E1E1F0F0F07878783C3C3C1E1E1E1F0F0F0F0787878787C3C3C3C3C3E1E1E1E1E1E1E1F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F1E1E1E1E1E1E1E3C3C3C3C3C3878787878F0F0F0F1E1E1E1E3C3C3C78787870F0F0E1E1E3C3C3C787870F0F1E1E1C3C387878F0F1E1E3C3C7878F0F1E1E3C3C7878F0E1E1C3C7878F0E1E1C3C7870F1E1C3C3878F0E1E3C3878F1E1C3C7870F1E3C3878F1E1C3C78F0E1E3C78";

arriav_ram_block ram_block1a68(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a68_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a68.clk0_core_clock_enable = "ena0";
defparam ram_block1a68.clk0_input_clock_enable = "ena0";
defparam ram_block1a68.clk0_output_clock_enable = "ena0";
defparam ram_block1a68.data_interleave_offset_in_bits = 1;
defparam ram_block1a68.data_interleave_width_in_bits = 1;
defparam ram_block1a68.init_file = "DDS_48_v1_nco_ii_0_sin.hex";
defparam ram_block1a68.init_file_layout = "port_a";
defparam ram_block1a68.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_c8g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a68.operation_mode = "rom";
defparam ram_block1a68.port_a_address_clear = "none";
defparam ram_block1a68.port_a_address_width = 13;
defparam ram_block1a68.port_a_data_out_clear = "none";
defparam ram_block1a68.port_a_data_out_clock = "clock0";
defparam ram_block1a68.port_a_data_width = 1;
defparam ram_block1a68.port_a_first_address = 32768;
defparam ram_block1a68.port_a_first_bit_number = 4;
defparam ram_block1a68.port_a_last_address = 40959;
defparam ram_block1a68.port_a_logical_ram_depth = 65536;
defparam ram_block1a68.port_a_logical_ram_width = 16;
defparam ram_block1a68.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a68.ram_block_type = "auto";
defparam ram_block1a68.mem_init3 = "01FC03F80FE03FC07F01FC07F00FE03F80FE03F80FF01FC07F01FC07F01FC07F01FC07F01FC07F01FC07F01FC07F01FC07F01FC07F01FC0FE03F80FE03F80FE07F01FC07F01F80FE03F80FC07F01FC0FE03F80FC07F01FC0FE03F81FC07F03F80FC07F01F80FE07F01F80FE07F01F80FE07F01F80FE07F01F80FC07F03F81FC07E03F01F80FE07F03F81FC0FE03F01F80FC07E03F01F80FC07E03F01F80FC07E07F03F81FC0FE07E03F01F80FC0FE07F03F01F80FC0FE07E03F01F81FC0FC07E07F03F01F81FC0FC07E07F03F03F81F80FC0FC07E07E03F03F81F81F80FC0FC07E07E03F03F03F81F81F80FC0FC0FE07E07E07F03F03F03F81F81F81F80FC0FC";
defparam ram_block1a68.mem_init2 = "0FC0FC07E07E07E07E07E03F03F03F03F03F03F03F81F81F81F81F81F81F81F81F81F81F81F81F81F81F81F81F81F81F81F81F81F81F81F81F81F81F81F81F03F03F03F03F03F03F03E07E07E07E07E07C0FC0FC0FC0FC1F81F81F81F83F03F03F03E07E07E07C0FC0FC0F81F81F83F03F03F07E07E07C0FC0FC1F81F83F03F03E07E07C0FC0F81F81F83F03E07E07C0FC0F81F81F03F03E07E0FC0FC1F81F03F07E07E0FC0F81F83F03E07E0FC0F81F83F03E07E0FC0F81F83F03E07E0FC1F81F03F07E07C0F81F83F07E07C0FC1F83F03E07C0FC1F83F07E07C0F81F83F07E0FC0F81F03E07C0FC1F83F07E0FC0F81F03E07C0F81F03E07E0FC1F83F07E0FC";
defparam ram_block1a68.mem_init1 = "1F83F07E0FC1F83F07E0FC1F83F07E0FC1F83F07E0FC1F83E07C0F81F03E07C0F83F07E0FC1F83F07C0F81F03E07C1F83F07E0F81F03E07C1F83F07C0F81F03E0FC1F83E07C0F83F07E0F81F03E0FC1F03E07C1F83F07C0F83F07E0F81F07E0F81F03E0FC1F03E0FC1F03E07C1F83E07C1F83E07C1F83E07C1F83E07C1F83E07C1F83E07C1F03E0FC1F03E0FC1F07E0F81F07E0F81F07C0F83F07C1F83E07C1F03E0FC1F07E0F81F07C0F83E07C1F83E0FC1F07E0F83F07C1F83E07C1F03E0F81F07C0F83E07C1F07E0F83F07C1F83E0FC1F07E0F83E07C1F03E0F83F07C1F83E0F81F07C0F83E0FC1F07C0F83E07C1F07E0F83E07C1F07E0F83E07C1F07E0F8";
defparam ram_block1a68.mem_init0 = "3E0FC1F07C0F83E0FC1F07C1F83E0F81F07C1F03E0F83F07C1F07E0F83E0FC1F07C1F83E0F83F07C1F07E0F83E0FC1F07C1F83E0F83E07C1F07C0F83E0F83F07C1F07C0F83E0F83F07C1F07E0F83E0F83F07C1F07C0F83E0F83F07C1F07C1F83E0F83E07C1F07C1F03E0F83E0F81F07C1F07C0F83E0F83E07C1F07C1F03E0F83E0F83F07C1F07C1F03E0F83E0F81F07C1F07C1F83E0F83E0F81F07C1F07C1F03E0F83E0F83F07C1F07C1F07E0F83E0F83E07C1F07C1F07C0F83E0F83E0F81F07C1F07C1F03E0F83E0F83E0FC1F07C1F07C1F83E0F83E0F83F07C1F07C1F07C0F83E0F83E0F81F07C1F07C1F07E0F83E0F83E0F81F07C1F07C1F03E0F83E0F83E";

arriav_ram_block ram_block1a84(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a84_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a84.clk0_core_clock_enable = "ena0";
defparam ram_block1a84.clk0_input_clock_enable = "ena0";
defparam ram_block1a84.clk0_output_clock_enable = "ena0";
defparam ram_block1a84.data_interleave_offset_in_bits = 1;
defparam ram_block1a84.data_interleave_width_in_bits = 1;
defparam ram_block1a84.init_file = "DDS_48_v1_nco_ii_0_sin.hex";
defparam ram_block1a84.init_file_layout = "port_a";
defparam ram_block1a84.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_c8g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a84.operation_mode = "rom";
defparam ram_block1a84.port_a_address_clear = "none";
defparam ram_block1a84.port_a_address_width = 13;
defparam ram_block1a84.port_a_data_out_clear = "none";
defparam ram_block1a84.port_a_data_out_clock = "clock0";
defparam ram_block1a84.port_a_data_width = 1;
defparam ram_block1a84.port_a_first_address = 40960;
defparam ram_block1a84.port_a_first_bit_number = 4;
defparam ram_block1a84.port_a_last_address = 49151;
defparam ram_block1a84.port_a_logical_ram_depth = 65536;
defparam ram_block1a84.port_a_logical_ram_width = 16;
defparam ram_block1a84.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a84.ram_block_type = "auto";
defparam ram_block1a84.mem_init3 = "000000000000000000000000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000001FFFFFFFFFFFFFFFFFFFFFF00000000000000000003FFFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFF000000000000007FFFFFFFFFFFFC000000000000FFFFFFFFFFFF800000000001FFFFFFFFFFF00000000001FFFFFFFFFF00000000007FFFFFFFFF0000000003FFFFFFFFE000000001FFFFFFFFC000000007FFFFFFFE00000000FFFFFFFF00000000FFFFFFFE00000003FFFFFFF00000003FFFFFFE0000000FFFFFFF0000000FFFFFFF0000001FFFFFF8000000FFF";
defparam ram_block1a84.mem_init2 = "FFFC000000FFFFFF8000003FFFFFE000000FFFFFF000000FFFFFF000000FFFFFE000003FFFFF800000FFFFFC00000FFFFFC00000FFFFFC00001FFFFF800003FFFFE00001FFFFF000007FFFF800007FFFF800007FFFF80000FFFFF00001FFFFC00007FFFF00001FFFFC0000FFFFE00007FFFE00003FFFF00007FFFE00007FFFE0000FFFFC0001FFFF00007FFFC0001FFFF00007FFFC0003FFFE0001FFFF0000FFFF0000FFFF80007FFF0000FFFF0000FFFF0001FFFE0003FFF80007FFF0001FFFC0007FFF0001FFFC0007FFF0001FFF8000FFFE0007FFE0003FFF0001FFF8001FFF8001FFF8001FFF8001FFF8001FFF8003FFF0003FFE0007FFC000FFF8003FFF";
defparam ram_block1a84.mem_init1 = "0007FFC001FFF8003FFE000FFF8003FFE000FFF8007FFC001FFF000FFF8003FFC001FFE000FFF0007FF8007FFC003FFC003FFE001FFE001FFE001FFE001FFE001FFE001FFC003FFC003FF8007FF8007FF000FFE001FFC003FF8007FF001FFE003FF8007FF001FFC003FF800FFE003FF800FFE003FF800FFE003FF800FFE003FF001FFC007FE003FF800FFC007FE003FF801FFC00FFE007FF003FF001FF800FFC00FFE007FE007FF003FF003FF001FF801FF801FF801FF801FF801FF801FF801FF801FF801FF003FF003FF007FE007FE00FFC00FF801FF803FF007FE007FC00FF801FF003FE007FC01FF803FF007FC00FF803FF007FC00FF803FE007FC01FF007";
defparam ram_block1a84.mem_init0 = "FE00FF803FE00FF803FE00FFC01FF007FC01FF007F803FE00FF803FE00FF803FC01FF007FC01FE00FF803FC01FF00FF803FE01FF007F803FC01FF00FF807FC01FE00FF007F803FC01FE00FF00FF807FC03FE01FE00FF00FF807F803FC03FE01FE00FF00FF007F807F807FC03FC03FC03FE01FE01FE01FE01FE00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FE01FE01FE01FE01FE03FC03FC03FC07F807F807F00FF00FE01FE01FC03FC03F807F80FF00FE01FE03FC03F807F00FF01FE03FC03F807F00FE01FC03F807F80FF01FC03F807F00FE01FC03F80FF01FE03F807F00FE03FC07F00FE03FC07F00FE03FC07F01FE03F807F01FC03F80FE03FC07F";

arriav_ram_block ram_block1a100(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a100_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a100.clk0_core_clock_enable = "ena0";
defparam ram_block1a100.clk0_input_clock_enable = "ena0";
defparam ram_block1a100.clk0_output_clock_enable = "ena0";
defparam ram_block1a100.data_interleave_offset_in_bits = 1;
defparam ram_block1a100.data_interleave_width_in_bits = 1;
defparam ram_block1a100.init_file = "DDS_48_v1_nco_ii_0_sin.hex";
defparam ram_block1a100.init_file_layout = "port_a";
defparam ram_block1a100.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_c8g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a100.operation_mode = "rom";
defparam ram_block1a100.port_a_address_clear = "none";
defparam ram_block1a100.port_a_address_width = 13;
defparam ram_block1a100.port_a_data_out_clear = "none";
defparam ram_block1a100.port_a_data_out_clock = "clock0";
defparam ram_block1a100.port_a_data_width = 1;
defparam ram_block1a100.port_a_first_address = 49152;
defparam ram_block1a100.port_a_first_bit_number = 4;
defparam ram_block1a100.port_a_last_address = 57343;
defparam ram_block1a100.port_a_logical_ram_depth = 65536;
defparam ram_block1a100.port_a_logical_ram_width = 16;
defparam ram_block1a100.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a100.ram_block_type = "auto";
defparam ram_block1a100.mem_init3 = "FC07F80FE03F807F01FC03F80FF01FC07F80FE01FC07F80FE01FC07F80FE01FC03F80FF01FE03F807F00FE01FC03F807F01FE03FC03F807F00FE01FC03F807F80FF01FE01FC03F807F80FF00FE01FE03FC03F807F807F00FF00FE01FE01FC03FC03FC07F807F807F80FF00FF00FF00FF00FE01FE01FE01FE01FE01FE01FE01FE01FE01FE01FE00FF00FF00FF00FF00FF807F807F807FC03FC03FC01FE01FE00FF00FF807F803FC03FE01FE00FF00FF807FC03FE01FE00FF007F803FC01FE00FF007FC03FE01FF007F803FC01FF00FF803FE01FF007F803FE00FF007FC01FF007F803FE00FF803FE00FF803FC01FF007FC01FF007FE00FF803FE00FF803FE00FF";
defparam ram_block1a100.mem_init2 = "C01FF007FC00FF803FE007FC01FF803FE007FC01FF803FF007FC00FF801FF003FE007FC00FFC01FF803FF003FE007FE00FFC00FFC01FF801FF801FF003FF003FF003FF003FF003FF003FF003FF003FF003FF001FF801FF801FFC00FFC00FFE007FE003FF001FF801FFC00FFE007FF003FF800FFC007FE003FF800FFC007FF001FF800FFE003FF800FFE003FF800FFE003FF800FFE003FF8007FF001FFC003FF800FFF001FFC003FF8007FF000FFE001FFC003FFC003FF8007FF8007FF000FFF000FFF000FFF000FFF000FFF000FFF8007FF8007FFC003FFC001FFE000FFF0007FF8003FFE001FFF0007FFC003FFE000FFF8003FFE000FFF8003FFF0007FFC001";
defparam ram_block1a100.mem_init1 = "FFF8003FFE0007FFC000FFF8001FFF8003FFF0003FFF0003FFF0003FFF0003FFF0003FFF0001FFF8000FFFC000FFFE0003FFF0001FFFC0007FFF0001FFFC0007FFF0001FFFC0003FFF8000FFFF0001FFFE0001FFFE0001FFFC0003FFFE0001FFFE0001FFFF0000FFFF80007FFFC0001FFFF00007FFFC0001FFFF00007FFFE0000FFFFC0000FFFFC0001FFFF80000FFFFC0000FFFFE00007FFFF00001FFFFC00007FFFF00001FFFFE00003FFFFC00003FFFFC00003FFFFC00001FFFFF00000FFFFF800003FFFFF000007FFFFE000007FFFFE000007FFFFE000003FFFFF800000FFFFFE000001FFFFFE000001FFFFFE000000FFFFFF8000003FFFFFE0000007FFF";
defparam ram_block1a100.mem_init0 = "FFE0000003FFFFFF0000001FFFFFFE0000001FFFFFFE0000000FFFFFFF80000001FFFFFFF80000000FFFFFFFE00000001FFFFFFFE00000000FFFFFFFFC000000007FFFFFFFF000000000FFFFFFFFF8000000001FFFFFFFFFC0000000001FFFFFFFFFF00000000001FFFFFFFFFFF000000000003FFFFFFFFFFFE0000000000007FFFFFFFFFFFFC00000000000001FFFFFFFFFFFFFFE0000000000000001FFFFFFFFFFFFFFFFF80000000000000000001FFFFFFFFFFFFFFFFFFFFFF000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000000000000000000000000000000000000000000000000000";

arriav_ram_block ram_block1a116(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a116_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a116.clk0_core_clock_enable = "ena0";
defparam ram_block1a116.clk0_input_clock_enable = "ena0";
defparam ram_block1a116.clk0_output_clock_enable = "ena0";
defparam ram_block1a116.data_interleave_offset_in_bits = 1;
defparam ram_block1a116.data_interleave_width_in_bits = 1;
defparam ram_block1a116.init_file = "DDS_48_v1_nco_ii_0_sin.hex";
defparam ram_block1a116.init_file_layout = "port_a";
defparam ram_block1a116.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_c8g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a116.operation_mode = "rom";
defparam ram_block1a116.port_a_address_clear = "none";
defparam ram_block1a116.port_a_address_width = 13;
defparam ram_block1a116.port_a_data_out_clear = "none";
defparam ram_block1a116.port_a_data_out_clock = "clock0";
defparam ram_block1a116.port_a_data_width = 1;
defparam ram_block1a116.port_a_first_address = 57344;
defparam ram_block1a116.port_a_first_bit_number = 4;
defparam ram_block1a116.port_a_last_address = 65535;
defparam ram_block1a116.port_a_logical_ram_depth = 65536;
defparam ram_block1a116.port_a_logical_ram_width = 16;
defparam ram_block1a116.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a116.ram_block_type = "auto";
defparam ram_block1a116.mem_init3 = "F83E0F83E0F81F07C1F07C1F03E0F83E0F83E0FC1F07C1F07C1F03E0F83E0F83E07C1F07C1F07C1F83E0F83E0F83F07C1F07C1F07E0F83E0F83E0F81F07C1F07C1F03E0F83E0F83E07C1F07C1F07C0F83E0F83E0FC1F07C1F07C1F83E0F83E0F81F07C1F07C1F03E0F83E0F83F07C1F07C1F03E0F83E0F81F07C1F07C1F83E0F83E0F81F07C1F07C0F83E0F83E07C1F07C1F03E0F83E0F81F07C1F07C0F83E0F83F07C1F07C1F83E0F83E07C1F07C1F83E0F83E0FC1F07C1F83E0F83E07C1F07C1F83E0F83E07C1F07C0F83E0F83F07C1F07E0F83E0FC1F07C1F83E0F83F07C1F07E0F83E0FC1F07C1F83E0F81F07C1F03E0F83F07C1F07E0F83E07C1F07E0F8";
defparam ram_block1a116.mem_init2 = "3E0FC1F07C0F83E0FC1F07C0F83E0FC1F07C0F83E07C1F07E0F83E07C1F03E0F83F07C1F83E0F81F07C0F83E0FC1F07E0F83F07C1F83E0FC1F07C0F83E07C1F03E0F81F07C0F83F07C1F83E0FC1F07E0F83F07C0F83E07C1F03E0FC1F07E0F81F07C0F83F07C1F83E07C1F03E0FC1F03E0FC1F07E0F81F07E0F81F07C0F83F07C0F83F07C0F83F07C0F83F07C0F83F07C0F83F07C0F81F07E0F81F07E0F81F03E0FC1F03E0FC1F83E07C1F83F07C0F81F07E0F81F03E0FC1F83E07C0F83F07E0F81F03E07C1F83F07C0F81F03E0FC1F83F07C0F81F03E07C1F83F07E0FC1F83E07C0F81F03E07C0F83F07E0FC1F83F07E0FC1F83F07E0FC1F83F07E0FC1F83F0";
defparam ram_block1a116.mem_init1 = "7E0FC1F83F07E0FC0F81F03E07C0F81F03E07E0FC1F83F07E07C0F81F03E07E0FC1F83F03E07C0FC1F83F07E07C0F81F83F07E07C0FC1F83F03E07C0FC1F81F03F07E0FC0F81F83F03E07E0FC0F81F83F03E07E0FC0F81F83F03E07E0FC0FC1F81F03F07E07E0FC0F81F81F03F03E07E07C0FC0F81F83F03F03E07E07C0FC0F81F81F83F03F07E07E07C0FC0FC1F81F81F83F03F03E07E07E07C0FC0FC0F81F81F81F83F03F03F03F07E07E07E07E07C0FC0FC0FC0FC0F81F81F81F81F81F81F81F03F03F03F03F03F03F03F03F03F03F03F03F03F03F03F03F03F03F03F03F03F03F03F03F03F03F03F03F81F81F81F81F81F81F80FC0FC0FC0FC0FC07E07E0";
defparam ram_block1a116.mem_init0 = "7E07E03F03F03F03F81F81F81FC0FC0FC0FE07E07E03F03F03F81F81F80FC0FC07E07E03F03F03F81F80FC0FC07E07E03F03F81F81FC0FC07E07F03F01F81FC0FC07E07F03F01F80FC0FE07E03F01F81FC0FE07E03F01F80FC0FE07F03F81FC0FC07E03F01F80FC07E03F01F80FC07E03F01F80FE07F03F81FC0FE03F01F80FC07F03F81FC07E03F01FC0FE03F01FC0FE03F01FC0FE03F01FC0FE03F01FC07E03F81FC07F03F80FE07F01FC07E03F80FE07F01FC07E03F80FE03F01FC07F01FC0FE03F80FE03F80FE07F01FC07F01FC07F01FC07F01FC07F01FC07F01FC07F01FC07F01FC07F01FC07F01FE03F80FE03F80FE01FC07F01FC07F80FE03F807F01";

arriav_ram_block ram_block1a36(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a36_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a36.clk0_core_clock_enable = "ena0";
defparam ram_block1a36.clk0_input_clock_enable = "ena0";
defparam ram_block1a36.clk0_output_clock_enable = "ena0";
defparam ram_block1a36.data_interleave_offset_in_bits = 1;
defparam ram_block1a36.data_interleave_width_in_bits = 1;
defparam ram_block1a36.init_file = "DDS_48_v1_nco_ii_0_sin.hex";
defparam ram_block1a36.init_file_layout = "port_a";
defparam ram_block1a36.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_c8g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a36.operation_mode = "rom";
defparam ram_block1a36.port_a_address_clear = "none";
defparam ram_block1a36.port_a_address_width = 13;
defparam ram_block1a36.port_a_data_out_clear = "none";
defparam ram_block1a36.port_a_data_out_clock = "clock0";
defparam ram_block1a36.port_a_data_width = 1;
defparam ram_block1a36.port_a_first_address = 16384;
defparam ram_block1a36.port_a_first_bit_number = 4;
defparam ram_block1a36.port_a_last_address = 24575;
defparam ram_block1a36.port_a_logical_ram_depth = 65536;
defparam ram_block1a36.port_a_logical_ram_width = 16;
defparam ram_block1a36.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a36.ram_block_type = "auto";
defparam ram_block1a36.mem_init3 = "03F80FE01FC07F00FE03F807F01FC03F80FF01FC07F80FE01FC07F80FF01FC03F80FF01FE03FC07F00FE01FC03F807F00FE01FC03F807F00FE01FC03F807F00FF01FE03FC03F807F80FF01FE01FC03FC03F807F80FF00FF01FE01FE03FC03FC07F807F807F80FF00FF00FF00FE01FE01FE01FE01FE01FE01FE01FE01FE01FE01FE01FE01FE01FE01FE01FE00FF00FF00FF00FF807F807F803FC03FC03FE01FE00FF00FF007F807FC03FC01FE00FF00FF807FC03FC01FE00FF007F803FC01FE00FF007FC03FE01FF007F803FE01FF007F803FE01FF007FC03FE00FF803FC01FF007FC01FE00FF803FE00FF803FE00FF803FE00FF803FE00FF803FE00FFC01FF00";
defparam ram_block1a36.mem_init2 = "7FC01FF803FE00FFC01FF007FE00FF801FF007FE00FFC01FF003FE007FC00FF801FF003FE007FE00FFC01FF801FF003FF003FE007FE007FC00FFC00FFC00FFC01FF801FF801FF801FF801FF801FF800FFC00FFC00FFC00FFE007FE007FF003FF001FF801FFC00FFE007FF003FF801FFC00FFE007FF001FF800FFE003FF001FFC007FF003FF800FFE003FF800FFE003FF800FFE003FF8007FF001FFC003FF800FFE001FFC003FF800FFF001FFE001FFC003FF8007FF800FFF000FFF000FFF001FFE001FFE001FFE001FFE000FFF000FFF000FFF8007FF8003FFC001FFE001FFF0007FF8003FFE001FFF0007FFC003FFE000FFF8003FFE000FFFC001FFF0007FFC";
defparam ram_block1a36.mem_init1 = "000FFF8001FFF0003FFE0007FFC000FFFC001FFF8001FFF8001FFF8001FFF8001FFF8000FFFC000FFFE0007FFF0003FFF8001FFFC0007FFF0001FFFC0007FFF0001FFFC0007FFF8000FFFE0001FFFC0003FFFC0003FFFC0007FFF80003FFFC0003FFFC0001FFFE0000FFFF00007FFFC0001FFFF00007FFFC0001FFFF00003FFFE00007FFFE0000FFFFC0000FFFFC00007FFFE00003FFFF00001FFFFC00007FFFF00001FFFFC00003FFFF800007FFFF800007FFFF800007FFFFC00003FFFFE00000FFFFF800003FFFFF000003FFFFE000007FFFFF000003FFFFF800000FFFFFE000003FFFFFC000007FFFFF8000003FFFFFC000001FFFFFF0000003FFFFFE0000";
defparam ram_block1a36.mem_init0 = "007FFFFFF0000001FFFFFFC0000007FFFFFF80000007FFFFFFC0000001FFFFFFF80000001FFFFFFFC00000007FFFFFFF800000007FFFFFFFC00000000FFFFFFFFC000000003FFFFFFFFC000000001FFFFFFFFF8000000000FFFFFFFFFF00000000003FFFFFFFFFF800000000007FFFFFFFFFFE000000000001FFFFFFFFFFFFC0000000000001FFFFFFFFFFFFFE000000000000001FFFFFFFFFFFFFFFE000000000000000007FFFFFFFFFFFFFFFFFFC0000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

arriav_ram_block ram_block1a52(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a52_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a52.clk0_core_clock_enable = "ena0";
defparam ram_block1a52.clk0_input_clock_enable = "ena0";
defparam ram_block1a52.clk0_output_clock_enable = "ena0";
defparam ram_block1a52.data_interleave_offset_in_bits = 1;
defparam ram_block1a52.data_interleave_width_in_bits = 1;
defparam ram_block1a52.init_file = "DDS_48_v1_nco_ii_0_sin.hex";
defparam ram_block1a52.init_file_layout = "port_a";
defparam ram_block1a52.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_c8g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a52.operation_mode = "rom";
defparam ram_block1a52.port_a_address_clear = "none";
defparam ram_block1a52.port_a_address_width = 13;
defparam ram_block1a52.port_a_data_out_clear = "none";
defparam ram_block1a52.port_a_data_out_clock = "clock0";
defparam ram_block1a52.port_a_data_width = 1;
defparam ram_block1a52.port_a_first_address = 24576;
defparam ram_block1a52.port_a_first_bit_number = 4;
defparam ram_block1a52.port_a_last_address = 32767;
defparam ram_block1a52.port_a_logical_ram_depth = 65536;
defparam ram_block1a52.port_a_logical_ram_width = 16;
defparam ram_block1a52.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a52.ram_block_type = "auto";
defparam ram_block1a52.mem_init3 = "0FC1F07C1F07C1F03E0F83E0F83E0FC1F07C1F07C1F83E0F83E0F83E07C1F07C1F07C1F83E0F83E0F83F07C1F07C1F07E0F83E0F83E0F81F07C1F07C1F03E0F83E0F83E07C1F07C1F07C0F83E0F83E0F81F07C1F07C1F83E0F83E0F83F07C1F07C1F03E0F83E0F83F07C1F07C1F03E0F83E0F83F07C1F07C1F03E0F83E0F83F07C1F07C1F83E0F83E0FC1F07C1F07C0F83E0F83E07C1F07C1F83E0F83E0FC1F07C1F07E0F83E0F81F07C1F07C0F83E0F83F07C1F07C0F83E0F83F07C1F07C0F83E0F81F07C1F07E0F83E0FC1F07C1F03E0F83E07C1F07C0F83E0F81F07C1F03E0F83E07C1F07C0F83E0F81F07C1F83E0F83F07C1F03E0F83E07C1F07E0F83E07";
defparam ram_block1a52.mem_init2 = "C1F07E0F83E07C1F07E0F83E07C1F07E0F83E07C1F07E0F83E07C1F03E0F83F07C1F83E0F81F07C0F83E0FC1F07E0F83F07C1F83E0F81F07C0F83E07C1F03E0F81F07C0F83E07C1F03E0F81F07E0F83F07C1F83E0FC1F03E0F81F07E0F83F07C0F83E07C1F83E0FC1F03E0F81F07E0F81F07C0F83F07C0F83F07C0F83E07C1F83E07C1F83E07C1F83E07C1F83E07C1F83E07C1F83E07C0F83F07C0F83F07C0F81F07E0F81F07E0FC1F03E0FC1F83E07C0F83F07E0F81F07E0FC1F03E07C1F83F07E0F81F03E0FC1F83F07C0F81F03E0FC1F83F07C0F81F03E07C1F83F07E0FC1F83E07C0F81F03E07C0F81F03E0FC1F83F07E0FC1F83F07E0FC1F83F07E0FC1F";
defparam ram_block1a52.mem_init1 = "83F07E0FC0F81F03E07C0F81F03E07E0FC1F83F07E0FC0F81F03E07C0FC1F83F07E07C0F81F03F07E0FC0F81F03F07E0FC0F81F03F07E0FC0F81F83F07E07C0FC1F83F03E07E0FC0F81F83F03E07E0FC0F81F83F03E07E0FC0F81F83F03E07E07C0FC1F81F83F03E07E07C0FC1F81F83F03F07E07E0FC0FC1F81F83F03F03E07E07C0FC0FC1F81F83F03F03E07E07E07C0FC0FC1F81F81F83F03F03F07E07E07E07C0FC0FC0FC1F81F81F81F83F03F03F03F03F07E07E07E07E07E07E0FC0FC0FC0FC0FC0FC0FC0FC0FC0FC1F81F81F81F81F81F81F81F81F81F81F81F81F81F80FC0FC0FC0FC0FC0FC0FC0FC0FC0FE07E07E07E07E07E07F03F03F03F03F01F";
defparam ram_block1a52.mem_init0 = "81F81F81F80FC0FC0FC07E07E07E03F03F03F01F81F81FC0FC0FC07E07E07F03F03F81F81FC0FC0FE07E07F03F03F81F80FC0FC07E07F03F01F81FC0FC07E07F03F01F81FC0FC07E03F03F81F80FC07E07F03F81F80FC07E03F03F81FC0FE07F03F81F80FC07E03F01F80FC07E03F01F80FC07F03F81FC0FE07F01F80FC07E03F81FC0FE03F01F80FE07F01F80FC07F03F80FC07F03F80FE07F01F80FE07F01FC0FE03F81FC07F03F80FE07F01FC07E03F80FE07F01FC07E03F80FE03F81FC07F01FC07F03F80FE03F80FE03F80FE03F01FC07F01FC07F01FC07F01FC07F01FC07F01FC03F80FE03F80FE03F80FE01FC07F01FC07F00FE03F80FE01FC07F01FC";

arriav_ram_block ram_block1a4(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a4_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.clk0_input_clock_enable = "ena0";
defparam ram_block1a4.clk0_output_clock_enable = "ena0";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.init_file = "DDS_48_v1_nco_ii_0_sin.hex";
defparam ram_block1a4.init_file_layout = "port_a";
defparam ram_block1a4.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_c8g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.operation_mode = "rom";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 13;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "clock0";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 8191;
defparam ram_block1a4.port_a_logical_ram_depth = 65536;
defparam ram_block1a4.port_a_logical_ram_width = 16;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.ram_block_type = "auto";
defparam ram_block1a4.mem_init3 = "7F01FC07F00FE03F80FE01FC07F01FC07F00FE03F80FE03F80FE03F807F01FC07F01FC07F01FC07F01FC07F01FC07F01F80FE03F80FE03F80FE03F81FC07F01FC07F03F80FE03F80FC07F01FC0FE03F80FC07F01FC0FE03F81FC07F03F80FE07F01FC0FE03F01FC0FE03F81FC07E03F81FC07E03F01FC0FE03F01F80FE07F03F80FC07E03F01FC0FE07F03F81FC07E03F01F80FC07E03F01F80FC07E03F03F81FC0FE07F03F81F80FC07E03F03F81FC0FC07E03F03F81F80FC07E07F03F01F81FC0FC07E07F03F01F81FC0FC07E07E03F03F81F81FC0FC0FE07E07F03F03F81F81FC0FC0FC07E07E07F03F03F01F81F81F80FC0FC0FC07E07E07E03F03F03F03";
defparam ram_block1a4.mem_init2 = "F01F81F81F81F81FC0FC0FC0FC0FC0FC0FE07E07E07E07E07E07E07E07E07E03F03F03F03F03F03F03F03F03F03F03F03F03F03F07E07E07E07E07E07E07E07E07E07E0FC0FC0FC0FC0FC0FC1F81F81F81F81F83F03F03F03F07E07E07E07C0FC0FC0FC1F81F81F83F03F03F07E07E07C0FC0FC0F81F81F83F03F07E07E07C0FC0F81F81F83F03F07E07E0FC0FC1F81F83F03F07E07C0FC0F81F83F03F07E07C0FC0F81F83F03E07E0FC0F81F83F03E07E0FC0F81F83F03E07E0FC0F81F83F07E07C0FC1F83F03E07E0FC1F81F03E07E0FC1F81F03E07E0FC1F81F03E07C0FC1F83F07E07C0F81F03E07E0FC1F83F07E0FC0F81F03E07C0F81F03E07E0FC1F83";
defparam ram_block1a4.mem_init1 = "F07E0FC1F83F07E0FC1F83F07E0FC1F83F07E0F81F03E07C0F81F03E07C0F83F07E0FC1F83F07C0F81F03E07C1F83F07E0F81F03E07C1F83F07E0F81F03E0FC1F83F07C0F81F07E0FC1F03E0FC1F83E07C0F83F07E0F81F07E0FC1F03E0FC1F03E07C1F83E07C1F83E07C0F83F07C0F83F07C0F83F07C0F83F07C0F83F07C0F83F07C0F83E07C1F83E07C1F83E07C1F03E0FC1F03E0F81F07E0F83F07C0F83E07C1F83E0FC1F03E0F81F07E0F83F07C1F83E0FC1F03E0F81F07C0F83E07C1F03E0F81F07C0F83E07C1F03E0F83F07C1F83E0FC1F07E0F83E07C1F03E0F83F07C1F83E0F81F07C0F83E0FC1F07C0F83E0FC1F07C0F83E0FC1F07C0F83E0FC1F07";
defparam ram_block1a4.mem_init0 = "C0F83E0FC1F07C0F83E0F81F07C1F83E0F83F07C1F03E0F83E07C1F07C0F83E0F81F07C1F03E0F83E07C1F07C0F83E0F81F07C1F07E0F83E0FC1F07C1F03E0F83E07C1F07C1F83E0F83E07C1F07C1F83E0F83E07C1F07C1F03E0F83E0FC1F07C1F07E0F83E0F83F07C1F07C0F83E0F83E07C1F07C1F07E0F83E0F83F07C1F07C1F83E0F83E0F81F07C1F07C1F83E0F83E0F81F07C1F07C1F83E0F83E0F81F07C1F07C1F83E0F83E0F83F07C1F07C1F03E0F83E0F83E07C1F07C1F07C0F83E0F83E0F81F07C1F07C1F03E0F83E0F83E0FC1F07C1F07C1F83E0F83E0F83F07C1F07C1F07C0F83E0F83E0F83F07C1F07C1F07E0F83E0F83E0F81F07C1F07C1F07E0";

arriav_ram_block ram_block1a20(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a20_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a20.clk0_core_clock_enable = "ena0";
defparam ram_block1a20.clk0_input_clock_enable = "ena0";
defparam ram_block1a20.clk0_output_clock_enable = "ena0";
defparam ram_block1a20.data_interleave_offset_in_bits = 1;
defparam ram_block1a20.data_interleave_width_in_bits = 1;
defparam ram_block1a20.init_file = "DDS_48_v1_nco_ii_0_sin.hex";
defparam ram_block1a20.init_file_layout = "port_a";
defparam ram_block1a20.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_c8g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a20.operation_mode = "rom";
defparam ram_block1a20.port_a_address_clear = "none";
defparam ram_block1a20.port_a_address_width = 13;
defparam ram_block1a20.port_a_data_out_clear = "none";
defparam ram_block1a20.port_a_data_out_clock = "clock0";
defparam ram_block1a20.port_a_data_width = 1;
defparam ram_block1a20.port_a_first_address = 8192;
defparam ram_block1a20.port_a_first_bit_number = 4;
defparam ram_block1a20.port_a_last_address = 16383;
defparam ram_block1a20.port_a_logical_ram_depth = 65536;
defparam ram_block1a20.port_a_logical_ram_width = 16;
defparam ram_block1a20.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a20.ram_block_type = "auto";
defparam ram_block1a20.mem_init3 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000007FFFFFFFFFFFFFFFFFFC00000000000000000FFFFFFFFFFFFFFFF000000000000000FFFFFFFFFFFFFF00000000000007FFFFFFFFFFFF000000000000FFFFFFFFFFFC00000000003FFFFFFFFFF80000000001FFFFFFFFFE0000000003FFFFFFFFF0000000007FFFFFFFF8000000007FFFFFFFE000000007FFFFFFFC00000003FFFFFFFC00000007FFFFFFF00000003FFFFFFF00000007FFFFFFC0000003FFFFFFC0000007FFFFFF0000001FFFFFFC00";
defparam ram_block1a20.mem_init2 = "0000FFFFFF8000001FFFFFF0000007FFFFF8000003FFFFFC000007FFFFF800000FFFFFE000003FFFFF800001FFFFFC00000FFFFF800001FFFFF800003FFFFE00000FFFFF800007FFFFC00003FFFFC00003FFFFC00003FFFF800007FFFF00001FFFFC00007FFFF00001FFFF80000FFFFC00007FFFE00007FFFE0000FFFFC0000FFFF80001FFFF00007FFFC0001FFFF00007FFFC0001FFFE0000FFFF00007FFF80007FFF80003FFFC0007FFF80007FFF80007FFF0000FFFE0003FFFC0007FFF0001FFFC0007FFF0001FFFC0007FFF0003FFF8001FFFC000FFFE0007FFE0003FFF0003FFF0003FFF0003FFF0003FFF0007FFE0007FFC000FFF8001FFF0003FFE000";
defparam ram_block1a20.mem_init1 = "7FFC001FFF0007FFE000FFF8003FFE000FFF8007FFC001FFF000FFF8003FFC001FFF000FFF0007FF8003FFC003FFE001FFE001FFE000FFF000FFF000FFF000FFF001FFE001FFE001FFE003FFC003FF8007FF000FFF001FFE003FF8007FF000FFE003FF8007FF001FFC003FF800FFE003FF800FFE003FF800FFE003FF801FFC007FF001FF800FFE003FF001FFC00FFE007FF003FF801FFC00FFE007FF003FF001FF801FFC00FFC00FFE007FE007FE007FE003FF003FF003FF003FF003FF003FF007FE007FE007FE007FC00FFC00FF801FF801FF003FF007FE00FFC00FF801FF003FE007FC00FF801FF007FE00FFC01FF003FE00FFC01FF007FE00FF803FF007FC";
defparam ram_block1a20.mem_init0 = "01FF007FE00FF803FE00FF803FE00FF803FE00FF803FE00FF803FE00FF007FC01FF007F803FE00FF807FC01FF00FF803FC01FF00FF803FC01FF00FF807FC01FE00FF007F803FC01FE00FF007F807FC03FE01FE00FF007F807FC03FC01FE01FE00FF00FF807F807F803FC03FC03FE01FE01FE01FE00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FE01FE01FE01FE03FC03FC03FC07F807F80FF00FF01FE01FE03FC03F807F807F00FF01FE03FC03F807F80FF01FE01FC03F807F00FE01FC03F807F00FE01FC03F807F00FE01FC07F80FF01FE03F807F01FE03FC07F00FE03FC07F01FE03F807F01FC03F80FE01FC07F00FE03F80";

arriav_ram_block ram_block1a69(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a69_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a69.clk0_core_clock_enable = "ena0";
defparam ram_block1a69.clk0_input_clock_enable = "ena0";
defparam ram_block1a69.clk0_output_clock_enable = "ena0";
defparam ram_block1a69.data_interleave_offset_in_bits = 1;
defparam ram_block1a69.data_interleave_width_in_bits = 1;
defparam ram_block1a69.init_file = "DDS_48_v1_nco_ii_0_sin.hex";
defparam ram_block1a69.init_file_layout = "port_a";
defparam ram_block1a69.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_c8g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a69.operation_mode = "rom";
defparam ram_block1a69.port_a_address_clear = "none";
defparam ram_block1a69.port_a_address_width = 13;
defparam ram_block1a69.port_a_data_out_clear = "none";
defparam ram_block1a69.port_a_data_out_clock = "clock0";
defparam ram_block1a69.port_a_data_width = 1;
defparam ram_block1a69.port_a_first_address = 32768;
defparam ram_block1a69.port_a_first_bit_number = 5;
defparam ram_block1a69.port_a_last_address = 40959;
defparam ram_block1a69.port_a_logical_ram_depth = 65536;
defparam ram_block1a69.port_a_logical_ram_width = 16;
defparam ram_block1a69.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a69.ram_block_type = "auto";
defparam ram_block1a69.mem_init3 = "0003FFF8001FFFC000FFFC000FFFE0007FFE0007FFF0003FFF0003FFF0003FFF0003FFF0003FFF0003FFF0003FFF0003FFF0003FFF0003FFE0007FFE0007FFE000FFFC000FFF8001FFF8003FFF0003FFE0007FFC000FFFC001FFF8003FFF0007FFC000FFF8001FFF0007FFE000FFF8001FFF0007FFE000FFF8003FFF0007FFC001FFF0007FFE000FFF8003FFE000FFF8003FFE000FFF8003FFE000FFF8003FFE000FFF8003FFE001FFF0007FFC001FFF000FFF8003FFE001FFF0007FFC003FFE000FFF0007FFC003FFE000FFF0007FF8003FFC001FFE000FFF8007FF8003FFC001FFE000FFF0007FF8007FFC003FFE001FFE000FFF000FFF8007FF8007FFC003";
defparam ram_block1a69.mem_init2 = "FFC003FFE001FFE001FFE000FFF000FFF000FFF0007FF8007FF8007FF8007FF8007FF8007FF8007FF8007FF8007FF8007FF8007FF8007FF8007FF8007FF800FFF000FFF000FFF000FFE001FFE001FFE003FFC003FFC003FF8007FF8007FF000FFF001FFE001FFC003FFC007FF8007FF000FFF001FFE003FFC003FF8007FF000FFE001FFC003FF8007FF800FFE001FFC003FF8007FF000FFE001FFC003FF800FFF001FFE003FF8007FF001FFE003FF8007FF001FFE003FF8007FF001FFE003FF800FFF001FFC007FF800FFE003FFC007FF001FFC003FF800FFE003FF8007FF001FFC007FF001FFC003FF800FFE003FF800FFE003FF800FFE001FFC007FF001FFC";
defparam ram_block1a69.mem_init1 = "007FF001FFC007FF001FFC007FF001FFC007FF001FFC007FE003FF800FFE003FF800FFE003FF800FFC007FF001FFC007FF001FF800FFE003FF800FFC007FF001FFC007FE003FF800FFE007FF001FFC00FFE003FF800FFC007FF001FF800FFE007FF001FFC00FFE003FF001FFC007FE003FF801FFC007FE003FF801FFC007FE003FF801FFC00FFE003FF001FFC00FFE007FF001FF800FFC007FF003FF801FFC00FFE003FF001FF800FFC007FE003FF801FFC00FFE007FF003FF801FFC00FFE007FF003FF801FFC00FFE007FF003FF801FFC00FFE007FE003FF001FF800FFC007FE007FF003FF801FFC00FFC007FE003FF001FF801FFC00FFE007FE003FF001FF8";
defparam ram_block1a69.mem_init0 = "01FFC00FFC007FE003FF003FF801FF800FFC00FFE007FF003FF001FF801FFC00FFC007FE007FF003FF001FF801FFC00FFC007FE007FE003FF003FF801FF800FFC00FFC007FE007FF003FF001FF801FF800FFC00FFC007FE007FF003FF003FF801FF801FFC00FFC00FFE007FE007FF003FF003FF801FF801FFC00FFC00FFE007FE007FF003FF003FF001FF801FF800FFC00FFC007FE007FE007FF003FF003FF001FF801FF800FFC00FFC00FFE007FE007FE003FF003FF003FF801FF801FF800FFC00FFC00FFE007FE007FE003FF003FF003FF801FF801FF800FFC00FFC00FFC007FE007FE007FF003FF003FF001FF801FF801FF800FFC00FFC00FFE007FE007FE";

arriav_ram_block ram_block1a85(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a85_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a85.clk0_core_clock_enable = "ena0";
defparam ram_block1a85.clk0_input_clock_enable = "ena0";
defparam ram_block1a85.clk0_output_clock_enable = "ena0";
defparam ram_block1a85.data_interleave_offset_in_bits = 1;
defparam ram_block1a85.data_interleave_width_in_bits = 1;
defparam ram_block1a85.init_file = "DDS_48_v1_nco_ii_0_sin.hex";
defparam ram_block1a85.init_file_layout = "port_a";
defparam ram_block1a85.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_c8g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a85.operation_mode = "rom";
defparam ram_block1a85.port_a_address_clear = "none";
defparam ram_block1a85.port_a_address_width = 13;
defparam ram_block1a85.port_a_data_out_clear = "none";
defparam ram_block1a85.port_a_data_out_clock = "clock0";
defparam ram_block1a85.port_a_data_width = 1;
defparam ram_block1a85.port_a_first_address = 40960;
defparam ram_block1a85.port_a_first_bit_number = 5;
defparam ram_block1a85.port_a_last_address = 49151;
defparam ram_block1a85.port_a_logical_ram_depth = 65536;
defparam ram_block1a85.port_a_logical_ram_width = 16;
defparam ram_block1a85.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a85.ram_block_type = "auto";
defparam ram_block1a85.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000FFFFFFFFFFFFFFFFFFFFF00000000000000000000FFFFFFFFFFFFFFFFFFE000000000000000003FFFFFFFFFFFFFFFFE0000000000000000FFFFFFFFFFFFFFFE000000000000000FFFFFFFFFFFFFFE00000000000000FFFFFFFFFFFFFF00000000000007FFFFFFFFF";
defparam ram_block1a85.mem_init2 = "FFFC0000000000007FFFFFFFFFFFE000000000000FFFFFFFFFFFF000000000001FFFFFFFFFFF800000000003FFFFFFFFFFC00000000003FFFFFFFFFF80000000001FFFFFFFFFF00000000007FFFFFFFFF80000000007FFFFFFFFF0000000003FFFFFFFFF0000000003FFFFFFFFE000000001FFFFFFFFF000000001FFFFFFFFE000000003FFFFFFFF000000003FFFFFFFF000000003FFFFFFFE00000000FFFFFFFF000000007FFFFFFF00000000FFFFFFFF00000001FFFFFFF80000000FFFFFFFC0000000FFFFFFFC0000000FFFFFFF80000001FFFFFFE0000000FFFFFFF80000007FFFFFF80000007FFFFFF80000007FFFFFF0000001FFFFFFC0000007FFFFFF";
defparam ram_block1a85.mem_init1 = "0000003FFFFFF8000001FFFFFF8000001FFFFFF8000003FFFFFF0000007FFFFFC000001FFFFFF0000007FFFFFC000003FFFFFE000001FFFFFE000001FFFFFE000001FFFFFC000003FFFFF8000007FFFFF000001FFFFFC000007FFFFF000001FFFFF800000FFFFFC000007FFFFE000007FFFFE000007FFFFE000007FFFFE00000FFFFFC00001FFFFF800003FFFFE000007FFFFC00001FFFFF00000FFFFF800003FFFFE00001FFFFF00000FFFFF000007FFFF800007FFFF800007FFFF800007FFFF800007FFFF00000FFFFF00001FFFFE00003FFFF800007FFFF00001FFFFC00007FFFF00001FFFFC00007FFFF00003FFFF80000FFFFC00007FFFE00003FFFF000";
defparam ram_block1a85.mem_init0 = "01FFFF80001FFFF80001FFFFC0000FFFFC0000FFFF80001FFFF80001FFFF80003FFFF00003FFFE00007FFFC0000FFFF80001FFFF00007FFFC0000FFFF80003FFFE0000FFFF80003FFFE0000FFFF80003FFFE0001FFFF00007FFF80003FFFE0001FFFF0000FFFF80007FFFC0003FFFC0001FFFE0001FFFE0001FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFE0001FFFE0001FFFE0003FFFC0003FFF80007FFF0000FFFE0001FFFC0003FFF80007FFF0001FFFE0003FFF8000FFFF0001FFFC0007FFF0001FFFC0007FFF8000FFFC0007FFF0001FFFC0007FFF0001FFF8000FFFE0003FFF0001FFFC000FFFE0003FFF0001FFF8000FFFC0007FFE0003FFF";

arriav_ram_block ram_block1a101(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a101_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a101.clk0_core_clock_enable = "ena0";
defparam ram_block1a101.clk0_input_clock_enable = "ena0";
defparam ram_block1a101.clk0_output_clock_enable = "ena0";
defparam ram_block1a101.data_interleave_offset_in_bits = 1;
defparam ram_block1a101.data_interleave_width_in_bits = 1;
defparam ram_block1a101.init_file = "DDS_48_v1_nco_ii_0_sin.hex";
defparam ram_block1a101.init_file_layout = "port_a";
defparam ram_block1a101.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_c8g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a101.operation_mode = "rom";
defparam ram_block1a101.port_a_address_clear = "none";
defparam ram_block1a101.port_a_address_width = 13;
defparam ram_block1a101.port_a_data_out_clear = "none";
defparam ram_block1a101.port_a_data_out_clock = "clock0";
defparam ram_block1a101.port_a_data_width = 1;
defparam ram_block1a101.port_a_first_address = 49152;
defparam ram_block1a101.port_a_first_bit_number = 5;
defparam ram_block1a101.port_a_last_address = 57343;
defparam ram_block1a101.port_a_logical_ram_depth = 65536;
defparam ram_block1a101.port_a_logical_ram_width = 16;
defparam ram_block1a101.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a101.ram_block_type = "auto";
defparam ram_block1a101.mem_init3 = "FFF8000FFFC0007FFE0003FFF0001FFF8000FFFE0007FFF0001FFF8000FFFE0003FFF0001FFFC0007FFF0001FFFC0007FFE0003FFFC0007FFF0001FFFC0007FFF0001FFFE0003FFF8000FFFF0001FFFC0003FFF80007FFF0000FFFE0001FFFC0003FFF80007FFF8000FFFF0000FFFF0000FFFE0001FFFE0001FFFE0001FFFE0001FFFE0001FFFF0000FFFF0000FFFF00007FFF80007FFFC0003FFFE0001FFFF0000FFFF80003FFFC0001FFFF0000FFFF80003FFFE0000FFFF80003FFFE0000FFFF80003FFFE00007FFFC0001FFFF00003FFFE00007FFFC0000FFFF80001FFFF80003FFFF00003FFFF00003FFFE00007FFFE00007FFFF00003FFFF00003FFFF00";
defparam ram_block1a101.mem_init2 = "001FFFF80000FFFFC00007FFFE00003FFFF80001FFFFC00007FFFF00001FFFFC00007FFFF00001FFFFC00003FFFF80000FFFFF00001FFFFE00001FFFFC00003FFFFC00003FFFFC00003FFFFC00003FFFFC00001FFFFE00001FFFFF00000FFFFF800003FFFFE00001FFFFF000007FFFFC00000FFFFF800003FFFFF000007FFFFE00000FFFFFC00000FFFFFC00000FFFFFC00000FFFFFC000007FFFFE000003FFFFF000001FFFFFC000007FFFFF000001FFFFFC000003FFFFF8000007FFFFF000000FFFFFF000000FFFFFF000000FFFFFF8000007FFFFFC000001FFFFFF0000007FFFFFC000001FFFFFF8000003FFFFFF0000003FFFFFF0000003FFFFFF8000001";
defparam ram_block1a101.mem_init1 = "FFFFFFC0000007FFFFFF0000001FFFFFFC0000003FFFFFFC0000003FFFFFFC0000003FFFFFFE0000000FFFFFFF00000003FFFFFFE00000007FFFFFFE00000007FFFFFFE00000003FFFFFFF00000001FFFFFFFE00000001FFFFFFFC00000001FFFFFFFE00000000FFFFFFFF800000001FFFFFFFF800000001FFFFFFFF800000000FFFFFFFFF000000001FFFFFFFFF000000000FFFFFFFFF8000000001FFFFFFFFF8000000001FFFFFFFFFC0000000003FFFFFFFFFC0000000001FFFFFFFFFF00000000003FFFFFFFFFF800000000007FFFFFFFFFF800000000003FFFFFFFFFFF000000000001FFFFFFFFFFFE000000000000FFFFFFFFFFFFC0000000000007FFF";
defparam ram_block1a101.mem_init0 = "FFFFFFFFFC0000000000001FFFFFFFFFFFFFE00000000000000FFFFFFFFFFFFFFE000000000000000FFFFFFFFFFFFFFFE0000000000000000FFFFFFFFFFFFFFFFF800000000000000000FFFFFFFFFFFFFFFFFFE00000000000000000001FFFFFFFFFFFFFFFFFFFFE00000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

arriav_ram_block ram_block1a117(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a117_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a117.clk0_core_clock_enable = "ena0";
defparam ram_block1a117.clk0_input_clock_enable = "ena0";
defparam ram_block1a117.clk0_output_clock_enable = "ena0";
defparam ram_block1a117.data_interleave_offset_in_bits = 1;
defparam ram_block1a117.data_interleave_width_in_bits = 1;
defparam ram_block1a117.init_file = "DDS_48_v1_nco_ii_0_sin.hex";
defparam ram_block1a117.init_file_layout = "port_a";
defparam ram_block1a117.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_c8g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a117.operation_mode = "rom";
defparam ram_block1a117.port_a_address_clear = "none";
defparam ram_block1a117.port_a_address_width = 13;
defparam ram_block1a117.port_a_data_out_clear = "none";
defparam ram_block1a117.port_a_data_out_clock = "clock0";
defparam ram_block1a117.port_a_data_width = 1;
defparam ram_block1a117.port_a_first_address = 57344;
defparam ram_block1a117.port_a_first_bit_number = 5;
defparam ram_block1a117.port_a_last_address = 65535;
defparam ram_block1a117.port_a_logical_ram_depth = 65536;
defparam ram_block1a117.port_a_logical_ram_width = 16;
defparam ram_block1a117.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a117.ram_block_type = "auto";
defparam ram_block1a117.mem_init3 = "FFC00FFC00FFE007FE007FE003FF003FF003FF001FF801FF801FFC00FFC00FFC007FE007FE007FE003FF003FF003FF801FF801FF800FFC00FFC00FFE007FE007FE003FF003FF003FF801FF801FF800FFC00FFC00FFE007FE007FE003FF003FF001FF801FF801FFC00FFC00FFC007FE007FE003FF003FF001FF801FF801FFC00FFC00FFE007FE007FF003FF003FF801FF801FFC00FFC00FFE007FE007FF003FF003FF801FF801FFC00FFC007FE007FE003FF003FF001FF801FFC00FFC007FE007FE003FF003FF801FF800FFC00FFC007FE007FF003FF001FF801FFC00FFC007FE007FF003FF001FF801FFC00FFE007FE003FF003FF801FF800FFC007FE007FF00";
defparam ram_block1a117.mem_init2 = "3FF001FF800FFC00FFE007FF003FF001FF800FFC007FE007FF003FF801FFC00FFC007FE003FF001FF800FFC00FFE007FF003FF801FFC00FFE007FF003FF801FFC00FFE007FF003FF801FFC00FFE007FF003FF800FFC007FE003FF001FF800FFE007FF003FF801FFC007FE003FF001FFC00FFE007FF001FF800FFE007FF003FF800FFC007FF003FF800FFC007FF003FF800FFC007FF001FF800FFE007FF001FFC00FFE003FF001FFC007FE003FF800FFE007FF001FFC00FFE003FF800FFC007FF001FFC007FE003FF800FFE003FF001FFC007FF001FFC007FE003FF800FFE003FF800FFE003FF800FFC007FF001FFC007FF001FFC007FF001FFC007FF001FFC00";
defparam ram_block1a117.mem_init1 = "7FF001FFC007FF000FFE003FF800FFE003FF800FFE003FF8007FF001FFC007FF001FFC003FF800FFE003FF8007FF001FFC007FF800FFE003FFC007FF001FFE003FF800FFF001FFC003FF800FFF001FFC003FF800FFF001FFC003FF800FFF001FFE003FF8007FF000FFE001FFC003FF8007FF000FFE003FFC003FF8007FF000FFE001FFC003FF8007FF800FFF001FFE001FFC003FFC007FF8007FF000FFF001FFE001FFC003FFC003FF8007FF8007FF800FFF000FFF000FFE001FFE001FFE001FFE003FFC003FFC003FFC003FFC003FFC003FFC003FFC003FFC003FFC003FFC003FFC003FFC003FFC003FFC001FFE001FFE001FFE000FFF000FFF000FFF8007FF";
defparam ram_block1a117.mem_init0 = "8007FFC003FFC003FFE001FFE000FFF000FFF8007FFC003FFC001FFE000FFF0007FF8003FFC003FFE000FFF0007FF8003FFC001FFE000FFF8007FFC001FFE000FFF8007FFC001FFF000FFF8003FFE001FFF0007FFC001FFF000FFF8003FFE000FFF8003FFE000FFF8003FFE000FFF8003FFE000FFF8003FFE000FFFC001FFF0007FFC001FFF8003FFE000FFFC001FFF0003FFE000FFFC001FFF0003FFE0007FFC001FFF8003FFF0007FFE0007FFC000FFF8001FFF8003FFF0003FFE0007FFE000FFFC000FFFC000FFF8001FFF8001FFF8001FFF8001FFF8001FFF8001FFF8001FFF8001FFF8001FFF8001FFFC000FFFC000FFFE0007FFE0007FFF0003FFF8001";

arriav_ram_block ram_block1a37(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a37_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a37.clk0_core_clock_enable = "ena0";
defparam ram_block1a37.clk0_input_clock_enable = "ena0";
defparam ram_block1a37.clk0_output_clock_enable = "ena0";
defparam ram_block1a37.data_interleave_offset_in_bits = 1;
defparam ram_block1a37.data_interleave_width_in_bits = 1;
defparam ram_block1a37.init_file = "DDS_48_v1_nco_ii_0_sin.hex";
defparam ram_block1a37.init_file_layout = "port_a";
defparam ram_block1a37.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_c8g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a37.operation_mode = "rom";
defparam ram_block1a37.port_a_address_clear = "none";
defparam ram_block1a37.port_a_address_width = 13;
defparam ram_block1a37.port_a_data_out_clear = "none";
defparam ram_block1a37.port_a_data_out_clock = "clock0";
defparam ram_block1a37.port_a_data_width = 1;
defparam ram_block1a37.port_a_first_address = 16384;
defparam ram_block1a37.port_a_first_bit_number = 5;
defparam ram_block1a37.port_a_last_address = 24575;
defparam ram_block1a37.port_a_logical_ram_depth = 65536;
defparam ram_block1a37.port_a_logical_ram_width = 16;
defparam ram_block1a37.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a37.ram_block_type = "auto";
defparam ram_block1a37.mem_init3 = "0007FFE0003FFF0001FFF8000FFFC0007FFF0003FFF8001FFFC0007FFF0003FFF8000FFFE0003FFF0001FFFC0007FFF0001FFFC0007FFF0001FFFC0007FFF0000FFFE0003FFF80007FFF0001FFFC0003FFF80007FFF0000FFFE0001FFFC0003FFF80007FFF8000FFFF0000FFFE0001FFFE0001FFFE0001FFFE0001FFFE0001FFFE0001FFFE0001FFFE0001FFFF0000FFFF00007FFF80007FFFC0003FFFE0001FFFF0000FFFF80003FFFC0001FFFF00007FFFC0003FFFE0000FFFF80003FFFE0000FFFFC0001FFFF00007FFFE0000FFFF80001FFFF00003FFFE00007FFFC0000FFFFC0001FFFF80001FFFF80001FFFF80001FFFF80001FFFF80001FFFFC0000FF";
defparam ram_block1a37.mem_init2 = "FFC00007FFFE00003FFFF00001FFFF80000FFFFE00003FFFF00001FFFFC00007FFFF00001FFFFE00003FFFF80000FFFFF00001FFFFE00003FFFFC00003FFFFC00007FFFF800007FFFF800007FFFF800003FFFFC00003FFFFE00001FFFFF00000FFFFF800003FFFFE00000FFFFF800003FFFFE00000FFFFF800001FFFFF000003FFFFF000007FFFFE000007FFFFE000007FFFFE000007FFFFF000003FFFFF800001FFFFFC000007FFFFF000001FFFFFC000007FFFFF800000FFFFFF000000FFFFFE000001FFFFFE000001FFFFFF000000FFFFFF8000007FFFFFC000001FFFFFF0000007FFFFFE000000FFFFFFC000001FFFFFF8000001FFFFFFC000000FFFFFFC";
defparam ram_block1a37.mem_init1 = "0000007FFFFFF0000001FFFFFFC0000003FFFFFF80000007FFFFFF80000007FFFFFF80000003FFFFFFE0000000FFFFFFF80000003FFFFFFF00000003FFFFFFF00000003FFFFFFF80000001FFFFFFFC00000003FFFFFFFC00000007FFFFFFFC00000003FFFFFFFE00000000FFFFFFFFC00000000FFFFFFFFC00000000FFFFFFFFE000000001FFFFFFFFC000000003FFFFFFFFE000000000FFFFFFFFFC000000000FFFFFFFFFC0000000007FFFFFFFFF80000000007FFFFFFFFFC0000000001FFFFFFFFFF80000000000FFFFFFFFFFE00000000000FFFFFFFFFFF800000000001FFFFFFFFFFFC000000000007FFFFFFFFFFFC000000000000FFFFFFFFFFFFE0000";
defparam ram_block1a37.mem_init0 = "000000000FFFFFFFFFFFFFC00000000000007FFFFFFFFFFFFFC000000000000007FFFFFFFFFFFFFFC0000000000000007FFFFFFFFFFFFFFFC00000000000000003FFFFFFFFFFFFFFFFFC0000000000000000007FFFFFFFFFFFFFFFFFFF0000000000000000000007FFFFFFFFFFFFFFFFFFFFFE0000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

arriav_ram_block ram_block1a53(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a53_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a53.clk0_core_clock_enable = "ena0";
defparam ram_block1a53.clk0_input_clock_enable = "ena0";
defparam ram_block1a53.clk0_output_clock_enable = "ena0";
defparam ram_block1a53.data_interleave_offset_in_bits = 1;
defparam ram_block1a53.data_interleave_width_in_bits = 1;
defparam ram_block1a53.init_file = "DDS_48_v1_nco_ii_0_sin.hex";
defparam ram_block1a53.init_file_layout = "port_a";
defparam ram_block1a53.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_c8g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a53.operation_mode = "rom";
defparam ram_block1a53.port_a_address_clear = "none";
defparam ram_block1a53.port_a_address_width = 13;
defparam ram_block1a53.port_a_data_out_clear = "none";
defparam ram_block1a53.port_a_data_out_clock = "clock0";
defparam ram_block1a53.port_a_data_width = 1;
defparam ram_block1a53.port_a_first_address = 24576;
defparam ram_block1a53.port_a_first_bit_number = 5;
defparam ram_block1a53.port_a_last_address = 32767;
defparam ram_block1a53.port_a_logical_ram_depth = 65536;
defparam ram_block1a53.port_a_logical_ram_width = 16;
defparam ram_block1a53.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a53.ram_block_type = "auto";
defparam ram_block1a53.mem_init3 = "003FF003FF003FF001FF801FF801FFC00FFC00FFC007FE007FE007FE003FF003FF003FF801FF801FF800FFC00FFC00FFE007FE007FE007FF003FF003FF001FF801FF801FFC00FFC00FFC007FE007FE007FF003FF003FF801FF801FF800FFC00FFC00FFE007FE007FF003FF003FF001FF801FF800FFC00FFC00FFE007FE007FF003FF003FF801FF801FFC00FFC00FFC007FE007FE003FF003FF801FF801FFC00FFC00FFE007FE007FF003FF003FF801FF800FFC00FFC007FE007FF003FF003FF801FF800FFC00FFE007FE003FF003FF001FF801FFC00FFC007FE007FF003FF001FF801FFC00FFC007FE007FF003FF801FF800FFC00FFE007FE003FF001FF801FF";
defparam ram_block1a53.mem_init2 = "C00FFE007FE003FF001FF801FFC00FFE007FE003FF001FF801FFC00FFE007FF003FF801FF800FFC007FE003FF001FF800FFC007FE007FF003FF801FFC00FFE007FF003FF801FFC00FFE007FF001FF800FFC007FE003FF001FF800FFE007FF003FF801FFC007FE003FF001FF800FFE007FF003FF800FFC007FF003FF801FFC007FE003FF801FFC007FE003FF801FFC007FE003FF801FFC007FF003FF800FFC007FF001FF800FFE003FF001FFC007FE003FF800FFE007FF001FFC00FFE003FF800FFE007FF001FFC007FF003FF800FFE003FF800FFC007FF001FFC007FF001FFC007FE003FF800FFE003FF800FFE003FF800FFE003FF800FFE003FF800FFE003FF";
defparam ram_block1a53.mem_init1 = "800FFE003FF800FFE003FF800FFE001FFC007FF001FFC007FF001FFC003FF800FFE003FF800FFF001FFC007FF000FFE003FF800FFF001FFC007FF800FFE003FFC007FF001FFE003FF8007FF001FFE003FF8007FF001FFE003FF8007FF001FFE003FFC007FF800FFE001FFC003FF8007FF000FFE001FFC003FF8007FF000FFE001FFC003FFC007FF800FFF001FFE001FFC003FFC007FF8007FF000FFF001FFE001FFC003FFC003FF8007FF8007FF000FFF000FFF001FFE001FFE001FFE003FFC003FFC003FFC003FFC003FFC007FF8007FF8007FF8007FF8007FF8007FF8007FF8003FFC003FFC003FFC003FFC003FFE001FFE001FFE001FFF000FFF000FFF000";
defparam ram_block1a53.mem_init0 = "7FF8007FF8003FFC003FFE001FFE000FFF000FFF8007FFC003FFC001FFE000FFF0007FF8003FFC001FFE000FFF0007FF8003FFC001FFF000FFF8003FFC001FFF000FFF8003FFC001FFF0007FF8003FFE000FFF8007FFC001FFF0007FFC001FFF0007FF8003FFE000FFF8003FFE000FFF8003FFF0007FFC001FFF0007FFC001FFF8003FFE000FFF8001FFF0007FFC000FFF8003FFF0007FFE000FFF8001FFF0003FFE0007FFC000FFF8001FFF0003FFE0007FFE000FFFC001FFF8001FFF8003FFF0003FFF0007FFE0007FFE0007FFE000FFFC000FFFC000FFFC000FFFC000FFFC000FFFC0007FFE0007FFE0007FFE0003FFF0003FFF0001FFF8001FFFC000FFFC";

arriav_ram_block ram_block1a5(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a5_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.clk0_input_clock_enable = "ena0";
defparam ram_block1a5.clk0_output_clock_enable = "ena0";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.init_file = "DDS_48_v1_nco_ii_0_sin.hex";
defparam ram_block1a5.init_file_layout = "port_a";
defparam ram_block1a5.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_c8g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.operation_mode = "rom";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 13;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "clock0";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 8191;
defparam ram_block1a5.port_a_logical_ram_depth = 65536;
defparam ram_block1a5.port_a_logical_ram_width = 16;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.ram_block_type = "auto";
defparam ram_block1a5.mem_init3 = "7FFE0007FFF0003FFF0001FFF8001FFF8000FFFC000FFFC000FFFC0007FFE0007FFE0007FFE0007FFE0007FFE0007FFE000FFFC000FFFC000FFFC001FFF8001FFF8003FFF0003FFF0007FFE000FFFC000FFF8001FFF0003FFE0007FFC000FFF8001FFF0003FFE000FFFC001FFF8003FFE0007FFC001FFF0003FFE000FFF8003FFF0007FFC001FFF0007FFC001FFF8003FFE000FFF8003FFE000FFF8003FFC001FFF0007FFC001FFF0007FFC003FFE000FFF8003FFC001FFF0007FF8003FFE001FFF0007FF8003FFE001FFF0007FF8003FFC001FFE000FFF0007FF8003FFC001FFE000FFF0007FF8007FFC003FFE001FFE000FFF000FFF8007FF8003FFC003FFC";
defparam ram_block1a5.mem_init2 = "001FFE001FFE001FFF000FFF000FFF000FFF8007FF8007FF8007FF8007FF8003FFC003FFC003FFC003FFC003FFC003FFC003FFC007FF8007FF8007FF8007FF8007FF800FFF000FFF000FFF001FFE001FFE001FFC003FFC003FF8007FF8007FF000FFF001FFE001FFC003FFC007FF8007FF000FFF001FFE003FFC007FF8007FF000FFE001FFC003FF8007FF000FFE001FFC003FF8007FF000FFE003FFC007FF800FFF001FFC003FF800FFF001FFC003FF800FFF001FFC003FF800FFF001FFC007FF800FFE003FFC007FF001FFE003FF800FFE001FFC007FF001FFE003FF800FFE003FF8007FF001FFC007FF001FFC007FF000FFE003FF800FFE003FF800FFE003";
defparam ram_block1a5.mem_init1 = "FF800FFE003FF800FFE003FF800FFE003FF800FFE003FF800FFE003FF800FFC007FF001FFC007FF001FFC007FE003FF800FFE003FF801FFC007FF001FFC00FFE003FF800FFE007FF001FFC00FFE003FF800FFC007FF001FF800FFE003FF001FFC007FE003FF801FFC007FF003FF800FFC007FF003FF800FFC007FF003FF800FFC007FF003FF801FFC007FE003FF801FFC00FFE003FF001FF800FFC007FF003FF801FFC00FFE003FF001FF800FFC007FE003FF001FFC00FFE007FF003FF801FFC00FFE007FF003FF801FFC00FFC007FE003FF001FF800FFC007FE003FF003FF801FFC00FFE007FF003FF001FF800FFC00FFE007FF003FF001FF800FFC00FFE007";
defparam ram_block1a5.mem_init0 = "FF003FF001FF800FFC00FFE007FE003FF003FF801FFC00FFC007FE007FF003FF001FF801FFC00FFC007FE007FF003FF001FF801FF800FFC00FFE007FE003FF003FF801FF801FFC00FFC007FE007FE003FF003FF801FF801FFC00FFC00FFE007FE007FF003FF003FF801FF800FFC00FFC007FE007FE007FF003FF003FF801FF801FFC00FFC00FFE007FE007FE003FF003FF001FF801FF801FFC00FFC00FFE007FE007FE003FF003FF003FF801FF801FFC00FFC00FFC007FE007FE007FF003FF003FF001FF801FF801FFC00FFC00FFC00FFE007FE007FE003FF003FF003FF801FF801FF800FFC00FFC00FFC007FE007FE007FF003FF003FF001FF801FF801FF800";

arriav_ram_block ram_block1a21(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a21_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a21.clk0_core_clock_enable = "ena0";
defparam ram_block1a21.clk0_input_clock_enable = "ena0";
defparam ram_block1a21.clk0_output_clock_enable = "ena0";
defparam ram_block1a21.data_interleave_offset_in_bits = 1;
defparam ram_block1a21.data_interleave_width_in_bits = 1;
defparam ram_block1a21.init_file = "DDS_48_v1_nco_ii_0_sin.hex";
defparam ram_block1a21.init_file_layout = "port_a";
defparam ram_block1a21.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_c8g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a21.operation_mode = "rom";
defparam ram_block1a21.port_a_address_clear = "none";
defparam ram_block1a21.port_a_address_width = 13;
defparam ram_block1a21.port_a_data_out_clear = "none";
defparam ram_block1a21.port_a_data_out_clock = "clock0";
defparam ram_block1a21.port_a_data_width = 1;
defparam ram_block1a21.port_a_first_address = 8192;
defparam ram_block1a21.port_a_first_bit_number = 5;
defparam ram_block1a21.port_a_last_address = 16383;
defparam ram_block1a21.port_a_logical_ram_depth = 65536;
defparam ram_block1a21.port_a_logical_ram_width = 16;
defparam ram_block1a21.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a21.ram_block_type = "auto";
defparam ram_block1a21.mem_init3 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFC000000000000000000001FFFFFFFFFFFFFFFFFFFC0000000000000000007FFFFFFFFFFFFFFFFF800000000000000007FFFFFFFFFFFFFFFC0000000000000007FFFFFFFFFFFFFFC000000000000007FFFFFFFFFFFFFC00000000000007FFFFFFFFFFFFE000000000";
defparam ram_block1a21.mem_init2 = "0000FFFFFFFFFFFFE0000000000007FFFFFFFFFFFC000000000007FFFFFFFFFFF000000000003FFFFFFFFFFE00000000000FFFFFFFFFFE00000000003FFFFFFFFFF00000000007FFFFFFFFFC0000000003FFFFFFFFFC0000000007FFFFFFFFE0000000007FFFFFFFFE000000000FFFFFFFFF8000000007FFFFFFFF000000000FFFFFFFFE000000007FFFFFFFE000000007FFFFFFFE00000000FFFFFFFF800000007FFFFFFFC00000007FFFFFFF800000007FFFFFFF00000003FFFFFFF80000001FFFFFFF80000001FFFFFFF80000003FFFFFFE0000000FFFFFFF80000003FFFFFFC0000003FFFFFFC0000003FFFFFF80000007FFFFFF0000001FFFFFFC000000";
defparam ram_block1a21.mem_init1 = "7FFFFFE0000007FFFFFF0000003FFFFFF0000007FFFFFE000000FFFFFFC000001FFFFFF0000007FFFFFC000003FFFFFE000001FFFFFF000000FFFFFF000000FFFFFE000001FFFFFE000003FFFFFC000007FFFFF000001FFFFFC000007FFFFF000003FFFFF800001FFFFFC00000FFFFFC00000FFFFFC00000FFFFFC00001FFFFF800001FFFFF000003FFFFE00000FFFFF800003FFFFE00000FFFFF800003FFFFE00001FFFFF00000FFFFF800007FFFF800003FFFFC00003FFFFC00003FFFFC00007FFFF800007FFFF80000FFFFF00001FFFFE00003FFFF80000FFFFF00001FFFFC00007FFFF00001FFFF80000FFFFE00003FFFF00001FFFF80000FFFFC00007FF";
defparam ram_block1a21.mem_init0 = "FE00007FFFF00003FFFF00003FFFF00003FFFF00003FFFF00003FFFF00007FFFE00007FFFC0000FFFF80001FFFF00003FFFE0000FFFFC0001FFFF00007FFFE0000FFFF80003FFFE0000FFFF80007FFFC0001FFFF00007FFF80003FFFE0001FFFF0000FFFF80007FFFC0003FFFC0001FFFE0001FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFE0001FFFE0003FFFC0003FFF80007FFF0000FFFE0001FFFC0003FFF80007FFF0001FFFC0003FFF8000FFFE0001FFFC0007FFF0001FFFC0007FFF0001FFFC0007FFF0001FFF8000FFFE0003FFF8001FFFC0007FFF0003FFF8001FFFC0007FFE0003FFF0001FFF8000FFFC000";

arriav_ram_block ram_block1a70(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a70_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a70.clk0_core_clock_enable = "ena0";
defparam ram_block1a70.clk0_input_clock_enable = "ena0";
defparam ram_block1a70.clk0_output_clock_enable = "ena0";
defparam ram_block1a70.data_interleave_offset_in_bits = 1;
defparam ram_block1a70.data_interleave_width_in_bits = 1;
defparam ram_block1a70.init_file = "DDS_48_v1_nco_ii_0_sin.hex";
defparam ram_block1a70.init_file_layout = "port_a";
defparam ram_block1a70.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_c8g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a70.operation_mode = "rom";
defparam ram_block1a70.port_a_address_clear = "none";
defparam ram_block1a70.port_a_address_width = 13;
defparam ram_block1a70.port_a_data_out_clear = "none";
defparam ram_block1a70.port_a_data_out_clock = "clock0";
defparam ram_block1a70.port_a_data_width = 1;
defparam ram_block1a70.port_a_first_address = 32768;
defparam ram_block1a70.port_a_first_bit_number = 6;
defparam ram_block1a70.port_a_last_address = 40959;
defparam ram_block1a70.port_a_logical_ram_depth = 65536;
defparam ram_block1a70.port_a_logical_ram_width = 16;
defparam ram_block1a70.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a70.ram_block_type = "auto";
defparam ram_block1a70.mem_init3 = "00000007FFFFFFC0000003FFFFFFE0000001FFFFFFF0000000FFFFFFF0000000FFFFFFF0000000FFFFFFF0000000FFFFFFF0000000FFFFFFE0000001FFFFFFE0000003FFFFFF80000007FFFFFF0000001FFFFFFC0000003FFFFFF8000000FFFFFFC0000007FFFFFF0000001FFFFFF8000000FFFFFFE0000007FFFFFF0000003FFFFFF0000001FFFFFF8000001FFFFFF8000001FFFFFF8000001FFFFFF8000001FFFFFF8000001FFFFFF0000003FFFFFF0000007FFFFFE000000FFFFFFC000001FFFFFF0000003FFFFFE000000FFFFFF8000003FFFFFE0000007FFFFF8000003FFFFFE000000FFFFFF8000003FFFFFE000001FFFFFF0000007FFFFF8000003FFF";
defparam ram_block1a70.mem_init2 = "FFC000001FFFFFE000001FFFFFF000000FFFFFF0000007FFFFF8000007FFFFF8000007FFFFF8000007FFFFF8000007FFFFF8000007FFFFF8000007FFFFF800000FFFFFF000000FFFFFE000001FFFFFE000003FFFFFC000007FFFFF800000FFFFFF000001FFFFFC000003FFFFF800000FFFFFF000001FFFFFC000007FFFFF000001FFFFFC000007FFFFF800001FFFFFC000007FFFFF000001FFFFFC000007FFFFF000001FFFFF800000FFFFFE000007FFFFF000001FFFFF800000FFFFFE000007FFFFF000003FFFFF800001FFFFFC00000FFFFFC000007FFFFE000007FFFFF000003FFFFF000003FFFFF800001FFFFF800001FFFFF800001FFFFFC00000FFFFFC";
defparam ram_block1a70.mem_init1 = "00000FFFFFC00000FFFFFC00000FFFFFC00000FFFFFC00001FFFFF800001FFFFF800001FFFFF800003FFFFF000003FFFFF000007FFFFE000007FFFFC00000FFFFFC00001FFFFF800001FFFFF000003FFFFE000007FFFFC00000FFFFF800001FFFFF000003FFFFE00000FFFFFC00001FFFFF800003FFFFE000007FFFFC00001FFFFF800003FFFFE00000FFFFFC00001FFFFF000007FFFFC00000FFFFF800003FFFFE00000FFFFF800003FFFFE000007FFFFC00001FFFFF000007FFFFC00001FFFFF000007FFFFC00001FFFFF000007FFFFC00001FFFFE00000FFFFF800003FFFFE00000FFFFF800003FFFFC00001FFFFF000007FFFFC00001FFFFE00000FFFFF8";
defparam ram_block1a70.mem_init0 = "00003FFFFC00001FFFFF000007FFFF800003FFFFE00000FFFFF000007FFFFC00003FFFFE00000FFFFF000007FFFFC00003FFFFE00001FFFFF000007FFFF800003FFFFC00001FFFFF00000FFFFF800007FFFFC00003FFFFE00000FFFFF000007FFFF800003FFFFC00001FFFFE00000FFFFF000007FFFF800003FFFFC00001FFFFE00000FFFFF00000FFFFF800007FFFFC00003FFFFE00001FFFFF00000FFFFF000007FFFF800003FFFFC00001FFFFE00001FFFFF00000FFFFF800007FFFF800003FFFFC00001FFFFE00001FFFFF00000FFFFF800007FFFF800003FFFFC00003FFFFE00001FFFFF00000FFFFF000007FFFF800007FFFFC00003FFFFE00001FFFFE";

arriav_ram_block ram_block1a86(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a86_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a86.clk0_core_clock_enable = "ena0";
defparam ram_block1a86.clk0_input_clock_enable = "ena0";
defparam ram_block1a86.clk0_output_clock_enable = "ena0";
defparam ram_block1a86.data_interleave_offset_in_bits = 1;
defparam ram_block1a86.data_interleave_width_in_bits = 1;
defparam ram_block1a86.init_file = "DDS_48_v1_nco_ii_0_sin.hex";
defparam ram_block1a86.init_file_layout = "port_a";
defparam ram_block1a86.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_c8g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a86.operation_mode = "rom";
defparam ram_block1a86.port_a_address_clear = "none";
defparam ram_block1a86.port_a_address_width = 13;
defparam ram_block1a86.port_a_data_out_clear = "none";
defparam ram_block1a86.port_a_data_out_clock = "clock0";
defparam ram_block1a86.port_a_data_width = 1;
defparam ram_block1a86.port_a_first_address = 40960;
defparam ram_block1a86.port_a_first_bit_number = 6;
defparam ram_block1a86.port_a_last_address = 49151;
defparam ram_block1a86.port_a_logical_ram_depth = 65536;
defparam ram_block1a86.port_a_logical_ram_width = 16;
defparam ram_block1a86.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a86.ram_block_type = "auto";
defparam ram_block1a86.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a86.mem_init2 = "FFFC0000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000007FFFFFFFFFFFFFFFFFFFFFC0000000000000000000007FFFFFFFFFFFFFFFFFFFF000000000000000000007FFFFFFFFFFFFFFFFFFF0000000000000000000FFFFFFFFFFFFFFFFFFE000000000000000000FFFFFFFFFFFFFFFFFE00000000000000000FFFFFFFFFFFFFFFFF00000000000000001FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF0000000000000007FFFFFFFFFFFFFFC000000000000003FFFFFFFFFFFFFF800000000000001FFFFFFFFFFFFFF800000000000007FFFFFFFFFFFFF80000000000000FFFFFFFFFFFFFC0000000000000";
defparam ram_block1a86.mem_init1 = "FFFFFFFFFFFFF80000000000007FFFFFFFFFFFF8000000000000FFFFFFFFFFFFC000000000000FFFFFFFFFFFFC000000000001FFFFFFFFFFFE000000000001FFFFFFFFFFFC000000000007FFFFFFFFFFF000000000003FFFFFFFFFFF000000000007FFFFFFFFFFC00000000001FFFFFFFFFFE00000000001FFFFFFFFFFE00000000003FFFFFFFFFF80000000001FFFFFFFFFFC0000000000FFFFFFFFFF80000000001FFFFFFFFFF0000000000FFFFFFFFFF80000000007FFFFFFFFF80000000007FFFFFFFFF0000000000FFFFFFFFFE0000000007FFFFFFFFF0000000003FFFFFFFFF0000000003FFFFFFFFF0000000007FFFFFFFFC000000001FFFFFFFFF000";
defparam ram_block1a86.mem_init0 = "0000007FFFFFFFF8000000003FFFFFFFFC000000007FFFFFFFF8000000007FFFFFFFF000000001FFFFFFFFC000000007FFFFFFFF000000003FFFFFFFF800000001FFFFFFFF800000001FFFFFFFF800000001FFFFFFFF000000007FFFFFFFE00000000FFFFFFFF800000003FFFFFFFC00000001FFFFFFFE00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFE00000001FFFFFFFE00000003FFFFFFF80000000FFFFFFFE00000003FFFFFFF80000000FFFFFFFE00000007FFFFFFF00000003FFFFFFF00000003FFFFFFF80000003FFFFFFF00000003FFFFFFF00000007FFFFFFE0000000FFFFFFFC0000001FFFFFFF00000007FFFFFFC0000001FFFFFFF";

arriav_ram_block ram_block1a102(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a102_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a102.clk0_core_clock_enable = "ena0";
defparam ram_block1a102.clk0_input_clock_enable = "ena0";
defparam ram_block1a102.clk0_output_clock_enable = "ena0";
defparam ram_block1a102.data_interleave_offset_in_bits = 1;
defparam ram_block1a102.data_interleave_width_in_bits = 1;
defparam ram_block1a102.init_file = "DDS_48_v1_nco_ii_0_sin.hex";
defparam ram_block1a102.init_file_layout = "port_a";
defparam ram_block1a102.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_c8g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a102.operation_mode = "rom";
defparam ram_block1a102.port_a_address_clear = "none";
defparam ram_block1a102.port_a_address_width = 13;
defparam ram_block1a102.port_a_data_out_clear = "none";
defparam ram_block1a102.port_a_data_out_clock = "clock0";
defparam ram_block1a102.port_a_data_width = 1;
defparam ram_block1a102.port_a_first_address = 49152;
defparam ram_block1a102.port_a_first_bit_number = 6;
defparam ram_block1a102.port_a_last_address = 57343;
defparam ram_block1a102.port_a_logical_ram_depth = 65536;
defparam ram_block1a102.port_a_logical_ram_width = 16;
defparam ram_block1a102.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a102.ram_block_type = "auto";
defparam ram_block1a102.mem_init3 = "FFFFFFF00000007FFFFFFC0000001FFFFFFF00000007FFFFFFE0000000FFFFFFFC0000001FFFFFFF80000001FFFFFFF80000003FFFFFFF80000001FFFFFFF80000001FFFFFFFC0000000FFFFFFFE00000003FFFFFFF80000000FFFFFFFE00000003FFFFFFF80000000FFFFFFFF00000000FFFFFFFE00000001FFFFFFFE00000001FFFFFFFE00000000FFFFFFFF000000007FFFFFFF800000003FFFFFFFE00000000FFFFFFFFC00000001FFFFFFFF000000003FFFFFFFF000000003FFFFFFFF000000003FFFFFFFF800000001FFFFFFFFC000000007FFFFFFFF000000001FFFFFFFFC000000003FFFFFFFFC000000007FFFFFFFF8000000003FFFFFFFFC000000";
defparam ram_block1a102.mem_init2 = "001FFFFFFFFF0000000007FFFFFFFFC000000001FFFFFFFFF8000000001FFFFFFFFF8000000001FFFFFFFFFC000000000FFFFFFFFFE0000000001FFFFFFFFFC0000000003FFFFFFFFFC0000000003FFFFFFFFFE0000000001FFFFFFFFFF00000000003FFFFFFFFFE00000000007FFFFFFFFFF00000000003FFFFFFFFFF80000000000FFFFFFFFFFF00000000000FFFFFFFFFFF000000000007FFFFFFFFFFC00000000001FFFFFFFFFFF800000000001FFFFFFFFFFFC000000000007FFFFFFFFFFF000000000000FFFFFFFFFFFF0000000000007FFFFFFFFFFFE0000000000007FFFFFFFFFFFE0000000000003FFFFFFFFFFFFC0000000000003FFFFFFFFFFFFE";
defparam ram_block1a102.mem_init1 = "00000000000007FFFFFFFFFFFFE00000000000003FFFFFFFFFFFFFC00000000000003FFFFFFFFFFFFFF000000000000003FFFFFFFFFFFFFF8000000000000007FFFFFFFFFFFFFFC000000000000001FFFFFFFFFFFFFFFE0000000000000001FFFFFFFFFFFFFFFF00000000000000001FFFFFFFFFFFFFFFFE00000000000000000FFFFFFFFFFFFFFFFFE000000000000000000FFFFFFFFFFFFFFFFFFE0000000000000000001FFFFFFFFFFFFFFFFFFFC00000000000000000001FFFFFFFFFFFFFFFFFFFFC0000000000000000000007FFFFFFFFFFFFFFFFFFFFFC00000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000007FFF";
defparam ram_block1a102.mem_init0 = "FFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

arriav_ram_block ram_block1a118(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a118_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a118.clk0_core_clock_enable = "ena0";
defparam ram_block1a118.clk0_input_clock_enable = "ena0";
defparam ram_block1a118.clk0_output_clock_enable = "ena0";
defparam ram_block1a118.data_interleave_offset_in_bits = 1;
defparam ram_block1a118.data_interleave_width_in_bits = 1;
defparam ram_block1a118.init_file = "DDS_48_v1_nco_ii_0_sin.hex";
defparam ram_block1a118.init_file_layout = "port_a";
defparam ram_block1a118.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_c8g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a118.operation_mode = "rom";
defparam ram_block1a118.port_a_address_clear = "none";
defparam ram_block1a118.port_a_address_width = 13;
defparam ram_block1a118.port_a_data_out_clear = "none";
defparam ram_block1a118.port_a_data_out_clock = "clock0";
defparam ram_block1a118.port_a_data_width = 1;
defparam ram_block1a118.port_a_first_address = 57344;
defparam ram_block1a118.port_a_first_bit_number = 6;
defparam ram_block1a118.port_a_last_address = 65535;
defparam ram_block1a118.port_a_logical_ram_depth = 65536;
defparam ram_block1a118.port_a_logical_ram_width = 16;
defparam ram_block1a118.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a118.ram_block_type = "auto";
defparam ram_block1a118.mem_init3 = "FFFFF00000FFFFF800007FFFFC00003FFFFC00001FFFFE00001FFFFF00000FFFFF800007FFFF800003FFFFC00003FFFFE00001FFFFF00000FFFFF000007FFFF800003FFFFC00003FFFFE00001FFFFF00000FFFFF000007FFFF800003FFFFC00001FFFFE00001FFFFF00000FFFFF800007FFFFC00003FFFFE00001FFFFE00000FFFFF000007FFFF800003FFFFC00001FFFFE00000FFFFF000007FFFF800003FFFFC00001FFFFE00000FFFFF800007FFFFC00003FFFFE00001FFFFF000007FFFF800003FFFFC00001FFFFF00000FFFFF800007FFFFC00001FFFFE00000FFFFF800007FFFFC00001FFFFE00000FFFFF800003FFFFC00001FFFFF000007FFFF80000";
defparam ram_block1a118.mem_init2 = "3FFFFE00000FFFFF000007FFFFC00001FFFFF000007FFFF800003FFFFE00000FFFFF800003FFFFE00000FFFFF000007FFFFC00001FFFFF000007FFFFC00001FFFFF000007FFFFC00001FFFFF000007FFFFC00000FFFFF800003FFFFE00000FFFFF800003FFFFE000007FFFFC00001FFFFF000007FFFFE00000FFFFF800003FFFFF000007FFFFC00000FFFFF800003FFFFF000007FFFFE00000FFFFF800001FFFFF000003FFFFE000007FFFFC00000FFFFF800001FFFFF000003FFFFF000007FFFFE000007FFFFC00000FFFFFC00001FFFFF800001FFFFF800003FFFFF000003FFFFF000003FFFFF000007FFFFE000007FFFFE000007FFFFE000007FFFFE00000";
defparam ram_block1a118.mem_init1 = "7FFFFE000007FFFFF000003FFFFF000003FFFFF000003FFFFF800001FFFFF800001FFFFFC00000FFFFFC000007FFFFE000007FFFFF000003FFFFF800001FFFFFC00000FFFFFE000003FFFFF000001FFFFFC00000FFFFFE000003FFFFF000001FFFFFC000007FFFFF000001FFFFFC000007FFFFF000003FFFFFC000007FFFFF000001FFFFFC000007FFFFF000001FFFFFE000003FFFFF8000007FFFFF000001FFFFFE000003FFFFFC000007FFFFF800000FFFFFF000000FFFFFE000001FFFFFE000003FFFFFC000003FFFFFC000003FFFFFC000003FFFFFC000003FFFFFC000003FFFFFC000003FFFFFC000001FFFFFE000001FFFFFF000000FFFFFF0000007FF";
defparam ram_block1a118.mem_init0 = "FFF8000003FFFFFC000001FFFFFF000000FFFFFF8000003FFFFFE000000FFFFFF8000003FFFFFC000000FFFFFF8000003FFFFFE000000FFFFFF8000001FFFFFF0000007FFFFFE000000FFFFFFC000001FFFFFF8000001FFFFFF0000003FFFFFF0000003FFFFFF0000003FFFFFF0000003FFFFFF0000003FFFFFF0000001FFFFFF8000001FFFFFFC000000FFFFFFE0000003FFFFFF0000001FFFFFFC0000007FFFFFE0000003FFFFFF80000007FFFFFF0000001FFFFFFC0000003FFFFFF8000000FFFFFFF0000000FFFFFFE0000001FFFFFFE0000001FFFFFFE0000001FFFFFFE0000001FFFFFFE0000001FFFFFFF0000000FFFFFFF80000007FFFFFFC0000001";

arriav_ram_block ram_block1a38(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a38_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a38.clk0_core_clock_enable = "ena0";
defparam ram_block1a38.clk0_input_clock_enable = "ena0";
defparam ram_block1a38.clk0_output_clock_enable = "ena0";
defparam ram_block1a38.data_interleave_offset_in_bits = 1;
defparam ram_block1a38.data_interleave_width_in_bits = 1;
defparam ram_block1a38.init_file = "DDS_48_v1_nco_ii_0_sin.hex";
defparam ram_block1a38.init_file_layout = "port_a";
defparam ram_block1a38.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_c8g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a38.operation_mode = "rom";
defparam ram_block1a38.port_a_address_clear = "none";
defparam ram_block1a38.port_a_address_width = 13;
defparam ram_block1a38.port_a_data_out_clear = "none";
defparam ram_block1a38.port_a_data_out_clock = "clock0";
defparam ram_block1a38.port_a_data_width = 1;
defparam ram_block1a38.port_a_first_address = 16384;
defparam ram_block1a38.port_a_first_bit_number = 6;
defparam ram_block1a38.port_a_last_address = 24575;
defparam ram_block1a38.port_a_logical_ram_depth = 65536;
defparam ram_block1a38.port_a_logical_ram_width = 16;
defparam ram_block1a38.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a38.ram_block_type = "auto";
defparam ram_block1a38.mem_init3 = "0000001FFFFFFF00000007FFFFFFC0000000FFFFFFF80000003FFFFFFF00000007FFFFFFE0000000FFFFFFFC0000000FFFFFFFC0000000FFFFFFFC0000000FFFFFFFE00000007FFFFFFF00000003FFFFFFF80000000FFFFFFFE00000003FFFFFFF800000007FFFFFFF00000001FFFFFFFE00000001FFFFFFFE00000001FFFFFFFE00000001FFFFFFFE00000000FFFFFFFF000000007FFFFFFFC00000001FFFFFFFF000000007FFFFFFFC00000000FFFFFFFFC00000001FFFFFFFF800000001FFFFFFFFC00000000FFFFFFFFE000000007FFFFFFFF000000001FFFFFFFFC000000003FFFFFFFF8000000007FFFFFFFF8000000007FFFFFFFF8000000003FFFFFF";
defparam ram_block1a38.mem_init2 = "FFC000000001FFFFFFFFF0000000007FFFFFFFFE000000000FFFFFFFFFC000000000FFFFFFFFFE0000000007FFFFFFFFF0000000001FFFFFFFFFC0000000003FFFFFFFFF80000000007FFFFFFFFF80000000003FFFFFFFFFE0000000000FFFFFFFFFF80000000001FFFFFFFFFF80000000001FFFFFFFFFF80000000000FFFFFFFFFFF00000000001FFFFFFFFFFE00000000001FFFFFFFFFFF000000000007FFFFFFFFFFC00000000000FFFFFFFFFFFC000000000007FFFFFFFFFFF000000000001FFFFFFFFFFFE000000000000FFFFFFFFFFFF8000000000003FFFFFFFFFFFF0000000000001FFFFFFFFFFFFC0000000000007FFFFFFFFFFFFC0000000000003";
defparam ram_block1a38.mem_init1 = "FFFFFFFFFFFFF00000000000003FFFFFFFFFFFFF800000000000007FFFFFFFFFFFFF800000000000001FFFFFFFFFFFFFF800000000000000FFFFFFFFFFFFFFF0000000000000007FFFFFFFFFFFFFFC0000000000000003FFFFFFFFFFFFFFFC0000000000000001FFFFFFFFFFFFFFFFC00000000000000003FFFFFFFFFFFFFFFFE000000000000000003FFFFFFFFFFFFFFFFFE0000000000000000003FFFFFFFFFFFFFFFFFFC00000000000000000007FFFFFFFFFFFFFFFFFFFC000000000000000000007FFFFFFFFFFFFFFFFFFFFE00000000000000000000007FFFFFFFFFFFFFFFFFFFFFFC000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFE0000";
defparam ram_block1a38.mem_init0 = "00000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

arriav_ram_block ram_block1a54(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a54_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a54.clk0_core_clock_enable = "ena0";
defparam ram_block1a54.clk0_input_clock_enable = "ena0";
defparam ram_block1a54.clk0_output_clock_enable = "ena0";
defparam ram_block1a54.data_interleave_offset_in_bits = 1;
defparam ram_block1a54.data_interleave_width_in_bits = 1;
defparam ram_block1a54.init_file = "DDS_48_v1_nco_ii_0_sin.hex";
defparam ram_block1a54.init_file_layout = "port_a";
defparam ram_block1a54.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_c8g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a54.operation_mode = "rom";
defparam ram_block1a54.port_a_address_clear = "none";
defparam ram_block1a54.port_a_address_width = 13;
defparam ram_block1a54.port_a_data_out_clear = "none";
defparam ram_block1a54.port_a_data_out_clock = "clock0";
defparam ram_block1a54.port_a_data_width = 1;
defparam ram_block1a54.port_a_first_address = 24576;
defparam ram_block1a54.port_a_first_bit_number = 6;
defparam ram_block1a54.port_a_last_address = 32767;
defparam ram_block1a54.port_a_logical_ram_depth = 65536;
defparam ram_block1a54.port_a_logical_ram_width = 16;
defparam ram_block1a54.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a54.ram_block_type = "auto";
defparam ram_block1a54.mem_init3 = "00000FFFFF00000FFFFF800007FFFFC00003FFFFC00001FFFFE00001FFFFF00000FFFFF800007FFFF800003FFFFC00001FFFFE00001FFFFF00000FFFFF000007FFFF800003FFFFC00003FFFFE00001FFFFF00000FFFFF800007FFFF800003FFFFC00001FFFFE00000FFFFF00000FFFFF800007FFFFC00003FFFFE00001FFFFF00000FFFFF800007FFFFC00003FFFFC00001FFFFE00000FFFFF800007FFFFC00003FFFFE00001FFFFF00000FFFFF800007FFFFC00003FFFFE00000FFFFF000007FFFF800003FFFFE00001FFFFF00000FFFFF800003FFFFC00001FFFFF00000FFFFF800003FFFFC00001FFFFF000007FFFF800003FFFFE00001FFFFF000007FFFF";
defparam ram_block1a54.mem_init2 = "C00001FFFFE00000FFFFF800003FFFFE00001FFFFF000007FFFFC00001FFFFF000007FFFF800003FFFFE00000FFFFF800003FFFFE00000FFFFF800003FFFFE00000FFFFF800003FFFFE00000FFFFF800003FFFFE00000FFFFF800001FFFFF000007FFFFC00001FFFFF000007FFFFE00000FFFFF800003FFFFF000007FFFFC00001FFFFF800003FFFFE000007FFFFC00001FFFFF800003FFFFF000007FFFFC00000FFFFF800001FFFFF000003FFFFE000007FFFFE00000FFFFFC00001FFFFF800001FFFFF000003FFFFF000007FFFFE000007FFFFC00000FFFFFC00000FFFFFC00001FFFFF800001FFFFF800001FFFFF800001FFFFF800001FFFFF800001FFFFF";
defparam ram_block1a54.mem_init1 = "800001FFFFF800001FFFFF800001FFFFFC00000FFFFFC00000FFFFFC000007FFFFE000007FFFFF000003FFFFF000001FFFFF800000FFFFFC000007FFFFE000003FFFFF000001FFFFF800000FFFFFE000007FFFFF000001FFFFF800000FFFFFE000003FFFFF800001FFFFFC000007FFFFF000001FFFFFC000007FFFFF000001FFFFFC000003FFFFF800000FFFFFE000003FFFFFC000007FFFFF000000FFFFFE000003FFFFFC000007FFFFF800000FFFFFF000000FFFFFE000001FFFFFE000003FFFFFC000003FFFFFC000003FFFFF8000007FFFFF8000007FFFFF8000007FFFFF8000003FFFFFC000003FFFFFC000001FFFFFE000001FFFFFF000000FFFFFF000";
defparam ram_block1a54.mem_init0 = "0007FFFFF8000003FFFFFE000001FFFFFF0000007FFFFFC000003FFFFFE000000FFFFFF8000003FFFFFE000000FFFFFF8000003FFFFFF0000007FFFFFC000000FFFFFF8000003FFFFFF0000007FFFFFE0000007FFFFFC000000FFFFFFC000000FFFFFF8000001FFFFFF8000001FFFFFF8000000FFFFFFC000000FFFFFFC0000007FFFFFE0000007FFFFFF0000003FFFFFF8000000FFFFFFE0000007FFFFFF0000001FFFFFFC0000007FFFFFF0000001FFFFFFE0000003FFFFFF80000007FFFFFF0000000FFFFFFE0000001FFFFFFE0000003FFFFFFC0000003FFFFFFC0000003FFFFFFC0000001FFFFFFE0000001FFFFFFF0000000FFFFFFF80000003FFFFFFC";

arriav_ram_block ram_block1a6(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a6_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.clk0_input_clock_enable = "ena0";
defparam ram_block1a6.clk0_output_clock_enable = "ena0";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.init_file = "DDS_48_v1_nco_ii_0_sin.hex";
defparam ram_block1a6.init_file_layout = "port_a";
defparam ram_block1a6.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_c8g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.operation_mode = "rom";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 13;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "clock0";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 8191;
defparam ram_block1a6.port_a_logical_ram_depth = 65536;
defparam ram_block1a6.port_a_logical_ram_width = 16;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.ram_block_type = "auto";
defparam ram_block1a6.mem_init3 = "7FFFFFF80000003FFFFFFE0000001FFFFFFF0000000FFFFFFF00000007FFFFFF80000007FFFFFF80000007FFFFFF8000000FFFFFFF0000000FFFFFFE0000001FFFFFFC0000003FFFFFF8000000FFFFFFF0000001FFFFFFC0000007FFFFFF0000001FFFFFFC000000FFFFFFE0000003FFFFFF8000001FFFFFFC000000FFFFFFC0000007FFFFFE0000007FFFFFE0000003FFFFFF0000003FFFFFF0000003FFFFFE0000007FFFFFE0000007FFFFFC000000FFFFFFC000001FFFFFF8000003FFFFFE0000007FFFFFC000001FFFFFF8000003FFFFFE000000FFFFFF8000003FFFFFE000000FFFFFF8000007FFFFFC000001FFFFFF000000FFFFFF8000003FFFFFC000";
defparam ram_block1a6.mem_init2 = "001FFFFFE000001FFFFFF000000FFFFFF0000007FFFFF8000007FFFFF8000003FFFFFC000003FFFFFC000003FFFFFC000003FFFFF8000007FFFFF8000007FFFFF800000FFFFFF000000FFFFFE000001FFFFFE000003FFFFFC000007FFFFF800000FFFFFE000001FFFFFC000007FFFFF800000FFFFFE000003FFFFF8000007FFFFF000001FFFFFC000007FFFFF000001FFFFFC000007FFFFF000003FFFFF800000FFFFFE000003FFFFF000001FFFFFC00000FFFFFE000003FFFFF000001FFFFF800000FFFFFC000007FFFFE000003FFFFF000001FFFFF800001FFFFFC00000FFFFFC000007FFFFE000007FFFFE000007FFFFF000003FFFFF000003FFFFF000003";
defparam ram_block1a6.mem_init1 = "FFFFF000003FFFFF000003FFFFF000003FFFFF000003FFFFF000003FFFFF000007FFFFE000007FFFFE000007FFFFC00000FFFFFC00001FFFFF800001FFFFF000003FFFFF000007FFFFE00000FFFFFC00000FFFFF800001FFFFF000003FFFFE000007FFFFC00001FFFFF800003FFFFF000007FFFFC00000FFFFF800003FFFFF000007FFFFC00001FFFFF800003FFFFE00000FFFFFC00001FFFFF000007FFFFC00001FFFFF000003FFFFE00000FFFFF800003FFFFE00000FFFFF800003FFFFE00000FFFFF800003FFFFE00000FFFFF800003FFFFE00000FFFFF800003FFFFC00001FFFFF000007FFFFC00001FFFFF00000FFFFF800003FFFFE00000FFFFF000007";
defparam ram_block1a6.mem_init0 = "FFFFC00001FFFFF00000FFFFF800003FFFFC00001FFFFF000007FFFF800003FFFFE00001FFFFF000007FFFF800003FFFFE00001FFFFF00000FFFFF800003FFFFC00001FFFFE00000FFFFF800007FFFFC00003FFFFE00001FFFFF00000FFFFF800007FFFFC00003FFFFE00000FFFFF000007FFFF800007FFFFC00003FFFFE00001FFFFF00000FFFFF800007FFFFC00003FFFFE00001FFFFE00000FFFFF000007FFFF800003FFFFC00003FFFFE00001FFFFF00000FFFFF800007FFFF800003FFFFC00001FFFFE00001FFFFF00000FFFFF000007FFFF800003FFFFC00003FFFFE00001FFFFF00000FFFFF000007FFFF800007FFFFC00003FFFFE00001FFFFE00000";

arriav_ram_block ram_block1a22(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a22_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a22.clk0_core_clock_enable = "ena0";
defparam ram_block1a22.clk0_input_clock_enable = "ena0";
defparam ram_block1a22.clk0_output_clock_enable = "ena0";
defparam ram_block1a22.data_interleave_offset_in_bits = 1;
defparam ram_block1a22.data_interleave_width_in_bits = 1;
defparam ram_block1a22.init_file = "DDS_48_v1_nco_ii_0_sin.hex";
defparam ram_block1a22.init_file_layout = "port_a";
defparam ram_block1a22.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_c8g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a22.operation_mode = "rom";
defparam ram_block1a22.port_a_address_clear = "none";
defparam ram_block1a22.port_a_address_width = 13;
defparam ram_block1a22.port_a_data_out_clear = "none";
defparam ram_block1a22.port_a_data_out_clock = "clock0";
defparam ram_block1a22.port_a_data_width = 1;
defparam ram_block1a22.port_a_first_address = 8192;
defparam ram_block1a22.port_a_first_bit_number = 6;
defparam ram_block1a22.port_a_last_address = 16383;
defparam ram_block1a22.port_a_logical_ram_depth = 65536;
defparam ram_block1a22.port_a_logical_ram_width = 16;
defparam ram_block1a22.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a22.ram_block_type = "auto";
defparam ram_block1a22.mem_init3 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000";
defparam ram_block1a22.mem_init2 = "0000FFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000FFFFFFFFFFFFFFFFFFFFFC000000000000000000007FFFFFFFFFFFFFFFFFFFC00000000000000000007FFFFFFFFFFFFFFFFFF8000000000000000000FFFFFFFFFFFFFFFFFF800000000000000000FFFFFFFFFFFFFFFFF800000000000000007FFFFFFFFFFFFFFFF00000000000000007FFFFFFFFFFFFFFF80000000000000007FFFFFFFFFFFFFFC000000000000001FFFFFFFFFFFFFFE000000000000003FFFFFFFFFFFFFF000000000000003FFFFFFFFFFFFFC00000000000003FFFFFFFFFFFFF80000000000001FFFFFFFFFFFFF";
defparam ram_block1a22.mem_init1 = "80000000000007FFFFFFFFFFFFC0000000000007FFFFFFFFFFFF0000000000001FFFFFFFFFFFF8000000000003FFFFFFFFFFFE000000000000FFFFFFFFFFFF000000000001FFFFFFFFFFFC000000000007FFFFFFFFFFE000000000007FFFFFFFFFFC00000000001FFFFFFFFFFF00000000000FFFFFFFFFFF00000000001FFFFFFFFFFE00000000003FFFFFFFFFF00000000003FFFFFFFFFF00000000003FFFFFFFFFE0000000000FFFFFFFFFF80000000003FFFFFFFFFC0000000003FFFFFFFFF80000000007FFFFFFFFF0000000001FFFFFFFFFC000000000FFFFFFFFFE0000000007FFFFFFFFE000000000FFFFFFFFFC000000001FFFFFFFFF0000000007FF";
defparam ram_block1a22.mem_init0 = "FFFFFF8000000003FFFFFFFFC000000003FFFFFFFFC000000003FFFFFFFF8000000007FFFFFFFF000000001FFFFFFFFC00000000FFFFFFFFE000000007FFFFFFFF000000003FFFFFFFF000000007FFFFFFFE000000007FFFFFFFC00000001FFFFFFFF000000007FFFFFFFC00000001FFFFFFFE00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000001FFFFFFFC00000003FFFFFFF80000000FFFFFFFE00000003FFFFFFF80000001FFFFFFFC0000000FFFFFFFE00000007FFFFFFE00000007FFFFFFE00000007FFFFFFE0000000FFFFFFFC0000001FFFFFFF80000003FFFFFFE00000007FFFFFFC0000001FFFFFFF0000000";

arriav_ram_block ram_block1a71(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a71_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a71.clk0_core_clock_enable = "ena0";
defparam ram_block1a71.clk0_input_clock_enable = "ena0";
defparam ram_block1a71.clk0_output_clock_enable = "ena0";
defparam ram_block1a71.data_interleave_offset_in_bits = 1;
defparam ram_block1a71.data_interleave_width_in_bits = 1;
defparam ram_block1a71.init_file = "DDS_48_v1_nco_ii_0_sin.hex";
defparam ram_block1a71.init_file_layout = "port_a";
defparam ram_block1a71.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_c8g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a71.operation_mode = "rom";
defparam ram_block1a71.port_a_address_clear = "none";
defparam ram_block1a71.port_a_address_width = 13;
defparam ram_block1a71.port_a_data_out_clear = "none";
defparam ram_block1a71.port_a_data_out_clock = "clock0";
defparam ram_block1a71.port_a_data_width = 1;
defparam ram_block1a71.port_a_first_address = 32768;
defparam ram_block1a71.port_a_first_bit_number = 7;
defparam ram_block1a71.port_a_last_address = 40959;
defparam ram_block1a71.port_a_logical_ram_depth = 65536;
defparam ram_block1a71.port_a_logical_ram_width = 16;
defparam ram_block1a71.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a71.ram_block_type = "auto";
defparam ram_block1a71.mem_init3 = "FFFFFFFFFFFFFFC00000000000001FFFFFFFFFFFFFF00000000000000FFFFFFFFFFFFFF00000000000000FFFFFFFFFFFFFF00000000000001FFFFFFFFFFFFFE00000000000007FFFFFFFFFFFFF00000000000003FFFFFFFFFFFFF80000000000003FFFFFFFFFFFFF00000000000007FFFFFFFFFFFFE0000000000000FFFFFFFFFFFFF00000000000007FFFFFFFFFFFF80000000000007FFFFFFFFFFFF80000000000007FFFFFFFFFFFF0000000000000FFFFFFFFFFFFE0000000000003FFFFFFFFFFFF0000000000001FFFFFFFFFFFF8000000000001FFFFFFFFFFFF8000000000001FFFFFFFFFFFF8000000000001FFFFFFFFFFFF0000000000007FFFFFFFFF";
defparam ram_block1a71.mem_init2 = "FFC000000000001FFFFFFFFFFFF000000000000FFFFFFFFFFFF8000000000007FFFFFFFFFFF8000000000007FFFFFFFFFFF8000000000007FFFFFFFFFFF800000000000FFFFFFFFFFFE000000000001FFFFFFFFFFFC000000000007FFFFFFFFFFF000000000003FFFFFFFFFFF800000000000FFFFFFFFFFFC00000000000FFFFFFFFFFFC000000000007FFFFFFFFFFC00000000000FFFFFFFFFFFC00000000000FFFFFFFFFFF800000000001FFFFFFFFFFF000000000007FFFFFFFFFFE00000000000FFFFFFFFFFF800000000003FFFFFFFFFFC00000000001FFFFFFFFFFF00000000000FFFFFFFFFFF800000000007FFFFFFFFFF800000000003FFFFFFFFFFC";
defparam ram_block1a71.mem_init1 = "00000000003FFFFFFFFFFC00000000003FFFFFFFFFFC00000000007FFFFFFFFFF800000000007FFFFFFFFFF00000000000FFFFFFFFFFE00000000003FFFFFFFFFFC00000000007FFFFFFFFFF00000000001FFFFFFFFFFC00000000007FFFFFFFFFF00000000001FFFFFFFFFFC00000000007FFFFFFFFFE00000000003FFFFFFFFFF80000000001FFFFFFFFFFC0000000000FFFFFFFFFFC00000000007FFFFFFFFFE00000000007FFFFFFFFFE00000000003FFFFFFFFFF00000000003FFFFFFFFFF00000000003FFFFFFFFFF00000000003FFFFFFFFFE00000000007FFFFFFFFFE00000000007FFFFFFFFFC0000000000FFFFFFFFFFC0000000001FFFFFFFFFF8";
defparam ram_block1a71.mem_init0 = "0000000003FFFFFFFFFF00000000007FFFFFFFFFE0000000000FFFFFFFFFFC0000000001FFFFFFFFFF00000000003FFFFFFFFFE0000000000FFFFFFFFFF80000000003FFFFFFFFFF00000000007FFFFFFFFFC0000000001FFFFFFFFFF00000000007FFFFFFFFFC0000000001FFFFFFFFFF00000000007FFFFFFFFFC0000000001FFFFFFFFFF00000000007FFFFFFFFFC0000000001FFFFFFFFFF0000000000FFFFFFFFFF80000000003FFFFFFFFFE0000000000FFFFFFFFFF80000000007FFFFFFFFFC0000000001FFFFFFFFFF00000000007FFFFFFFFF80000000003FFFFFFFFFE0000000000FFFFFFFFFF00000000007FFFFFFFFFC0000000001FFFFFFFFFE";

arriav_ram_block ram_block1a87(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a87_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a87.clk0_core_clock_enable = "ena0";
defparam ram_block1a87.clk0_input_clock_enable = "ena0";
defparam ram_block1a87.clk0_output_clock_enable = "ena0";
defparam ram_block1a87.data_interleave_offset_in_bits = 1;
defparam ram_block1a87.data_interleave_width_in_bits = 1;
defparam ram_block1a87.init_file = "DDS_48_v1_nco_ii_0_sin.hex";
defparam ram_block1a87.init_file_layout = "port_a";
defparam ram_block1a87.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_c8g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a87.operation_mode = "rom";
defparam ram_block1a87.port_a_address_clear = "none";
defparam ram_block1a87.port_a_address_width = 13;
defparam ram_block1a87.port_a_data_out_clear = "none";
defparam ram_block1a87.port_a_data_out_clock = "clock0";
defparam ram_block1a87.port_a_data_width = 1;
defparam ram_block1a87.port_a_first_address = 40960;
defparam ram_block1a87.port_a_first_bit_number = 7;
defparam ram_block1a87.port_a_last_address = 49151;
defparam ram_block1a87.port_a_logical_ram_depth = 65536;
defparam ram_block1a87.port_a_logical_ram_width = 16;
defparam ram_block1a87.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a87.ram_block_type = "auto";
defparam ram_block1a87.mem_init3 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000000000000000000000000000000";
defparam ram_block1a87.mem_init2 = "0003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000003FFFFFFFFFFFFF";
defparam ram_block1a87.mem_init1 = "FFFFFFFFFFFFF800000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000FFFFFFFFFFFFFFFFFFFFFFC0000000000000000000001FFFFFFFFFFFFFFFFFFFFFE0000000000000000000007FFFFFFFFFFFFFFFFFFFFC000000000000000000007FFFFFFFFFFFFFFFFFFFF000000000000000000007FFFFFFFFFFFFFFFFFFF80000000000000000000FFFFFFFFFFFFFFFFFFFE0000000000000000000FFFFFFFFFFFFFFFFFFF0000000000000000000FFFFFFFFFFFFFFFFFFC000000000000000000FFF";
defparam ram_block1a87.mem_init0 = "FFFFFFFFFFFFFFF8000000000000000003FFFFFFFFFFFFFFFFF800000000000000000FFFFFFFFFFFFFFFFFC00000000000000000FFFFFFFFFFFFFFFFF800000000000000007FFFFFFFFFFFFFFFF80000000000000000FFFFFFFFFFFFFFFFE00000000000000007FFFFFFFFFFFFFFFC0000000000000001FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFE0000000000000001FFFFFFFFFFFFFFF8000000000000001FFFFFFFFFFFFFFF8000000000000001FFFFFFFFFFFFFFF000000000000000FFFFFFFFFFFFFFF800000000000000FFFFFFFFFFFFFFF000000000000001FFFFFFFFFFFFFFC00000000000000FFFFFFFFFFFFFFC00000000000000";

arriav_ram_block ram_block1a103(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a103_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a103.clk0_core_clock_enable = "ena0";
defparam ram_block1a103.clk0_input_clock_enable = "ena0";
defparam ram_block1a103.clk0_output_clock_enable = "ena0";
defparam ram_block1a103.data_interleave_offset_in_bits = 1;
defparam ram_block1a103.data_interleave_width_in_bits = 1;
defparam ram_block1a103.init_file = "DDS_48_v1_nco_ii_0_sin.hex";
defparam ram_block1a103.init_file_layout = "port_a";
defparam ram_block1a103.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_c8g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a103.operation_mode = "rom";
defparam ram_block1a103.port_a_address_clear = "none";
defparam ram_block1a103.port_a_address_width = 13;
defparam ram_block1a103.port_a_data_out_clear = "none";
defparam ram_block1a103.port_a_data_out_clock = "clock0";
defparam ram_block1a103.port_a_data_width = 1;
defparam ram_block1a103.port_a_first_address = 49152;
defparam ram_block1a103.port_a_first_bit_number = 7;
defparam ram_block1a103.port_a_last_address = 57343;
defparam ram_block1a103.port_a_logical_ram_depth = 65536;
defparam ram_block1a103.port_a_logical_ram_width = 16;
defparam ram_block1a103.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a103.ram_block_type = "auto";
defparam ram_block1a103.mem_init3 = "000000000000007FFFFFFFFFFFFFE000000000000007FFFFFFFFFFFFFF000000000000001FFFFFFFFFFFFFFE000000000000003FFFFFFFFFFFFFFE000000000000001FFFFFFFFFFFFFFF0000000000000003FFFFFFFFFFFFFFF0000000000000003FFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFE0000000000000001FFFFFFFFFFFFFFFF00000000000000007FFFFFFFFFFFFFFFC0000000000000000FFFFFFFFFFFFFFFFE00000000000000003FFFFFFFFFFFFFFFFC00000000000000003FFFFFFFFFFFFFFFFE000000000000000007FFFFFFFFFFFFFFFFE000000000000000003FFFFFFFFFFFFFFFFF8000000000000000003FFFFFFFFFFFFFFF";
defparam ram_block1a103.mem_init2 = "FFE0000000000000000007FFFFFFFFFFFFFFFFFE0000000000000000001FFFFFFFFFFFFFFFFFFE0000000000000000000FFFFFFFFFFFFFFFFFFFE00000000000000000003FFFFFFFFFFFFFFFFFFFC00000000000000000001FFFFFFFFFFFFFFFFFFFFC000000000000000000007FFFFFFFFFFFFFFFFFFFFC000000000000000000000FFFFFFFFFFFFFFFFFFFFFF00000000000000000000007FFFFFFFFFFFFFFFFFFFFFE00000000000000000000001FFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000003FFFFFFFFFFFFF";
defparam ram_block1a103.mem_init1 = "FFFFFFFFFFFFF8000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000";
defparam ram_block1a103.mem_init0 = "000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

arriav_ram_block ram_block1a119(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a119_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a119.clk0_core_clock_enable = "ena0";
defparam ram_block1a119.clk0_input_clock_enable = "ena0";
defparam ram_block1a119.clk0_output_clock_enable = "ena0";
defparam ram_block1a119.data_interleave_offset_in_bits = 1;
defparam ram_block1a119.data_interleave_width_in_bits = 1;
defparam ram_block1a119.init_file = "DDS_48_v1_nco_ii_0_sin.hex";
defparam ram_block1a119.init_file_layout = "port_a";
defparam ram_block1a119.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_c8g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a119.operation_mode = "rom";
defparam ram_block1a119.port_a_address_clear = "none";
defparam ram_block1a119.port_a_address_width = 13;
defparam ram_block1a119.port_a_data_out_clear = "none";
defparam ram_block1a119.port_a_data_out_clock = "clock0";
defparam ram_block1a119.port_a_data_width = 1;
defparam ram_block1a119.port_a_first_address = 57344;
defparam ram_block1a119.port_a_first_bit_number = 7;
defparam ram_block1a119.port_a_last_address = 65535;
defparam ram_block1a119.port_a_logical_ram_depth = 65536;
defparam ram_block1a119.port_a_logical_ram_width = 16;
defparam ram_block1a119.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a119.ram_block_type = "auto";
defparam ram_block1a119.mem_init3 = "FFFFFFFFFF00000000007FFFFFFFFFC0000000001FFFFFFFFFE0000000000FFFFFFFFFF80000000003FFFFFFFFFC0000000001FFFFFFFFFF00000000007FFFFFFFFFC0000000003FFFFFFFFFE0000000000FFFFFFFFFF80000000003FFFFFFFFFE0000000001FFFFFFFFFF00000000007FFFFFFFFFC0000000001FFFFFFFFFF00000000007FFFFFFFFFC0000000001FFFFFFFFFF00000000007FFFFFFFFFC0000000001FFFFFFFFFF00000000007FFFFFFFFFC0000000001FFFFFFFFFF80000000003FFFFFFFFFE0000000000FFFFFFFFFF80000000001FFFFFFFFFF00000000007FFFFFFFFFE0000000000FFFFFFFFFFC0000000001FFFFFFFFFF8000000000";
defparam ram_block1a119.mem_init2 = "3FFFFFFFFFF00000000007FFFFFFFFFE00000000007FFFFFFFFFC0000000000FFFFFFFFFFC0000000000FFFFFFFFFF80000000001FFFFFFFFFF80000000001FFFFFFFFFF80000000001FFFFFFFFFF80000000000FFFFFFFFFFC0000000000FFFFFFFFFFC00000000007FFFFFFFFFE00000000007FFFFFFFFFF00000000003FFFFFFFFFF80000000000FFFFFFFFFFC00000000007FFFFFFFFFF00000000001FFFFFFFFFFC00000000007FFFFFFFFFF00000000001FFFFFFFFFFC00000000007FFFFFFFFFF80000000000FFFFFFFFFFE00000000001FFFFFFFFFFC00000000003FFFFFFFFFFC00000000007FFFFFFFFFF800000000007FFFFFFFFFF80000000000";
defparam ram_block1a119.mem_init1 = "7FFFFFFFFFF800000000003FFFFFFFFFFC00000000003FFFFFFFFFFE00000000001FFFFFFFFFFF000000000007FFFFFFFFFF800000000003FFFFFFFFFFE00000000000FFFFFFFFFFFC00000000001FFFFFFFFFFF000000000003FFFFFFFFFFE000000000007FFFFFFFFFFE000000000007FFFFFFFFFFC000000000007FFFFFFFFFFE000000000007FFFFFFFFFFE000000000003FFFFFFFFFFF800000000001FFFFFFFFFFFC000000000007FFFFFFFFFFF000000000000FFFFFFFFFFFE000000000003FFFFFFFFFFFC000000000003FFFFFFFFFFFC000000000003FFFFFFFFFFFC000000000003FFFFFFFFFFFE000000000001FFFFFFFFFFFF0000000000007FF";
defparam ram_block1a119.mem_init0 = "FFFFFFFFFC000000000001FFFFFFFFFFFF0000000000003FFFFFFFFFFFF0000000000003FFFFFFFFFFFF0000000000003FFFFFFFFFFFF0000000000001FFFFFFFFFFFF8000000000000FFFFFFFFFFFFE0000000000001FFFFFFFFFFFFC0000000000003FFFFFFFFFFFFC0000000000003FFFFFFFFFFFFC0000000000001FFFFFFFFFFFFE0000000000000FFFFFFFFFFFFFC0000000000001FFFFFFFFFFFFF80000000000003FFFFFFFFFFFFF80000000000001FFFFFFFFFFFFFC0000000000000FFFFFFFFFFFFFF00000000000001FFFFFFFFFFFFFE00000000000001FFFFFFFFFFFFFE00000000000001FFFFFFFFFFFFFF000000000000007FFFFFFFFFFFFFE";

arriav_ram_block ram_block1a39(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a39_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a39.clk0_core_clock_enable = "ena0";
defparam ram_block1a39.clk0_input_clock_enable = "ena0";
defparam ram_block1a39.clk0_output_clock_enable = "ena0";
defparam ram_block1a39.data_interleave_offset_in_bits = 1;
defparam ram_block1a39.data_interleave_width_in_bits = 1;
defparam ram_block1a39.init_file = "DDS_48_v1_nco_ii_0_sin.hex";
defparam ram_block1a39.init_file_layout = "port_a";
defparam ram_block1a39.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_c8g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a39.operation_mode = "rom";
defparam ram_block1a39.port_a_address_clear = "none";
defparam ram_block1a39.port_a_address_width = 13;
defparam ram_block1a39.port_a_data_out_clear = "none";
defparam ram_block1a39.port_a_data_out_clock = "clock0";
defparam ram_block1a39.port_a_data_width = 1;
defparam ram_block1a39.port_a_first_address = 16384;
defparam ram_block1a39.port_a_first_bit_number = 7;
defparam ram_block1a39.port_a_last_address = 24575;
defparam ram_block1a39.port_a_logical_ram_depth = 65536;
defparam ram_block1a39.port_a_logical_ram_width = 16;
defparam ram_block1a39.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a39.ram_block_type = "auto";
defparam ram_block1a39.mem_init3 = "FFFFFFFFFFFFFF000000000000003FFFFFFFFFFFFFF800000000000000FFFFFFFFFFFFFFE000000000000003FFFFFFFFFFFFFFC000000000000003FFFFFFFFFFFFFFE000000000000000FFFFFFFFFFFFFFF8000000000000001FFFFFFFFFFFFFFF8000000000000000FFFFFFFFFFFFFFFE0000000000000001FFFFFFFFFFFFFFFE0000000000000001FFFFFFFFFFFFFFFF00000000000000003FFFFFFFFFFFFFFFF00000000000000003FFFFFFFFFFFFFFFFC00000000000000007FFFFFFFFFFFFFFFFC00000000000000001FFFFFFFFFFFFFFFFF000000000000000003FFFFFFFFFFFFFFFFF8000000000000000007FFFFFFFFFFFFFFFFF8000000000000000";
defparam ram_block1a39.mem_init2 = "003FFFFFFFFFFFFFFFFFF0000000000000000001FFFFFFFFFFFFFFFFFFC0000000000000000001FFFFFFFFFFFFFFFFFFF00000000000000000003FFFFFFFFFFFFFFFFFFF800000000000000000007FFFFFFFFFFFFFFFFFFFE000000000000000000007FFFFFFFFFFFFFFFFFFFF8000000000000000000007FFFFFFFFFFFFFFFFFFFFF0000000000000000000001FFFFFFFFFFFFFFFFFFFFFF00000000000000000000003FFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000";
defparam ram_block1a39.mem_init1 = "0000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000000000000000000000000001FFFF";
defparam ram_block1a39.mem_init0 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

arriav_ram_block ram_block1a55(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a55_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a55.clk0_core_clock_enable = "ena0";
defparam ram_block1a55.clk0_input_clock_enable = "ena0";
defparam ram_block1a55.clk0_output_clock_enable = "ena0";
defparam ram_block1a55.data_interleave_offset_in_bits = 1;
defparam ram_block1a55.data_interleave_width_in_bits = 1;
defparam ram_block1a55.init_file = "DDS_48_v1_nco_ii_0_sin.hex";
defparam ram_block1a55.init_file_layout = "port_a";
defparam ram_block1a55.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_c8g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a55.operation_mode = "rom";
defparam ram_block1a55.port_a_address_clear = "none";
defparam ram_block1a55.port_a_address_width = 13;
defparam ram_block1a55.port_a_data_out_clear = "none";
defparam ram_block1a55.port_a_data_out_clock = "clock0";
defparam ram_block1a55.port_a_data_width = 1;
defparam ram_block1a55.port_a_first_address = 24576;
defparam ram_block1a55.port_a_first_bit_number = 7;
defparam ram_block1a55.port_a_last_address = 32767;
defparam ram_block1a55.port_a_logical_ram_depth = 65536;
defparam ram_block1a55.port_a_logical_ram_width = 16;
defparam ram_block1a55.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a55.ram_block_type = "auto";
defparam ram_block1a55.mem_init3 = "0000000000FFFFFFFFFF80000000003FFFFFFFFFC0000000001FFFFFFFFFF00000000007FFFFFFFFF80000000003FFFFFFFFFE0000000000FFFFFFFFFF00000000007FFFFFFFFFC0000000001FFFFFFFFFF00000000007FFFFFFFFF80000000003FFFFFFFFFE0000000000FFFFFFFFFF80000000003FFFFFFFFFE0000000000FFFFFFFFFF80000000003FFFFFFFFFC0000000001FFFFFFFFFF80000000003FFFFFFFFFE0000000000FFFFFFFFFF80000000003FFFFFFFFFE0000000000FFFFFFFFFF80000000001FFFFFFFFFF00000000007FFFFFFFFFC0000000000FFFFFFFFFF80000000003FFFFFFFFFF00000000007FFFFFFFFFE0000000000FFFFFFFFFF";
defparam ram_block1a55.mem_init2 = "C0000000001FFFFFFFFFF80000000001FFFFFFFFFF00000000003FFFFFFFFFF00000000007FFFFFFFFFE00000000007FFFFFFFFFE00000000007FFFFFFFFFE00000000007FFFFFFFFFE00000000007FFFFFFFFFE00000000007FFFFFFFFFF00000000003FFFFFFFFFF00000000001FFFFFFFFFF80000000000FFFFFFFFFFC00000000007FFFFFFFFFE00000000003FFFFFFFFFF80000000000FFFFFFFFFFC00000000007FFFFFFFFFF00000000001FFFFFFFFFFE00000000003FFFFFFFFFF80000000000FFFFFFFFFFF00000000001FFFFFFFFFFC00000000003FFFFFFFFFFC00000000007FFFFFFFFFF800000000007FFFFFFFFFF800000000007FFFFFFFFFF";
defparam ram_block1a55.mem_init1 = "800000000007FFFFFFFFFF800000000003FFFFFFFFFFC00000000003FFFFFFFFFFE00000000000FFFFFFFFFFF000000000007FFFFFFFFFFC00000000001FFFFFFFFFFF000000000007FFFFFFFFFFE00000000000FFFFFFFFFFF800000000001FFFFFFFFFFF800000000003FFFFFFFFFFF000000000003FFFFFFFFFFF000000000003FFFFFFFFFFF800000000001FFFFFFFFFFFC00000000000FFFFFFFFFFFE000000000003FFFFFFFFFFF800000000000FFFFFFFFFFFE000000000001FFFFFFFFFFFC000000000003FFFFFFFFFFF8000000000007FFFFFFFFFFF8000000000007FFFFFFFFFFFC000000000003FFFFFFFFFFFE000000000000FFFFFFFFFFFF000";
defparam ram_block1a55.mem_init0 = "0000000007FFFFFFFFFFFE000000000000FFFFFFFFFFFFC000000000001FFFFFFFFFFFF8000000000001FFFFFFFFFFFF8000000000000FFFFFFFFFFFFC0000000000007FFFFFFFFFFFF0000000000001FFFFFFFFFFFFC0000000000003FFFFFFFFFFFF80000000000007FFFFFFFFFFFF80000000000003FFFFFFFFFFFFC0000000000001FFFFFFFFFFFFF00000000000007FFFFFFFFFFFFE0000000000000FFFFFFFFFFFFFC0000000000000FFFFFFFFFFFFFE00000000000007FFFFFFFFFFFFF00000000000001FFFFFFFFFFFFFE00000000000003FFFFFFFFFFFFFC00000000000003FFFFFFFFFFFFFE00000000000000FFFFFFFFFFFFFF800000000000003";

arriav_ram_block ram_block1a7(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a7_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.clk0_input_clock_enable = "ena0";
defparam ram_block1a7.clk0_output_clock_enable = "ena0";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.init_file = "DDS_48_v1_nco_ii_0_sin.hex";
defparam ram_block1a7.init_file_layout = "port_a";
defparam ram_block1a7.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_c8g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.operation_mode = "rom";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 13;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "clock0";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 8191;
defparam ram_block1a7.port_a_logical_ram_depth = 65536;
defparam ram_block1a7.port_a_logical_ram_width = 16;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.ram_block_type = "auto";
defparam ram_block1a7.mem_init3 = "800000000000003FFFFFFFFFFFFFE00000000000000FFFFFFFFFFFFFF800000000000007FFFFFFFFFFFFF80000000000000FFFFFFFFFFFFFF00000000000001FFFFFFFFFFFFFC0000000000000FFFFFFFFFFFFFE00000000000007FFFFFFFFFFFFE0000000000000FFFFFFFFFFFFFC0000000000001FFFFFFFFFFFFF00000000000007FFFFFFFFFFFF80000000000003FFFFFFFFFFFFC0000000000003FFFFFFFFFFFF80000000000007FFFFFFFFFFFF0000000000001FFFFFFFFFFFFC0000000000007FFFFFFFFFFFE0000000000003FFFFFFFFFFFF0000000000003FFFFFFFFFFFF0000000000007FFFFFFFFFFFE000000000000FFFFFFFFFFFFC000000000";
defparam ram_block1a7.mem_init2 = "001FFFFFFFFFFFE000000000000FFFFFFFFFFFF8000000000007FFFFFFFFFFFC000000000003FFFFFFFFFFFC000000000003FFFFFFFFFFF8000000000007FFFFFFFFFFF000000000000FFFFFFFFFFFE000000000003FFFFFFFFFFF800000000000FFFFFFFFFFFE000000000007FFFFFFFFFFF000000000003FFFFFFFFFFF800000000001FFFFFFFFFFF800000000001FFFFFFFFFFF800000000003FFFFFFFFFFF000000000003FFFFFFFFFFE00000000000FFFFFFFFFFFC00000000001FFFFFFFFFFF000000000007FFFFFFFFFFC00000000001FFFFFFFFFFE00000000000FFFFFFFFFFF800000000007FFFFFFFFFF800000000003FFFFFFFFFFC00000000003";
defparam ram_block1a7.mem_init1 = "FFFFFFFFFFC00000000003FFFFFFFFFFC00000000003FFFFFFFFFFC00000000007FFFFFFFFFF800000000007FFFFFFFFFF00000000001FFFFFFFFFFE00000000003FFFFFFFFFF80000000000FFFFFFFFFFF00000000001FFFFFFFFFFC00000000007FFFFFFFFFE00000000003FFFFFFFFFF80000000000FFFFFFFFFFC00000000007FFFFFFFFFE00000000003FFFFFFFFFF00000000001FFFFFFFFFF80000000001FFFFFFFFFFC0000000000FFFFFFFFFFC0000000000FFFFFFFFFFC0000000000FFFFFFFFFFC0000000000FFFFFFFFFFC0000000000FFFFFFFFFFC0000000001FFFFFFFFFF80000000001FFFFFFFFFF00000000003FFFFFFFFFF00000000007";
defparam ram_block1a7.mem_init0 = "FFFFFFFFFE0000000000FFFFFFFFFFC0000000001FFFFFFFFFF80000000003FFFFFFFFFE00000000007FFFFFFFFFC0000000001FFFFFFFFFF00000000003FFFFFFFFFE0000000000FFFFFFFFFF80000000003FFFFFFFFFE0000000000FFFFFFFFFF80000000003FFFFFFFFFF00000000007FFFFFFFFF80000000003FFFFFFFFFE0000000000FFFFFFFFFF80000000003FFFFFFFFFE0000000000FFFFFFFFFF80000000003FFFFFFFFFC0000000001FFFFFFFFFF00000000007FFFFFFFFFC0000000001FFFFFFFFFE0000000000FFFFFFFFFF80000000003FFFFFFFFFC0000000001FFFFFFFFFF00000000007FFFFFFFFF80000000003FFFFFFFFFE0000000000";

arriav_ram_block ram_block1a23(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a23_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a23.clk0_core_clock_enable = "ena0";
defparam ram_block1a23.clk0_input_clock_enable = "ena0";
defparam ram_block1a23.clk0_output_clock_enable = "ena0";
defparam ram_block1a23.data_interleave_offset_in_bits = 1;
defparam ram_block1a23.data_interleave_width_in_bits = 1;
defparam ram_block1a23.init_file = "DDS_48_v1_nco_ii_0_sin.hex";
defparam ram_block1a23.init_file_layout = "port_a";
defparam ram_block1a23.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_c8g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a23.operation_mode = "rom";
defparam ram_block1a23.port_a_address_clear = "none";
defparam ram_block1a23.port_a_address_width = 13;
defparam ram_block1a23.port_a_data_out_clear = "none";
defparam ram_block1a23.port_a_data_out_clock = "clock0";
defparam ram_block1a23.port_a_data_width = 1;
defparam ram_block1a23.port_a_first_address = 8192;
defparam ram_block1a23.port_a_first_bit_number = 7;
defparam ram_block1a23.port_a_last_address = 16383;
defparam ram_block1a23.port_a_logical_ram_depth = 65536;
defparam ram_block1a23.port_a_logical_ram_width = 16;
defparam ram_block1a23.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a23.ram_block_type = "auto";
defparam ram_block1a23.mem_init3 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a23.mem_init2 = "FFFF00000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000";
defparam ram_block1a23.mem_init1 = "00000000000007FFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000007FFFFFFFFFFFFFFFFFFFFFF80000000000000000000001FFFFFFFFFFFFFFFFFFFFFF0000000000000000000001FFFFFFFFFFFFFFFFFFFFFC000000000000000000003FFFFFFFFFFFFFFFFFFFFC00000000000000000000FFFFFFFFFFFFFFFFFFFFC00000000000000000003FFFFFFFFFFFFFFFFFFF80000000000000000001FFFFFFFFFFFFFFFFFFF00000000000000000007FFFFFFFFFFFFFFFFFF0000000000000000001FFFFFFFFFFFFFFFFFF800";
defparam ram_block1a23.mem_init0 = "0000000000000003FFFFFFFFFFFFFFFFFC000000000000000003FFFFFFFFFFFFFFFFF800000000000000001FFFFFFFFFFFFFFFFF000000000000000007FFFFFFFFFFFFFFFFC00000000000000007FFFFFFFFFFFFFFFF80000000000000001FFFFFFFFFFFFFFFF80000000000000001FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFE0000000000000003FFFFFFFFFFFFFFF0000000000000003FFFFFFFFFFFFFFE000000000000000FFFFFFFFFFFFFFF8000000000000007FFFFFFFFFFFFFF800000000000000FFFFFFFFFFFFFFE000000000000003FFFFFFFFFFFFFF800000000000001FFFFFFFFFFFFFF";

arriav_ram_block ram_block1a72(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a72_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a72.clk0_core_clock_enable = "ena0";
defparam ram_block1a72.clk0_input_clock_enable = "ena0";
defparam ram_block1a72.clk0_output_clock_enable = "ena0";
defparam ram_block1a72.data_interleave_offset_in_bits = 1;
defparam ram_block1a72.data_interleave_width_in_bits = 1;
defparam ram_block1a72.init_file = "DDS_48_v1_nco_ii_0_sin.hex";
defparam ram_block1a72.init_file_layout = "port_a";
defparam ram_block1a72.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_c8g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a72.operation_mode = "rom";
defparam ram_block1a72.port_a_address_clear = "none";
defparam ram_block1a72.port_a_address_width = 13;
defparam ram_block1a72.port_a_data_out_clear = "none";
defparam ram_block1a72.port_a_data_out_clock = "clock0";
defparam ram_block1a72.port_a_data_width = 1;
defparam ram_block1a72.port_a_first_address = 32768;
defparam ram_block1a72.port_a_first_bit_number = 8;
defparam ram_block1a72.port_a_last_address = 40959;
defparam ram_block1a72.port_a_logical_ram_depth = 65536;
defparam ram_block1a72.port_a_logical_ram_width = 16;
defparam ram_block1a72.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a72.ram_block_type = "auto";
defparam ram_block1a72.mem_init3 = "FFFFFFFFFFFFFFC0000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000";
defparam ram_block1a72.mem_init2 = "003FFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFF800000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000FFFFFFFFFFFFFFFFFFFFFFF800000000000000000000003FFFFFFFFFFFFFFFFFFFFFFC00000000000000000000003FFFFFFFFFFFFFFFFFFFFFFC00000000000000000000007FFFFFFFFFFFFFFFFFFFFFF00000000000000000000001FFFFFFFFFFFFFFFFFFFFFF80000000000000000000003FFFFFFFFFFFFFFFFFFFFFF00000000000000000000007FFFFFFFFFFFFFFFFFFFFF80000000000000000000003";
defparam ram_block1a72.mem_init1 = "FFFFFFFFFFFFFFFFFFFFFC0000000000000000000003FFFFFFFFFFFFFFFFFFFFF8000000000000000000000FFFFFFFFFFFFFFFFFFFFFE0000000000000000000003FFFFFFFFFFFFFFFFFFFFF0000000000000000000003FFFFFFFFFFFFFFFFFFFFF0000000000000000000003FFFFFFFFFFFFFFFFFFFFE0000000000000000000007FFFFFFFFFFFFFFFFFFFFC000000000000000000003FFFFFFFFFFFFFFFFFFFFE000000000000000000001FFFFFFFFFFFFFFFFFFFFF000000000000000000000FFFFFFFFFFFFFFFFFFFFF000000000000000000001FFFFFFFFFFFFFFFFFFFFE000000000000000000003FFFFFFFFFFFFFFFFFFFFC000000000000000000007";
defparam ram_block1a72.mem_init0 = "FFFFFFFFFFFFFFFFFFFF000000000000000000001FFFFFFFFFFFFFFFFFFFFC00000000000000000000FFFFFFFFFFFFFFFFFFFFE000000000000000000007FFFFFFFFFFFFFFFFFFFF000000000000000000003FFFFFFFFFFFFFFFFFFFF000000000000000000003FFFFFFFFFFFFFFFFFFFF000000000000000000003FFFFFFFFFFFFFFFFFFFF000000000000000000003FFFFFFFFFFFFFFFFFFFF000000000000000000007FFFFFFFFFFFFFFFFFFFE000000000000000000007FFFFFFFFFFFFFFFFFFFC00000000000000000000FFFFFFFFFFFFFFFFFFFF800000000000000000001FFFFFFFFFFFFFFFFFFFF000000000000000000003FFFFFFFFFFFFFFFFFFFE";

arriav_ram_block ram_block1a88(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a88_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a88.clk0_core_clock_enable = "ena0";
defparam ram_block1a88.clk0_input_clock_enable = "ena0";
defparam ram_block1a88.clk0_output_clock_enable = "ena0";
defparam ram_block1a88.data_interleave_offset_in_bits = 1;
defparam ram_block1a88.data_interleave_width_in_bits = 1;
defparam ram_block1a88.init_file = "DDS_48_v1_nco_ii_0_sin.hex";
defparam ram_block1a88.init_file_layout = "port_a";
defparam ram_block1a88.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_c8g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a88.operation_mode = "rom";
defparam ram_block1a88.port_a_address_clear = "none";
defparam ram_block1a88.port_a_address_width = 13;
defparam ram_block1a88.port_a_data_out_clear = "none";
defparam ram_block1a88.port_a_data_out_clock = "clock0";
defparam ram_block1a88.port_a_data_width = 1;
defparam ram_block1a88.port_a_first_address = 40960;
defparam ram_block1a88.port_a_first_bit_number = 8;
defparam ram_block1a88.port_a_last_address = 49151;
defparam ram_block1a88.port_a_logical_ram_depth = 65536;
defparam ram_block1a88.port_a_logical_ram_width = 16;
defparam ram_block1a88.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a88.ram_block_type = "auto";
defparam ram_block1a88.mem_init3 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000000000000000000000000000000";
defparam ram_block1a88.mem_init2 = "00000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a88.mem_init1 = "FFFFFFFFFFFFF8000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a88.mem_init0 = "FFFFFFFFFFFFFFF8000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000003FFFFFFFFFFFFFF";

arriav_ram_block ram_block1a104(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a104_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a104.clk0_core_clock_enable = "ena0";
defparam ram_block1a104.clk0_input_clock_enable = "ena0";
defparam ram_block1a104.clk0_output_clock_enable = "ena0";
defparam ram_block1a104.data_interleave_offset_in_bits = 1;
defparam ram_block1a104.data_interleave_width_in_bits = 1;
defparam ram_block1a104.init_file = "DDS_48_v1_nco_ii_0_sin.hex";
defparam ram_block1a104.init_file_layout = "port_a";
defparam ram_block1a104.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_c8g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a104.operation_mode = "rom";
defparam ram_block1a104.port_a_address_clear = "none";
defparam ram_block1a104.port_a_address_width = 13;
defparam ram_block1a104.port_a_data_out_clear = "none";
defparam ram_block1a104.port_a_data_out_clock = "clock0";
defparam ram_block1a104.port_a_data_width = 1;
defparam ram_block1a104.port_a_first_address = 49152;
defparam ram_block1a104.port_a_first_bit_number = 8;
defparam ram_block1a104.port_a_last_address = 57343;
defparam ram_block1a104.port_a_logical_ram_depth = 65536;
defparam ram_block1a104.port_a_logical_ram_width = 16;
defparam ram_block1a104.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a104.ram_block_type = "auto";
defparam ram_block1a104.mem_init3 = "FFFFFFFFFFFFFF800000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000000000003FFFFFFFFFFFFFFF";
defparam ram_block1a104.mem_init2 = "FFFFFFFFFFFFFFFFFFFFF80000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000000003FFFFFFFFFFFFF";
defparam ram_block1a104.mem_init1 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000000000000000000000";
defparam ram_block1a104.mem_init0 = "000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

arriav_ram_block ram_block1a120(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a120_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a120.clk0_core_clock_enable = "ena0";
defparam ram_block1a120.clk0_input_clock_enable = "ena0";
defparam ram_block1a120.clk0_output_clock_enable = "ena0";
defparam ram_block1a120.data_interleave_offset_in_bits = 1;
defparam ram_block1a120.data_interleave_width_in_bits = 1;
defparam ram_block1a120.init_file = "DDS_48_v1_nco_ii_0_sin.hex";
defparam ram_block1a120.init_file_layout = "port_a";
defparam ram_block1a120.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_c8g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a120.operation_mode = "rom";
defparam ram_block1a120.port_a_address_clear = "none";
defparam ram_block1a120.port_a_address_width = 13;
defparam ram_block1a120.port_a_data_out_clear = "none";
defparam ram_block1a120.port_a_data_out_clock = "clock0";
defparam ram_block1a120.port_a_data_width = 1;
defparam ram_block1a120.port_a_first_address = 57344;
defparam ram_block1a120.port_a_first_bit_number = 8;
defparam ram_block1a120.port_a_last_address = 65535;
defparam ram_block1a120.port_a_logical_ram_depth = 65536;
defparam ram_block1a120.port_a_logical_ram_width = 16;
defparam ram_block1a120.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a120.ram_block_type = "auto";
defparam ram_block1a120.mem_init3 = "FFFFFFFFFFFFFFFFFFFF800000000000000000001FFFFFFFFFFFFFFFFFFFF000000000000000000003FFFFFFFFFFFFFFFFFFFE000000000000000000007FFFFFFFFFFFFFFFFFFFC00000000000000000000FFFFFFFFFFFFFFFFFFFFC00000000000000000001FFFFFFFFFFFFFFFFFFFF800000000000000000001FFFFFFFFFFFFFFFFFFFF800000000000000000001FFFFFFFFFFFFFFFFFFFF800000000000000000001FFFFFFFFFFFFFFFFFFFF800000000000000000001FFFFFFFFFFFFFFFFFFFFC00000000000000000000FFFFFFFFFFFFFFFFFFFFE000000000000000000007FFFFFFFFFFFFFFFFFFFF000000000000000000001FFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a120.mem_init2 = "C000000000000000000007FFFFFFFFFFFFFFFFFFFF800000000000000000000FFFFFFFFFFFFFFFFFFFFF000000000000000000001FFFFFFFFFFFFFFFFFFFFE000000000000000000001FFFFFFFFFFFFFFFFFFFFF000000000000000000000FFFFFFFFFFFFFFFFFFFFF8000000000000000000007FFFFFFFFFFFFFFFFFFFFC000000000000000000000FFFFFFFFFFFFFFFFFFFFF8000000000000000000001FFFFFFFFFFFFFFFFFFFFF8000000000000000000001FFFFFFFFFFFFFFFFFFFFF8000000000000000000000FFFFFFFFFFFFFFFFFFFFFE0000000000000000000003FFFFFFFFFFFFFFFFFFFFF80000000000000000000007FFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a120.mem_init1 = "80000000000000000000003FFFFFFFFFFFFFFFFFFFFFC0000000000000000000001FFFFFFFFFFFFFFFFFFFFFF80000000000000000000003FFFFFFFFFFFFFFFFFFFFFF00000000000000000000001FFFFFFFFFFFFFFFFFFFFFFC00000000000000000000007FFFFFFFFFFFFFFFFFFFFFF800000000000000000000007FFFFFFFFFFFFFFFFFFFFFF800000000000000000000003FFFFFFFFFFFFFFFFFFFFFFE000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFF000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFF800";
defparam ram_block1a120.mem_init0 = "0000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000007FFFFFFFFFFFFFF";

arriav_ram_block ram_block1a40(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a40_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a40.clk0_core_clock_enable = "ena0";
defparam ram_block1a40.clk0_input_clock_enable = "ena0";
defparam ram_block1a40.clk0_output_clock_enable = "ena0";
defparam ram_block1a40.data_interleave_offset_in_bits = 1;
defparam ram_block1a40.data_interleave_width_in_bits = 1;
defparam ram_block1a40.init_file = "DDS_48_v1_nco_ii_0_sin.hex";
defparam ram_block1a40.init_file_layout = "port_a";
defparam ram_block1a40.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_c8g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a40.operation_mode = "rom";
defparam ram_block1a40.port_a_address_clear = "none";
defparam ram_block1a40.port_a_address_width = 13;
defparam ram_block1a40.port_a_data_out_clear = "none";
defparam ram_block1a40.port_a_data_out_clock = "clock0";
defparam ram_block1a40.port_a_data_width = 1;
defparam ram_block1a40.port_a_first_address = 16384;
defparam ram_block1a40.port_a_first_bit_number = 8;
defparam ram_block1a40.port_a_last_address = 24575;
defparam ram_block1a40.port_a_logical_ram_depth = 65536;
defparam ram_block1a40.port_a_logical_ram_width = 16;
defparam ram_block1a40.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a40.ram_block_type = "auto";
defparam ram_block1a40.mem_init3 = "00000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000";
defparam ram_block1a40.mem_init2 = "000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000";
defparam ram_block1a40.mem_init1 = "00000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000000000000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a40.mem_init0 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

arriav_ram_block ram_block1a56(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a56_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a56.clk0_core_clock_enable = "ena0";
defparam ram_block1a56.clk0_input_clock_enable = "ena0";
defparam ram_block1a56.clk0_output_clock_enable = "ena0";
defparam ram_block1a56.data_interleave_offset_in_bits = 1;
defparam ram_block1a56.data_interleave_width_in_bits = 1;
defparam ram_block1a56.init_file = "DDS_48_v1_nco_ii_0_sin.hex";
defparam ram_block1a56.init_file_layout = "port_a";
defparam ram_block1a56.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_c8g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a56.operation_mode = "rom";
defparam ram_block1a56.port_a_address_clear = "none";
defparam ram_block1a56.port_a_address_width = 13;
defparam ram_block1a56.port_a_data_out_clear = "none";
defparam ram_block1a56.port_a_data_out_clock = "clock0";
defparam ram_block1a56.port_a_data_width = 1;
defparam ram_block1a56.port_a_first_address = 24576;
defparam ram_block1a56.port_a_first_bit_number = 8;
defparam ram_block1a56.port_a_last_address = 32767;
defparam ram_block1a56.port_a_logical_ram_depth = 65536;
defparam ram_block1a56.port_a_logical_ram_width = 16;
defparam ram_block1a56.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a56.ram_block_type = "auto";
defparam ram_block1a56.mem_init3 = "000000000000000000007FFFFFFFFFFFFFFFFFFFC00000000000000000000FFFFFFFFFFFFFFFFFFFF800000000000000000001FFFFFFFFFFFFFFFFFFFF000000000000000000003FFFFFFFFFFFFFFFFFFFF000000000000000000007FFFFFFFFFFFFFFFFFFFE000000000000000000007FFFFFFFFFFFFFFFFFFFE000000000000000000007FFFFFFFFFFFFFFFFFFFC000000000000000000007FFFFFFFFFFFFFFFFFFFE000000000000000000007FFFFFFFFFFFFFFFFFFFE000000000000000000007FFFFFFFFFFFFFFFFFFFF000000000000000000003FFFFFFFFFFFFFFFFFFFF800000000000000000000FFFFFFFFFFFFFFFFFFFFE00000000000000000000";
defparam ram_block1a56.mem_init2 = "3FFFFFFFFFFFFFFFFFFFF800000000000000000000FFFFFFFFFFFFFFFFFFFFF000000000000000000001FFFFFFFFFFFFFFFFFFFFE000000000000000000001FFFFFFFFFFFFFFFFFFFFE000000000000000000001FFFFFFFFFFFFFFFFFFFFF000000000000000000000FFFFFFFFFFFFFFFFFFFFF8000000000000000000003FFFFFFFFFFFFFFFFFFFFE0000000000000000000007FFFFFFFFFFFFFFFFFFFFC000000000000000000000FFFFFFFFFFFFFFFFFFFFFE0000000000000000000007FFFFFFFFFFFFFFFFFFFFF0000000000000000000003FFFFFFFFFFFFFFFFFFFFFC0000000000000000000007FFFFFFFFFFFFFFFFFFFFF8000000000000000000000";
defparam ram_block1a56.mem_init1 = "7FFFFFFFFFFFFFFFFFFFFF80000000000000000000003FFFFFFFFFFFFFFFFFFFFFE0000000000000000000000FFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000FFFFFFFFFFFFFFFFFFFFFFE00000000000000000000007FFFFFFFFFFFFFFFFFFFFFF80000000000000000000000FFFFFFFFFFFFFFFFFFFFFFF000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFC00000000000000000000001FFFFFFFFFFFFFFFFFFFFFFF800000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000FFF";
defparam ram_block1a56.mem_init0 = "FFFFFFFFFFFFFFFFFFFFFE0000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000";

arriav_ram_block ram_block1a8(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a8_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a8.clk0_core_clock_enable = "ena0";
defparam ram_block1a8.clk0_input_clock_enable = "ena0";
defparam ram_block1a8.clk0_output_clock_enable = "ena0";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.init_file = "DDS_48_v1_nco_ii_0_sin.hex";
defparam ram_block1a8.init_file_layout = "port_a";
defparam ram_block1a8.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_c8g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a8.operation_mode = "rom";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 13;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "clock0";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 8191;
defparam ram_block1a8.port_a_logical_ram_depth = 65536;
defparam ram_block1a8.port_a_logical_ram_width = 16;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a8.ram_block_type = "auto";
defparam ram_block1a8.mem_init3 = "000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000FFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a8.mem_init2 = "FFE000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFF000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFF000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFC00000000000000000000001FFFFFFFFFFFFFFFFFFFFFFE00000000000000000000003FFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000FFFFFFFFFFFFFFFFFFFFFFE00000000000000000000007FFFFFFFFFFFFFFFFFFFFFE0000000000000000000000FFFFFFFFFFFFFFFFFFFFFF80000000000000000000003FFFFFFFFFFFFFFFFFFFFFC";
defparam ram_block1a8.mem_init1 = "0000000000000000000003FFFFFFFFFFFFFFFFFFFFFC0000000000000000000007FFFFFFFFFFFFFFFFFFFFF8000000000000000000001FFFFFFFFFFFFFFFFFFFFFC000000000000000000000FFFFFFFFFFFFFFFFFFFFFE0000000000000000000007FFFFFFFFFFFFFFFFFFFFC000000000000000000000FFFFFFFFFFFFFFFFFFFFF8000000000000000000003FFFFFFFFFFFFFFFFFFFFE000000000000000000001FFFFFFFFFFFFFFFFFFFFF000000000000000000000FFFFFFFFFFFFFFFFFFFFF000000000000000000000FFFFFFFFFFFFFFFFFFFFF000000000000000000001FFFFFFFFFFFFFFFFFFFFE000000000000000000003FFFFFFFFFFFFFFFFFFFF8";
defparam ram_block1a8.mem_init0 = "00000000000000000000FFFFFFFFFFFFFFFFFFFFE000000000000000000003FFFFFFFFFFFFFFFFFFFF800000000000000000001FFFFFFFFFFFFFFFFFFFFC00000000000000000000FFFFFFFFFFFFFFFFFFFFC00000000000000000000FFFFFFFFFFFFFFFFFFFFC000000000000000000007FFFFFFFFFFFFFFFFFFFC00000000000000000000FFFFFFFFFFFFFFFFFFFFC00000000000000000000FFFFFFFFFFFFFFFFFFFFC00000000000000000001FFFFFFFFFFFFFFFFFFFF800000000000000000001FFFFFFFFFFFFFFFFFFFF000000000000000000003FFFFFFFFFFFFFFFFFFFE000000000000000000007FFFFFFFFFFFFFFFFFFFC00000000000000000000";

arriav_ram_block ram_block1a24(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a24_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a24.clk0_core_clock_enable = "ena0";
defparam ram_block1a24.clk0_input_clock_enable = "ena0";
defparam ram_block1a24.clk0_output_clock_enable = "ena0";
defparam ram_block1a24.data_interleave_offset_in_bits = 1;
defparam ram_block1a24.data_interleave_width_in_bits = 1;
defparam ram_block1a24.init_file = "DDS_48_v1_nco_ii_0_sin.hex";
defparam ram_block1a24.init_file_layout = "port_a";
defparam ram_block1a24.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_c8g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a24.operation_mode = "rom";
defparam ram_block1a24.port_a_address_clear = "none";
defparam ram_block1a24.port_a_address_width = 13;
defparam ram_block1a24.port_a_data_out_clear = "none";
defparam ram_block1a24.port_a_data_out_clock = "clock0";
defparam ram_block1a24.port_a_data_width = 1;
defparam ram_block1a24.port_a_first_address = 8192;
defparam ram_block1a24.port_a_first_bit_number = 8;
defparam ram_block1a24.port_a_last_address = 16383;
defparam ram_block1a24.port_a_logical_ram_depth = 65536;
defparam ram_block1a24.port_a_logical_ram_width = 16;
defparam ram_block1a24.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a24.ram_block_type = "auto";
defparam ram_block1a24.mem_init3 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a24.mem_init2 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000000000000000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000000000000000000";
defparam ram_block1a24.mem_init1 = "00000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000";
defparam ram_block1a24.mem_init0 = "0000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000";

arriav_ram_block ram_block1a73(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a73_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a73.clk0_core_clock_enable = "ena0";
defparam ram_block1a73.clk0_input_clock_enable = "ena0";
defparam ram_block1a73.clk0_output_clock_enable = "ena0";
defparam ram_block1a73.data_interleave_offset_in_bits = 1;
defparam ram_block1a73.data_interleave_width_in_bits = 1;
defparam ram_block1a73.init_file = "DDS_48_v1_nco_ii_0_sin.hex";
defparam ram_block1a73.init_file_layout = "port_a";
defparam ram_block1a73.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_c8g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a73.operation_mode = "rom";
defparam ram_block1a73.port_a_address_clear = "none";
defparam ram_block1a73.port_a_address_width = 13;
defparam ram_block1a73.port_a_data_out_clear = "none";
defparam ram_block1a73.port_a_data_out_clock = "clock0";
defparam ram_block1a73.port_a_data_width = 1;
defparam ram_block1a73.port_a_first_address = 32768;
defparam ram_block1a73.port_a_first_bit_number = 9;
defparam ram_block1a73.port_a_last_address = 40959;
defparam ram_block1a73.port_a_logical_ram_depth = 65536;
defparam ram_block1a73.port_a_logical_ram_width = 16;
defparam ram_block1a73.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a73.ram_block_type = "auto";
defparam ram_block1a73.mem_init3 = "000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000";
defparam ram_block1a73.mem_init2 = "000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a73.mem_init1 = "FFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a73.mem_init0 = "FFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE";

arriav_ram_block ram_block1a89(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a89_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a89.clk0_core_clock_enable = "ena0";
defparam ram_block1a89.clk0_input_clock_enable = "ena0";
defparam ram_block1a89.clk0_output_clock_enable = "ena0";
defparam ram_block1a89.data_interleave_offset_in_bits = 1;
defparam ram_block1a89.data_interleave_width_in_bits = 1;
defparam ram_block1a89.init_file = "DDS_48_v1_nco_ii_0_sin.hex";
defparam ram_block1a89.init_file_layout = "port_a";
defparam ram_block1a89.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_c8g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a89.operation_mode = "rom";
defparam ram_block1a89.port_a_address_clear = "none";
defparam ram_block1a89.port_a_address_width = 13;
defparam ram_block1a89.port_a_data_out_clear = "none";
defparam ram_block1a89.port_a_data_out_clock = "clock0";
defparam ram_block1a89.port_a_data_width = 1;
defparam ram_block1a89.port_a_first_address = 40960;
defparam ram_block1a89.port_a_first_bit_number = 9;
defparam ram_block1a89.port_a_last_address = 49151;
defparam ram_block1a89.port_a_logical_ram_depth = 65536;
defparam ram_block1a89.port_a_logical_ram_width = 16;
defparam ram_block1a89.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a89.ram_block_type = "auto";
defparam ram_block1a89.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a89.mem_init2 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a89.mem_init1 = "00000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000000000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a89.mem_init0 = "0000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000000000000000000000";

arriav_ram_block ram_block1a105(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a105_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a105.clk0_core_clock_enable = "ena0";
defparam ram_block1a105.clk0_input_clock_enable = "ena0";
defparam ram_block1a105.clk0_output_clock_enable = "ena0";
defparam ram_block1a105.data_interleave_offset_in_bits = 1;
defparam ram_block1a105.data_interleave_width_in_bits = 1;
defparam ram_block1a105.init_file = "DDS_48_v1_nco_ii_0_sin.hex";
defparam ram_block1a105.init_file_layout = "port_a";
defparam ram_block1a105.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_c8g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a105.operation_mode = "rom";
defparam ram_block1a105.port_a_address_clear = "none";
defparam ram_block1a105.port_a_address_width = 13;
defparam ram_block1a105.port_a_data_out_clear = "none";
defparam ram_block1a105.port_a_data_out_clock = "clock0";
defparam ram_block1a105.port_a_data_width = 1;
defparam ram_block1a105.port_a_first_address = 49152;
defparam ram_block1a105.port_a_first_bit_number = 9;
defparam ram_block1a105.port_a_last_address = 57343;
defparam ram_block1a105.port_a_logical_ram_depth = 65536;
defparam ram_block1a105.port_a_logical_ram_width = 16;
defparam ram_block1a105.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a105.ram_block_type = "auto";
defparam ram_block1a105.mem_init3 = "00000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000";
defparam ram_block1a105.mem_init2 = "00000000000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000000000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000";
defparam ram_block1a105.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a105.mem_init0 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

arriav_ram_block ram_block1a121(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a121_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a121.clk0_core_clock_enable = "ena0";
defparam ram_block1a121.clk0_input_clock_enable = "ena0";
defparam ram_block1a121.clk0_output_clock_enable = "ena0";
defparam ram_block1a121.data_interleave_offset_in_bits = 1;
defparam ram_block1a121.data_interleave_width_in_bits = 1;
defparam ram_block1a121.init_file = "DDS_48_v1_nco_ii_0_sin.hex";
defparam ram_block1a121.init_file_layout = "port_a";
defparam ram_block1a121.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_c8g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a121.operation_mode = "rom";
defparam ram_block1a121.port_a_address_clear = "none";
defparam ram_block1a121.port_a_address_width = 13;
defparam ram_block1a121.port_a_data_out_clear = "none";
defparam ram_block1a121.port_a_data_out_clock = "clock0";
defparam ram_block1a121.port_a_data_width = 1;
defparam ram_block1a121.port_a_first_address = 57344;
defparam ram_block1a121.port_a_first_bit_number = 9;
defparam ram_block1a121.port_a_last_address = 65535;
defparam ram_block1a121.port_a_logical_ram_depth = 65536;
defparam ram_block1a121.port_a_logical_ram_width = 16;
defparam ram_block1a121.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a121.ram_block_type = "auto";
defparam ram_block1a121.mem_init3 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a121.mem_init2 = "FFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a121.mem_init1 = "FFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000000";
defparam ram_block1a121.mem_init0 = "0000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000";

arriav_ram_block ram_block1a41(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a41_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a41.clk0_core_clock_enable = "ena0";
defparam ram_block1a41.clk0_input_clock_enable = "ena0";
defparam ram_block1a41.clk0_output_clock_enable = "ena0";
defparam ram_block1a41.data_interleave_offset_in_bits = 1;
defparam ram_block1a41.data_interleave_width_in_bits = 1;
defparam ram_block1a41.init_file = "DDS_48_v1_nco_ii_0_sin.hex";
defparam ram_block1a41.init_file_layout = "port_a";
defparam ram_block1a41.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_c8g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a41.operation_mode = "rom";
defparam ram_block1a41.port_a_address_clear = "none";
defparam ram_block1a41.port_a_address_width = 13;
defparam ram_block1a41.port_a_data_out_clear = "none";
defparam ram_block1a41.port_a_data_out_clock = "clock0";
defparam ram_block1a41.port_a_data_width = 1;
defparam ram_block1a41.port_a_first_address = 16384;
defparam ram_block1a41.port_a_first_bit_number = 9;
defparam ram_block1a41.port_a_last_address = 24575;
defparam ram_block1a41.port_a_logical_ram_depth = 65536;
defparam ram_block1a41.port_a_logical_ram_width = 16;
defparam ram_block1a41.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a41.ram_block_type = "auto";
defparam ram_block1a41.mem_init3 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFF";
defparam ram_block1a41.mem_init2 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFF";
defparam ram_block1a41.mem_init1 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a41.mem_init0 = "000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

arriav_ram_block ram_block1a57(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a57_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a57.clk0_core_clock_enable = "ena0";
defparam ram_block1a57.clk0_input_clock_enable = "ena0";
defparam ram_block1a57.clk0_output_clock_enable = "ena0";
defparam ram_block1a57.data_interleave_offset_in_bits = 1;
defparam ram_block1a57.data_interleave_width_in_bits = 1;
defparam ram_block1a57.init_file = "DDS_48_v1_nco_ii_0_sin.hex";
defparam ram_block1a57.init_file_layout = "port_a";
defparam ram_block1a57.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_c8g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a57.operation_mode = "rom";
defparam ram_block1a57.port_a_address_clear = "none";
defparam ram_block1a57.port_a_address_width = 13;
defparam ram_block1a57.port_a_data_out_clear = "none";
defparam ram_block1a57.port_a_data_out_clock = "clock0";
defparam ram_block1a57.port_a_data_width = 1;
defparam ram_block1a57.port_a_first_address = 24576;
defparam ram_block1a57.port_a_first_bit_number = 9;
defparam ram_block1a57.port_a_last_address = 32767;
defparam ram_block1a57.port_a_logical_ram_depth = 65536;
defparam ram_block1a57.port_a_logical_ram_width = 16;
defparam ram_block1a57.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a57.ram_block_type = "auto";
defparam ram_block1a57.mem_init3 = "00000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000";
defparam ram_block1a57.mem_init2 = "0000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000";
defparam ram_block1a57.mem_init1 = "00000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a57.mem_init0 = "FFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFF";

arriav_ram_block ram_block1a9(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a9_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a9.clk0_core_clock_enable = "ena0";
defparam ram_block1a9.clk0_input_clock_enable = "ena0";
defparam ram_block1a9.clk0_output_clock_enable = "ena0";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.init_file = "DDS_48_v1_nco_ii_0_sin.hex";
defparam ram_block1a9.init_file_layout = "port_a";
defparam ram_block1a9.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_c8g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a9.operation_mode = "rom";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 13;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "clock0";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 8191;
defparam ram_block1a9.port_a_logical_ram_depth = 65536;
defparam ram_block1a9.port_a_logical_ram_width = 16;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a9.ram_block_type = "auto";
defparam ram_block1a9.mem_init3 = "FFFFFFFFFFFFFFC000000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a9.mem_init2 = "FFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000";
defparam ram_block1a9.mem_init1 = "0000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000";
defparam ram_block1a9.mem_init0 = "00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000000000000000000";

arriav_ram_block ram_block1a25(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a25_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a25.clk0_core_clock_enable = "ena0";
defparam ram_block1a25.clk0_input_clock_enable = "ena0";
defparam ram_block1a25.clk0_output_clock_enable = "ena0";
defparam ram_block1a25.data_interleave_offset_in_bits = 1;
defparam ram_block1a25.data_interleave_width_in_bits = 1;
defparam ram_block1a25.init_file = "DDS_48_v1_nco_ii_0_sin.hex";
defparam ram_block1a25.init_file_layout = "port_a";
defparam ram_block1a25.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_c8g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a25.operation_mode = "rom";
defparam ram_block1a25.port_a_address_clear = "none";
defparam ram_block1a25.port_a_address_width = 13;
defparam ram_block1a25.port_a_data_out_clear = "none";
defparam ram_block1a25.port_a_data_out_clock = "clock0";
defparam ram_block1a25.port_a_data_width = 1;
defparam ram_block1a25.port_a_first_address = 8192;
defparam ram_block1a25.port_a_first_bit_number = 9;
defparam ram_block1a25.port_a_last_address = 16383;
defparam ram_block1a25.port_a_logical_ram_depth = 65536;
defparam ram_block1a25.port_a_logical_ram_width = 16;
defparam ram_block1a25.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a25.ram_block_type = "auto";
defparam ram_block1a25.mem_init3 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000000000000000000000000";
defparam ram_block1a25.mem_init2 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a25.mem_init1 = "FFFFFFFFFFFFF80000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000000000000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a25.mem_init0 = "FFFFFFFFFFFFFFFC00000000000000000000000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

arriav_ram_block ram_block1a74(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a74_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a74.clk0_core_clock_enable = "ena0";
defparam ram_block1a74.clk0_input_clock_enable = "ena0";
defparam ram_block1a74.clk0_output_clock_enable = "ena0";
defparam ram_block1a74.data_interleave_offset_in_bits = 1;
defparam ram_block1a74.data_interleave_width_in_bits = 1;
defparam ram_block1a74.init_file = "DDS_48_v1_nco_ii_0_sin.hex";
defparam ram_block1a74.init_file_layout = "port_a";
defparam ram_block1a74.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_c8g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a74.operation_mode = "rom";
defparam ram_block1a74.port_a_address_clear = "none";
defparam ram_block1a74.port_a_address_width = 13;
defparam ram_block1a74.port_a_data_out_clear = "none";
defparam ram_block1a74.port_a_data_out_clock = "clock0";
defparam ram_block1a74.port_a_data_width = 1;
defparam ram_block1a74.port_a_first_address = 32768;
defparam ram_block1a74.port_a_first_bit_number = 10;
defparam ram_block1a74.port_a_last_address = 40959;
defparam ram_block1a74.port_a_logical_ram_depth = 65536;
defparam ram_block1a74.port_a_logical_ram_width = 16;
defparam ram_block1a74.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a74.ram_block_type = "auto";
defparam ram_block1a74.mem_init3 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000";
defparam ram_block1a74.mem_init2 = "0000000000000000000000000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a74.mem_init1 = "FFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000000000000000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a74.mem_init0 = "FFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE";

arriav_ram_block ram_block1a90(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a90_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a90.clk0_core_clock_enable = "ena0";
defparam ram_block1a90.clk0_input_clock_enable = "ena0";
defparam ram_block1a90.clk0_output_clock_enable = "ena0";
defparam ram_block1a90.data_interleave_offset_in_bits = 1;
defparam ram_block1a90.data_interleave_width_in_bits = 1;
defparam ram_block1a90.init_file = "DDS_48_v1_nco_ii_0_sin.hex";
defparam ram_block1a90.init_file_layout = "port_a";
defparam ram_block1a90.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_c8g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a90.operation_mode = "rom";
defparam ram_block1a90.port_a_address_clear = "none";
defparam ram_block1a90.port_a_address_width = 13;
defparam ram_block1a90.port_a_data_out_clear = "none";
defparam ram_block1a90.port_a_data_out_clock = "clock0";
defparam ram_block1a90.port_a_data_width = 1;
defparam ram_block1a90.port_a_first_address = 40960;
defparam ram_block1a90.port_a_first_bit_number = 10;
defparam ram_block1a90.port_a_last_address = 49151;
defparam ram_block1a90.port_a_logical_ram_depth = 65536;
defparam ram_block1a90.port_a_logical_ram_width = 16;
defparam ram_block1a90.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a90.ram_block_type = "auto";
defparam ram_block1a90.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a90.mem_init2 = "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a90.mem_init1 = "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a90.mem_init0 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

arriav_ram_block ram_block1a106(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a106_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a106.clk0_core_clock_enable = "ena0";
defparam ram_block1a106.clk0_input_clock_enable = "ena0";
defparam ram_block1a106.clk0_output_clock_enable = "ena0";
defparam ram_block1a106.data_interleave_offset_in_bits = 1;
defparam ram_block1a106.data_interleave_width_in_bits = 1;
defparam ram_block1a106.init_file = "DDS_48_v1_nco_ii_0_sin.hex";
defparam ram_block1a106.init_file_layout = "port_a";
defparam ram_block1a106.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_c8g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a106.operation_mode = "rom";
defparam ram_block1a106.port_a_address_clear = "none";
defparam ram_block1a106.port_a_address_width = 13;
defparam ram_block1a106.port_a_data_out_clear = "none";
defparam ram_block1a106.port_a_data_out_clock = "clock0";
defparam ram_block1a106.port_a_data_width = 1;
defparam ram_block1a106.port_a_first_address = 49152;
defparam ram_block1a106.port_a_first_bit_number = 10;
defparam ram_block1a106.port_a_last_address = 57343;
defparam ram_block1a106.port_a_logical_ram_depth = 65536;
defparam ram_block1a106.port_a_logical_ram_width = 16;
defparam ram_block1a106.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a106.ram_block_type = "auto";
defparam ram_block1a106.mem_init3 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a106.mem_init2 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a106.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a106.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

arriav_ram_block ram_block1a122(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a122_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a122.clk0_core_clock_enable = "ena0";
defparam ram_block1a122.clk0_input_clock_enable = "ena0";
defparam ram_block1a122.clk0_output_clock_enable = "ena0";
defparam ram_block1a122.data_interleave_offset_in_bits = 1;
defparam ram_block1a122.data_interleave_width_in_bits = 1;
defparam ram_block1a122.init_file = "DDS_48_v1_nco_ii_0_sin.hex";
defparam ram_block1a122.init_file_layout = "port_a";
defparam ram_block1a122.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_c8g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a122.operation_mode = "rom";
defparam ram_block1a122.port_a_address_clear = "none";
defparam ram_block1a122.port_a_address_width = 13;
defparam ram_block1a122.port_a_data_out_clear = "none";
defparam ram_block1a122.port_a_data_out_clock = "clock0";
defparam ram_block1a122.port_a_data_width = 1;
defparam ram_block1a122.port_a_first_address = 57344;
defparam ram_block1a122.port_a_first_bit_number = 10;
defparam ram_block1a122.port_a_last_address = 65535;
defparam ram_block1a122.port_a_logical_ram_depth = 65536;
defparam ram_block1a122.port_a_logical_ram_width = 16;
defparam ram_block1a122.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a122.ram_block_type = "auto";
defparam ram_block1a122.mem_init3 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000000000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a122.mem_init2 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000000000000000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000000000000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a122.mem_init1 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a122.mem_init0 = "0000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

arriav_ram_block ram_block1a42(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a42_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a42.clk0_core_clock_enable = "ena0";
defparam ram_block1a42.clk0_input_clock_enable = "ena0";
defparam ram_block1a42.clk0_output_clock_enable = "ena0";
defparam ram_block1a42.data_interleave_offset_in_bits = 1;
defparam ram_block1a42.data_interleave_width_in_bits = 1;
defparam ram_block1a42.init_file = "DDS_48_v1_nco_ii_0_sin.hex";
defparam ram_block1a42.init_file_layout = "port_a";
defparam ram_block1a42.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_c8g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a42.operation_mode = "rom";
defparam ram_block1a42.port_a_address_clear = "none";
defparam ram_block1a42.port_a_address_width = 13;
defparam ram_block1a42.port_a_data_out_clear = "none";
defparam ram_block1a42.port_a_data_out_clock = "clock0";
defparam ram_block1a42.port_a_data_width = 1;
defparam ram_block1a42.port_a_first_address = 16384;
defparam ram_block1a42.port_a_first_bit_number = 10;
defparam ram_block1a42.port_a_last_address = 24575;
defparam ram_block1a42.port_a_logical_ram_depth = 65536;
defparam ram_block1a42.port_a_logical_ram_width = 16;
defparam ram_block1a42.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a42.ram_block_type = "auto";
defparam ram_block1a42.mem_init3 = "00000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a42.mem_init2 = "00000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a42.mem_init1 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a42.mem_init0 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

arriav_ram_block ram_block1a58(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a58_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a58.clk0_core_clock_enable = "ena0";
defparam ram_block1a58.clk0_input_clock_enable = "ena0";
defparam ram_block1a58.clk0_output_clock_enable = "ena0";
defparam ram_block1a58.data_interleave_offset_in_bits = 1;
defparam ram_block1a58.data_interleave_width_in_bits = 1;
defparam ram_block1a58.init_file = "DDS_48_v1_nco_ii_0_sin.hex";
defparam ram_block1a58.init_file_layout = "port_a";
defparam ram_block1a58.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_c8g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a58.operation_mode = "rom";
defparam ram_block1a58.port_a_address_clear = "none";
defparam ram_block1a58.port_a_address_width = 13;
defparam ram_block1a58.port_a_data_out_clear = "none";
defparam ram_block1a58.port_a_data_out_clock = "clock0";
defparam ram_block1a58.port_a_data_width = 1;
defparam ram_block1a58.port_a_first_address = 24576;
defparam ram_block1a58.port_a_first_bit_number = 10;
defparam ram_block1a58.port_a_last_address = 32767;
defparam ram_block1a58.port_a_logical_ram_depth = 65536;
defparam ram_block1a58.port_a_logical_ram_width = 16;
defparam ram_block1a58.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a58.ram_block_type = "auto";
defparam ram_block1a58.mem_init3 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000000000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000";
defparam ram_block1a58.mem_init2 = "000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000000000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000";
defparam ram_block1a58.mem_init1 = "0000000000000000000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a58.mem_init0 = "FFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000000000000000000000000000000000000000000000";

arriav_ram_block ram_block1a10(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a10_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a10.clk0_core_clock_enable = "ena0";
defparam ram_block1a10.clk0_input_clock_enable = "ena0";
defparam ram_block1a10.clk0_output_clock_enable = "ena0";
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.init_file = "DDS_48_v1_nco_ii_0_sin.hex";
defparam ram_block1a10.init_file_layout = "port_a";
defparam ram_block1a10.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_c8g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a10.operation_mode = "rom";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 13;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "clock0";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 8191;
defparam ram_block1a10.port_a_logical_ram_depth = 65536;
defparam ram_block1a10.port_a_logical_ram_width = 16;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a10.ram_block_type = "auto";
defparam ram_block1a10.mem_init3 = "000000000000000000000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a10.mem_init2 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a10.mem_init1 = "0000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000000000000000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a10.mem_init0 = "00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000000000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000000000000000000000000000000000000000000000000000000000";

arriav_ram_block ram_block1a26(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a26_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a26.clk0_core_clock_enable = "ena0";
defparam ram_block1a26.clk0_input_clock_enable = "ena0";
defparam ram_block1a26.clk0_output_clock_enable = "ena0";
defparam ram_block1a26.data_interleave_offset_in_bits = 1;
defparam ram_block1a26.data_interleave_width_in_bits = 1;
defparam ram_block1a26.init_file = "DDS_48_v1_nco_ii_0_sin.hex";
defparam ram_block1a26.init_file_layout = "port_a";
defparam ram_block1a26.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_c8g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a26.operation_mode = "rom";
defparam ram_block1a26.port_a_address_clear = "none";
defparam ram_block1a26.port_a_address_width = 13;
defparam ram_block1a26.port_a_data_out_clear = "none";
defparam ram_block1a26.port_a_data_out_clock = "clock0";
defparam ram_block1a26.port_a_data_width = 1;
defparam ram_block1a26.port_a_first_address = 8192;
defparam ram_block1a26.port_a_first_bit_number = 10;
defparam ram_block1a26.port_a_last_address = 16383;
defparam ram_block1a26.port_a_logical_ram_depth = 65536;
defparam ram_block1a26.port_a_logical_ram_width = 16;
defparam ram_block1a26.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a26.ram_block_type = "auto";
defparam ram_block1a26.mem_init3 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a26.mem_init2 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a26.mem_init1 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a26.mem_init0 = "000000000000000000000000000000000000000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000000000000000000000";

arriav_ram_block ram_block1a75(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a75_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a75.clk0_core_clock_enable = "ena0";
defparam ram_block1a75.clk0_input_clock_enable = "ena0";
defparam ram_block1a75.clk0_output_clock_enable = "ena0";
defparam ram_block1a75.data_interleave_offset_in_bits = 1;
defparam ram_block1a75.data_interleave_width_in_bits = 1;
defparam ram_block1a75.init_file = "DDS_48_v1_nco_ii_0_sin.hex";
defparam ram_block1a75.init_file_layout = "port_a";
defparam ram_block1a75.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_c8g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a75.operation_mode = "rom";
defparam ram_block1a75.port_a_address_clear = "none";
defparam ram_block1a75.port_a_address_width = 13;
defparam ram_block1a75.port_a_data_out_clear = "none";
defparam ram_block1a75.port_a_data_out_clock = "clock0";
defparam ram_block1a75.port_a_data_width = 1;
defparam ram_block1a75.port_a_first_address = 32768;
defparam ram_block1a75.port_a_first_bit_number = 11;
defparam ram_block1a75.port_a_last_address = 40959;
defparam ram_block1a75.port_a_logical_ram_depth = 65536;
defparam ram_block1a75.port_a_logical_ram_width = 16;
defparam ram_block1a75.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a75.ram_block_type = "auto";
defparam ram_block1a75.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a75.mem_init2 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a75.mem_init1 = "FFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a75.mem_init0 = "00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE";

arriav_ram_block ram_block1a91(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a91_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a91.clk0_core_clock_enable = "ena0";
defparam ram_block1a91.clk0_input_clock_enable = "ena0";
defparam ram_block1a91.clk0_output_clock_enable = "ena0";
defparam ram_block1a91.data_interleave_offset_in_bits = 1;
defparam ram_block1a91.data_interleave_width_in_bits = 1;
defparam ram_block1a91.init_file = "DDS_48_v1_nco_ii_0_sin.hex";
defparam ram_block1a91.init_file_layout = "port_a";
defparam ram_block1a91.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_c8g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a91.operation_mode = "rom";
defparam ram_block1a91.port_a_address_clear = "none";
defparam ram_block1a91.port_a_address_width = 13;
defparam ram_block1a91.port_a_data_out_clear = "none";
defparam ram_block1a91.port_a_data_out_clock = "clock0";
defparam ram_block1a91.port_a_data_width = 1;
defparam ram_block1a91.port_a_first_address = 40960;
defparam ram_block1a91.port_a_first_bit_number = 11;
defparam ram_block1a91.port_a_last_address = 49151;
defparam ram_block1a91.port_a_logical_ram_depth = 65536;
defparam ram_block1a91.port_a_logical_ram_width = 16;
defparam ram_block1a91.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a91.ram_block_type = "auto";
defparam ram_block1a91.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a91.mem_init2 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a91.mem_init1 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a91.mem_init0 = "000000000000000000000000000000000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

arriav_ram_block ram_block1a107(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a107_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a107.clk0_core_clock_enable = "ena0";
defparam ram_block1a107.clk0_input_clock_enable = "ena0";
defparam ram_block1a107.clk0_output_clock_enable = "ena0";
defparam ram_block1a107.data_interleave_offset_in_bits = 1;
defparam ram_block1a107.data_interleave_width_in_bits = 1;
defparam ram_block1a107.init_file = "DDS_48_v1_nco_ii_0_sin.hex";
defparam ram_block1a107.init_file_layout = "port_a";
defparam ram_block1a107.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_c8g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a107.operation_mode = "rom";
defparam ram_block1a107.port_a_address_clear = "none";
defparam ram_block1a107.port_a_address_width = 13;
defparam ram_block1a107.port_a_data_out_clear = "none";
defparam ram_block1a107.port_a_data_out_clock = "clock0";
defparam ram_block1a107.port_a_data_width = 1;
defparam ram_block1a107.port_a_first_address = 49152;
defparam ram_block1a107.port_a_first_bit_number = 11;
defparam ram_block1a107.port_a_last_address = 57343;
defparam ram_block1a107.port_a_logical_ram_depth = 65536;
defparam ram_block1a107.port_a_logical_ram_width = 16;
defparam ram_block1a107.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a107.ram_block_type = "auto";
defparam ram_block1a107.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a107.mem_init2 = "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a107.mem_init1 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a107.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

arriav_ram_block ram_block1a123(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a123_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a123.clk0_core_clock_enable = "ena0";
defparam ram_block1a123.clk0_input_clock_enable = "ena0";
defparam ram_block1a123.clk0_output_clock_enable = "ena0";
defparam ram_block1a123.data_interleave_offset_in_bits = 1;
defparam ram_block1a123.data_interleave_width_in_bits = 1;
defparam ram_block1a123.init_file = "DDS_48_v1_nco_ii_0_sin.hex";
defparam ram_block1a123.init_file_layout = "port_a";
defparam ram_block1a123.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_c8g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a123.operation_mode = "rom";
defparam ram_block1a123.port_a_address_clear = "none";
defparam ram_block1a123.port_a_address_width = 13;
defparam ram_block1a123.port_a_data_out_clear = "none";
defparam ram_block1a123.port_a_data_out_clock = "clock0";
defparam ram_block1a123.port_a_data_width = 1;
defparam ram_block1a123.port_a_first_address = 57344;
defparam ram_block1a123.port_a_first_bit_number = 11;
defparam ram_block1a123.port_a_last_address = 65535;
defparam ram_block1a123.port_a_logical_ram_depth = 65536;
defparam ram_block1a123.port_a_logical_ram_width = 16;
defparam ram_block1a123.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a123.ram_block_type = "auto";
defparam ram_block1a123.mem_init3 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000";
defparam ram_block1a123.mem_init2 = "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a123.mem_init1 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a123.mem_init0 = "FFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000000000000000000000000000000000000000";

arriav_ram_block ram_block1a43(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a43_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a43.clk0_core_clock_enable = "ena0";
defparam ram_block1a43.clk0_input_clock_enable = "ena0";
defparam ram_block1a43.clk0_output_clock_enable = "ena0";
defparam ram_block1a43.data_interleave_offset_in_bits = 1;
defparam ram_block1a43.data_interleave_width_in_bits = 1;
defparam ram_block1a43.init_file = "DDS_48_v1_nco_ii_0_sin.hex";
defparam ram_block1a43.init_file_layout = "port_a";
defparam ram_block1a43.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_c8g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a43.operation_mode = "rom";
defparam ram_block1a43.port_a_address_clear = "none";
defparam ram_block1a43.port_a_address_width = 13;
defparam ram_block1a43.port_a_data_out_clear = "none";
defparam ram_block1a43.port_a_data_out_clock = "clock0";
defparam ram_block1a43.port_a_data_width = 1;
defparam ram_block1a43.port_a_first_address = 16384;
defparam ram_block1a43.port_a_first_bit_number = 11;
defparam ram_block1a43.port_a_last_address = 24575;
defparam ram_block1a43.port_a_logical_ram_depth = 65536;
defparam ram_block1a43.port_a_logical_ram_width = 16;
defparam ram_block1a43.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a43.ram_block_type = "auto";
defparam ram_block1a43.mem_init3 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a43.mem_init2 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a43.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a43.mem_init0 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

arriav_ram_block ram_block1a59(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a59_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a59.clk0_core_clock_enable = "ena0";
defparam ram_block1a59.clk0_input_clock_enable = "ena0";
defparam ram_block1a59.clk0_output_clock_enable = "ena0";
defparam ram_block1a59.data_interleave_offset_in_bits = 1;
defparam ram_block1a59.data_interleave_width_in_bits = 1;
defparam ram_block1a59.init_file = "DDS_48_v1_nco_ii_0_sin.hex";
defparam ram_block1a59.init_file_layout = "port_a";
defparam ram_block1a59.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_c8g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a59.operation_mode = "rom";
defparam ram_block1a59.port_a_address_clear = "none";
defparam ram_block1a59.port_a_address_width = 13;
defparam ram_block1a59.port_a_data_out_clear = "none";
defparam ram_block1a59.port_a_data_out_clock = "clock0";
defparam ram_block1a59.port_a_data_width = 1;
defparam ram_block1a59.port_a_first_address = 24576;
defparam ram_block1a59.port_a_first_bit_number = 11;
defparam ram_block1a59.port_a_last_address = 32767;
defparam ram_block1a59.port_a_logical_ram_depth = 65536;
defparam ram_block1a59.port_a_logical_ram_width = 16;
defparam ram_block1a59.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a59.ram_block_type = "auto";
defparam ram_block1a59.mem_init3 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a59.mem_init2 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000";
defparam ram_block1a59.mem_init1 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a59.mem_init0 = "0000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

arriav_ram_block ram_block1a11(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a11_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a11.clk0_core_clock_enable = "ena0";
defparam ram_block1a11.clk0_input_clock_enable = "ena0";
defparam ram_block1a11.clk0_output_clock_enable = "ena0";
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.init_file = "DDS_48_v1_nco_ii_0_sin.hex";
defparam ram_block1a11.init_file_layout = "port_a";
defparam ram_block1a11.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_c8g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a11.operation_mode = "rom";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 13;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "clock0";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 8191;
defparam ram_block1a11.port_a_logical_ram_depth = 65536;
defparam ram_block1a11.port_a_logical_ram_width = 16;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a11.ram_block_type = "auto";
defparam ram_block1a11.mem_init3 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000";
defparam ram_block1a11.mem_init2 = "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a11.mem_init1 = "0000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a11.mem_init0 = "FFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

arriav_ram_block ram_block1a27(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a27_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a27.clk0_core_clock_enable = "ena0";
defparam ram_block1a27.clk0_input_clock_enable = "ena0";
defparam ram_block1a27.clk0_output_clock_enable = "ena0";
defparam ram_block1a27.data_interleave_offset_in_bits = 1;
defparam ram_block1a27.data_interleave_width_in_bits = 1;
defparam ram_block1a27.init_file = "DDS_48_v1_nco_ii_0_sin.hex";
defparam ram_block1a27.init_file_layout = "port_a";
defparam ram_block1a27.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_c8g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a27.operation_mode = "rom";
defparam ram_block1a27.port_a_address_clear = "none";
defparam ram_block1a27.port_a_address_width = 13;
defparam ram_block1a27.port_a_data_out_clear = "none";
defparam ram_block1a27.port_a_data_out_clock = "clock0";
defparam ram_block1a27.port_a_data_width = 1;
defparam ram_block1a27.port_a_first_address = 8192;
defparam ram_block1a27.port_a_first_bit_number = 11;
defparam ram_block1a27.port_a_last_address = 16383;
defparam ram_block1a27.port_a_logical_ram_depth = 65536;
defparam ram_block1a27.port_a_logical_ram_width = 16;
defparam ram_block1a27.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a27.ram_block_type = "auto";
defparam ram_block1a27.mem_init3 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a27.mem_init2 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a27.mem_init1 = "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a27.mem_init0 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

arriav_ram_block ram_block1a76(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a76_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a76.clk0_core_clock_enable = "ena0";
defparam ram_block1a76.clk0_input_clock_enable = "ena0";
defparam ram_block1a76.clk0_output_clock_enable = "ena0";
defparam ram_block1a76.data_interleave_offset_in_bits = 1;
defparam ram_block1a76.data_interleave_width_in_bits = 1;
defparam ram_block1a76.init_file = "DDS_48_v1_nco_ii_0_sin.hex";
defparam ram_block1a76.init_file_layout = "port_a";
defparam ram_block1a76.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_c8g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a76.operation_mode = "rom";
defparam ram_block1a76.port_a_address_clear = "none";
defparam ram_block1a76.port_a_address_width = 13;
defparam ram_block1a76.port_a_data_out_clear = "none";
defparam ram_block1a76.port_a_data_out_clock = "clock0";
defparam ram_block1a76.port_a_data_width = 1;
defparam ram_block1a76.port_a_first_address = 32768;
defparam ram_block1a76.port_a_first_bit_number = 12;
defparam ram_block1a76.port_a_last_address = 40959;
defparam ram_block1a76.port_a_logical_ram_depth = 65536;
defparam ram_block1a76.port_a_logical_ram_width = 16;
defparam ram_block1a76.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a76.ram_block_type = "auto";
defparam ram_block1a76.mem_init3 = "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a76.mem_init2 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a76.mem_init1 = "0000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a76.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE";

arriav_ram_block ram_block1a92(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a92_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a92.clk0_core_clock_enable = "ena0";
defparam ram_block1a92.clk0_input_clock_enable = "ena0";
defparam ram_block1a92.clk0_output_clock_enable = "ena0";
defparam ram_block1a92.data_interleave_offset_in_bits = 1;
defparam ram_block1a92.data_interleave_width_in_bits = 1;
defparam ram_block1a92.init_file = "DDS_48_v1_nco_ii_0_sin.hex";
defparam ram_block1a92.init_file_layout = "port_a";
defparam ram_block1a92.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_c8g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a92.operation_mode = "rom";
defparam ram_block1a92.port_a_address_clear = "none";
defparam ram_block1a92.port_a_address_width = 13;
defparam ram_block1a92.port_a_data_out_clear = "none";
defparam ram_block1a92.port_a_data_out_clock = "clock0";
defparam ram_block1a92.port_a_data_width = 1;
defparam ram_block1a92.port_a_first_address = 40960;
defparam ram_block1a92.port_a_first_bit_number = 12;
defparam ram_block1a92.port_a_last_address = 49151;
defparam ram_block1a92.port_a_logical_ram_depth = 65536;
defparam ram_block1a92.port_a_logical_ram_width = 16;
defparam ram_block1a92.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a92.ram_block_type = "auto";
defparam ram_block1a92.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a92.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a92.mem_init1 = "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a92.mem_init0 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

arriav_ram_block ram_block1a108(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a108_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a108.clk0_core_clock_enable = "ena0";
defparam ram_block1a108.clk0_input_clock_enable = "ena0";
defparam ram_block1a108.clk0_output_clock_enable = "ena0";
defparam ram_block1a108.data_interleave_offset_in_bits = 1;
defparam ram_block1a108.data_interleave_width_in_bits = 1;
defparam ram_block1a108.init_file = "DDS_48_v1_nco_ii_0_sin.hex";
defparam ram_block1a108.init_file_layout = "port_a";
defparam ram_block1a108.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_c8g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a108.operation_mode = "rom";
defparam ram_block1a108.port_a_address_clear = "none";
defparam ram_block1a108.port_a_address_width = 13;
defparam ram_block1a108.port_a_data_out_clear = "none";
defparam ram_block1a108.port_a_data_out_clock = "clock0";
defparam ram_block1a108.port_a_data_width = 1;
defparam ram_block1a108.port_a_first_address = 49152;
defparam ram_block1a108.port_a_first_bit_number = 12;
defparam ram_block1a108.port_a_last_address = 57343;
defparam ram_block1a108.port_a_logical_ram_depth = 65536;
defparam ram_block1a108.port_a_logical_ram_width = 16;
defparam ram_block1a108.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a108.ram_block_type = "auto";
defparam ram_block1a108.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a108.mem_init2 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a108.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a108.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

arriav_ram_block ram_block1a124(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a124_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a124.clk0_core_clock_enable = "ena0";
defparam ram_block1a124.clk0_input_clock_enable = "ena0";
defparam ram_block1a124.clk0_output_clock_enable = "ena0";
defparam ram_block1a124.data_interleave_offset_in_bits = 1;
defparam ram_block1a124.data_interleave_width_in_bits = 1;
defparam ram_block1a124.init_file = "DDS_48_v1_nco_ii_0_sin.hex";
defparam ram_block1a124.init_file_layout = "port_a";
defparam ram_block1a124.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_c8g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a124.operation_mode = "rom";
defparam ram_block1a124.port_a_address_clear = "none";
defparam ram_block1a124.port_a_address_width = 13;
defparam ram_block1a124.port_a_data_out_clear = "none";
defparam ram_block1a124.port_a_data_out_clock = "clock0";
defparam ram_block1a124.port_a_data_width = 1;
defparam ram_block1a124.port_a_first_address = 57344;
defparam ram_block1a124.port_a_first_bit_number = 12;
defparam ram_block1a124.port_a_last_address = 65535;
defparam ram_block1a124.port_a_logical_ram_depth = 65536;
defparam ram_block1a124.port_a_logical_ram_width = 16;
defparam ram_block1a124.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a124.ram_block_type = "auto";
defparam ram_block1a124.mem_init3 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a124.mem_init2 = "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000";
defparam ram_block1a124.mem_init1 = "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a124.mem_init0 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

arriav_ram_block ram_block1a44(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a44_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a44.clk0_core_clock_enable = "ena0";
defparam ram_block1a44.clk0_input_clock_enable = "ena0";
defparam ram_block1a44.clk0_output_clock_enable = "ena0";
defparam ram_block1a44.data_interleave_offset_in_bits = 1;
defparam ram_block1a44.data_interleave_width_in_bits = 1;
defparam ram_block1a44.init_file = "DDS_48_v1_nco_ii_0_sin.hex";
defparam ram_block1a44.init_file_layout = "port_a";
defparam ram_block1a44.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_c8g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a44.operation_mode = "rom";
defparam ram_block1a44.port_a_address_clear = "none";
defparam ram_block1a44.port_a_address_width = 13;
defparam ram_block1a44.port_a_data_out_clear = "none";
defparam ram_block1a44.port_a_data_out_clock = "clock0";
defparam ram_block1a44.port_a_data_width = 1;
defparam ram_block1a44.port_a_first_address = 16384;
defparam ram_block1a44.port_a_first_bit_number = 12;
defparam ram_block1a44.port_a_last_address = 24575;
defparam ram_block1a44.port_a_logical_ram_depth = 65536;
defparam ram_block1a44.port_a_logical_ram_width = 16;
defparam ram_block1a44.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a44.ram_block_type = "auto";
defparam ram_block1a44.mem_init3 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a44.mem_init2 = "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a44.mem_init1 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a44.mem_init0 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

arriav_ram_block ram_block1a60(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a60_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a60.clk0_core_clock_enable = "ena0";
defparam ram_block1a60.clk0_input_clock_enable = "ena0";
defparam ram_block1a60.clk0_output_clock_enable = "ena0";
defparam ram_block1a60.data_interleave_offset_in_bits = 1;
defparam ram_block1a60.data_interleave_width_in_bits = 1;
defparam ram_block1a60.init_file = "DDS_48_v1_nco_ii_0_sin.hex";
defparam ram_block1a60.init_file_layout = "port_a";
defparam ram_block1a60.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_c8g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a60.operation_mode = "rom";
defparam ram_block1a60.port_a_address_clear = "none";
defparam ram_block1a60.port_a_address_width = 13;
defparam ram_block1a60.port_a_data_out_clear = "none";
defparam ram_block1a60.port_a_data_out_clock = "clock0";
defparam ram_block1a60.port_a_data_width = 1;
defparam ram_block1a60.port_a_first_address = 24576;
defparam ram_block1a60.port_a_first_bit_number = 12;
defparam ram_block1a60.port_a_last_address = 32767;
defparam ram_block1a60.port_a_logical_ram_depth = 65536;
defparam ram_block1a60.port_a_logical_ram_width = 16;
defparam ram_block1a60.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a60.ram_block_type = "auto";
defparam ram_block1a60.mem_init3 = "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a60.mem_init2 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a60.mem_init1 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a60.mem_init0 = "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

arriav_ram_block ram_block1a12(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a12_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a12.clk0_core_clock_enable = "ena0";
defparam ram_block1a12.clk0_input_clock_enable = "ena0";
defparam ram_block1a12.clk0_output_clock_enable = "ena0";
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.init_file = "DDS_48_v1_nco_ii_0_sin.hex";
defparam ram_block1a12.init_file_layout = "port_a";
defparam ram_block1a12.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_c8g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a12.operation_mode = "rom";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 13;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "clock0";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 8191;
defparam ram_block1a12.port_a_logical_ram_depth = 65536;
defparam ram_block1a12.port_a_logical_ram_width = 16;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a12.ram_block_type = "auto";
defparam ram_block1a12.mem_init3 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a12.mem_init2 = "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a12.mem_init1 = "FFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a12.mem_init0 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

arriav_ram_block ram_block1a28(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a28_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a28.clk0_core_clock_enable = "ena0";
defparam ram_block1a28.clk0_input_clock_enable = "ena0";
defparam ram_block1a28.clk0_output_clock_enable = "ena0";
defparam ram_block1a28.data_interleave_offset_in_bits = 1;
defparam ram_block1a28.data_interleave_width_in_bits = 1;
defparam ram_block1a28.init_file = "DDS_48_v1_nco_ii_0_sin.hex";
defparam ram_block1a28.init_file_layout = "port_a";
defparam ram_block1a28.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_c8g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a28.operation_mode = "rom";
defparam ram_block1a28.port_a_address_clear = "none";
defparam ram_block1a28.port_a_address_width = 13;
defparam ram_block1a28.port_a_data_out_clear = "none";
defparam ram_block1a28.port_a_data_out_clock = "clock0";
defparam ram_block1a28.port_a_data_width = 1;
defparam ram_block1a28.port_a_first_address = 8192;
defparam ram_block1a28.port_a_first_bit_number = 12;
defparam ram_block1a28.port_a_last_address = 16383;
defparam ram_block1a28.port_a_logical_ram_depth = 65536;
defparam ram_block1a28.port_a_logical_ram_width = 16;
defparam ram_block1a28.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a28.ram_block_type = "auto";
defparam ram_block1a28.mem_init3 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a28.mem_init2 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a28.mem_init1 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a28.mem_init0 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

arriav_ram_block ram_block1a77(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a77_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a77.clk0_core_clock_enable = "ena0";
defparam ram_block1a77.clk0_input_clock_enable = "ena0";
defparam ram_block1a77.clk0_output_clock_enable = "ena0";
defparam ram_block1a77.data_interleave_offset_in_bits = 1;
defparam ram_block1a77.data_interleave_width_in_bits = 1;
defparam ram_block1a77.init_file = "DDS_48_v1_nco_ii_0_sin.hex";
defparam ram_block1a77.init_file_layout = "port_a";
defparam ram_block1a77.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_c8g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a77.operation_mode = "rom";
defparam ram_block1a77.port_a_address_clear = "none";
defparam ram_block1a77.port_a_address_width = 13;
defparam ram_block1a77.port_a_data_out_clear = "none";
defparam ram_block1a77.port_a_data_out_clock = "clock0";
defparam ram_block1a77.port_a_data_width = 1;
defparam ram_block1a77.port_a_first_address = 32768;
defparam ram_block1a77.port_a_first_bit_number = 13;
defparam ram_block1a77.port_a_last_address = 40959;
defparam ram_block1a77.port_a_logical_ram_depth = 65536;
defparam ram_block1a77.port_a_logical_ram_width = 16;
defparam ram_block1a77.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a77.ram_block_type = "auto";
defparam ram_block1a77.mem_init3 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a77.mem_init2 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a77.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a77.mem_init0 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE";

arriav_ram_block ram_block1a93(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a93_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a93.clk0_core_clock_enable = "ena0";
defparam ram_block1a93.clk0_input_clock_enable = "ena0";
defparam ram_block1a93.clk0_output_clock_enable = "ena0";
defparam ram_block1a93.data_interleave_offset_in_bits = 1;
defparam ram_block1a93.data_interleave_width_in_bits = 1;
defparam ram_block1a93.init_file = "DDS_48_v1_nco_ii_0_sin.hex";
defparam ram_block1a93.init_file_layout = "port_a";
defparam ram_block1a93.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_c8g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a93.operation_mode = "rom";
defparam ram_block1a93.port_a_address_clear = "none";
defparam ram_block1a93.port_a_address_width = 13;
defparam ram_block1a93.port_a_data_out_clear = "none";
defparam ram_block1a93.port_a_data_out_clock = "clock0";
defparam ram_block1a93.port_a_data_width = 1;
defparam ram_block1a93.port_a_first_address = 40960;
defparam ram_block1a93.port_a_first_bit_number = 13;
defparam ram_block1a93.port_a_last_address = 49151;
defparam ram_block1a93.port_a_logical_ram_depth = 65536;
defparam ram_block1a93.port_a_logical_ram_width = 16;
defparam ram_block1a93.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a93.ram_block_type = "auto";
defparam ram_block1a93.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a93.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a93.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a93.mem_init0 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

arriav_ram_block ram_block1a109(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a109_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a109.clk0_core_clock_enable = "ena0";
defparam ram_block1a109.clk0_input_clock_enable = "ena0";
defparam ram_block1a109.clk0_output_clock_enable = "ena0";
defparam ram_block1a109.data_interleave_offset_in_bits = 1;
defparam ram_block1a109.data_interleave_width_in_bits = 1;
defparam ram_block1a109.init_file = "DDS_48_v1_nco_ii_0_sin.hex";
defparam ram_block1a109.init_file_layout = "port_a";
defparam ram_block1a109.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_c8g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a109.operation_mode = "rom";
defparam ram_block1a109.port_a_address_clear = "none";
defparam ram_block1a109.port_a_address_width = 13;
defparam ram_block1a109.port_a_data_out_clear = "none";
defparam ram_block1a109.port_a_data_out_clock = "clock0";
defparam ram_block1a109.port_a_data_width = 1;
defparam ram_block1a109.port_a_first_address = 49152;
defparam ram_block1a109.port_a_first_bit_number = 13;
defparam ram_block1a109.port_a_last_address = 57343;
defparam ram_block1a109.port_a_logical_ram_depth = 65536;
defparam ram_block1a109.port_a_logical_ram_width = 16;
defparam ram_block1a109.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a109.ram_block_type = "auto";
defparam ram_block1a109.mem_init3 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a109.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a109.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a109.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

arriav_ram_block ram_block1a125(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a125_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a125.clk0_core_clock_enable = "ena0";
defparam ram_block1a125.clk0_input_clock_enable = "ena0";
defparam ram_block1a125.clk0_output_clock_enable = "ena0";
defparam ram_block1a125.data_interleave_offset_in_bits = 1;
defparam ram_block1a125.data_interleave_width_in_bits = 1;
defparam ram_block1a125.init_file = "DDS_48_v1_nco_ii_0_sin.hex";
defparam ram_block1a125.init_file_layout = "port_a";
defparam ram_block1a125.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_c8g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a125.operation_mode = "rom";
defparam ram_block1a125.port_a_address_clear = "none";
defparam ram_block1a125.port_a_address_width = 13;
defparam ram_block1a125.port_a_data_out_clear = "none";
defparam ram_block1a125.port_a_data_out_clock = "clock0";
defparam ram_block1a125.port_a_data_width = 1;
defparam ram_block1a125.port_a_first_address = 57344;
defparam ram_block1a125.port_a_first_bit_number = 13;
defparam ram_block1a125.port_a_last_address = 65535;
defparam ram_block1a125.port_a_logical_ram_depth = 65536;
defparam ram_block1a125.port_a_logical_ram_width = 16;
defparam ram_block1a125.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a125.ram_block_type = "auto";
defparam ram_block1a125.mem_init3 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a125.mem_init2 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a125.mem_init1 = "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a125.mem_init0 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

arriav_ram_block ram_block1a45(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a45_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a45.clk0_core_clock_enable = "ena0";
defparam ram_block1a45.clk0_input_clock_enable = "ena0";
defparam ram_block1a45.clk0_output_clock_enable = "ena0";
defparam ram_block1a45.data_interleave_offset_in_bits = 1;
defparam ram_block1a45.data_interleave_width_in_bits = 1;
defparam ram_block1a45.init_file = "DDS_48_v1_nco_ii_0_sin.hex";
defparam ram_block1a45.init_file_layout = "port_a";
defparam ram_block1a45.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_c8g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a45.operation_mode = "rom";
defparam ram_block1a45.port_a_address_clear = "none";
defparam ram_block1a45.port_a_address_width = 13;
defparam ram_block1a45.port_a_data_out_clear = "none";
defparam ram_block1a45.port_a_data_out_clock = "clock0";
defparam ram_block1a45.port_a_data_width = 1;
defparam ram_block1a45.port_a_first_address = 16384;
defparam ram_block1a45.port_a_first_bit_number = 13;
defparam ram_block1a45.port_a_last_address = 24575;
defparam ram_block1a45.port_a_logical_ram_depth = 65536;
defparam ram_block1a45.port_a_logical_ram_width = 16;
defparam ram_block1a45.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a45.ram_block_type = "auto";
defparam ram_block1a45.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a45.mem_init2 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a45.mem_init1 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a45.mem_init0 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

arriav_ram_block ram_block1a61(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a61_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a61.clk0_core_clock_enable = "ena0";
defparam ram_block1a61.clk0_input_clock_enable = "ena0";
defparam ram_block1a61.clk0_output_clock_enable = "ena0";
defparam ram_block1a61.data_interleave_offset_in_bits = 1;
defparam ram_block1a61.data_interleave_width_in_bits = 1;
defparam ram_block1a61.init_file = "DDS_48_v1_nco_ii_0_sin.hex";
defparam ram_block1a61.init_file_layout = "port_a";
defparam ram_block1a61.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_c8g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a61.operation_mode = "rom";
defparam ram_block1a61.port_a_address_clear = "none";
defparam ram_block1a61.port_a_address_width = 13;
defparam ram_block1a61.port_a_data_out_clear = "none";
defparam ram_block1a61.port_a_data_out_clock = "clock0";
defparam ram_block1a61.port_a_data_width = 1;
defparam ram_block1a61.port_a_first_address = 24576;
defparam ram_block1a61.port_a_first_bit_number = 13;
defparam ram_block1a61.port_a_last_address = 32767;
defparam ram_block1a61.port_a_logical_ram_depth = 65536;
defparam ram_block1a61.port_a_logical_ram_width = 16;
defparam ram_block1a61.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a61.ram_block_type = "auto";
defparam ram_block1a61.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a61.mem_init2 = "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a61.mem_init1 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a61.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

arriav_ram_block ram_block1a13(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a13_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a13.clk0_core_clock_enable = "ena0";
defparam ram_block1a13.clk0_input_clock_enable = "ena0";
defparam ram_block1a13.clk0_output_clock_enable = "ena0";
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.init_file = "DDS_48_v1_nco_ii_0_sin.hex";
defparam ram_block1a13.init_file_layout = "port_a";
defparam ram_block1a13.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_c8g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a13.operation_mode = "rom";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 13;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "clock0";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 8191;
defparam ram_block1a13.port_a_logical_ram_depth = 65536;
defparam ram_block1a13.port_a_logical_ram_width = 16;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a13.ram_block_type = "auto";
defparam ram_block1a13.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a13.mem_init2 = "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a13.mem_init1 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a13.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

arriav_ram_block ram_block1a29(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a29_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a29.clk0_core_clock_enable = "ena0";
defparam ram_block1a29.clk0_input_clock_enable = "ena0";
defparam ram_block1a29.clk0_output_clock_enable = "ena0";
defparam ram_block1a29.data_interleave_offset_in_bits = 1;
defparam ram_block1a29.data_interleave_width_in_bits = 1;
defparam ram_block1a29.init_file = "DDS_48_v1_nco_ii_0_sin.hex";
defparam ram_block1a29.init_file_layout = "port_a";
defparam ram_block1a29.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_c8g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a29.operation_mode = "rom";
defparam ram_block1a29.port_a_address_clear = "none";
defparam ram_block1a29.port_a_address_width = 13;
defparam ram_block1a29.port_a_data_out_clear = "none";
defparam ram_block1a29.port_a_data_out_clock = "clock0";
defparam ram_block1a29.port_a_data_width = 1;
defparam ram_block1a29.port_a_first_address = 8192;
defparam ram_block1a29.port_a_first_bit_number = 13;
defparam ram_block1a29.port_a_last_address = 16383;
defparam ram_block1a29.port_a_logical_ram_depth = 65536;
defparam ram_block1a29.port_a_logical_ram_width = 16;
defparam ram_block1a29.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a29.ram_block_type = "auto";
defparam ram_block1a29.mem_init3 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a29.mem_init2 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a29.mem_init1 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a29.mem_init0 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

arriav_ram_block ram_block1a78(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a78_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a78.clk0_core_clock_enable = "ena0";
defparam ram_block1a78.clk0_input_clock_enable = "ena0";
defparam ram_block1a78.clk0_output_clock_enable = "ena0";
defparam ram_block1a78.data_interleave_offset_in_bits = 1;
defparam ram_block1a78.data_interleave_width_in_bits = 1;
defparam ram_block1a78.init_file = "DDS_48_v1_nco_ii_0_sin.hex";
defparam ram_block1a78.init_file_layout = "port_a";
defparam ram_block1a78.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_c8g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a78.operation_mode = "rom";
defparam ram_block1a78.port_a_address_clear = "none";
defparam ram_block1a78.port_a_address_width = 13;
defparam ram_block1a78.port_a_data_out_clear = "none";
defparam ram_block1a78.port_a_data_out_clock = "clock0";
defparam ram_block1a78.port_a_data_width = 1;
defparam ram_block1a78.port_a_first_address = 32768;
defparam ram_block1a78.port_a_first_bit_number = 14;
defparam ram_block1a78.port_a_last_address = 40959;
defparam ram_block1a78.port_a_logical_ram_depth = 65536;
defparam ram_block1a78.port_a_logical_ram_width = 16;
defparam ram_block1a78.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a78.ram_block_type = "auto";
defparam ram_block1a78.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a78.mem_init2 = "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a78.mem_init1 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a78.mem_init0 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE";

arriav_ram_block ram_block1a94(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a94_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a94.clk0_core_clock_enable = "ena0";
defparam ram_block1a94.clk0_input_clock_enable = "ena0";
defparam ram_block1a94.clk0_output_clock_enable = "ena0";
defparam ram_block1a94.data_interleave_offset_in_bits = 1;
defparam ram_block1a94.data_interleave_width_in_bits = 1;
defparam ram_block1a94.init_file = "DDS_48_v1_nco_ii_0_sin.hex";
defparam ram_block1a94.init_file_layout = "port_a";
defparam ram_block1a94.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_c8g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a94.operation_mode = "rom";
defparam ram_block1a94.port_a_address_clear = "none";
defparam ram_block1a94.port_a_address_width = 13;
defparam ram_block1a94.port_a_data_out_clear = "none";
defparam ram_block1a94.port_a_data_out_clock = "clock0";
defparam ram_block1a94.port_a_data_width = 1;
defparam ram_block1a94.port_a_first_address = 40960;
defparam ram_block1a94.port_a_first_bit_number = 14;
defparam ram_block1a94.port_a_last_address = 49151;
defparam ram_block1a94.port_a_logical_ram_depth = 65536;
defparam ram_block1a94.port_a_logical_ram_width = 16;
defparam ram_block1a94.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a94.ram_block_type = "auto";
defparam ram_block1a94.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a94.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a94.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a94.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

arriav_ram_block ram_block1a110(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a110_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a110.clk0_core_clock_enable = "ena0";
defparam ram_block1a110.clk0_input_clock_enable = "ena0";
defparam ram_block1a110.clk0_output_clock_enable = "ena0";
defparam ram_block1a110.data_interleave_offset_in_bits = 1;
defparam ram_block1a110.data_interleave_width_in_bits = 1;
defparam ram_block1a110.init_file = "DDS_48_v1_nco_ii_0_sin.hex";
defparam ram_block1a110.init_file_layout = "port_a";
defparam ram_block1a110.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_c8g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a110.operation_mode = "rom";
defparam ram_block1a110.port_a_address_clear = "none";
defparam ram_block1a110.port_a_address_width = 13;
defparam ram_block1a110.port_a_data_out_clear = "none";
defparam ram_block1a110.port_a_data_out_clock = "clock0";
defparam ram_block1a110.port_a_data_width = 1;
defparam ram_block1a110.port_a_first_address = 49152;
defparam ram_block1a110.port_a_first_bit_number = 14;
defparam ram_block1a110.port_a_last_address = 57343;
defparam ram_block1a110.port_a_logical_ram_depth = 65536;
defparam ram_block1a110.port_a_logical_ram_width = 16;
defparam ram_block1a110.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a110.ram_block_type = "auto";
defparam ram_block1a110.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a110.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a110.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a110.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

arriav_ram_block ram_block1a126(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a126_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a126.clk0_core_clock_enable = "ena0";
defparam ram_block1a126.clk0_input_clock_enable = "ena0";
defparam ram_block1a126.clk0_output_clock_enable = "ena0";
defparam ram_block1a126.data_interleave_offset_in_bits = 1;
defparam ram_block1a126.data_interleave_width_in_bits = 1;
defparam ram_block1a126.init_file = "DDS_48_v1_nco_ii_0_sin.hex";
defparam ram_block1a126.init_file_layout = "port_a";
defparam ram_block1a126.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_c8g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a126.operation_mode = "rom";
defparam ram_block1a126.port_a_address_clear = "none";
defparam ram_block1a126.port_a_address_width = 13;
defparam ram_block1a126.port_a_data_out_clear = "none";
defparam ram_block1a126.port_a_data_out_clock = "clock0";
defparam ram_block1a126.port_a_data_width = 1;
defparam ram_block1a126.port_a_first_address = 57344;
defparam ram_block1a126.port_a_first_bit_number = 14;
defparam ram_block1a126.port_a_last_address = 65535;
defparam ram_block1a126.port_a_logical_ram_depth = 65536;
defparam ram_block1a126.port_a_logical_ram_width = 16;
defparam ram_block1a126.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a126.ram_block_type = "auto";
defparam ram_block1a126.mem_init3 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a126.mem_init2 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a126.mem_init1 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a126.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

arriav_ram_block ram_block1a46(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a46_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a46.clk0_core_clock_enable = "ena0";
defparam ram_block1a46.clk0_input_clock_enable = "ena0";
defparam ram_block1a46.clk0_output_clock_enable = "ena0";
defparam ram_block1a46.data_interleave_offset_in_bits = 1;
defparam ram_block1a46.data_interleave_width_in_bits = 1;
defparam ram_block1a46.init_file = "DDS_48_v1_nco_ii_0_sin.hex";
defparam ram_block1a46.init_file_layout = "port_a";
defparam ram_block1a46.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_c8g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a46.operation_mode = "rom";
defparam ram_block1a46.port_a_address_clear = "none";
defparam ram_block1a46.port_a_address_width = 13;
defparam ram_block1a46.port_a_data_out_clear = "none";
defparam ram_block1a46.port_a_data_out_clock = "clock0";
defparam ram_block1a46.port_a_data_width = 1;
defparam ram_block1a46.port_a_first_address = 16384;
defparam ram_block1a46.port_a_first_bit_number = 14;
defparam ram_block1a46.port_a_last_address = 24575;
defparam ram_block1a46.port_a_logical_ram_depth = 65536;
defparam ram_block1a46.port_a_logical_ram_width = 16;
defparam ram_block1a46.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a46.ram_block_type = "auto";
defparam ram_block1a46.mem_init3 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a46.mem_init2 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a46.mem_init1 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a46.mem_init0 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

arriav_ram_block ram_block1a62(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a62_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a62.clk0_core_clock_enable = "ena0";
defparam ram_block1a62.clk0_input_clock_enable = "ena0";
defparam ram_block1a62.clk0_output_clock_enable = "ena0";
defparam ram_block1a62.data_interleave_offset_in_bits = 1;
defparam ram_block1a62.data_interleave_width_in_bits = 1;
defparam ram_block1a62.init_file = "DDS_48_v1_nco_ii_0_sin.hex";
defparam ram_block1a62.init_file_layout = "port_a";
defparam ram_block1a62.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_c8g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a62.operation_mode = "rom";
defparam ram_block1a62.port_a_address_clear = "none";
defparam ram_block1a62.port_a_address_width = 13;
defparam ram_block1a62.port_a_data_out_clear = "none";
defparam ram_block1a62.port_a_data_out_clock = "clock0";
defparam ram_block1a62.port_a_data_width = 1;
defparam ram_block1a62.port_a_first_address = 24576;
defparam ram_block1a62.port_a_first_bit_number = 14;
defparam ram_block1a62.port_a_last_address = 32767;
defparam ram_block1a62.port_a_logical_ram_depth = 65536;
defparam ram_block1a62.port_a_logical_ram_width = 16;
defparam ram_block1a62.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a62.ram_block_type = "auto";
defparam ram_block1a62.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a62.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a62.mem_init1 = "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a62.mem_init0 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

arriav_ram_block ram_block1a14(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a14_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a14.clk0_core_clock_enable = "ena0";
defparam ram_block1a14.clk0_input_clock_enable = "ena0";
defparam ram_block1a14.clk0_output_clock_enable = "ena0";
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.init_file = "DDS_48_v1_nco_ii_0_sin.hex";
defparam ram_block1a14.init_file_layout = "port_a";
defparam ram_block1a14.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_c8g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a14.operation_mode = "rom";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 13;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "clock0";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 8191;
defparam ram_block1a14.port_a_logical_ram_depth = 65536;
defparam ram_block1a14.port_a_logical_ram_width = 16;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a14.ram_block_type = "auto";
defparam ram_block1a14.mem_init3 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a14.mem_init2 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a14.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a14.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

arriav_ram_block ram_block1a30(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a30_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a30.clk0_core_clock_enable = "ena0";
defparam ram_block1a30.clk0_input_clock_enable = "ena0";
defparam ram_block1a30.clk0_output_clock_enable = "ena0";
defparam ram_block1a30.data_interleave_offset_in_bits = 1;
defparam ram_block1a30.data_interleave_width_in_bits = 1;
defparam ram_block1a30.init_file = "DDS_48_v1_nco_ii_0_sin.hex";
defparam ram_block1a30.init_file_layout = "port_a";
defparam ram_block1a30.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_c8g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a30.operation_mode = "rom";
defparam ram_block1a30.port_a_address_clear = "none";
defparam ram_block1a30.port_a_address_width = 13;
defparam ram_block1a30.port_a_data_out_clear = "none";
defparam ram_block1a30.port_a_data_out_clock = "clock0";
defparam ram_block1a30.port_a_data_width = 1;
defparam ram_block1a30.port_a_first_address = 8192;
defparam ram_block1a30.port_a_first_bit_number = 14;
defparam ram_block1a30.port_a_last_address = 16383;
defparam ram_block1a30.port_a_logical_ram_depth = 65536;
defparam ram_block1a30.port_a_logical_ram_width = 16;
defparam ram_block1a30.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a30.ram_block_type = "auto";
defparam ram_block1a30.mem_init3 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a30.mem_init2 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a30.mem_init1 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a30.mem_init0 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

arriav_ram_block ram_block1a79(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a79_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a79.clk0_core_clock_enable = "ena0";
defparam ram_block1a79.clk0_input_clock_enable = "ena0";
defparam ram_block1a79.clk0_output_clock_enable = "ena0";
defparam ram_block1a79.data_interleave_offset_in_bits = 1;
defparam ram_block1a79.data_interleave_width_in_bits = 1;
defparam ram_block1a79.init_file = "DDS_48_v1_nco_ii_0_sin.hex";
defparam ram_block1a79.init_file_layout = "port_a";
defparam ram_block1a79.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_c8g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a79.operation_mode = "rom";
defparam ram_block1a79.port_a_address_clear = "none";
defparam ram_block1a79.port_a_address_width = 13;
defparam ram_block1a79.port_a_data_out_clear = "none";
defparam ram_block1a79.port_a_data_out_clock = "clock0";
defparam ram_block1a79.port_a_data_width = 1;
defparam ram_block1a79.port_a_first_address = 32768;
defparam ram_block1a79.port_a_first_bit_number = 15;
defparam ram_block1a79.port_a_last_address = 40959;
defparam ram_block1a79.port_a_logical_ram_depth = 65536;
defparam ram_block1a79.port_a_logical_ram_width = 16;
defparam ram_block1a79.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a79.ram_block_type = "auto";
defparam ram_block1a79.mem_init3 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a79.mem_init2 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a79.mem_init1 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a79.mem_init0 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE";

arriav_ram_block ram_block1a95(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a95_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a95.clk0_core_clock_enable = "ena0";
defparam ram_block1a95.clk0_input_clock_enable = "ena0";
defparam ram_block1a95.clk0_output_clock_enable = "ena0";
defparam ram_block1a95.data_interleave_offset_in_bits = 1;
defparam ram_block1a95.data_interleave_width_in_bits = 1;
defparam ram_block1a95.init_file = "DDS_48_v1_nco_ii_0_sin.hex";
defparam ram_block1a95.init_file_layout = "port_a";
defparam ram_block1a95.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_c8g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a95.operation_mode = "rom";
defparam ram_block1a95.port_a_address_clear = "none";
defparam ram_block1a95.port_a_address_width = 13;
defparam ram_block1a95.port_a_data_out_clear = "none";
defparam ram_block1a95.port_a_data_out_clock = "clock0";
defparam ram_block1a95.port_a_data_width = 1;
defparam ram_block1a95.port_a_first_address = 40960;
defparam ram_block1a95.port_a_first_bit_number = 15;
defparam ram_block1a95.port_a_last_address = 49151;
defparam ram_block1a95.port_a_logical_ram_depth = 65536;
defparam ram_block1a95.port_a_logical_ram_width = 16;
defparam ram_block1a95.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a95.ram_block_type = "auto";
defparam ram_block1a95.mem_init3 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a95.mem_init2 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a95.mem_init1 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a95.mem_init0 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

arriav_ram_block ram_block1a111(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a111_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a111.clk0_core_clock_enable = "ena0";
defparam ram_block1a111.clk0_input_clock_enable = "ena0";
defparam ram_block1a111.clk0_output_clock_enable = "ena0";
defparam ram_block1a111.data_interleave_offset_in_bits = 1;
defparam ram_block1a111.data_interleave_width_in_bits = 1;
defparam ram_block1a111.init_file = "DDS_48_v1_nco_ii_0_sin.hex";
defparam ram_block1a111.init_file_layout = "port_a";
defparam ram_block1a111.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_c8g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a111.operation_mode = "rom";
defparam ram_block1a111.port_a_address_clear = "none";
defparam ram_block1a111.port_a_address_width = 13;
defparam ram_block1a111.port_a_data_out_clear = "none";
defparam ram_block1a111.port_a_data_out_clock = "clock0";
defparam ram_block1a111.port_a_data_width = 1;
defparam ram_block1a111.port_a_first_address = 49152;
defparam ram_block1a111.port_a_first_bit_number = 15;
defparam ram_block1a111.port_a_last_address = 57343;
defparam ram_block1a111.port_a_logical_ram_depth = 65536;
defparam ram_block1a111.port_a_logical_ram_width = 16;
defparam ram_block1a111.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a111.ram_block_type = "auto";
defparam ram_block1a111.mem_init3 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a111.mem_init2 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a111.mem_init1 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a111.mem_init0 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

arriav_ram_block ram_block1a127(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a127_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a127.clk0_core_clock_enable = "ena0";
defparam ram_block1a127.clk0_input_clock_enable = "ena0";
defparam ram_block1a127.clk0_output_clock_enable = "ena0";
defparam ram_block1a127.data_interleave_offset_in_bits = 1;
defparam ram_block1a127.data_interleave_width_in_bits = 1;
defparam ram_block1a127.init_file = "DDS_48_v1_nco_ii_0_sin.hex";
defparam ram_block1a127.init_file_layout = "port_a";
defparam ram_block1a127.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_c8g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a127.operation_mode = "rom";
defparam ram_block1a127.port_a_address_clear = "none";
defparam ram_block1a127.port_a_address_width = 13;
defparam ram_block1a127.port_a_data_out_clear = "none";
defparam ram_block1a127.port_a_data_out_clock = "clock0";
defparam ram_block1a127.port_a_data_width = 1;
defparam ram_block1a127.port_a_first_address = 57344;
defparam ram_block1a127.port_a_first_bit_number = 15;
defparam ram_block1a127.port_a_last_address = 65535;
defparam ram_block1a127.port_a_logical_ram_depth = 65536;
defparam ram_block1a127.port_a_logical_ram_width = 16;
defparam ram_block1a127.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a127.ram_block_type = "auto";
defparam ram_block1a127.mem_init3 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a127.mem_init2 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a127.mem_init1 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a127.mem_init0 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

arriav_ram_block ram_block1a47(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a47_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a47.clk0_core_clock_enable = "ena0";
defparam ram_block1a47.clk0_input_clock_enable = "ena0";
defparam ram_block1a47.clk0_output_clock_enable = "ena0";
defparam ram_block1a47.data_interleave_offset_in_bits = 1;
defparam ram_block1a47.data_interleave_width_in_bits = 1;
defparam ram_block1a47.init_file = "DDS_48_v1_nco_ii_0_sin.hex";
defparam ram_block1a47.init_file_layout = "port_a";
defparam ram_block1a47.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_c8g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a47.operation_mode = "rom";
defparam ram_block1a47.port_a_address_clear = "none";
defparam ram_block1a47.port_a_address_width = 13;
defparam ram_block1a47.port_a_data_out_clear = "none";
defparam ram_block1a47.port_a_data_out_clock = "clock0";
defparam ram_block1a47.port_a_data_width = 1;
defparam ram_block1a47.port_a_first_address = 16384;
defparam ram_block1a47.port_a_first_bit_number = 15;
defparam ram_block1a47.port_a_last_address = 24575;
defparam ram_block1a47.port_a_logical_ram_depth = 65536;
defparam ram_block1a47.port_a_logical_ram_width = 16;
defparam ram_block1a47.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a47.ram_block_type = "auto";
defparam ram_block1a47.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a47.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a47.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a47.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

arriav_ram_block ram_block1a63(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a63_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a63.clk0_core_clock_enable = "ena0";
defparam ram_block1a63.clk0_input_clock_enable = "ena0";
defparam ram_block1a63.clk0_output_clock_enable = "ena0";
defparam ram_block1a63.data_interleave_offset_in_bits = 1;
defparam ram_block1a63.data_interleave_width_in_bits = 1;
defparam ram_block1a63.init_file = "DDS_48_v1_nco_ii_0_sin.hex";
defparam ram_block1a63.init_file_layout = "port_a";
defparam ram_block1a63.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_c8g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a63.operation_mode = "rom";
defparam ram_block1a63.port_a_address_clear = "none";
defparam ram_block1a63.port_a_address_width = 13;
defparam ram_block1a63.port_a_data_out_clear = "none";
defparam ram_block1a63.port_a_data_out_clock = "clock0";
defparam ram_block1a63.port_a_data_width = 1;
defparam ram_block1a63.port_a_first_address = 24576;
defparam ram_block1a63.port_a_first_bit_number = 15;
defparam ram_block1a63.port_a_last_address = 32767;
defparam ram_block1a63.port_a_logical_ram_depth = 65536;
defparam ram_block1a63.port_a_logical_ram_width = 16;
defparam ram_block1a63.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a63.ram_block_type = "auto";
defparam ram_block1a63.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a63.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a63.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a63.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

arriav_ram_block ram_block1a15(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a15_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a15.clk0_core_clock_enable = "ena0";
defparam ram_block1a15.clk0_input_clock_enable = "ena0";
defparam ram_block1a15.clk0_output_clock_enable = "ena0";
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.init_file = "DDS_48_v1_nco_ii_0_sin.hex";
defparam ram_block1a15.init_file_layout = "port_a";
defparam ram_block1a15.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_c8g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a15.operation_mode = "rom";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 13;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "clock0";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 8191;
defparam ram_block1a15.port_a_logical_ram_depth = 65536;
defparam ram_block1a15.port_a_logical_ram_width = 16;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a15.ram_block_type = "auto";
defparam ram_block1a15.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a15.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a15.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a15.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

arriav_ram_block ram_block1a31(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a31_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a31.clk0_core_clock_enable = "ena0";
defparam ram_block1a31.clk0_input_clock_enable = "ena0";
defparam ram_block1a31.clk0_output_clock_enable = "ena0";
defparam ram_block1a31.data_interleave_offset_in_bits = 1;
defparam ram_block1a31.data_interleave_width_in_bits = 1;
defparam ram_block1a31.init_file = "DDS_48_v1_nco_ii_0_sin.hex";
defparam ram_block1a31.init_file_layout = "port_a";
defparam ram_block1a31.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_c8g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a31.operation_mode = "rom";
defparam ram_block1a31.port_a_address_clear = "none";
defparam ram_block1a31.port_a_address_width = 13;
defparam ram_block1a31.port_a_data_out_clear = "none";
defparam ram_block1a31.port_a_data_out_clock = "clock0";
defparam ram_block1a31.port_a_data_width = 1;
defparam ram_block1a31.port_a_first_address = 8192;
defparam ram_block1a31.port_a_first_bit_number = 15;
defparam ram_block1a31.port_a_last_address = 16383;
defparam ram_block1a31.port_a_logical_ram_depth = 65536;
defparam ram_block1a31.port_a_logical_ram_width = 16;
defparam ram_block1a31.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a31.ram_block_type = "auto";
defparam ram_block1a31.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a31.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a31.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a31.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

dffeas \out_address_reg_a[2] (
	.clk(clock0),
	.d(\address_reg_a[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clocken0),
	.q(out_address_reg_a_2),
	.prn(vcc));
defparam \out_address_reg_a[2] .is_wysiwyg = "true";
defparam \out_address_reg_a[2] .power_up = "low";

dffeas \out_address_reg_a[0] (
	.clk(clock0),
	.d(\address_reg_a[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clocken0),
	.q(out_address_reg_a_0),
	.prn(vcc));
defparam \out_address_reg_a[0] .is_wysiwyg = "true";
defparam \out_address_reg_a[0] .power_up = "low";

dffeas \out_address_reg_a[1] (
	.clk(clock0),
	.d(\address_reg_a[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clocken0),
	.q(out_address_reg_a_1),
	.prn(vcc));
defparam \out_address_reg_a[1] .is_wysiwyg = "true";
defparam \out_address_reg_a[1] .power_up = "low";

dffeas \address_reg_a[2] (
	.clk(clock0),
	.d(address_a[15]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clocken0),
	.q(\address_reg_a[2]~q ),
	.prn(vcc));
defparam \address_reg_a[2] .is_wysiwyg = "true";
defparam \address_reg_a[2] .power_up = "low";

dffeas \address_reg_a[0] (
	.clk(clock0),
	.d(address_a[13]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clocken0),
	.q(\address_reg_a[0]~q ),
	.prn(vcc));
defparam \address_reg_a[0] .is_wysiwyg = "true";
defparam \address_reg_a[0] .power_up = "low";

dffeas \address_reg_a[1] (
	.clk(clock0),
	.d(address_a[14]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clocken0),
	.q(\address_reg_a[1]~q ),
	.prn(vcc));
defparam \address_reg_a[1] .is_wysiwyg = "true";
defparam \address_reg_a[1] .power_up = "low";

endmodule

module DDS_48_v1_asj_nco_as_m_cen_1 (
	ram_block1a64,
	ram_block1a80,
	ram_block1a96,
	ram_block1a112,
	ram_block1a32,
	ram_block1a48,
	ram_block1a0,
	ram_block1a16,
	ram_block1a65,
	ram_block1a81,
	ram_block1a97,
	ram_block1a113,
	ram_block1a33,
	ram_block1a49,
	ram_block1a1,
	ram_block1a17,
	ram_block1a66,
	ram_block1a82,
	ram_block1a98,
	ram_block1a114,
	ram_block1a34,
	ram_block1a50,
	ram_block1a2,
	ram_block1a18,
	ram_block1a67,
	ram_block1a83,
	ram_block1a99,
	ram_block1a115,
	ram_block1a35,
	ram_block1a51,
	ram_block1a3,
	ram_block1a19,
	ram_block1a68,
	ram_block1a84,
	ram_block1a100,
	ram_block1a116,
	ram_block1a36,
	ram_block1a52,
	ram_block1a4,
	ram_block1a20,
	ram_block1a69,
	ram_block1a85,
	ram_block1a101,
	ram_block1a117,
	ram_block1a37,
	ram_block1a53,
	ram_block1a5,
	ram_block1a21,
	ram_block1a70,
	ram_block1a86,
	ram_block1a102,
	ram_block1a118,
	ram_block1a38,
	ram_block1a54,
	ram_block1a6,
	ram_block1a22,
	ram_block1a71,
	ram_block1a87,
	ram_block1a103,
	ram_block1a119,
	ram_block1a39,
	ram_block1a55,
	ram_block1a7,
	ram_block1a23,
	ram_block1a72,
	ram_block1a88,
	ram_block1a104,
	ram_block1a120,
	ram_block1a40,
	ram_block1a56,
	ram_block1a8,
	ram_block1a24,
	ram_block1a73,
	ram_block1a89,
	ram_block1a105,
	ram_block1a121,
	ram_block1a41,
	ram_block1a57,
	ram_block1a9,
	ram_block1a25,
	ram_block1a74,
	ram_block1a90,
	ram_block1a106,
	ram_block1a122,
	ram_block1a42,
	ram_block1a58,
	ram_block1a10,
	ram_block1a26,
	ram_block1a75,
	ram_block1a91,
	ram_block1a107,
	ram_block1a123,
	ram_block1a43,
	ram_block1a59,
	ram_block1a11,
	ram_block1a27,
	ram_block1a76,
	ram_block1a92,
	ram_block1a108,
	ram_block1a124,
	ram_block1a44,
	ram_block1a60,
	ram_block1a12,
	ram_block1a28,
	ram_block1a77,
	ram_block1a93,
	ram_block1a109,
	ram_block1a125,
	ram_block1a45,
	ram_block1a61,
	ram_block1a13,
	ram_block1a29,
	ram_block1a78,
	ram_block1a94,
	ram_block1a110,
	ram_block1a126,
	ram_block1a46,
	ram_block1a62,
	ram_block1a14,
	ram_block1a30,
	ram_block1a79,
	ram_block1a95,
	ram_block1a111,
	ram_block1a127,
	ram_block1a47,
	ram_block1a63,
	ram_block1a15,
	ram_block1a31,
	rom_add_0,
	rom_add_1,
	rom_add_2,
	rom_add_3,
	rom_add_4,
	rom_add_5,
	rom_add_6,
	rom_add_7,
	rom_add_8,
	rom_add_9,
	rom_add_10,
	rom_add_11,
	rom_add_12,
	clk,
	clken)/* synthesis synthesis_greybox=1 */;
output 	ram_block1a64;
output 	ram_block1a80;
output 	ram_block1a96;
output 	ram_block1a112;
output 	ram_block1a32;
output 	ram_block1a48;
output 	ram_block1a0;
output 	ram_block1a16;
output 	ram_block1a65;
output 	ram_block1a81;
output 	ram_block1a97;
output 	ram_block1a113;
output 	ram_block1a33;
output 	ram_block1a49;
output 	ram_block1a1;
output 	ram_block1a17;
output 	ram_block1a66;
output 	ram_block1a82;
output 	ram_block1a98;
output 	ram_block1a114;
output 	ram_block1a34;
output 	ram_block1a50;
output 	ram_block1a2;
output 	ram_block1a18;
output 	ram_block1a67;
output 	ram_block1a83;
output 	ram_block1a99;
output 	ram_block1a115;
output 	ram_block1a35;
output 	ram_block1a51;
output 	ram_block1a3;
output 	ram_block1a19;
output 	ram_block1a68;
output 	ram_block1a84;
output 	ram_block1a100;
output 	ram_block1a116;
output 	ram_block1a36;
output 	ram_block1a52;
output 	ram_block1a4;
output 	ram_block1a20;
output 	ram_block1a69;
output 	ram_block1a85;
output 	ram_block1a101;
output 	ram_block1a117;
output 	ram_block1a37;
output 	ram_block1a53;
output 	ram_block1a5;
output 	ram_block1a21;
output 	ram_block1a70;
output 	ram_block1a86;
output 	ram_block1a102;
output 	ram_block1a118;
output 	ram_block1a38;
output 	ram_block1a54;
output 	ram_block1a6;
output 	ram_block1a22;
output 	ram_block1a71;
output 	ram_block1a87;
output 	ram_block1a103;
output 	ram_block1a119;
output 	ram_block1a39;
output 	ram_block1a55;
output 	ram_block1a7;
output 	ram_block1a23;
output 	ram_block1a72;
output 	ram_block1a88;
output 	ram_block1a104;
output 	ram_block1a120;
output 	ram_block1a40;
output 	ram_block1a56;
output 	ram_block1a8;
output 	ram_block1a24;
output 	ram_block1a73;
output 	ram_block1a89;
output 	ram_block1a105;
output 	ram_block1a121;
output 	ram_block1a41;
output 	ram_block1a57;
output 	ram_block1a9;
output 	ram_block1a25;
output 	ram_block1a74;
output 	ram_block1a90;
output 	ram_block1a106;
output 	ram_block1a122;
output 	ram_block1a42;
output 	ram_block1a58;
output 	ram_block1a10;
output 	ram_block1a26;
output 	ram_block1a75;
output 	ram_block1a91;
output 	ram_block1a107;
output 	ram_block1a123;
output 	ram_block1a43;
output 	ram_block1a59;
output 	ram_block1a11;
output 	ram_block1a27;
output 	ram_block1a76;
output 	ram_block1a92;
output 	ram_block1a108;
output 	ram_block1a124;
output 	ram_block1a44;
output 	ram_block1a60;
output 	ram_block1a12;
output 	ram_block1a28;
output 	ram_block1a77;
output 	ram_block1a93;
output 	ram_block1a109;
output 	ram_block1a125;
output 	ram_block1a45;
output 	ram_block1a61;
output 	ram_block1a13;
output 	ram_block1a29;
output 	ram_block1a78;
output 	ram_block1a94;
output 	ram_block1a110;
output 	ram_block1a126;
output 	ram_block1a46;
output 	ram_block1a62;
output 	ram_block1a14;
output 	ram_block1a30;
output 	ram_block1a79;
output 	ram_block1a95;
output 	ram_block1a111;
output 	ram_block1a127;
output 	ram_block1a47;
output 	ram_block1a63;
output 	ram_block1a15;
output 	ram_block1a31;
input 	rom_add_0;
input 	rom_add_1;
input 	rom_add_2;
input 	rom_add_3;
input 	rom_add_4;
input 	rom_add_5;
input 	rom_add_6;
input 	rom_add_7;
input 	rom_add_8;
input 	rom_add_9;
input 	rom_add_10;
input 	rom_add_11;
input 	rom_add_12;
input 	clk;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



DDS_48_v1_altsyncram_2 altsyncram_component0(
	.ram_block1a64(ram_block1a64),
	.ram_block1a80(ram_block1a80),
	.ram_block1a96(ram_block1a96),
	.ram_block1a112(ram_block1a112),
	.ram_block1a32(ram_block1a32),
	.ram_block1a48(ram_block1a48),
	.ram_block1a0(ram_block1a0),
	.ram_block1a16(ram_block1a16),
	.ram_block1a65(ram_block1a65),
	.ram_block1a81(ram_block1a81),
	.ram_block1a97(ram_block1a97),
	.ram_block1a113(ram_block1a113),
	.ram_block1a33(ram_block1a33),
	.ram_block1a49(ram_block1a49),
	.ram_block1a1(ram_block1a1),
	.ram_block1a17(ram_block1a17),
	.ram_block1a66(ram_block1a66),
	.ram_block1a82(ram_block1a82),
	.ram_block1a98(ram_block1a98),
	.ram_block1a114(ram_block1a114),
	.ram_block1a34(ram_block1a34),
	.ram_block1a50(ram_block1a50),
	.ram_block1a2(ram_block1a2),
	.ram_block1a18(ram_block1a18),
	.ram_block1a67(ram_block1a67),
	.ram_block1a83(ram_block1a83),
	.ram_block1a99(ram_block1a99),
	.ram_block1a115(ram_block1a115),
	.ram_block1a35(ram_block1a35),
	.ram_block1a51(ram_block1a51),
	.ram_block1a3(ram_block1a3),
	.ram_block1a19(ram_block1a19),
	.ram_block1a68(ram_block1a68),
	.ram_block1a84(ram_block1a84),
	.ram_block1a100(ram_block1a100),
	.ram_block1a116(ram_block1a116),
	.ram_block1a36(ram_block1a36),
	.ram_block1a52(ram_block1a52),
	.ram_block1a4(ram_block1a4),
	.ram_block1a20(ram_block1a20),
	.ram_block1a69(ram_block1a69),
	.ram_block1a85(ram_block1a85),
	.ram_block1a101(ram_block1a101),
	.ram_block1a117(ram_block1a117),
	.ram_block1a37(ram_block1a37),
	.ram_block1a53(ram_block1a53),
	.ram_block1a5(ram_block1a5),
	.ram_block1a21(ram_block1a21),
	.ram_block1a70(ram_block1a70),
	.ram_block1a86(ram_block1a86),
	.ram_block1a102(ram_block1a102),
	.ram_block1a118(ram_block1a118),
	.ram_block1a38(ram_block1a38),
	.ram_block1a54(ram_block1a54),
	.ram_block1a6(ram_block1a6),
	.ram_block1a22(ram_block1a22),
	.ram_block1a71(ram_block1a71),
	.ram_block1a87(ram_block1a87),
	.ram_block1a103(ram_block1a103),
	.ram_block1a119(ram_block1a119),
	.ram_block1a39(ram_block1a39),
	.ram_block1a55(ram_block1a55),
	.ram_block1a7(ram_block1a7),
	.ram_block1a23(ram_block1a23),
	.ram_block1a72(ram_block1a72),
	.ram_block1a88(ram_block1a88),
	.ram_block1a104(ram_block1a104),
	.ram_block1a120(ram_block1a120),
	.ram_block1a40(ram_block1a40),
	.ram_block1a56(ram_block1a56),
	.ram_block1a8(ram_block1a8),
	.ram_block1a24(ram_block1a24),
	.ram_block1a73(ram_block1a73),
	.ram_block1a89(ram_block1a89),
	.ram_block1a105(ram_block1a105),
	.ram_block1a121(ram_block1a121),
	.ram_block1a41(ram_block1a41),
	.ram_block1a57(ram_block1a57),
	.ram_block1a9(ram_block1a9),
	.ram_block1a25(ram_block1a25),
	.ram_block1a74(ram_block1a74),
	.ram_block1a90(ram_block1a90),
	.ram_block1a106(ram_block1a106),
	.ram_block1a122(ram_block1a122),
	.ram_block1a42(ram_block1a42),
	.ram_block1a58(ram_block1a58),
	.ram_block1a10(ram_block1a10),
	.ram_block1a26(ram_block1a26),
	.ram_block1a75(ram_block1a75),
	.ram_block1a91(ram_block1a91),
	.ram_block1a107(ram_block1a107),
	.ram_block1a123(ram_block1a123),
	.ram_block1a43(ram_block1a43),
	.ram_block1a59(ram_block1a59),
	.ram_block1a11(ram_block1a11),
	.ram_block1a27(ram_block1a27),
	.ram_block1a76(ram_block1a76),
	.ram_block1a92(ram_block1a92),
	.ram_block1a108(ram_block1a108),
	.ram_block1a124(ram_block1a124),
	.ram_block1a44(ram_block1a44),
	.ram_block1a60(ram_block1a60),
	.ram_block1a12(ram_block1a12),
	.ram_block1a28(ram_block1a28),
	.ram_block1a77(ram_block1a77),
	.ram_block1a93(ram_block1a93),
	.ram_block1a109(ram_block1a109),
	.ram_block1a125(ram_block1a125),
	.ram_block1a45(ram_block1a45),
	.ram_block1a61(ram_block1a61),
	.ram_block1a13(ram_block1a13),
	.ram_block1a29(ram_block1a29),
	.ram_block1a78(ram_block1a78),
	.ram_block1a94(ram_block1a94),
	.ram_block1a110(ram_block1a110),
	.ram_block1a126(ram_block1a126),
	.ram_block1a46(ram_block1a46),
	.ram_block1a62(ram_block1a62),
	.ram_block1a14(ram_block1a14),
	.ram_block1a30(ram_block1a30),
	.ram_block1a79(ram_block1a79),
	.ram_block1a95(ram_block1a95),
	.ram_block1a111(ram_block1a111),
	.ram_block1a127(ram_block1a127),
	.ram_block1a47(ram_block1a47),
	.ram_block1a63(ram_block1a63),
	.ram_block1a15(ram_block1a15),
	.ram_block1a31(ram_block1a31),
	.address_a({gnd,gnd,gnd,rom_add_12,rom_add_11,rom_add_10,rom_add_9,rom_add_8,rom_add_7,rom_add_6,rom_add_5,rom_add_4,rom_add_3,rom_add_2,rom_add_1,rom_add_0}),
	.clock0(clk),
	.clocken0(clken));

endmodule

module DDS_48_v1_altsyncram_2 (
	ram_block1a64,
	ram_block1a80,
	ram_block1a96,
	ram_block1a112,
	ram_block1a32,
	ram_block1a48,
	ram_block1a0,
	ram_block1a16,
	ram_block1a65,
	ram_block1a81,
	ram_block1a97,
	ram_block1a113,
	ram_block1a33,
	ram_block1a49,
	ram_block1a1,
	ram_block1a17,
	ram_block1a66,
	ram_block1a82,
	ram_block1a98,
	ram_block1a114,
	ram_block1a34,
	ram_block1a50,
	ram_block1a2,
	ram_block1a18,
	ram_block1a67,
	ram_block1a83,
	ram_block1a99,
	ram_block1a115,
	ram_block1a35,
	ram_block1a51,
	ram_block1a3,
	ram_block1a19,
	ram_block1a68,
	ram_block1a84,
	ram_block1a100,
	ram_block1a116,
	ram_block1a36,
	ram_block1a52,
	ram_block1a4,
	ram_block1a20,
	ram_block1a69,
	ram_block1a85,
	ram_block1a101,
	ram_block1a117,
	ram_block1a37,
	ram_block1a53,
	ram_block1a5,
	ram_block1a21,
	ram_block1a70,
	ram_block1a86,
	ram_block1a102,
	ram_block1a118,
	ram_block1a38,
	ram_block1a54,
	ram_block1a6,
	ram_block1a22,
	ram_block1a71,
	ram_block1a87,
	ram_block1a103,
	ram_block1a119,
	ram_block1a39,
	ram_block1a55,
	ram_block1a7,
	ram_block1a23,
	ram_block1a72,
	ram_block1a88,
	ram_block1a104,
	ram_block1a120,
	ram_block1a40,
	ram_block1a56,
	ram_block1a8,
	ram_block1a24,
	ram_block1a73,
	ram_block1a89,
	ram_block1a105,
	ram_block1a121,
	ram_block1a41,
	ram_block1a57,
	ram_block1a9,
	ram_block1a25,
	ram_block1a74,
	ram_block1a90,
	ram_block1a106,
	ram_block1a122,
	ram_block1a42,
	ram_block1a58,
	ram_block1a10,
	ram_block1a26,
	ram_block1a75,
	ram_block1a91,
	ram_block1a107,
	ram_block1a123,
	ram_block1a43,
	ram_block1a59,
	ram_block1a11,
	ram_block1a27,
	ram_block1a76,
	ram_block1a92,
	ram_block1a108,
	ram_block1a124,
	ram_block1a44,
	ram_block1a60,
	ram_block1a12,
	ram_block1a28,
	ram_block1a77,
	ram_block1a93,
	ram_block1a109,
	ram_block1a125,
	ram_block1a45,
	ram_block1a61,
	ram_block1a13,
	ram_block1a29,
	ram_block1a78,
	ram_block1a94,
	ram_block1a110,
	ram_block1a126,
	ram_block1a46,
	ram_block1a62,
	ram_block1a14,
	ram_block1a30,
	ram_block1a79,
	ram_block1a95,
	ram_block1a111,
	ram_block1a127,
	ram_block1a47,
	ram_block1a63,
	ram_block1a15,
	ram_block1a31,
	address_a,
	clock0,
	clocken0)/* synthesis synthesis_greybox=1 */;
output 	ram_block1a64;
output 	ram_block1a80;
output 	ram_block1a96;
output 	ram_block1a112;
output 	ram_block1a32;
output 	ram_block1a48;
output 	ram_block1a0;
output 	ram_block1a16;
output 	ram_block1a65;
output 	ram_block1a81;
output 	ram_block1a97;
output 	ram_block1a113;
output 	ram_block1a33;
output 	ram_block1a49;
output 	ram_block1a1;
output 	ram_block1a17;
output 	ram_block1a66;
output 	ram_block1a82;
output 	ram_block1a98;
output 	ram_block1a114;
output 	ram_block1a34;
output 	ram_block1a50;
output 	ram_block1a2;
output 	ram_block1a18;
output 	ram_block1a67;
output 	ram_block1a83;
output 	ram_block1a99;
output 	ram_block1a115;
output 	ram_block1a35;
output 	ram_block1a51;
output 	ram_block1a3;
output 	ram_block1a19;
output 	ram_block1a68;
output 	ram_block1a84;
output 	ram_block1a100;
output 	ram_block1a116;
output 	ram_block1a36;
output 	ram_block1a52;
output 	ram_block1a4;
output 	ram_block1a20;
output 	ram_block1a69;
output 	ram_block1a85;
output 	ram_block1a101;
output 	ram_block1a117;
output 	ram_block1a37;
output 	ram_block1a53;
output 	ram_block1a5;
output 	ram_block1a21;
output 	ram_block1a70;
output 	ram_block1a86;
output 	ram_block1a102;
output 	ram_block1a118;
output 	ram_block1a38;
output 	ram_block1a54;
output 	ram_block1a6;
output 	ram_block1a22;
output 	ram_block1a71;
output 	ram_block1a87;
output 	ram_block1a103;
output 	ram_block1a119;
output 	ram_block1a39;
output 	ram_block1a55;
output 	ram_block1a7;
output 	ram_block1a23;
output 	ram_block1a72;
output 	ram_block1a88;
output 	ram_block1a104;
output 	ram_block1a120;
output 	ram_block1a40;
output 	ram_block1a56;
output 	ram_block1a8;
output 	ram_block1a24;
output 	ram_block1a73;
output 	ram_block1a89;
output 	ram_block1a105;
output 	ram_block1a121;
output 	ram_block1a41;
output 	ram_block1a57;
output 	ram_block1a9;
output 	ram_block1a25;
output 	ram_block1a74;
output 	ram_block1a90;
output 	ram_block1a106;
output 	ram_block1a122;
output 	ram_block1a42;
output 	ram_block1a58;
output 	ram_block1a10;
output 	ram_block1a26;
output 	ram_block1a75;
output 	ram_block1a91;
output 	ram_block1a107;
output 	ram_block1a123;
output 	ram_block1a43;
output 	ram_block1a59;
output 	ram_block1a11;
output 	ram_block1a27;
output 	ram_block1a76;
output 	ram_block1a92;
output 	ram_block1a108;
output 	ram_block1a124;
output 	ram_block1a44;
output 	ram_block1a60;
output 	ram_block1a12;
output 	ram_block1a28;
output 	ram_block1a77;
output 	ram_block1a93;
output 	ram_block1a109;
output 	ram_block1a125;
output 	ram_block1a45;
output 	ram_block1a61;
output 	ram_block1a13;
output 	ram_block1a29;
output 	ram_block1a78;
output 	ram_block1a94;
output 	ram_block1a110;
output 	ram_block1a126;
output 	ram_block1a46;
output 	ram_block1a62;
output 	ram_block1a14;
output 	ram_block1a30;
output 	ram_block1a79;
output 	ram_block1a95;
output 	ram_block1a111;
output 	ram_block1a127;
output 	ram_block1a47;
output 	ram_block1a63;
output 	ram_block1a15;
output 	ram_block1a31;
input 	[15:0] address_a;
input 	clock0;
input 	clocken0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



DDS_48_v1_altsyncram_78g1 auto_generated(
	.ram_block1a641(ram_block1a64),
	.ram_block1a801(ram_block1a80),
	.ram_block1a961(ram_block1a96),
	.ram_block1a1121(ram_block1a112),
	.ram_block1a321(ram_block1a32),
	.ram_block1a481(ram_block1a48),
	.ram_block1a01(ram_block1a0),
	.ram_block1a161(ram_block1a16),
	.ram_block1a651(ram_block1a65),
	.ram_block1a811(ram_block1a81),
	.ram_block1a971(ram_block1a97),
	.ram_block1a1131(ram_block1a113),
	.ram_block1a331(ram_block1a33),
	.ram_block1a491(ram_block1a49),
	.ram_block1a128(ram_block1a1),
	.ram_block1a171(ram_block1a17),
	.ram_block1a661(ram_block1a66),
	.ram_block1a821(ram_block1a82),
	.ram_block1a981(ram_block1a98),
	.ram_block1a1141(ram_block1a114),
	.ram_block1a341(ram_block1a34),
	.ram_block1a501(ram_block1a50),
	.ram_block1a210(ram_block1a2),
	.ram_block1a181(ram_block1a18),
	.ram_block1a671(ram_block1a67),
	.ram_block1a831(ram_block1a83),
	.ram_block1a991(ram_block1a99),
	.ram_block1a1151(ram_block1a115),
	.ram_block1a351(ram_block1a35),
	.ram_block1a511(ram_block1a51),
	.ram_block1a310(ram_block1a3),
	.ram_block1a191(ram_block1a19),
	.ram_block1a681(ram_block1a68),
	.ram_block1a841(ram_block1a84),
	.ram_block1a1001(ram_block1a100),
	.ram_block1a1161(ram_block1a116),
	.ram_block1a361(ram_block1a36),
	.ram_block1a521(ram_block1a52),
	.ram_block1a410(ram_block1a4),
	.ram_block1a201(ram_block1a20),
	.ram_block1a691(ram_block1a69),
	.ram_block1a851(ram_block1a85),
	.ram_block1a1011(ram_block1a101),
	.ram_block1a1171(ram_block1a117),
	.ram_block1a371(ram_block1a37),
	.ram_block1a531(ram_block1a53),
	.ram_block1a510(ram_block1a5),
	.ram_block1a211(ram_block1a21),
	.ram_block1a701(ram_block1a70),
	.ram_block1a861(ram_block1a86),
	.ram_block1a1021(ram_block1a102),
	.ram_block1a1181(ram_block1a118),
	.ram_block1a381(ram_block1a38),
	.ram_block1a541(ram_block1a54),
	.ram_block1a610(ram_block1a6),
	.ram_block1a221(ram_block1a22),
	.ram_block1a711(ram_block1a71),
	.ram_block1a871(ram_block1a87),
	.ram_block1a1031(ram_block1a103),
	.ram_block1a1191(ram_block1a119),
	.ram_block1a391(ram_block1a39),
	.ram_block1a551(ram_block1a55),
	.ram_block1a710(ram_block1a7),
	.ram_block1a231(ram_block1a23),
	.ram_block1a721(ram_block1a72),
	.ram_block1a881(ram_block1a88),
	.ram_block1a1041(ram_block1a104),
	.ram_block1a1201(ram_block1a120),
	.ram_block1a401(ram_block1a40),
	.ram_block1a561(ram_block1a56),
	.ram_block1a810(ram_block1a8),
	.ram_block1a241(ram_block1a24),
	.ram_block1a731(ram_block1a73),
	.ram_block1a891(ram_block1a89),
	.ram_block1a1051(ram_block1a105),
	.ram_block1a1211(ram_block1a121),
	.ram_block1a411(ram_block1a41),
	.ram_block1a571(ram_block1a57),
	.ram_block1a910(ram_block1a9),
	.ram_block1a251(ram_block1a25),
	.ram_block1a741(ram_block1a74),
	.ram_block1a901(ram_block1a90),
	.ram_block1a1061(ram_block1a106),
	.ram_block1a1221(ram_block1a122),
	.ram_block1a421(ram_block1a42),
	.ram_block1a581(ram_block1a58),
	.ram_block1a1010(ram_block1a10),
	.ram_block1a261(ram_block1a26),
	.ram_block1a751(ram_block1a75),
	.ram_block1a911(ram_block1a91),
	.ram_block1a1071(ram_block1a107),
	.ram_block1a1231(ram_block1a123),
	.ram_block1a431(ram_block1a43),
	.ram_block1a591(ram_block1a59),
	.ram_block1a1110(ram_block1a11),
	.ram_block1a271(ram_block1a27),
	.ram_block1a761(ram_block1a76),
	.ram_block1a921(ram_block1a92),
	.ram_block1a1081(ram_block1a108),
	.ram_block1a1241(ram_block1a124),
	.ram_block1a441(ram_block1a44),
	.ram_block1a601(ram_block1a60),
	.ram_block1a129(ram_block1a12),
	.ram_block1a281(ram_block1a28),
	.ram_block1a771(ram_block1a77),
	.ram_block1a931(ram_block1a93),
	.ram_block1a1091(ram_block1a109),
	.ram_block1a1251(ram_block1a125),
	.ram_block1a451(ram_block1a45),
	.ram_block1a611(ram_block1a61),
	.ram_block1a131(ram_block1a13),
	.ram_block1a291(ram_block1a29),
	.ram_block1a781(ram_block1a78),
	.ram_block1a941(ram_block1a94),
	.ram_block1a1101(ram_block1a110),
	.ram_block1a1261(ram_block1a126),
	.ram_block1a461(ram_block1a46),
	.ram_block1a621(ram_block1a62),
	.ram_block1a141(ram_block1a14),
	.ram_block1a301(ram_block1a30),
	.ram_block1a791(ram_block1a79),
	.ram_block1a951(ram_block1a95),
	.ram_block1a1111(ram_block1a111),
	.ram_block1a1271(ram_block1a127),
	.ram_block1a471(ram_block1a47),
	.ram_block1a631(ram_block1a63),
	.ram_block1a151(ram_block1a15),
	.ram_block1a311(ram_block1a31),
	.address_a({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.clock0(clock0),
	.clocken0(clocken0));

endmodule

module DDS_48_v1_altsyncram_78g1 (
	ram_block1a641,
	ram_block1a801,
	ram_block1a961,
	ram_block1a1121,
	ram_block1a321,
	ram_block1a481,
	ram_block1a01,
	ram_block1a161,
	ram_block1a651,
	ram_block1a811,
	ram_block1a971,
	ram_block1a1131,
	ram_block1a331,
	ram_block1a491,
	ram_block1a128,
	ram_block1a171,
	ram_block1a661,
	ram_block1a821,
	ram_block1a981,
	ram_block1a1141,
	ram_block1a341,
	ram_block1a501,
	ram_block1a210,
	ram_block1a181,
	ram_block1a671,
	ram_block1a831,
	ram_block1a991,
	ram_block1a1151,
	ram_block1a351,
	ram_block1a511,
	ram_block1a310,
	ram_block1a191,
	ram_block1a681,
	ram_block1a841,
	ram_block1a1001,
	ram_block1a1161,
	ram_block1a361,
	ram_block1a521,
	ram_block1a410,
	ram_block1a201,
	ram_block1a691,
	ram_block1a851,
	ram_block1a1011,
	ram_block1a1171,
	ram_block1a371,
	ram_block1a531,
	ram_block1a510,
	ram_block1a211,
	ram_block1a701,
	ram_block1a861,
	ram_block1a1021,
	ram_block1a1181,
	ram_block1a381,
	ram_block1a541,
	ram_block1a610,
	ram_block1a221,
	ram_block1a711,
	ram_block1a871,
	ram_block1a1031,
	ram_block1a1191,
	ram_block1a391,
	ram_block1a551,
	ram_block1a710,
	ram_block1a231,
	ram_block1a721,
	ram_block1a881,
	ram_block1a1041,
	ram_block1a1201,
	ram_block1a401,
	ram_block1a561,
	ram_block1a810,
	ram_block1a241,
	ram_block1a731,
	ram_block1a891,
	ram_block1a1051,
	ram_block1a1211,
	ram_block1a411,
	ram_block1a571,
	ram_block1a910,
	ram_block1a251,
	ram_block1a741,
	ram_block1a901,
	ram_block1a1061,
	ram_block1a1221,
	ram_block1a421,
	ram_block1a581,
	ram_block1a1010,
	ram_block1a261,
	ram_block1a751,
	ram_block1a911,
	ram_block1a1071,
	ram_block1a1231,
	ram_block1a431,
	ram_block1a591,
	ram_block1a1110,
	ram_block1a271,
	ram_block1a761,
	ram_block1a921,
	ram_block1a1081,
	ram_block1a1241,
	ram_block1a441,
	ram_block1a601,
	ram_block1a129,
	ram_block1a281,
	ram_block1a771,
	ram_block1a931,
	ram_block1a1091,
	ram_block1a1251,
	ram_block1a451,
	ram_block1a611,
	ram_block1a131,
	ram_block1a291,
	ram_block1a781,
	ram_block1a941,
	ram_block1a1101,
	ram_block1a1261,
	ram_block1a461,
	ram_block1a621,
	ram_block1a141,
	ram_block1a301,
	ram_block1a791,
	ram_block1a951,
	ram_block1a1111,
	ram_block1a1271,
	ram_block1a471,
	ram_block1a631,
	ram_block1a151,
	ram_block1a311,
	address_a,
	clock0,
	clocken0)/* synthesis synthesis_greybox=1 */;
output 	ram_block1a641;
output 	ram_block1a801;
output 	ram_block1a961;
output 	ram_block1a1121;
output 	ram_block1a321;
output 	ram_block1a481;
output 	ram_block1a01;
output 	ram_block1a161;
output 	ram_block1a651;
output 	ram_block1a811;
output 	ram_block1a971;
output 	ram_block1a1131;
output 	ram_block1a331;
output 	ram_block1a491;
output 	ram_block1a128;
output 	ram_block1a171;
output 	ram_block1a661;
output 	ram_block1a821;
output 	ram_block1a981;
output 	ram_block1a1141;
output 	ram_block1a341;
output 	ram_block1a501;
output 	ram_block1a210;
output 	ram_block1a181;
output 	ram_block1a671;
output 	ram_block1a831;
output 	ram_block1a991;
output 	ram_block1a1151;
output 	ram_block1a351;
output 	ram_block1a511;
output 	ram_block1a310;
output 	ram_block1a191;
output 	ram_block1a681;
output 	ram_block1a841;
output 	ram_block1a1001;
output 	ram_block1a1161;
output 	ram_block1a361;
output 	ram_block1a521;
output 	ram_block1a410;
output 	ram_block1a201;
output 	ram_block1a691;
output 	ram_block1a851;
output 	ram_block1a1011;
output 	ram_block1a1171;
output 	ram_block1a371;
output 	ram_block1a531;
output 	ram_block1a510;
output 	ram_block1a211;
output 	ram_block1a701;
output 	ram_block1a861;
output 	ram_block1a1021;
output 	ram_block1a1181;
output 	ram_block1a381;
output 	ram_block1a541;
output 	ram_block1a610;
output 	ram_block1a221;
output 	ram_block1a711;
output 	ram_block1a871;
output 	ram_block1a1031;
output 	ram_block1a1191;
output 	ram_block1a391;
output 	ram_block1a551;
output 	ram_block1a710;
output 	ram_block1a231;
output 	ram_block1a721;
output 	ram_block1a881;
output 	ram_block1a1041;
output 	ram_block1a1201;
output 	ram_block1a401;
output 	ram_block1a561;
output 	ram_block1a810;
output 	ram_block1a241;
output 	ram_block1a731;
output 	ram_block1a891;
output 	ram_block1a1051;
output 	ram_block1a1211;
output 	ram_block1a411;
output 	ram_block1a571;
output 	ram_block1a910;
output 	ram_block1a251;
output 	ram_block1a741;
output 	ram_block1a901;
output 	ram_block1a1061;
output 	ram_block1a1221;
output 	ram_block1a421;
output 	ram_block1a581;
output 	ram_block1a1010;
output 	ram_block1a261;
output 	ram_block1a751;
output 	ram_block1a911;
output 	ram_block1a1071;
output 	ram_block1a1231;
output 	ram_block1a431;
output 	ram_block1a591;
output 	ram_block1a1110;
output 	ram_block1a271;
output 	ram_block1a761;
output 	ram_block1a921;
output 	ram_block1a1081;
output 	ram_block1a1241;
output 	ram_block1a441;
output 	ram_block1a601;
output 	ram_block1a129;
output 	ram_block1a281;
output 	ram_block1a771;
output 	ram_block1a931;
output 	ram_block1a1091;
output 	ram_block1a1251;
output 	ram_block1a451;
output 	ram_block1a611;
output 	ram_block1a131;
output 	ram_block1a291;
output 	ram_block1a781;
output 	ram_block1a941;
output 	ram_block1a1101;
output 	ram_block1a1261;
output 	ram_block1a461;
output 	ram_block1a621;
output 	ram_block1a141;
output 	ram_block1a301;
output 	ram_block1a791;
output 	ram_block1a951;
output 	ram_block1a1111;
output 	ram_block1a1271;
output 	ram_block1a471;
output 	ram_block1a631;
output 	ram_block1a151;
output 	ram_block1a311;
input 	[15:0] address_a;
input 	clock0;
input 	clocken0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a64_PORTADATAOUT_bus;
wire [143:0] ram_block1a80_PORTADATAOUT_bus;
wire [143:0] ram_block1a96_PORTADATAOUT_bus;
wire [143:0] ram_block1a112_PORTADATAOUT_bus;
wire [143:0] ram_block1a32_PORTADATAOUT_bus;
wire [143:0] ram_block1a48_PORTADATAOUT_bus;
wire [143:0] ram_block1a0_PORTADATAOUT_bus;
wire [143:0] ram_block1a16_PORTADATAOUT_bus;
wire [143:0] ram_block1a65_PORTADATAOUT_bus;
wire [143:0] ram_block1a81_PORTADATAOUT_bus;
wire [143:0] ram_block1a97_PORTADATAOUT_bus;
wire [143:0] ram_block1a113_PORTADATAOUT_bus;
wire [143:0] ram_block1a33_PORTADATAOUT_bus;
wire [143:0] ram_block1a49_PORTADATAOUT_bus;
wire [143:0] ram_block1a1_PORTADATAOUT_bus;
wire [143:0] ram_block1a17_PORTADATAOUT_bus;
wire [143:0] ram_block1a66_PORTADATAOUT_bus;
wire [143:0] ram_block1a82_PORTADATAOUT_bus;
wire [143:0] ram_block1a98_PORTADATAOUT_bus;
wire [143:0] ram_block1a114_PORTADATAOUT_bus;
wire [143:0] ram_block1a34_PORTADATAOUT_bus;
wire [143:0] ram_block1a50_PORTADATAOUT_bus;
wire [143:0] ram_block1a2_PORTADATAOUT_bus;
wire [143:0] ram_block1a18_PORTADATAOUT_bus;
wire [143:0] ram_block1a67_PORTADATAOUT_bus;
wire [143:0] ram_block1a83_PORTADATAOUT_bus;
wire [143:0] ram_block1a99_PORTADATAOUT_bus;
wire [143:0] ram_block1a115_PORTADATAOUT_bus;
wire [143:0] ram_block1a35_PORTADATAOUT_bus;
wire [143:0] ram_block1a51_PORTADATAOUT_bus;
wire [143:0] ram_block1a3_PORTADATAOUT_bus;
wire [143:0] ram_block1a19_PORTADATAOUT_bus;
wire [143:0] ram_block1a68_PORTADATAOUT_bus;
wire [143:0] ram_block1a84_PORTADATAOUT_bus;
wire [143:0] ram_block1a100_PORTADATAOUT_bus;
wire [143:0] ram_block1a116_PORTADATAOUT_bus;
wire [143:0] ram_block1a36_PORTADATAOUT_bus;
wire [143:0] ram_block1a52_PORTADATAOUT_bus;
wire [143:0] ram_block1a4_PORTADATAOUT_bus;
wire [143:0] ram_block1a20_PORTADATAOUT_bus;
wire [143:0] ram_block1a69_PORTADATAOUT_bus;
wire [143:0] ram_block1a85_PORTADATAOUT_bus;
wire [143:0] ram_block1a101_PORTADATAOUT_bus;
wire [143:0] ram_block1a117_PORTADATAOUT_bus;
wire [143:0] ram_block1a37_PORTADATAOUT_bus;
wire [143:0] ram_block1a53_PORTADATAOUT_bus;
wire [143:0] ram_block1a5_PORTADATAOUT_bus;
wire [143:0] ram_block1a21_PORTADATAOUT_bus;
wire [143:0] ram_block1a70_PORTADATAOUT_bus;
wire [143:0] ram_block1a86_PORTADATAOUT_bus;
wire [143:0] ram_block1a102_PORTADATAOUT_bus;
wire [143:0] ram_block1a118_PORTADATAOUT_bus;
wire [143:0] ram_block1a38_PORTADATAOUT_bus;
wire [143:0] ram_block1a54_PORTADATAOUT_bus;
wire [143:0] ram_block1a6_PORTADATAOUT_bus;
wire [143:0] ram_block1a22_PORTADATAOUT_bus;
wire [143:0] ram_block1a71_PORTADATAOUT_bus;
wire [143:0] ram_block1a87_PORTADATAOUT_bus;
wire [143:0] ram_block1a103_PORTADATAOUT_bus;
wire [143:0] ram_block1a119_PORTADATAOUT_bus;
wire [143:0] ram_block1a39_PORTADATAOUT_bus;
wire [143:0] ram_block1a55_PORTADATAOUT_bus;
wire [143:0] ram_block1a7_PORTADATAOUT_bus;
wire [143:0] ram_block1a23_PORTADATAOUT_bus;
wire [143:0] ram_block1a72_PORTADATAOUT_bus;
wire [143:0] ram_block1a88_PORTADATAOUT_bus;
wire [143:0] ram_block1a104_PORTADATAOUT_bus;
wire [143:0] ram_block1a120_PORTADATAOUT_bus;
wire [143:0] ram_block1a40_PORTADATAOUT_bus;
wire [143:0] ram_block1a56_PORTADATAOUT_bus;
wire [143:0] ram_block1a8_PORTADATAOUT_bus;
wire [143:0] ram_block1a24_PORTADATAOUT_bus;
wire [143:0] ram_block1a73_PORTADATAOUT_bus;
wire [143:0] ram_block1a89_PORTADATAOUT_bus;
wire [143:0] ram_block1a105_PORTADATAOUT_bus;
wire [143:0] ram_block1a121_PORTADATAOUT_bus;
wire [143:0] ram_block1a41_PORTADATAOUT_bus;
wire [143:0] ram_block1a57_PORTADATAOUT_bus;
wire [143:0] ram_block1a9_PORTADATAOUT_bus;
wire [143:0] ram_block1a25_PORTADATAOUT_bus;
wire [143:0] ram_block1a74_PORTADATAOUT_bus;
wire [143:0] ram_block1a90_PORTADATAOUT_bus;
wire [143:0] ram_block1a106_PORTADATAOUT_bus;
wire [143:0] ram_block1a122_PORTADATAOUT_bus;
wire [143:0] ram_block1a42_PORTADATAOUT_bus;
wire [143:0] ram_block1a58_PORTADATAOUT_bus;
wire [143:0] ram_block1a10_PORTADATAOUT_bus;
wire [143:0] ram_block1a26_PORTADATAOUT_bus;
wire [143:0] ram_block1a75_PORTADATAOUT_bus;
wire [143:0] ram_block1a91_PORTADATAOUT_bus;
wire [143:0] ram_block1a107_PORTADATAOUT_bus;
wire [143:0] ram_block1a123_PORTADATAOUT_bus;
wire [143:0] ram_block1a43_PORTADATAOUT_bus;
wire [143:0] ram_block1a59_PORTADATAOUT_bus;
wire [143:0] ram_block1a11_PORTADATAOUT_bus;
wire [143:0] ram_block1a27_PORTADATAOUT_bus;
wire [143:0] ram_block1a76_PORTADATAOUT_bus;
wire [143:0] ram_block1a92_PORTADATAOUT_bus;
wire [143:0] ram_block1a108_PORTADATAOUT_bus;
wire [143:0] ram_block1a124_PORTADATAOUT_bus;
wire [143:0] ram_block1a44_PORTADATAOUT_bus;
wire [143:0] ram_block1a60_PORTADATAOUT_bus;
wire [143:0] ram_block1a12_PORTADATAOUT_bus;
wire [143:0] ram_block1a28_PORTADATAOUT_bus;
wire [143:0] ram_block1a77_PORTADATAOUT_bus;
wire [143:0] ram_block1a93_PORTADATAOUT_bus;
wire [143:0] ram_block1a109_PORTADATAOUT_bus;
wire [143:0] ram_block1a125_PORTADATAOUT_bus;
wire [143:0] ram_block1a45_PORTADATAOUT_bus;
wire [143:0] ram_block1a61_PORTADATAOUT_bus;
wire [143:0] ram_block1a13_PORTADATAOUT_bus;
wire [143:0] ram_block1a29_PORTADATAOUT_bus;
wire [143:0] ram_block1a78_PORTADATAOUT_bus;
wire [143:0] ram_block1a94_PORTADATAOUT_bus;
wire [143:0] ram_block1a110_PORTADATAOUT_bus;
wire [143:0] ram_block1a126_PORTADATAOUT_bus;
wire [143:0] ram_block1a46_PORTADATAOUT_bus;
wire [143:0] ram_block1a62_PORTADATAOUT_bus;
wire [143:0] ram_block1a14_PORTADATAOUT_bus;
wire [143:0] ram_block1a30_PORTADATAOUT_bus;
wire [143:0] ram_block1a79_PORTADATAOUT_bus;
wire [143:0] ram_block1a95_PORTADATAOUT_bus;
wire [143:0] ram_block1a111_PORTADATAOUT_bus;
wire [143:0] ram_block1a127_PORTADATAOUT_bus;
wire [143:0] ram_block1a47_PORTADATAOUT_bus;
wire [143:0] ram_block1a63_PORTADATAOUT_bus;
wire [143:0] ram_block1a15_PORTADATAOUT_bus;
wire [143:0] ram_block1a31_PORTADATAOUT_bus;

assign ram_block1a641 = ram_block1a64_PORTADATAOUT_bus[0];

assign ram_block1a801 = ram_block1a80_PORTADATAOUT_bus[0];

assign ram_block1a961 = ram_block1a96_PORTADATAOUT_bus[0];

assign ram_block1a1121 = ram_block1a112_PORTADATAOUT_bus[0];

assign ram_block1a321 = ram_block1a32_PORTADATAOUT_bus[0];

assign ram_block1a481 = ram_block1a48_PORTADATAOUT_bus[0];

assign ram_block1a01 = ram_block1a0_PORTADATAOUT_bus[0];

assign ram_block1a161 = ram_block1a16_PORTADATAOUT_bus[0];

assign ram_block1a651 = ram_block1a65_PORTADATAOUT_bus[0];

assign ram_block1a811 = ram_block1a81_PORTADATAOUT_bus[0];

assign ram_block1a971 = ram_block1a97_PORTADATAOUT_bus[0];

assign ram_block1a1131 = ram_block1a113_PORTADATAOUT_bus[0];

assign ram_block1a331 = ram_block1a33_PORTADATAOUT_bus[0];

assign ram_block1a491 = ram_block1a49_PORTADATAOUT_bus[0];

assign ram_block1a128 = ram_block1a1_PORTADATAOUT_bus[0];

assign ram_block1a171 = ram_block1a17_PORTADATAOUT_bus[0];

assign ram_block1a661 = ram_block1a66_PORTADATAOUT_bus[0];

assign ram_block1a821 = ram_block1a82_PORTADATAOUT_bus[0];

assign ram_block1a981 = ram_block1a98_PORTADATAOUT_bus[0];

assign ram_block1a1141 = ram_block1a114_PORTADATAOUT_bus[0];

assign ram_block1a341 = ram_block1a34_PORTADATAOUT_bus[0];

assign ram_block1a501 = ram_block1a50_PORTADATAOUT_bus[0];

assign ram_block1a210 = ram_block1a2_PORTADATAOUT_bus[0];

assign ram_block1a181 = ram_block1a18_PORTADATAOUT_bus[0];

assign ram_block1a671 = ram_block1a67_PORTADATAOUT_bus[0];

assign ram_block1a831 = ram_block1a83_PORTADATAOUT_bus[0];

assign ram_block1a991 = ram_block1a99_PORTADATAOUT_bus[0];

assign ram_block1a1151 = ram_block1a115_PORTADATAOUT_bus[0];

assign ram_block1a351 = ram_block1a35_PORTADATAOUT_bus[0];

assign ram_block1a511 = ram_block1a51_PORTADATAOUT_bus[0];

assign ram_block1a310 = ram_block1a3_PORTADATAOUT_bus[0];

assign ram_block1a191 = ram_block1a19_PORTADATAOUT_bus[0];

assign ram_block1a681 = ram_block1a68_PORTADATAOUT_bus[0];

assign ram_block1a841 = ram_block1a84_PORTADATAOUT_bus[0];

assign ram_block1a1001 = ram_block1a100_PORTADATAOUT_bus[0];

assign ram_block1a1161 = ram_block1a116_PORTADATAOUT_bus[0];

assign ram_block1a361 = ram_block1a36_PORTADATAOUT_bus[0];

assign ram_block1a521 = ram_block1a52_PORTADATAOUT_bus[0];

assign ram_block1a410 = ram_block1a4_PORTADATAOUT_bus[0];

assign ram_block1a201 = ram_block1a20_PORTADATAOUT_bus[0];

assign ram_block1a691 = ram_block1a69_PORTADATAOUT_bus[0];

assign ram_block1a851 = ram_block1a85_PORTADATAOUT_bus[0];

assign ram_block1a1011 = ram_block1a101_PORTADATAOUT_bus[0];

assign ram_block1a1171 = ram_block1a117_PORTADATAOUT_bus[0];

assign ram_block1a371 = ram_block1a37_PORTADATAOUT_bus[0];

assign ram_block1a531 = ram_block1a53_PORTADATAOUT_bus[0];

assign ram_block1a510 = ram_block1a5_PORTADATAOUT_bus[0];

assign ram_block1a211 = ram_block1a21_PORTADATAOUT_bus[0];

assign ram_block1a701 = ram_block1a70_PORTADATAOUT_bus[0];

assign ram_block1a861 = ram_block1a86_PORTADATAOUT_bus[0];

assign ram_block1a1021 = ram_block1a102_PORTADATAOUT_bus[0];

assign ram_block1a1181 = ram_block1a118_PORTADATAOUT_bus[0];

assign ram_block1a381 = ram_block1a38_PORTADATAOUT_bus[0];

assign ram_block1a541 = ram_block1a54_PORTADATAOUT_bus[0];

assign ram_block1a610 = ram_block1a6_PORTADATAOUT_bus[0];

assign ram_block1a221 = ram_block1a22_PORTADATAOUT_bus[0];

assign ram_block1a711 = ram_block1a71_PORTADATAOUT_bus[0];

assign ram_block1a871 = ram_block1a87_PORTADATAOUT_bus[0];

assign ram_block1a1031 = ram_block1a103_PORTADATAOUT_bus[0];

assign ram_block1a1191 = ram_block1a119_PORTADATAOUT_bus[0];

assign ram_block1a391 = ram_block1a39_PORTADATAOUT_bus[0];

assign ram_block1a551 = ram_block1a55_PORTADATAOUT_bus[0];

assign ram_block1a710 = ram_block1a7_PORTADATAOUT_bus[0];

assign ram_block1a231 = ram_block1a23_PORTADATAOUT_bus[0];

assign ram_block1a721 = ram_block1a72_PORTADATAOUT_bus[0];

assign ram_block1a881 = ram_block1a88_PORTADATAOUT_bus[0];

assign ram_block1a1041 = ram_block1a104_PORTADATAOUT_bus[0];

assign ram_block1a1201 = ram_block1a120_PORTADATAOUT_bus[0];

assign ram_block1a401 = ram_block1a40_PORTADATAOUT_bus[0];

assign ram_block1a561 = ram_block1a56_PORTADATAOUT_bus[0];

assign ram_block1a810 = ram_block1a8_PORTADATAOUT_bus[0];

assign ram_block1a241 = ram_block1a24_PORTADATAOUT_bus[0];

assign ram_block1a731 = ram_block1a73_PORTADATAOUT_bus[0];

assign ram_block1a891 = ram_block1a89_PORTADATAOUT_bus[0];

assign ram_block1a1051 = ram_block1a105_PORTADATAOUT_bus[0];

assign ram_block1a1211 = ram_block1a121_PORTADATAOUT_bus[0];

assign ram_block1a411 = ram_block1a41_PORTADATAOUT_bus[0];

assign ram_block1a571 = ram_block1a57_PORTADATAOUT_bus[0];

assign ram_block1a910 = ram_block1a9_PORTADATAOUT_bus[0];

assign ram_block1a251 = ram_block1a25_PORTADATAOUT_bus[0];

assign ram_block1a741 = ram_block1a74_PORTADATAOUT_bus[0];

assign ram_block1a901 = ram_block1a90_PORTADATAOUT_bus[0];

assign ram_block1a1061 = ram_block1a106_PORTADATAOUT_bus[0];

assign ram_block1a1221 = ram_block1a122_PORTADATAOUT_bus[0];

assign ram_block1a421 = ram_block1a42_PORTADATAOUT_bus[0];

assign ram_block1a581 = ram_block1a58_PORTADATAOUT_bus[0];

assign ram_block1a1010 = ram_block1a10_PORTADATAOUT_bus[0];

assign ram_block1a261 = ram_block1a26_PORTADATAOUT_bus[0];

assign ram_block1a751 = ram_block1a75_PORTADATAOUT_bus[0];

assign ram_block1a911 = ram_block1a91_PORTADATAOUT_bus[0];

assign ram_block1a1071 = ram_block1a107_PORTADATAOUT_bus[0];

assign ram_block1a1231 = ram_block1a123_PORTADATAOUT_bus[0];

assign ram_block1a431 = ram_block1a43_PORTADATAOUT_bus[0];

assign ram_block1a591 = ram_block1a59_PORTADATAOUT_bus[0];

assign ram_block1a1110 = ram_block1a11_PORTADATAOUT_bus[0];

assign ram_block1a271 = ram_block1a27_PORTADATAOUT_bus[0];

assign ram_block1a761 = ram_block1a76_PORTADATAOUT_bus[0];

assign ram_block1a921 = ram_block1a92_PORTADATAOUT_bus[0];

assign ram_block1a1081 = ram_block1a108_PORTADATAOUT_bus[0];

assign ram_block1a1241 = ram_block1a124_PORTADATAOUT_bus[0];

assign ram_block1a441 = ram_block1a44_PORTADATAOUT_bus[0];

assign ram_block1a601 = ram_block1a60_PORTADATAOUT_bus[0];

assign ram_block1a129 = ram_block1a12_PORTADATAOUT_bus[0];

assign ram_block1a281 = ram_block1a28_PORTADATAOUT_bus[0];

assign ram_block1a771 = ram_block1a77_PORTADATAOUT_bus[0];

assign ram_block1a931 = ram_block1a93_PORTADATAOUT_bus[0];

assign ram_block1a1091 = ram_block1a109_PORTADATAOUT_bus[0];

assign ram_block1a1251 = ram_block1a125_PORTADATAOUT_bus[0];

assign ram_block1a451 = ram_block1a45_PORTADATAOUT_bus[0];

assign ram_block1a611 = ram_block1a61_PORTADATAOUT_bus[0];

assign ram_block1a131 = ram_block1a13_PORTADATAOUT_bus[0];

assign ram_block1a291 = ram_block1a29_PORTADATAOUT_bus[0];

assign ram_block1a781 = ram_block1a78_PORTADATAOUT_bus[0];

assign ram_block1a941 = ram_block1a94_PORTADATAOUT_bus[0];

assign ram_block1a1101 = ram_block1a110_PORTADATAOUT_bus[0];

assign ram_block1a1261 = ram_block1a126_PORTADATAOUT_bus[0];

assign ram_block1a461 = ram_block1a46_PORTADATAOUT_bus[0];

assign ram_block1a621 = ram_block1a62_PORTADATAOUT_bus[0];

assign ram_block1a141 = ram_block1a14_PORTADATAOUT_bus[0];

assign ram_block1a301 = ram_block1a30_PORTADATAOUT_bus[0];

assign ram_block1a791 = ram_block1a79_PORTADATAOUT_bus[0];

assign ram_block1a951 = ram_block1a95_PORTADATAOUT_bus[0];

assign ram_block1a1111 = ram_block1a111_PORTADATAOUT_bus[0];

assign ram_block1a1271 = ram_block1a127_PORTADATAOUT_bus[0];

assign ram_block1a471 = ram_block1a47_PORTADATAOUT_bus[0];

assign ram_block1a631 = ram_block1a63_PORTADATAOUT_bus[0];

assign ram_block1a151 = ram_block1a15_PORTADATAOUT_bus[0];

assign ram_block1a311 = ram_block1a31_PORTADATAOUT_bus[0];

arriav_ram_block ram_block1a64(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a64_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a64.clk0_core_clock_enable = "ena0";
defparam ram_block1a64.clk0_input_clock_enable = "ena0";
defparam ram_block1a64.clk0_output_clock_enable = "ena0";
defparam ram_block1a64.data_interleave_offset_in_bits = 1;
defparam ram_block1a64.data_interleave_width_in_bits = 1;
defparam ram_block1a64.init_file = "DDS_48_v1_nco_ii_0_cos.hex";
defparam ram_block1a64.init_file_layout = "port_a";
defparam ram_block1a64.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0121|altsyncram:altsyncram_component0|altsyncram_78g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a64.operation_mode = "rom";
defparam ram_block1a64.port_a_address_clear = "none";
defparam ram_block1a64.port_a_address_width = 13;
defparam ram_block1a64.port_a_data_out_clear = "none";
defparam ram_block1a64.port_a_data_out_clock = "clock0";
defparam ram_block1a64.port_a_data_width = 1;
defparam ram_block1a64.port_a_first_address = 32768;
defparam ram_block1a64.port_a_first_bit_number = 0;
defparam ram_block1a64.port_a_last_address = 40959;
defparam ram_block1a64.port_a_logical_ram_depth = 65536;
defparam ram_block1a64.port_a_logical_ram_width = 16;
defparam ram_block1a64.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a64.ram_block_type = "auto";
defparam ram_block1a64.mem_init3 = "1E0F07C3E0F07C1F0F83E0F83E0F83E0F81F07C0F81F07E0FC0F81F81F03F03F03F03F81F81FC0FE07F01FC07E03FC07F01FE03FC03F807F803FC03FE01FF007FC00FF801FF801FFC00FFE003FFC003FFC001FFF0003FFF8000FFFF00003FFFF00000FFFFFE000000FFFFFFFE0000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000001FFFFFFF8000001FFFFF800007FFFE0000FFFF0001FFF8001FFF0007FF8007FF001FFC00FFC00FFC00FF803FE00FF007F807F807F807F00FE01FC07F01FC0FE03F01F80FC0FC07E07E0FC0FC0F81F83F07E0F81F07C1F83E0F83E0F87C1F0783E1F0783C1E0F0F87C3C1E1E0F0F0F0F8787878787";
defparam ram_block1a64.mem_init2 = "8F0F0F0E1E1E3C387870E1E3C7870E1C3871E3C78E1C78E1C70E3C71C38E3871C71C38E38E38E38E38E38E39C71C718E38C71CE38C718E31CE31C639CE31CE718C739CE318C6318C6318C6739CE6319CE6339CC67319CC673398CC6633198CCE67331998CCC666333319999CCCCCC6666666666333333333333326666666666CCCCCD9999B3336666CCC999332664CD99B3264CD993264C993264C99366C99366C9B264D9364D93649B26C93649B24DB26D924DB249B64926DB24926DB6D924924924DB6DB6DA492492492DB6DA4925B6D2496DA496D24B692DA4B692DA4B49692D25A5B4B4B49696969696969694B4B4A5A5AD2D694B5A52D694A5AD6B5A529";
defparam ram_block1a64.mem_init1 = "4A5294A56B5AD4A56B5A95AD4AD4A56A56AD4AD4A95AB52A54A952A54A952AD5AA55AA55AAD52A954AA552A955AA955AAB556AA9552AA9554AAA5554AAA95556AAAA55555AAAAA9555555AAAAAAAA95555555555555555AAAAAAAAAAD5555555555555554AAAAAAAAD555554AAAAAD55552AAA95554AAA9555AAA9556AAB554AA9552AB556AA552AB55AAD56A954AB54AB54A956AD52A54A952B56AD4A95A952B52B52B52B5A95AD4A56B5A94A5295AD6B5A5294A52D6B4A5AD296B4A5A52D2D6969694B4B4B4B4B4969696D2D25A5B49692D25B496D25B692DB492DB4925B6D24925B6DB6D249249249249249B6DB6D924936DB24936C926D924DB26D926C93";
defparam ram_block1a64.mem_init0 = "649B26C9B26C9B26C9B364D9B264C9B366CD9B3664C99B3266CC99B33666CCC9999333266664CCCCCC99999999999999999999999999CCCCCCE666673331999CCC66633199CCE673399CC673398CE6319CC6339CC6318CE739CE739CE318C739C631CE31CE31CE39C738E71C638E31C71C738E38E38E38E38E1C71C70E38E1C70E3C71E3870E3C78F1E3C78F1E1C3C7870F0E1E1E1E3C3C3C3C3C1E1E1E0F0F0787C3E1F0F87C1E0F83C1F07C1F07C1F03E0F81F03E07E0FC0FC0FC0FC0FC07E03F01FC07F01FC07F80FF00FF00FF007FC01FF007FE00FFE007FF001FFE001FFF0003FFF0000FFFF00001FFFFE000001FFFFFFF00000000003FFFFFFFFFFFFFF";

arriav_ram_block ram_block1a80(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a80_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a80.clk0_core_clock_enable = "ena0";
defparam ram_block1a80.clk0_input_clock_enable = "ena0";
defparam ram_block1a80.clk0_output_clock_enable = "ena0";
defparam ram_block1a80.data_interleave_offset_in_bits = 1;
defparam ram_block1a80.data_interleave_width_in_bits = 1;
defparam ram_block1a80.init_file = "DDS_48_v1_nco_ii_0_cos.hex";
defparam ram_block1a80.init_file_layout = "port_a";
defparam ram_block1a80.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0121|altsyncram:altsyncram_component0|altsyncram_78g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a80.operation_mode = "rom";
defparam ram_block1a80.port_a_address_clear = "none";
defparam ram_block1a80.port_a_address_width = 13;
defparam ram_block1a80.port_a_data_out_clear = "none";
defparam ram_block1a80.port_a_data_out_clock = "clock0";
defparam ram_block1a80.port_a_data_width = 1;
defparam ram_block1a80.port_a_first_address = 40960;
defparam ram_block1a80.port_a_first_bit_number = 0;
defparam ram_block1a80.port_a_last_address = 49151;
defparam ram_block1a80.port_a_logical_ram_depth = 65536;
defparam ram_block1a80.port_a_logical_ram_width = 16;
defparam ram_block1a80.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a80.ram_block_type = "auto";
defparam ram_block1a80.mem_init3 = "B56AD5AB56AD52A54A952A54A952A54A952A55AB56AD5AB56AD5AB56A952A54A952A54AB56AD5AB56AD5AA54A952A54AB56AD5AB54A952A54AB56AD5AA54A952AD5AB56A952A55AB56A952A55AB56A952A55AB54A952AD5AA54AB56A952AD5AA54AB56A952AD5AA55AB54AB56A956AD52AD5AA55AA54AB54AB56A956A956A956A956AD52AD52AD52A956A956A956A956A954AB54AB55AA55AAD52AD56A954AB54AA552AD56A954AA55AAD56A954AA552A954AB55AAD56AB552A954AA552A955AAD56AA552AB55AA954AAD56AA556AA552AB552AB552AB552AA556AA556AAD54AA955AAB556AA554AA9552AA554AA9556AAD55AAA554AAB554AAB554AAB554AAB";
defparam ram_block1a80.mem_init2 = "555AAA5552AAD556AAB555AAA9554AAAD556AAA5556AAAD554AAA9555AAAB5554AAA95556AAA95556AAAB5555AAAAD5554AAAAD5555AAAA955556AAAA955554AAAAA555556AAAAAD555552AAAAA9555555AAAAAAA55555552AAAAAAAD55555555AAAAAAAAAB55555555554AAAAAAAAAAAAA955555555555555555556AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAD5555555555555555556AAAAAAAAAAAAB55555555552AAAAAAAA955555556AAAAAAA5555554AAAAAA555555AAAAAB55555AAAAAD55552AAAA55556AAAA55552AAAD5556AAAD5552AAA5556AAA5556AAA5552AAB554AAA5552AAD552AAD55AAA554AA9552AA554AA955AA9";
defparam ram_block1a80.mem_init1 = "552AB552A955AA954AAD56AB55AA956AB55AAD56A954AB54AA55AA55AA55AA55AA54AB54A956AD52A54A956AD5AB56AD5AB56AD4A952B56AD4A95AB52A56A56AD4AD4AD5A95A95A95AD4AD4AD4A56A52B5295AD4AD6B5295AD4A5295AD6A5294A5295AD6B5AD6B5AD694A5294A5AD6B4A52D6B4A52D6B4A5AD296B4A5A52D696B4B5A5AD2D29696B4B4B4A5A5A5A5A5A5A5A5A5A5A5A5A5A5B4B4B4B69696D2D25A5B4B696D2DA5B49692DA5B496D25B496D25B492DA496D24B6D25B6D24B6D2496DB4925B6DA4924B6DB6D2492492DB6DB6DB6DB6DB6DB6DB6DB6DB6D924924936DB6D924936DB64926DB24936D926DB249B649B649B649B649B64DB26D936C";
defparam ram_block1a80.mem_init0 = "9B24D93649B26C9B26C9B26C9B364D9366C9B364C9B364C9B366CD93264C993266CD9B3264CD9B3266CC99B33664CC999332664CCD99933326664CCC99999333336666666CCCCCCCCC9999999999999999999999999999CCCCCCCCC66666673333399998CCCE6663333999CCC66633399CCC6633199CC6633198CE63319CC67319CC67318CE6319CE6318CE739CC6318C6318C6318C6318E739C6318E738C739C639C639C638C738E71CE39C718E39C71CE38E31C71C738E38E38E38E38E38E38E38F1C71C70E38E1C71E38F1C78E3C70E3C70E3C78F1C3870E1C3870E1E3C7870F1E1C3C387870F0F0E1E1E1E1E1E1E1E1E1E1E1F0F0F078783C3E1F0F0783C";

arriav_ram_block ram_block1a96(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a96_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a96.clk0_core_clock_enable = "ena0";
defparam ram_block1a96.clk0_input_clock_enable = "ena0";
defparam ram_block1a96.clk0_output_clock_enable = "ena0";
defparam ram_block1a96.data_interleave_offset_in_bits = 1;
defparam ram_block1a96.data_interleave_width_in_bits = 1;
defparam ram_block1a96.init_file = "DDS_48_v1_nco_ii_0_cos.hex";
defparam ram_block1a96.init_file_layout = "port_a";
defparam ram_block1a96.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0121|altsyncram:altsyncram_component0|altsyncram_78g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a96.operation_mode = "rom";
defparam ram_block1a96.port_a_address_clear = "none";
defparam ram_block1a96.port_a_address_width = 13;
defparam ram_block1a96.port_a_data_out_clear = "none";
defparam ram_block1a96.port_a_data_out_clock = "clock0";
defparam ram_block1a96.port_a_data_width = 1;
defparam ram_block1a96.port_a_first_address = 49152;
defparam ram_block1a96.port_a_first_bit_number = 0;
defparam ram_block1a96.port_a_last_address = 57343;
defparam ram_block1a96.port_a_logical_ram_depth = 65536;
defparam ram_block1a96.port_a_logical_ram_width = 16;
defparam ram_block1a96.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a96.ram_block_type = "auto";
defparam ram_block1a96.mem_init3 = "783C1E1F0F8783C3C1E1E1F0F0F0F0F0F0F0F0F0F0F0E1E1E1C3C387870F1E1C3C78F0E1C3870E1C3871E3C78E1C78E1C78E3C71E38F1C70E38E1C71C71E38E38E38E38E38E38E38E39C71C718E38E71C738E31C738E71CE39C638C738C738C739C639CE318C739CE318C6318C6318C6318C6739CE6318CE7318CE6319CC67319CC673198CE633198CC6733198CC66733998CCC6673339998CCCE6663333399999CCCCCCC6666666673333333333333333333333333332666666666CCCCCCD99999333326664CCC99993336664CC999332664CD99B3266CC99B3664C99B366CC993264C99366CD9B264D9B264D9B26CD9364D9B26C9B26C9B26C9B24D93649B2";
defparam ram_block1a96.mem_init2 = "6D936C9B64DB24DB24DB24DB24DB249B6C936D9249B6C924DB6D924936DB6D924924936DB6DB6DB6DB6DB6DB6DB6DB6DB692492496DB6DA4924B6DB4925B6D2496DA496DB496DA496D24B6925B496D25B496D25B4B692D25B4B696D2DA5B4B49696D2D2DA5A5A5B4B4B4B4B4B4B4B4B4B4B4B4B4B4A5A5A5AD2D29696B4B5A5AD2D694B4A5AD296B4A5AD694A5AD694A5AD6B4A5294A52D6B5AD6B5AD6B5294A5294AD6B5294A56B5295AD6A56B5295A94AD4A56A56A56B52B52B52B56A56A56AD4AD4A95AB52A56AD5A952A56AD5AB56AD5AB56AD52A54A956AD52A55AA54AB54AB54AB54AB54AA55AA552AD56AB55AAD52AB55AAD56AA552AB552A955AA955";
defparam ram_block1a96.mem_init1 = "2AB552AA554AA9552AA554AAB556AA9556AA9554AAA555AAA9554AAAD554AAAD554AAA95556AAAD5556AAA95554AAAAD5554AAAA955556AAAAB55555AAAAAB555554AAAAAA5555554AAAAAAAD55555552AAAAAAAA95555555555AAAAAAAAAAAAAD5555555555555555556AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAD55555555555555555552AAAAAAAAAAAAA55555555555AAAAAAAAAB555555556AAAAAAA95555554AAAAAAB5555552AAAAA9555556AAAAAD55554AAAAA555552AAAAD55552AAAB55556AAAA55556AAAB5555AAAAD5552AAAD5552AAA5555AAAB5552AAA5556AAAD554AAAD556AAA5552AAB555AAAD556AA9554AAB555";
defparam ram_block1a96.mem_init0 = "AAA555AAA555AAA555AAA554AAB556AAD552AA554AA9552AA554AAD55AAB552AA556AAD54AAD54AA955AA955AA955AA954AAD54AAD56AA552AB55AA954AAD56AB552A954AA552A955AAD56AB55AA552A954AA552AD56AB54AA552AD56A954AA55AA552AD56A956AB54AB55AA55AA552AD52AD52AD52AD52A956A956A956AD52AD52AD52AD52AD5AA55AA54AB54AB56A956AD52AD5AA55AB54AB56A952AD5AA54AB56A952AD5AA54AB56A952A55AB54A952AD5AB54A952AD5AB54A952AD5AB56A952A54AB56AD5AA54A952A55AB56AD5AA54A952A54AB56AD5AB56AD5AA54A952A54A952AD5AB56AD5AB56AD5AB54A952A54A952A54A952A54A956AD5AB56AD5A";

arriav_ram_block ram_block1a112(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a112_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a112.clk0_core_clock_enable = "ena0";
defparam ram_block1a112.clk0_input_clock_enable = "ena0";
defparam ram_block1a112.clk0_output_clock_enable = "ena0";
defparam ram_block1a112.data_interleave_offset_in_bits = 1;
defparam ram_block1a112.data_interleave_width_in_bits = 1;
defparam ram_block1a112.init_file = "DDS_48_v1_nco_ii_0_cos.hex";
defparam ram_block1a112.init_file_layout = "port_a";
defparam ram_block1a112.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0121|altsyncram:altsyncram_component0|altsyncram_78g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a112.operation_mode = "rom";
defparam ram_block1a112.port_a_address_clear = "none";
defparam ram_block1a112.port_a_address_width = 13;
defparam ram_block1a112.port_a_data_out_clear = "none";
defparam ram_block1a112.port_a_data_out_clock = "clock0";
defparam ram_block1a112.port_a_data_width = 1;
defparam ram_block1a112.port_a_first_address = 57344;
defparam ram_block1a112.port_a_first_bit_number = 0;
defparam ram_block1a112.port_a_last_address = 65535;
defparam ram_block1a112.port_a_logical_ram_depth = 65536;
defparam ram_block1a112.port_a_logical_ram_width = 16;
defparam ram_block1a112.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a112.ram_block_type = "auto";
defparam ram_block1a112.mem_init3 = "FFFFFFFFFFFFFF80000000001FFFFFFF000000FFFFF00001FFFE0001FFF8001FFF000FFF001FFC00FFE00FFC01FF007FC01FE01FE01FE03FC07F01FC07F01F80FC07E07E07E07E07E0FC0F81F03E0F81F07C1F07C1F0783E0F07C3E1F0F87C3C1E1E0F0F0F07878787878F0F0F0E1E1C3C7870F1E3C78F1E3C78E1C38F1C78E1C70E38E1C71C70E38E38E38E38E39C71C718E38C71CE39C738E718E718E718C739C6318E739CE739CE6318C67398C67318CE63399CC673399CCE6733198CCC6673331999CCCCCE666667333333333333333333333333326666664CCCC99993332666CCD99B3266CC99B3264CD9B366CD9B264C9B364D9B26C9B26C9B26C9B24D";
defparam ram_block1a112.mem_init2 = "926C936C9B64936C926D9249B6D924936DB6DB2492492492492496DB6DB492496DB4925B6925B692DB496D25B49692D25B4B49696D2D2D25A5A5A5A5A52D2D2D69694B4A5AD296B4A5AD694A5294B5AD6B5294A52B5AD4A56B52B5A95A95A95A952B52A56AD5A952A54A956AD52A55AA55AA552AD56AB55AA954AAD55AA9552AA555AAAD552AAB5552AAA55552AAA955556AAAAA5555556AAAAAAAA55555555555555556AAAAAAAAAB55555555555555552AAAAAAAB5555552AAAAB55554AAAAD5552AAA5554AAA5552AA9552AAD55AAB552AB552A954AA552A956AB54AB54AB56A952A54A952A54A95AB52A56A56AD4AD4A56A56B52B5AD4A56B5AD4A5294A5";
defparam ram_block1a112.mem_init1 = "294B5AD6B4A52D694B5A52D696B4B4A5A5A52D2D2D2D2D2D2D25A5A5B4B49692D25A4B692DA4B692DA496D24B6D2496DB4924B6DB6924924924B6DB6DB64924924936DB6C9249B6C924DB249B64936C9B649B24D926C9B24D9364D9364C9B26CD9326CD93264C993264C9933664C99B33664CC999332666CCCD999B3333666666CCCCCCCCCC99999999999998CCCCCCCCCC666667333319998CCC666333199CCE6633198CC663399CC67319CC67398CE7318CE739CC6318C6318C6318E739C631CE718E738C718E718E31C638E71C638E31C71C738E38E38E38E38E38E3871C71C38E3871C78E1C70E3C70E3C78F1C3870E1C3C78F0E1C3C3878F0F0E1E1E1E3";
defparam ram_block1a112.mem_init0 = "C3C3C3C3C3E1E1E1E0F0F0787C3E1E0F0783C1F0F83C1F07C3E0F83E0F83F07C1F03E0FC1F83F03E07E07E0FC0FC07E07E03F01F80FE07F01FC07F00FE01FC03FC03FC03FC01FE00FF803FE007FE007FE007FF001FFC003FFC001FFF0003FFF0001FFFE0000FFFFC00003FFFFF0000003FFFFFFF00000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000FFFFFFFE000000FFFFFE00001FFFF80001FFFE0003FFF8001FFF0007FF8007FF800FFE007FF003FF003FE007FC01FF00FF807F803FC03F807F80FF01FC07F80FC07F01FC0FE07F03F03F81F81F81F81F03F03E07E0FC1F03E07C1F03E0F83E0F83E0F83E1F07C1E0F87C1E0F0";

arriav_ram_block ram_block1a32(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a32_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a32.clk0_core_clock_enable = "ena0";
defparam ram_block1a32.clk0_input_clock_enable = "ena0";
defparam ram_block1a32.clk0_output_clock_enable = "ena0";
defparam ram_block1a32.data_interleave_offset_in_bits = 1;
defparam ram_block1a32.data_interleave_width_in_bits = 1;
defparam ram_block1a32.init_file = "DDS_48_v1_nco_ii_0_cos.hex";
defparam ram_block1a32.init_file_layout = "port_a";
defparam ram_block1a32.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0121|altsyncram:altsyncram_component0|altsyncram_78g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a32.operation_mode = "rom";
defparam ram_block1a32.port_a_address_clear = "none";
defparam ram_block1a32.port_a_address_width = 13;
defparam ram_block1a32.port_a_data_out_clear = "none";
defparam ram_block1a32.port_a_data_out_clock = "clock0";
defparam ram_block1a32.port_a_data_width = 1;
defparam ram_block1a32.port_a_first_address = 16384;
defparam ram_block1a32.port_a_first_bit_number = 0;
defparam ram_block1a32.port_a_last_address = 24575;
defparam ram_block1a32.port_a_logical_ram_depth = 65536;
defparam ram_block1a32.port_a_logical_ram_width = 16;
defparam ram_block1a32.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a32.ram_block_type = "auto";
defparam ram_block1a32.mem_init3 = "783C1E1F0F8783C3C1E1E1F0F0F0F0F0F0F0F0F0F0F0E1E1E1C3C387870F1E1C3C78F0E1C3870E1C3871E3C78E1C78E1C78E3C71E38F1C70E38E1C71C71E38E38E38E38E38E38E38E39C71C718E38E71C738E31C738E71CE39C638C738C738C739C639CE318C739CE318C6318C6318C6318C6739CE6318CE7318CE6319CC67319CC673198CE633198CC6733198CC66733998CCC6673339998CCCE6663333399999CCCCCCC6666666673333333333333333333333333332666666666CCCCCCD99999333326664CCC99993336664CC999332664CD99B3266CC99B3664C99B366CC993264C99366CD9B264D9B264D9B26CD9364D9B26C9B26C9B26C9B24D93649B2";
defparam ram_block1a32.mem_init2 = "6D936C9B64DB24DB24DB24DB24DB249B6C936D9249B6C924DB6D924936DB6D924924936DB6DB6DB6DB6DB6DB6DB6DB6DB692492496DB6DA4924B6DB4925B6D2496DA496DB496DA496D24B6925B496D25B496D25B4B692D25B4B696D2DA5B4B49696D2D2DA5A5A5B4B4B4B4B4B4B4B4B4B4B4B4B4B4A5A5A5AD2D29696B4B5A5AD2D694B4A5AD296B4A5AD694A5AD694A5AD6B4A5294A52D6B5AD6B5AD6B5294A5294AD6B5294A56B5295AD6A56B5295A94AD4A56A56A56B52B52B52B56A56A56AD4AD4A95AB52A56AD5A952A56AD5AB56AD5AB56AD52A54A956AD52A55AA54AB54AB54AB54AB54AA55AA552AD56AB55AAD52AB55AAD56AA552AB552A955AA955";
defparam ram_block1a32.mem_init1 = "2AB552AA554AA9552AA554AAB556AA9556AA9554AAA555AAA9554AAAD554AAAD554AAA95556AAAD5556AAA95554AAAAD5554AAAA955556AAAAB55555AAAAAB555554AAAAAA5555554AAAAAAAD55555552AAAAAAAA95555555555AAAAAAAAAAAAAD5555555555555555556AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAD55555555555555555552AAAAAAAAAAAAA55555555555AAAAAAAAAB555555556AAAAAAA95555554AAAAAAB5555552AAAAA9555556AAAAAD55554AAAAA555552AAAAD55552AAAB55556AAAA55556AAAB5555AAAAD5552AAAD5552AAA5555AAAB5552AAA5556AAAD554AAAD556AAA5552AAB555AAAD556AA9554AAB555";
defparam ram_block1a32.mem_init0 = "AAA555AAA555AAA555AAA554AAB556AAD552AA554AA9552AA554AAD55AAB552AA556AAD54AAD54AA955AA955AA955AA954AAD54AAD56AA552AB55AA954AAD56AB552A954AA552A955AAD56AB55AA552A954AA552AD56AB54AA552AD56A954AA55AA552AD56A956AB54AB55AA55AA552AD52AD52AD52AD52A956A956A956AD52AD52AD52AD52AD5AA55AA54AB54AB56A956AD52AD5AA55AB54AB56A952AD5AA54AB56A952AD5AA54AB56A952A55AB54A952AD5AB54A952AD5AB54A952AD5AB56A952A54AB56AD5AA54A952A55AB56AD5AA54A952A54AB56AD5AB56AD5AA54A952A54A952AD5AB56AD5AB56AD5AB54A952A54A952A54A952A54A956AD5AB56AD5A";

arriav_ram_block ram_block1a48(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a48_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a48.clk0_core_clock_enable = "ena0";
defparam ram_block1a48.clk0_input_clock_enable = "ena0";
defparam ram_block1a48.clk0_output_clock_enable = "ena0";
defparam ram_block1a48.data_interleave_offset_in_bits = 1;
defparam ram_block1a48.data_interleave_width_in_bits = 1;
defparam ram_block1a48.init_file = "DDS_48_v1_nco_ii_0_cos.hex";
defparam ram_block1a48.init_file_layout = "port_a";
defparam ram_block1a48.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0121|altsyncram:altsyncram_component0|altsyncram_78g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a48.operation_mode = "rom";
defparam ram_block1a48.port_a_address_clear = "none";
defparam ram_block1a48.port_a_address_width = 13;
defparam ram_block1a48.port_a_data_out_clear = "none";
defparam ram_block1a48.port_a_data_out_clock = "clock0";
defparam ram_block1a48.port_a_data_width = 1;
defparam ram_block1a48.port_a_first_address = 24576;
defparam ram_block1a48.port_a_first_bit_number = 0;
defparam ram_block1a48.port_a_last_address = 32767;
defparam ram_block1a48.port_a_logical_ram_depth = 65536;
defparam ram_block1a48.port_a_logical_ram_width = 16;
defparam ram_block1a48.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a48.ram_block_type = "auto";
defparam ram_block1a48.mem_init3 = "FFFFFFFFFFFFFF80000000001FFFFFFF000000FFFFF00001FFFE0001FFF8001FFF000FFF001FFC00FFE00FFC01FF007FC01FE01FE01FE03FC07F01FC07F01F80FC07E07E07E07E07E0FC0F81F03E0F81F07C1F07C1F0783E0F07C3E1F0F87C3C1E1E0F0F0F07878787878F0F0F0E1E1C3C7870F1E3C78F1E3C78E1C38F1C78E1C70E38E1C71C70E38E38E38E38E39C71C718E38C71CE39C738E718E718E718C739C6318E739CE739CE6318C67398C67318CE63399CC673399CCE6733198CCC6673331999CCCCCE666667333333333333333333333333326666664CCCC99993332666CCD99B3266CC99B3264CD9B366CD9B264C9B364D9B26C9B26C9B26C9B24D";
defparam ram_block1a48.mem_init2 = "926C936C9B64936C926D9249B6D924936DB6DB2492492492492496DB6DB492496DB4925B6925B692DB496D25B49692D25B4B49696D2D2D25A5A5A5A5A52D2D2D69694B4A5AD296B4A5AD694A5294B5AD6B5294A52B5AD4A56B52B5A95A95A95A952B52A56AD5A952A54A956AD52A55AA55AA552AD56AB55AA954AAD55AA9552AA555AAAD552AAB5552AAA55552AAA955556AAAAA5555556AAAAAAAA55555555555555556AAAAAAAAAB55555555555555552AAAAAAAB5555552AAAAB55554AAAAD5552AAA5554AAA5552AA9552AAD55AAB552AB552A954AA552A956AB54AB54AB56A952A54A952A54A95AB52A56A56AD4AD4A56A56B52B5AD4A56B5AD4A5294A5";
defparam ram_block1a48.mem_init1 = "294B5AD6B4A52D694B5A52D696B4B4A5A5A52D2D2D2D2D2D2D25A5A5B4B49692D25A4B692DA4B692DA496D24B6D2496DB4924B6DB6924924924B6DB6DB64924924936DB6C9249B6C924DB249B64936C9B649B24D926C9B24D9364D9364C9B26CD9326CD93264C993264C9933664C99B33664CC999332666CCCD999B3333666666CCCCCCCCCC99999999999998CCCCCCCCCC666667333319998CCC666333199CCE6633198CC663399CC67319CC67398CE7318CE739CC6318C6318C6318E739C631CE718E738C718E718E31C638E71C638E31C71C738E38E38E38E38E38E3871C71C38E3871C78E1C70E3C70E3C78F1C3870E1C3C78F0E1C3C3878F0F0E1E1E1E3";
defparam ram_block1a48.mem_init0 = "C3C3C3C3C3E1E1E1E0F0F0787C3E1E0F0783C1F0F83C1F07C3E0F83E0F83F07C1F03E0FC1F83F03E07E07E0FC0FC07E07E03F01F80FE07F01FC07F00FE01FC03FC03FC03FC01FE00FF803FE007FE007FE007FF001FFC003FFC001FFF0003FFF0001FFFE0000FFFFC00003FFFFF0000003FFFFFFF00000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000FFFFFFFE000000FFFFFE00001FFFF80001FFFE0003FFF8001FFF0007FF8007FF800FFE007FF003FF003FE007FC01FF00FF807F803FC03F807F80FF01FC07F80FC07F01FC0FE07F03F03F81F81F81F81F03F03E07E0FC1F03E07C1F03E0F83E0F83E0F83E1F07C1E0F87C1E0F0";

arriav_ram_block ram_block1a0(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a0_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.clk0_input_clock_enable = "ena0";
defparam ram_block1a0.clk0_output_clock_enable = "ena0";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.init_file = "DDS_48_v1_nco_ii_0_cos.hex";
defparam ram_block1a0.init_file_layout = "port_a";
defparam ram_block1a0.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0121|altsyncram:altsyncram_component0|altsyncram_78g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.operation_mode = "rom";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 13;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "clock0";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 8191;
defparam ram_block1a0.port_a_logical_ram_depth = 65536;
defparam ram_block1a0.port_a_logical_ram_width = 16;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.ram_block_type = "auto";
defparam ram_block1a0.mem_init3 = "1E0F07C3E0F07C1F0F83E0F83E0F83E0F81F07C0F81F07E0FC0F81F81F03F03F03F03F81F81FC0FE07F01FC07E03FC07F01FE03FC03F807F803FC03FE01FF007FC00FF801FF801FFC00FFE003FFC003FFC001FFF0003FFF8000FFFF00003FFFF00000FFFFFE000000FFFFFFFE0000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000001FFFFFFF8000001FFFFF800007FFFE0000FFFF0001FFF8001FFF0007FF8007FF001FFC00FFC00FFC00FF803FE00FF007F807F807F807F00FE01FC07F01FC0FE03F01F80FC0FC07E07E0FC0FC0F81F83F07E0F81F07C1F83E0F83E0F87C1F0783E1F0783C1E0F0F87C3C1E1E0F0F0F0F8787878787";
defparam ram_block1a0.mem_init2 = "8F0F0F0E1E1E3C387870E1E3C7870E1C3871E3C78E1C78E1C70E3C71C38E3871C71C38E38E38E38E38E38E39C71C718E38C71CE38C718E31CE31C639CE31CE718C739CE318C6318C6318C6739CE6319CE6339CC67319CC673398CC6633198CCE67331998CCC666333319999CCCCCC6666666666333333333333326666666666CCCCCD9999B3336666CCC999332664CD99B3264CD993264C993264C99366C99366C9B264D9364D93649B26C93649B24DB26D924DB249B64926DB24926DB6D924924924DB6DB6DA492492492DB6DA4925B6D2496DA496D24B692DA4B692DA4B49692D25A5B4B4B49696969696969694B4B4A5A5AD2D694B5A52D694A5AD6B5A529";
defparam ram_block1a0.mem_init1 = "4A5294A56B5AD4A56B5A95AD4AD4A56A56AD4AD4A95AB52A54A952A54A952AD5AA55AA55AAD52A954AA552A955AA955AAB556AA9552AA9554AAA5554AAA95556AAAA55555AAAAA9555555AAAAAAAA95555555555555555AAAAAAAAAAD5555555555555554AAAAAAAAD555554AAAAAD55552AAA95554AAA9555AAA9556AAB554AA9552AB556AA552AB55AAD56A954AB54AB54A956AD52A54A952B56AD4A95A952B52B52B52B5A95AD4A56B5A94A5295AD6B5A5294A52D6B4A5AD296B4A5A52D2D6969694B4B4B4B4B4969696D2D25A5B49692D25B496D25B692DB492DB4925B6D24925B6DB6D249249249249249B6DB6D924936DB24936C926D924DB26D926C93";
defparam ram_block1a0.mem_init0 = "649B26C9B26C9B26C9B364D9B264C9B366CD9B3664C99B3266CC99B33666CCC9999333266664CCCCCC99999999999999999999999999CCCCCCE666673331999CCC66633199CCE673399CC673398CE6319CC6339CC6318CE739CE739CE318C739C631CE31CE31CE39C738E71C638E31C71C738E38E38E38E38E1C71C70E38E1C70E3C71E3870E3C78F1E3C78F1E1C3C7870F0E1E1E1E3C3C3C3C3C1E1E1E0F0F0787C3E1F0F87C1E0F83C1F07C1F07C1F03E0F81F03E07E0FC0FC0FC0FC0FC07E03F01FC07F01FC07F80FF00FF00FF007FC01FF007FE00FFE007FF001FFE001FFF0003FFF0000FFFF00001FFFFE000001FFFFFFF00000000003FFFFFFFFFFFFFF";

arriav_ram_block ram_block1a16(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a16_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a16.clk0_core_clock_enable = "ena0";
defparam ram_block1a16.clk0_input_clock_enable = "ena0";
defparam ram_block1a16.clk0_output_clock_enable = "ena0";
defparam ram_block1a16.data_interleave_offset_in_bits = 1;
defparam ram_block1a16.data_interleave_width_in_bits = 1;
defparam ram_block1a16.init_file = "DDS_48_v1_nco_ii_0_cos.hex";
defparam ram_block1a16.init_file_layout = "port_a";
defparam ram_block1a16.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0121|altsyncram:altsyncram_component0|altsyncram_78g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a16.operation_mode = "rom";
defparam ram_block1a16.port_a_address_clear = "none";
defparam ram_block1a16.port_a_address_width = 13;
defparam ram_block1a16.port_a_data_out_clear = "none";
defparam ram_block1a16.port_a_data_out_clock = "clock0";
defparam ram_block1a16.port_a_data_width = 1;
defparam ram_block1a16.port_a_first_address = 8192;
defparam ram_block1a16.port_a_first_bit_number = 0;
defparam ram_block1a16.port_a_last_address = 16383;
defparam ram_block1a16.port_a_logical_ram_depth = 65536;
defparam ram_block1a16.port_a_logical_ram_width = 16;
defparam ram_block1a16.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a16.ram_block_type = "auto";
defparam ram_block1a16.mem_init3 = "B56AD5AB56AD52A54A952A54A952A54A952A55AB56AD5AB56AD5AB56A952A54A952A54AB56AD5AB56AD5AA54A952A54AB56AD5AB54A952A54AB56AD5AA54A952AD5AB56A952A55AB56A952A55AB56A952A55AB54A952AD5AA54AB56A952AD5AA54AB56A952AD5AA55AB54AB56A956AD52AD5AA55AA54AB54AB56A956A956A956A956AD52AD52AD52A956A956A956A956A954AB54AB55AA55AAD52AD56A954AB54AA552AD56A954AA55AAD56A954AA552A954AB55AAD56AB552A954AA552A955AAD56AA552AB55AA954AAD56AA556AA552AB552AB552AB552AA556AA556AAD54AA955AAB556AA554AA9552AA554AA9556AAD55AAA554AAB554AAB554AAB554AAB";
defparam ram_block1a16.mem_init2 = "555AAA5552AAD556AAB555AAA9554AAAD556AAA5556AAAD554AAA9555AAAB5554AAA95556AAA95556AAAB5555AAAAD5554AAAAD5555AAAA955556AAAA955554AAAAA555556AAAAAD555552AAAAA9555555AAAAAAA55555552AAAAAAAD55555555AAAAAAAAAB55555555554AAAAAAAAAAAAA955555555555555555556AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAD5555555555555555556AAAAAAAAAAAAB55555555552AAAAAAAA955555556AAAAAAA5555554AAAAAA555555AAAAAB55555AAAAAD55552AAAA55556AAAA55552AAAD5556AAAD5552AAA5556AAA5556AAA5552AAB554AAA5552AAD552AAD55AAA554AA9552AA554AA955AA9";
defparam ram_block1a16.mem_init1 = "552AB552A955AA954AAD56AB55AA956AB55AAD56A954AB54AA55AA55AA55AA55AA54AB54A956AD52A54A956AD5AB56AD5AB56AD4A952B56AD4A95AB52A56A56AD4AD4AD5A95A95A95AD4AD4AD4A56A52B5295AD4AD6B5295AD4A5295AD6A5294A5295AD6B5AD6B5AD694A5294A5AD6B4A52D6B4A52D6B4A5AD296B4A5A52D696B4B5A5AD2D29696B4B4B4A5A5A5A5A5A5A5A5A5A5A5A5A5A5B4B4B4B69696D2D25A5B4B696D2DA5B49692DA5B496D25B496D25B492DA496D24B6D25B6D24B6D2496DB4925B6DA4924B6DB6D2492492DB6DB6DB6DB6DB6DB6DB6DB6DB6D924924936DB6D924936DB64926DB24936D926DB249B649B649B649B649B64DB26D936C";
defparam ram_block1a16.mem_init0 = "9B24D93649B26C9B26C9B26C9B364D9366C9B364C9B364C9B366CD93264C993266CD9B3264CD9B3266CC99B33664CC999332664CCD99933326664CCC99999333336666666CCCCCCCCC9999999999999999999999999999CCCCCCCCC66666673333399998CCCE6663333999CCC66633399CCC6633199CC6633198CE63319CC67319CC67318CE6319CE6318CE739CC6318C6318C6318C6318E739C6318E738C739C639C639C638C738E71CE39C718E39C71CE38E31C71C738E38E38E38E38E38E38E38F1C71C70E38E1C71E38F1C78E3C70E3C70E3C78F1C3870E1C3870E1E3C7870F1E1C3C387870F0F0E1E1E1E1E1E1E1E1E1E1E1F0F0F078783C3E1F0F0783C";

arriav_ram_block ram_block1a65(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a65_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a65.clk0_core_clock_enable = "ena0";
defparam ram_block1a65.clk0_input_clock_enable = "ena0";
defparam ram_block1a65.clk0_output_clock_enable = "ena0";
defparam ram_block1a65.data_interleave_offset_in_bits = 1;
defparam ram_block1a65.data_interleave_width_in_bits = 1;
defparam ram_block1a65.init_file = "DDS_48_v1_nco_ii_0_cos.hex";
defparam ram_block1a65.init_file_layout = "port_a";
defparam ram_block1a65.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0121|altsyncram:altsyncram_component0|altsyncram_78g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a65.operation_mode = "rom";
defparam ram_block1a65.port_a_address_clear = "none";
defparam ram_block1a65.port_a_address_width = 13;
defparam ram_block1a65.port_a_data_out_clear = "none";
defparam ram_block1a65.port_a_data_out_clock = "clock0";
defparam ram_block1a65.port_a_data_width = 1;
defparam ram_block1a65.port_a_first_address = 32768;
defparam ram_block1a65.port_a_first_bit_number = 1;
defparam ram_block1a65.port_a_last_address = 40959;
defparam ram_block1a65.port_a_logical_ram_depth = 65536;
defparam ram_block1a65.port_a_logical_ram_width = 16;
defparam ram_block1a65.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a65.ram_block_type = "auto";
defparam ram_block1a65.mem_init3 = "4AA552A955AAD54AA556AA556AA556AA554AAD55AAB552AA555AAB554AA9556AA9556AAB554AAA5552AAB5552AA95552AAB5556AAA95552AAA95556AAAB55552AAAA55554AAAAB55555AAAAA9555556AAAAAB5555556AAAAAAA555555556AAAAAAAAA555555555555AAAAAAAAAAAAAAAAAA5555555555555555555555555555555555555555556AAAAAAAAAAAAAAAAAD555555555552AAAAAAAAB55555555AAAAAAAD555555AAAAAAD55555AAAAA955556AAAA955552AAAB5555AAAAD5552AAAD555AAAB5556AAA5556AAB555AAAD556AA9554AAB556AA9552AAD55AAB552AA556AAD54AAD54AAD56AA552AB55AAD56AB55AAD56A954AB55AA55AAD52AD52AD5";
defparam ram_block1a65.mem_init2 = "2A55AA54AB54A952AD5AB54A952A54A952A54A952B56AD4A95AB56A56AD4AD5A95A952B52B52B52B52B52B5295A95AD4AD6A56B5295AD4A56B5A94AD6B5A94A5295AD6B5AD6B5AD6B5AD6B5AD6B4A5294B5AD694A5AD694A5AD296B4A5AD296B4A5A52D29694B4A5A5AD2D2969696B4B4B4B4B4A5A5A5A5A5A5A4B4B4B4B4B4969696D2D2DA5A4B4B696D2DA5B4B696D2DA4B696D25B496D25B496D25B492DA4B6D24B6925B6925B6D24B6DA492DB6924B6DB692492DB6DB4924924B6DB6DB6DB6DB6924924936DB6DB6DB6DB6C9249249B6DB6C9249B6DB24936DB24936D924DB64936D926D924DB24DB24DB24D926D936C93649B26D93649B26C9364D9364D";
defparam ram_block1a65.mem_init1 = "9364D9364D9366C9B26CD9366C99364C9B366C99326CD9B366CD9B366CD9B366CC993366CC99B3266CC99B3266CCD99332664CCD99B332666CCC999933326664CCCC99999333332666666CCCCCCCCD9999999999999999333333333319999999999999998CCCCCCCCE6666673333319999CCCCE66673331999CCCE667333998CCE66333998CC6633399CCE673198CC673398CE67319CC67319CC67318CE6319CC6339CC6339CE6318C6739CE739CE6318C639CE739CE738C631CE738C639CE318E718E738C738C738E718E71CE39C638E71CE39C718E39C71CE38E31C71C638E38E39C71C71C71C71C71C71C71C71C71E38E38E3C71C70E38E1C71C38E1C70E3";
defparam ram_block1a65.mem_init0 = "871C38F1C38F1C38F1C3871E3C78F1C3870E1C3878F1E3C3870F1E3C3878F0F1E1E3C3C787870F0F0F1E1E1E1E1E1E1E1E1E1E1E1E1E0F0F0F078787C3C1E1E0F0787C3E1E0F0783C1E0F87C3E0F07C1E0F83C1F07C1F0F83E0F83E0FC1F07C1F83E0FC1F03E0FC1F83F07E07C0FC1F81F83F03F03F03F03F01F81F80FC0FE07F03F81FC07F03F80FE03F80FE01FC07F80FF01FE01FC03FC03FC01FE01FF00FF807FC01FF007FE00FFC01FF801FF801FFC00FFE003FF800FFF000FFF000FFF8003FFE0007FFE0007FFF0000FFFF00007FFFE00007FFFF000007FFFFE000001FFFFFFC0000000FFFFFFFFE00000000001FFFFFFFFFFFFFFFFFC00000000000000";

arriav_ram_block ram_block1a81(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a81_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a81.clk0_core_clock_enable = "ena0";
defparam ram_block1a81.clk0_input_clock_enable = "ena0";
defparam ram_block1a81.clk0_output_clock_enable = "ena0";
defparam ram_block1a81.data_interleave_offset_in_bits = 1;
defparam ram_block1a81.data_interleave_width_in_bits = 1;
defparam ram_block1a81.init_file = "DDS_48_v1_nco_ii_0_cos.hex";
defparam ram_block1a81.init_file_layout = "port_a";
defparam ram_block1a81.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0121|altsyncram:altsyncram_component0|altsyncram_78g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a81.operation_mode = "rom";
defparam ram_block1a81.port_a_address_clear = "none";
defparam ram_block1a81.port_a_address_width = 13;
defparam ram_block1a81.port_a_data_out_clear = "none";
defparam ram_block1a81.port_a_data_out_clock = "clock0";
defparam ram_block1a81.port_a_data_width = 1;
defparam ram_block1a81.port_a_first_address = 40960;
defparam ram_block1a81.port_a_first_bit_number = 1;
defparam ram_block1a81.port_a_last_address = 49151;
defparam ram_block1a81.port_a_logical_ram_depth = 65536;
defparam ram_block1a81.port_a_logical_ram_width = 16;
defparam ram_block1a81.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a81.ram_block_type = "auto";
defparam ram_block1a81.mem_init3 = "7319CC67319CCE63398CE63398CE63398CE63398CE63398CE63398CE67319CC67319CC67319CC67319CC663398CE63398CE63398CC67319CC67319CC663398CE63398CE67319CC673198CE63398CE67319CC673398CE63399CC673198CE63399CC673198CE63399CC673398CE67319CCE63399CC663398CC673198CE673198CE67319CCE63319CCE673198CE673198CE673398CC673399CC663319CCE673398CC663319CCE673399CC6633198CC6633198CC673399CCE6733198CC6633198CC6633199CCE6733998CC6633199CCE6633198CCE6733198CCE6633199CCE66333998CC66733199CCC66733199CCC66733199CCC666333998CCC667333998CCC667";
defparam ram_block1a81.mem_init2 = "333999CCCE663331998CCC6667333999CCCE6663331999CCCC66673339998CCCC666733319998CCCE666733339999CCCCC66663333399998CCCCE666673333399999CCCCCE666663333331999998CCCCCC6666666333333319999999CCCCCCCCC66666666673333333333399999999999998CCCCCCCCCCCCCCCCCCCE6666666666666666666666666666666666666666666666666664CCCCCCCCCCCCCCCCCCD999999999999933333333336666666664CCCCCCCD99999993333332666666CCCCCC99999933333666664CCCC99999333326666CCCC9999B33326664CCC99993332666CCCD9993336666CCD9993336664CC999B33666CCD99B33666CCD99B33664";
defparam ram_block1a81.mem_init1 = "CC99933664CC99B32664CD9933664CD9933664CD9B3266CD993366CC993366CC993266CD9B3264C993264CD9B366CD9B366CD9B264C993264D9B366C99326CD9B264D9B364C9B364C9B264D9B26CD9366C9B364D9B26C9B364D9364C9B26C9B26C9B364D9364D9364DB26C9B26C9B26D9364D926C9B26D93649B26D936C9B24D926C93649B64DB26D926D936C936C936C936C936C936C936C926D926DB24DB64936C926DB249B6C924DB64936DB24936DB24936DB64924DB6D924936DB6D924924DB6DB6C924924926DB6DB6DB6DB64924924924924924924924924924B6DB6DB6DB6DB492492492DB6DB6924924B6DB692492DB6D2492DB6D2492DB6924B6DA";
defparam ram_block1a81.mem_init0 = "496DB492DB6925B6925B6925B692DB492DA496D25B692DA496D25B496D25B496D25B49692DA4B696D25A4B696D2DA5B4B696D2DA5B4B49696D2D25A5B4B4B69696D2D2D2DA5A5A5A5A4B4B4B4B4B4B4B4B4B4B4B4B4B4B5A5A5A5A52D2D2D2969694B4B5A5A52D29696B4B5A52D29694B5A52D694B4A52D694B5A5296B4A52D6B4A52D6B5A5294B5AD6B5A5294A5294A5294A5294A5294A5294AD6B5AD6A5294AD6B5294AD6A5295AD4A56B52B5A94AD4A56A56B52B5295A95A95A95A95A95A95A95AB52B52A56A54AD4A95AB52A56AD5A952A56AD5AB56AD5AB56AD5AB56AD52A54AB56A952AD5AA55AB54AB54AB54AB54AB54AB55AA552AD56A954AA552A95";

arriav_ram_block ram_block1a97(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a97_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a97.clk0_core_clock_enable = "ena0";
defparam ram_block1a97.clk0_input_clock_enable = "ena0";
defparam ram_block1a97.clk0_output_clock_enable = "ena0";
defparam ram_block1a97.data_interleave_offset_in_bits = 1;
defparam ram_block1a97.data_interleave_width_in_bits = 1;
defparam ram_block1a97.init_file = "DDS_48_v1_nco_ii_0_cos.hex";
defparam ram_block1a97.init_file_layout = "port_a";
defparam ram_block1a97.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0121|altsyncram:altsyncram_component0|altsyncram_78g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a97.operation_mode = "rom";
defparam ram_block1a97.port_a_address_clear = "none";
defparam ram_block1a97.port_a_address_width = 13;
defparam ram_block1a97.port_a_data_out_clear = "none";
defparam ram_block1a97.port_a_data_out_clock = "clock0";
defparam ram_block1a97.port_a_data_width = 1;
defparam ram_block1a97.port_a_first_address = 49152;
defparam ram_block1a97.port_a_first_bit_number = 1;
defparam ram_block1a97.port_a_last_address = 57343;
defparam ram_block1a97.port_a_logical_ram_depth = 65536;
defparam ram_block1a97.port_a_logical_ram_width = 16;
defparam ram_block1a97.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a97.ram_block_type = "auto";
defparam ram_block1a97.mem_init3 = "2A954AB55AAD56A954AB54AA55AA55AA55AA55AA55AA54AB54A956AD52A54AB56AD5AA54A952A54A952B56AD5AB52A54AD5A952B56A54AD5A95AB52B52B56A56A56A56A56A56A56A56B52B52B5A95AD4AD6A56B5295AD4A56B5295AD6A5295AD6B5294A56B5AD6B5A94A5294A5294A5294A52D6B5AD6B5A5294A5AD6B4A52D6B4A52D6B4A5AD694B5A52D694B5A52D296B4A5A52D29694B4A5A5AD2D69696B4B4B5A5A5A52D2D2D2D29696969696969696969696969696D2D2D2D2DA5A5A5B4B4B4969692D2DA5A4B4B696D2D25A4B49692D25B4B696D25A4B692D25B496D25A4B692DA4B6D25B496D24B692DB496DA4B6D24B6925B6925B6925B6924B6D2496";
defparam ram_block1a97.mem_init2 = "DB4925B6D2496DB692496DB692496DB6DA4924B6DB6DA4924924B6DB6DB6DB4924924924924924924924924924924924924924924DB6DB6DB6D924924936DB6DB24924DB6DB24924DB6D924936DB24936DB24936D9249B6C926DB249B6C926DB24DB649B6C936C926D926D926D926D926D926D926D936C93649B64DB26D936C9B64DB26D93649B26D9364DB26C9B24D9364D926C9B26C9B26C9B26C9B26C9B26C9B264D9364D9326C9B364D9326C9B364D9B26CD9326CD9366C99366CD9326CD9B264D9B366C993264C9B366CD9B366CD9B366CD9B366CD9B3264C993366CD993266CD993266CD993366CC99B3266CC99B3666CC99B3266CC99933664CC99B33";
defparam ram_block1a97.mem_init1 = "666CC999332664CC999332666CCD99B332664CCD9993336664CCD999B3326664CCD999B33326664CCCD999B333266664CCCD9999B3333266666CCCCC999999333332666666CCCCCCD9999999B33333336666666664CCCCCCCCCC9999999999999B33333333333333333326666666666666666666666666666666666666666666666666663333333333333333333319999999999999CCCCCCCCCCC666666666733333333199999998CCCCCCC66666673333331999998CCCCCE6666633333399999CCCCCE66663333319998CCCCE6666333319998CCCC666633331999CCCCE66633339998CCCE6663331999CCCC6663331999CCCE667333999CCCE667333998CCC";
defparam ram_block1a97.mem_init0 = "666333999CCC666333999CCC66733199CCCE66333998CCE6633399CCC66733199CCE6633399CCC66733998CC66733998CC6633399CCE6633198CC6673399CCE6733198CC6633198CC6633198CC6633198CC663319CCE673399CCE633198CC663399CCE633198CE673398CC663399CCE63319CCE63319CCE673198CE67319CCE63319CCE63319CC663399CC673398CE67319CCE63399CC673398CE67319CC663398CE67319CC663398CE67319CC673398CE63398CC67319CC673398CE63398CE67319CC67319CC663398CE63398CE63399CC67319CC67319CC67319CC663398CE63398CE63398CE63398CE63398CC67319CC67319CC67319CC67319CC67319CC6";

arriav_ram_block ram_block1a113(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a113_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a113.clk0_core_clock_enable = "ena0";
defparam ram_block1a113.clk0_input_clock_enable = "ena0";
defparam ram_block1a113.clk0_output_clock_enable = "ena0";
defparam ram_block1a113.data_interleave_offset_in_bits = 1;
defparam ram_block1a113.data_interleave_width_in_bits = 1;
defparam ram_block1a113.init_file = "DDS_48_v1_nco_ii_0_cos.hex";
defparam ram_block1a113.init_file_layout = "port_a";
defparam ram_block1a113.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0121|altsyncram:altsyncram_component0|altsyncram_78g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a113.operation_mode = "rom";
defparam ram_block1a113.port_a_address_clear = "none";
defparam ram_block1a113.port_a_address_width = 13;
defparam ram_block1a113.port_a_data_out_clear = "none";
defparam ram_block1a113.port_a_data_out_clock = "clock0";
defparam ram_block1a113.port_a_data_width = 1;
defparam ram_block1a113.port_a_first_address = 57344;
defparam ram_block1a113.port_a_first_bit_number = 1;
defparam ram_block1a113.port_a_last_address = 65535;
defparam ram_block1a113.port_a_logical_ram_depth = 65536;
defparam ram_block1a113.port_a_logical_ram_width = 16;
defparam ram_block1a113.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a113.ram_block_type = "auto";
defparam ram_block1a113.mem_init3 = "FFFFFFFFFFFFFFFFFFFFFFFFE0000000000000FFFFFFFFFE00000001FFFFFFE000000FFFFFE00000FFFFF00001FFFF80001FFFE0001FFFC0007FFE0007FFE000FFF8007FF8007FF800FFF001FFC00FFE007FE007FE007FC00FF803FE00FF803FE01FF00FF007F807F807F00FF00FE01FC07F80FE03F80FE03F80FE03F01F80FE07F03F01F81F80FC0FC0FC0FC0FC1F81F81F03F07E0FC1F83F07E0F81F07E0F83E07C1F07C1F07C1F07C1F0783E0F87C1F0F83C1E0F87C3E1F0F87C3E1F0F0787C3C1E1E0F0F0F878787C3C3C3C3C3C3C3C3C3C3C3C3C38787878F0F0E1E1C3C3878F0E1E3C3870F1E3C3870E1C3870E1C3870E3C78E1C38F1C38F1C38F1C38E";
defparam ram_block1a113.mem_init2 = "1C70E38F1C78E38F1C71E38E38E1C71C71C71C38E38E38E38E38E71C71C71C718E38E39C71C638E31C718E39C718E31C638C718E71CE31C639C639C639CE31CE718E738C631CE738C6318E739CE739CE739CE739CC6318C6739CC6319CE6319CE6339CC67319CE63398CE67319CC663399CC6633198CC6633198CCE6633199CCC666333199CCCC66633339999CCCCE66667333339999998CCCCCCCC66666666666666667333333333266666666666666664CCCCCCCD999999B3333266666CCCC9999B3336666CCC999B332664CC999332664CD99B3266CC99B3264CD993266CD9B3264C993264C99326CD9B364C9B366C99364C9B264D9366C9B26C99364D936";
defparam ram_block1a113.mem_init1 = "4D926C9B26C9B64D926C9B64DB26D936C93649B649B649B649B6C936D926DB249B6C924DB6C924DB6C9249B6DB64924926DB6DB6DB24924924924924924924924925B6DB6DB6D2492496DB6D24925B6D2492DB6924B6D2496DA496DA496D24B6925B496DA4B692DA4B692DA5B496D2DA5B49692D25A4B4B69692D2DA5A5B4B4B49696969696D2D2D2D2D2D2D29696969696B4B4B5A5A5AD2D29694B4A5A52D694B4A5AD296B4A52D694A5AD694A52D6B5A5294A5296B5AD6B5AD6B5AD4A5294A56B5AD4A5295AD4A52B5A94AD4A56B52B5A95A95AD4AD4AD4AD4AD4AD4AD5A95A952B52A56AD4A95AB56A54A952A56AD5AB56A952A54A956AD52A55AB54AB54A";
defparam ram_block1a113.mem_init0 = "956A956A954AB54AB55AA552A954AB55AAD56AA552A955AA954AAD54AAD55AA955AAB556AAD55AAB554AAB556AA9554AAB555AAAD554AAA5556AAA5554AAA95556AAA95556AAAB55552AAAB55554AAAAB55555AAAAA9555556AAAAAA5555555AAAAAAAB555555556AAAAAAAAAA55555555555555AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA55555555555555AAAAAAAAAAB555555554AAAAAAA95555554AAAAAAD555552AAAAA555552AAAA955556AAAAD5554AAAA55552AAA95556AAAD555AAAB5552AAA5552AAB555AAAD556AA9554AAB554AAB556AA9552AA554AA9552AB556AA556AA556AA556AB552AB55AAD54AA55";

arriav_ram_block ram_block1a33(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a33_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a33.clk0_core_clock_enable = "ena0";
defparam ram_block1a33.clk0_input_clock_enable = "ena0";
defparam ram_block1a33.clk0_output_clock_enable = "ena0";
defparam ram_block1a33.data_interleave_offset_in_bits = 1;
defparam ram_block1a33.data_interleave_width_in_bits = 1;
defparam ram_block1a33.init_file = "DDS_48_v1_nco_ii_0_cos.hex";
defparam ram_block1a33.init_file_layout = "port_a";
defparam ram_block1a33.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0121|altsyncram:altsyncram_component0|altsyncram_78g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a33.operation_mode = "rom";
defparam ram_block1a33.port_a_address_clear = "none";
defparam ram_block1a33.port_a_address_width = 13;
defparam ram_block1a33.port_a_data_out_clear = "none";
defparam ram_block1a33.port_a_data_out_clock = "clock0";
defparam ram_block1a33.port_a_data_width = 1;
defparam ram_block1a33.port_a_first_address = 16384;
defparam ram_block1a33.port_a_first_bit_number = 1;
defparam ram_block1a33.port_a_last_address = 24575;
defparam ram_block1a33.port_a_logical_ram_depth = 65536;
defparam ram_block1a33.port_a_logical_ram_width = 16;
defparam ram_block1a33.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a33.ram_block_type = "auto";
defparam ram_block1a33.mem_init3 = "52A954AA552AD56A954AB55AA55AA55AA55AA55AA55AB54AB56A952AD5AA54A956AD5AB56AD5AB56AD5AB56AD4A952B56AD4A95AB52A56A54AD4A95A95AB52B52B52B52B52B52B52B5295A95AD4AD4A56A52B5A95AD4A56B5294AD6A5295AD6A5294AD6B5AD6A5294A5294A5294A5294A5294A5294B5AD6B5A5294B5AD694A5AD694A5AD294B5A52D694A5A52D694B5A52D29694B5A5AD2D29694B4B5A5A52D2D296969694B4B4B4B5A5A5A5A5A5A5A5A5A5A5A5A5A5A4B4B4B4B4B6969696D2D2DA5A5B4B49696D2D25A5B4B696D2DA5B4B696D2DA4B496D2DA4B692D25B496D25B496D25B496D24B692DB496D24B6925B692DB492DB492DB492DB6925B6D24";
defparam ram_block1a33.mem_init2 = "B6DA492DB692496DB692496DB692492DB6DA492492DB6DB6924924925B6DB6DB6DB6DA4924924924924924924924924924DB6DB6DB6DB6C924924926DB6DB64924936DB6D924936DB64924DB6D9249B6D9249B6D924DB64926DB249B6C926D924DB649B6C936C926D926D926D926D926D926D926D936C936C9B64DB24D926C93649B26D936C9B24D936C9B26C9364D936C9B26C9B26C9B64D9364D9364D9B26C9B26C9B264D9364D9B26C9B364D9B26CD9366C9B364C9B264D9B264D9B364C9B366C99326CD9B364C993264C9B366CD9B366CD9B3664C993264C99B366CC993266CD993266CD993366CC99B3664CD9933664CD9933664CC99B32664CD9933266";
defparam ram_block1a33.mem_init1 = "4CD99B33666CCD99B33666CCD99B332664CCD999333666CCCD9993336666CCC999933326664CCC9999B33326666CCCC999993333266664CCCCD99999333332666666CCCCCC99999993333333666666664CCCCCCCCD9999999999333333333333366666666666666666664CCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCE66666666666666666663333333333333399999999999CCCCCCCCCC666666667333333319999998CCCCCCC6666663333331999998CCCCCE666673333399999CCCCCE66663333399998CCCC6666733339999CCCCE66633331999CCCC66663333999CCCC66673331998CCCE667333999CCCC6663331998CCE667333999";
defparam ram_block1a33.mem_init0 = "CCC666333999CCC666333998CCC66733199CCC66733199CCC66733199CCC66333998CCE6733198CCE6633199CCE6633198CCE6733198CC6633399CCE6733198CC6633198CC6633199CCE673399CC6633198CC6633198CC673399CCE673198CC663399CCE673198CC673399CC663399CCE63319CCE63319CCE673198CE67319CCE63319CCE63319CC663398CC673398CE67319CCE63399CC673398CE63319CC673398CE63319CC673398CE63399CC67319CCE63398CE63319CC67319CCE63398CE63398CC67319CC67319CC663398CE63398CE63398CC67319CC67319CC67319CC67319CCE63398CE63398CE63398CE63398CE63398CE63398CE67319CC67319C";

arriav_ram_block ram_block1a49(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a49_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a49.clk0_core_clock_enable = "ena0";
defparam ram_block1a49.clk0_input_clock_enable = "ena0";
defparam ram_block1a49.clk0_output_clock_enable = "ena0";
defparam ram_block1a49.data_interleave_offset_in_bits = 1;
defparam ram_block1a49.data_interleave_width_in_bits = 1;
defparam ram_block1a49.init_file = "DDS_48_v1_nco_ii_0_cos.hex";
defparam ram_block1a49.init_file_layout = "port_a";
defparam ram_block1a49.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0121|altsyncram:altsyncram_component0|altsyncram_78g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a49.operation_mode = "rom";
defparam ram_block1a49.port_a_address_clear = "none";
defparam ram_block1a49.port_a_address_width = 13;
defparam ram_block1a49.port_a_data_out_clear = "none";
defparam ram_block1a49.port_a_data_out_clock = "clock0";
defparam ram_block1a49.port_a_data_width = 1;
defparam ram_block1a49.port_a_first_address = 24576;
defparam ram_block1a49.port_a_first_bit_number = 1;
defparam ram_block1a49.port_a_last_address = 32767;
defparam ram_block1a49.port_a_logical_ram_depth = 65536;
defparam ram_block1a49.port_a_logical_ram_width = 16;
defparam ram_block1a49.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a49.ram_block_type = "auto";
defparam ram_block1a49.mem_init3 = "000000000000007FFFFFFFFFFFFFFFFF00000000000FFFFFFFFE00000007FFFFFF000000FFFFFC00001FFFFC0000FFFFC0001FFFE0001FFFC000FFFC000FFF8003FFE001FFE001FFE003FF800FFE007FF003FF003FF007FE00FFC01FF007FC03FE01FF00FF007F807F807F00FF01FE03FC07F00FE03F80FE03F81FC07F03F81FC0FE07E03F03F01F81F81F81F81F83F03F07E07C0FC1F83F07E0F81F07E0F83F07C1F07E0F83E0F83E1F07C1F0783E0F07C1E0F87C3E0F0783C1E0F0F87C3C1E0F0F0787C3C3C1E1E1E0F0F0F0F0F0F0F0F0F0F0F0F0F1E1E1E1C3C3C7878F0F1E1E3C3878F1E1C3878F1E3C3870E1C3871E3C78F1C3871E3871E3871E3871C3";
defparam ram_block1a49.mem_init2 = "8E1C70E3871C70E38E1C71C78E38E38F1C71C71C71C71C71C71C71C71C738E38E38C71C718E38E71C738E31C738E71CE38C738E71CE31CE39C639C639CE31CE318E738C639CE718C639CE739CE738C6318CE739CE739CC6318CE7398C67398C67318CE6319CC67319CC67319CCE63399CC663319CCE6733998CC66333998CCE66333999CCCE6673331999CCCCE66673333199999CCCCCCE666666663333333333333333199999999993333333333333333666666666CCCCCC9999993333266664CCC99993332666CCC999B336664CC99933666CC99B3266CC99B3266CD993266CD9B366CD9B366CD9B366C99326CD9B264D9326CD9366C9B26CD9364D9364D93";
defparam ram_block1a49.mem_init1 = "64D9364D926C9B24D936C9B24D926D936C93649B649B649B64936C936D924DB64936D9249B6D9249B6DB24926DB6DB24924926DB6DB6DB6DB6D92492492DB6DB6DB6DB6DA4924925B6DB692492DB6DA492DB6924B6DA496DB492DB492DA496DA4B6925B496D25B496D25B496D2DA4B696D2DA5B4B696D2DA5A4B4B69696D2D2D25A5A5A5A5A4B4B4B4B4B4B4A5A5A5A5A5AD2D2D29696B4B4A5A52D29694B4A5AD296B4A5AD296B4A52D6B4A52D6B5A5294A5AD6B5AD6B5AD6B5AD6B5AD6B5294A52B5AD6A52B5AD4A56B5295AD4AD6A56B52B5295A95A95A95A95A95A952B52B56A56AD4AD5AB52A56AD5A952A54A952A54A952A55AB56A952A55AA54AB54A9";
defparam ram_block1a49.mem_init0 = "56A956A956AB54AB55AA552AD56AB55AAD56AB55AA954AAD56AA556AA556AAD54AA955AAB556AA9552AAD55AAA5552AAD556AAB555AAAD554AAAD555AAAB5556AAA95556AAAB5555AAAA955552AAAAD55552AAAAB555556AAAAAB5555556AAAAAAB55555555AAAAAAAAA9555555555556AAAAAAAAAAAAAAAAAD555555555555555555555555555555555555555554AAAAAAAAAAAAAAAAAB555555555554AAAAAAAAAD55555554AAAAAAAD555555AAAAAAD555552AAAAB55555AAAAA55554AAAA95555AAAAD5552AAA95552AAAD555AAA95552AA9555AAA9554AAA555AAAD552AAD552AA555AAB554AA955AAB556AA554AAD54AAD54AAD54AA556AB552A954AA5";

arriav_ram_block ram_block1a1(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a1_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.clk0_input_clock_enable = "ena0";
defparam ram_block1a1.clk0_output_clock_enable = "ena0";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.init_file = "DDS_48_v1_nco_ii_0_cos.hex";
defparam ram_block1a1.init_file_layout = "port_a";
defparam ram_block1a1.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0121|altsyncram:altsyncram_component0|altsyncram_78g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.operation_mode = "rom";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 13;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "clock0";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 8191;
defparam ram_block1a1.port_a_logical_ram_depth = 65536;
defparam ram_block1a1.port_a_logical_ram_width = 16;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.ram_block_type = "auto";
defparam ram_block1a1.mem_init3 = "54AA556AB55AA955AAD54AAD54AAD54AAD55AA9552AA554AA9552AAD55AAA555AAA5552AAD556AAB555AAA9554AAA9555AAAB5556AAAD5552AAA95554AAAA55556AAAAD55552AAAA955554AAAAA9555556AAAAAA55555552AAAAAAA555555555AAAAAAAAAAB55555555555554AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAB55555555555554AAAAAAAAAAD55555555AAAAAAAB5555554AAAAAAD555552AAAAB55555AAAAA55555AAAA95555AAAAD5552AAAD5552AAA5554AAAD554AAA5556AAB555AAA5552AAD55AAA555AAB556AAD55AAB552AB556AA556AA552AB552A954AAD56AB55AA552A954AB55AA55AA552AD52AD52";
defparam ram_block1a1.mem_init2 = "A55AA55AB54A956AD52A54A952AD5AB56AD4A952A54AD5AB52A56AD4A95A952B52B56A56A56A56A56A56A56B52B52B5A95AD4A56A52B5A94A56B5294A56B5AD4A5294A56B5AD6B5AD6B5AD294A5294B5AD694A52D6B4A52D694A5AD296B4A5A52D694B4A5A52D29696B4B4B5A5A5AD2D2D2D2D296969696969696D2D2D2D2D25A5A5B4B4B69692D2DA5A4B49692D25B4B696D25B4B692DA4B692DA4B6D25B492DA496D24B6D24B6D2496DA492DB692496DB492496DB6D2492496DB6DB6DB49249249249249249249249249B6DB6DB6C924924DB6DB24926DB64926DB64926DB249B6C936D926DB24DB24DB24DB24D926D936C9B64DB26C9364DB26C9B26C9364";
defparam ram_block1a1.mem_init1 = "D9364D9326C9B26CD9364C9B264D9326CD9B264D9B366C993264C993264C99B366CC9933664C99B3266CC99B33664CC999332664CC999B332666CCCD999B33326666CCCCC99999B333333666666664CCCCCCCCCCCCCCCC9999999999CCCCCCCCCCCCCCCCC66666666333333399999CCCCCE666733339998CCC6667331998CCC66733198CCE6633198CC6633198CC673398CC67319CCE63398CE7319CC67398CE7318CE7318C6739CC6318C6739CE739CE739CE739CE318C639CE718C639CE31CE718E738C738C738C718E71CE31C638C718E31C738E31C718E38C71C738E38E31C71C71C71CE38E38E38E38E3871C71C71C70E38E38F1C71E38E3C71E38E1C70";
defparam ram_block1a1.mem_init0 = "E3871E3871E3871E3870E3C78E1C3870E1C3870E1C3878F1E1C3878F0E1E3C387870F0E1E1E3C3C3C387878787878787878787878787C3C3C3E1E1E0F0F0787C3C1E1F0F87C3E1F0F87C3E0F0783E1F07C3E0F83C1F07C1F07C1F07C1F07C0F83E0FC1F03E0FC1F83F07E0FC1F81F03F03F07E07E07E07E07E03F03F01F81FC0FE03F01F80FE03F80FE03F80FE03FC07F00FE01FE01FC03FC03FC01FE01FF00FF803FE00FF803FE007FC00FFC00FFC00FFE007FF001FFE003FFC003FFC003FFE000FFFC000FFFC0007FFF0000FFFF00003FFFF00001FFFFE00000FFFFFE000000FFFFFFF00000000FFFFFFFFFE0000000000000FFFFFFFFFFFFFFFFFFFFFFFFF";

arriav_ram_block ram_block1a17(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a17_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a17.clk0_core_clock_enable = "ena0";
defparam ram_block1a17.clk0_input_clock_enable = "ena0";
defparam ram_block1a17.clk0_output_clock_enable = "ena0";
defparam ram_block1a17.data_interleave_offset_in_bits = 1;
defparam ram_block1a17.data_interleave_width_in_bits = 1;
defparam ram_block1a17.init_file = "DDS_48_v1_nco_ii_0_cos.hex";
defparam ram_block1a17.init_file_layout = "port_a";
defparam ram_block1a17.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0121|altsyncram:altsyncram_component0|altsyncram_78g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a17.operation_mode = "rom";
defparam ram_block1a17.port_a_address_clear = "none";
defparam ram_block1a17.port_a_address_width = 13;
defparam ram_block1a17.port_a_data_out_clear = "none";
defparam ram_block1a17.port_a_data_out_clock = "clock0";
defparam ram_block1a17.port_a_data_width = 1;
defparam ram_block1a17.port_a_first_address = 8192;
defparam ram_block1a17.port_a_first_bit_number = 1;
defparam ram_block1a17.port_a_last_address = 16383;
defparam ram_block1a17.port_a_logical_ram_depth = 65536;
defparam ram_block1a17.port_a_logical_ram_width = 16;
defparam ram_block1a17.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a17.ram_block_type = "auto";
defparam ram_block1a17.mem_init3 = "C67319CC67319CC67319CC67319CC67319CC663398CE63398CE63398CE63398CE63398CC67319CC67319CC67319CC673398CE63398CE63398CC67319CC67319CCE63398CE63399CC67319CC663398CE63399CC67319CCE63398CC67319CCE63398CC67319CCE63399CC673398CE67319CCE63399CC673398CC673198CE673198CE67319CCE63319CCE673198CE673198CE673398CC663399CCE633198CE673398CC6633198CE673399CCE673198CC6633198CC6633198CC6633198CC6633199CCE673399CCC6633198CCE6733998CC6633399CCC6633399CCC66733998CCE6733199CCC66733998CCE66333998CCE66733199CCC667333998CCC667333998CCC";
defparam ram_block1a17.mem_init2 = "666333999CCCE667333999CCCE6673331998CCC66673331998CCCE66633339998CCCE666733319998CCCC6666333319998CCCCE66663333199998CCCCE6666733333999998CCCCCE666663333331999999CCCCCCC666666633333333199999999CCCCCCCCCC666666666673333333333333199999999999999999998CCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCC9999999999999999999B333333333333266666666664CCCCCCCCD9999999B33333336666666CCCCCC99999933333266666CCCCC99999B333366664CCCC9999B33366664CCC9999B3336664CCC999B3336664CCD9993336664CC999B33666CCC999332664CC99933266CCD";
defparam ram_block1a17.mem_init1 = "99B32664CD9933266CC99B3266CCD9B3266CC99B3266CD993366CC993366CC993366CD993264C99B366CD9B366CD9B366CD9B366CD9B264C99326CD9B364C9B366C99366CD9326CD9366C99366C9B364D9B26C99364D9B26C99364D9364C9B26C9B26C9B26C9B26C9B26C9B26C9364D93649B26C9B64D936C9B24D936C9B64DB26D936C9B64DB24D926D936C936C936C936C936C936C936C926D926DB24DB649B6C926DB249B6C926DB24936D9249B6D9249B6D924936DB649249B6DB649249B6DB6D924924936DB6DB6DB64924924924924924924924924924924924924924925B6DB6DB6DA4924924B6DB6DA4924B6DB6D2492DB6D2492DB6D2496DB4925B6";
defparam ram_block1a17.mem_init0 = "D2496DA492DB492DB492DB492DA496DA4B6D25B692DA496D25B496DA4B692DA4B496D25B49692DA4B496D2DA5B49692D25A4B49696D2DA5A4B4B69692D2D25A5A5B4B4B4B696969696D2D2D2D2D2D2D2D2D2D2D2D2D2D29696969694B4B4B5A5A5AD2D2D696B4B4A5A52D29694B4A5AD29694B5A52D694B5A52D6B4A5AD694A5AD694A5AD6B4A5294B5AD6B5AD694A5294A5294A5294A52B5AD6B5AD4A5295AD6B5294AD6B5295AD4A56B5295AD4AD6A56B52B5A95A95AD4AD4AD4AD4AD4AD4AD4AD5A95A95AB52B56A54AD5A952B56A54A95AB56AD5A952A54A952A54AB56AD5AA54A956AD52A55AA54AB54AB54AB54AB54AB54AA55AA552AD56AB55AA552A9";

arriav_ram_block ram_block1a66(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a66_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a66.clk0_core_clock_enable = "ena0";
defparam ram_block1a66.clk0_input_clock_enable = "ena0";
defparam ram_block1a66.clk0_output_clock_enable = "ena0";
defparam ram_block1a66.data_interleave_offset_in_bits = 1;
defparam ram_block1a66.data_interleave_width_in_bits = 1;
defparam ram_block1a66.init_file = "DDS_48_v1_nco_ii_0_cos.hex";
defparam ram_block1a66.init_file_layout = "port_a";
defparam ram_block1a66.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0121|altsyncram:altsyncram_component0|altsyncram_78g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a66.operation_mode = "rom";
defparam ram_block1a66.port_a_address_clear = "none";
defparam ram_block1a66.port_a_address_width = 13;
defparam ram_block1a66.port_a_data_out_clear = "none";
defparam ram_block1a66.port_a_data_out_clock = "clock0";
defparam ram_block1a66.port_a_data_width = 1;
defparam ram_block1a66.port_a_first_address = 32768;
defparam ram_block1a66.port_a_first_bit_number = 2;
defparam ram_block1a66.port_a_last_address = 40959;
defparam ram_block1a66.port_a_logical_ram_depth = 65536;
defparam ram_block1a66.port_a_logical_ram_width = 16;
defparam ram_block1a66.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a66.ram_block_type = "auto";
defparam ram_block1a66.mem_init3 = "933664CD9933666CC99B33664CC99B33666CC999332664CC999332666CCD99B332664CCD9993336664CCD999B3326664CCD999B33326664CCCD999B333266664CCCC999993333266666CCCCCD99999B3333326666664CCCCCCC99999999B333333333666666666666CCCCCCCCCCCCCCCCCC9999999999999999999999999999999999999999998CCCCCCCCCCCCCCCCCE66666666666333333333399999999CCCCCCCE666666333333199999CCCCCE66667333319999CCCCC666633331999CCCCE66633339998CCC6667333999CCCE667331998CCC66733199CCCE6633399CCC66733198CCE6733198CC6633399CCE673399CCE673198CC663399CCE63319CCE6";
defparam ram_block1a66.mem_init2 = "3399CC673398CE63319CC67319CC67319CC67319CC67318CE63398C67318CE6319CE6339CC6339CC6339CC6319CE6318CE7398C6319CE7398C6318CE739CE739CE6318C6318C6318C6318C6318C739CE739CE718C6318E739CE318C739CE318C739C631CE718C739C631CE318E718C738C738C739C639C639C638C738C738C718E718E31CE39C738C718E31C638C718E31C738E71C638E71C638E71C638E31C738E38C71C638E39C71C738E38E31C71C738E38E38E31C71C71C71C738E38E38E38E38E38E38E38E38E38E38E38F1C71C71C71C70E38E38E3C71C71C38E38E1C71C78E38E1C71E38E3C71C38E3C71E38E1C70E3871C38E1C78E3C70E3871E3871";
defparam ram_block1a66.mem_init1 = "E3871E3871E3870E3C70E1C78F1E3870E3C78F1E3C70E1C3870E1C3870E1C3870F1E3C78F0E1C3C78F0E1C3C78F0E1E3C3878F0E1E3C3C7870F0E1E1C3C387870F0F1E1E1C3C3C38787870F0F0F0F1E1E1E1E1E1E1E1E1C3C3C3C3C3E1E1E1E1E1E1E1E1F0F0F0F0F07878783C3C3E1E1E0F0F078783C3E1E1F0F0787C3C1E0F0F87C3C1E0F0783C3E1F0F87C1E0F0783C1F0F87C1E0F87C1E0F87C1F0F83E1F07C3E0F83C1F07C1F0783E0F83E0F83E0F83E0F83E0F83F07C1F07C0F83E0FC1F07E0F83F07C0F83F07E0F81F03E07C0F81F03E07E0FC1F81F03F03E07E07C0FC0FC1F81F81F81F81F81F81F81F81F81FC0FC0FC07E07F03F01F81FC0FE07F03";
defparam ram_block1a66.mem_init0 = "F81FC0FE03F01FC0FE03F81FC07F01FC07F01FC07F01FC03F80FE03FC07F00FE01FC03F807F80FF00FE01FE01FE01FE01FE01FE01FE00FF00FF807F803FE01FF007F803FE00FF803FE00FF803FF007FE00FFC01FF801FF003FF003FF001FF801FFC00FFE003FF001FFC007FF800FFE001FFC003FFC003FFC001FFE000FFF0007FFC001FFF8003FFF0003FFF0001FFF8000FFFE0001FFFC0003FFFE0001FFFF00007FFFE00007FFFF00001FFFFE00001FFFFF000003FFFFF000000FFFFFF0000003FFFFFF80000007FFFFFFF000000007FFFFFFFF80000000007FFFFFFFFFFE00000000000000FFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000";

arriav_ram_block ram_block1a82(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a82_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a82.clk0_core_clock_enable = "ena0";
defparam ram_block1a82.clk0_input_clock_enable = "ena0";
defparam ram_block1a82.clk0_output_clock_enable = "ena0";
defparam ram_block1a82.data_interleave_offset_in_bits = 1;
defparam ram_block1a82.data_interleave_width_in_bits = 1;
defparam ram_block1a82.init_file = "DDS_48_v1_nco_ii_0_cos.hex";
defparam ram_block1a82.init_file_layout = "port_a";
defparam ram_block1a82.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0121|altsyncram:altsyncram_component0|altsyncram_78g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a82.operation_mode = "rom";
defparam ram_block1a82.port_a_address_clear = "none";
defparam ram_block1a82.port_a_address_width = 13;
defparam ram_block1a82.port_a_data_out_clear = "none";
defparam ram_block1a82.port_a_data_out_clock = "clock0";
defparam ram_block1a82.port_a_data_width = 1;
defparam ram_block1a82.port_a_first_address = 40960;
defparam ram_block1a82.port_a_first_bit_number = 2;
defparam ram_block1a82.port_a_last_address = 49151;
defparam ram_block1a82.port_a_logical_ram_depth = 65536;
defparam ram_block1a82.port_a_logical_ram_width = 16;
defparam ram_block1a82.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a82.ram_block_type = "auto";
defparam ram_block1a82.mem_init3 = "A5AD694A5AD694B5AD294B5AD294B5AD294B5AD294B5AD294B5AD294B5A5296B5A5296B5A5296B5A5296B4A52D6B4A52D6B4A52D694A5AD694A5AD694B5AD294B5AD294B5A5296B5A52D6B4A52D6B4A5AD694A5AD294B5AD296B5A52D6B4A52D694A5AD294B5AD296B5A52D6B4A5AD694B5AD296B4A52D694A5AD294B5A52D6B4A5AD694B5A5296B4A5AD294B5A52D6B4A5AD296B5A52D694B5A5296B4A5AD296B4A5AD694B5A52D694B5A52D694B5A52D694A5AD296B4A5A52D694B5A52D694B5A52D694B5A52D296B4A5AD296B4B5A52D694B5A5AD296B4B5A52D694B4A5AD2D694B5A5AD29694B5A5AD29694B5A5AD29694B4A5AD2D696B4A5A52D29694B5";
defparam ram_block1a82.mem_init2 = "A5AD2D696B4B5A5AD2D696B4B5A5AD2D696B4B4A5A52D29696B4B5A5AD2D29696B4B5A5A52D2D696B4B4A5A5AD2D2969694B4B5A5A52D2D29696B4B4B5A5A5AD2D2D69696B4B4B4A5A5A5AD2D2D2969696B4B4B4B5A5A5A5AD2D2D2D696969696B4B4B4B4B5A5A5A5A5A5AD2D2D2D2D2D2D296969696969696969694B4B4B4B4B4B4B4B4B4B4B4B4B4B4B4B4B4B4B4B4B4B4B4B4B4B696969696969696969692D2D2D2D2D2D25A5A5A5A5A4B4B4B4B49696969692D2D2D25A5A5A4B4B4B4969696D2D2D25A5A5B4B4B69696D2D2DA5A5B4B4B69692D2D25A5B4B49696D2D25A5B4B49696D2DA5A4B4B696D2DA5A4B49692D2DA5B4B696D2DA5B4B696D2DA5B49";
defparam ram_block1a82.mem_init1 = "692D25A4B696D2DA4B49692DA5B49692DA5B49692DA4B496D25A4B692DA5B496D25B4B692DA4B692DA4B696D25B496D25B496D24B692DA4B692DA4B6D25B496D24B692DA496D25B692DB496D24B6925B492DA496D24B6D25B6925B692DB492DB492DA496DA496DA496DB492DB492DB4925B6924B6D24B6DA492DB4925B6D2496DB4925B6D2496DB4924B6DA4925B6DA4925B6DA4925B6DA4924B6DB492496DB6DA4924B6DB6D2492496DB6DA4924925B6DB6DA492492496DB6DB6DA492492492496DB6DB6DB6DB6DB4924924924924924924924924924924924924924924924924924926DB6DB6DB6DB6DB24924924924DB6DB6DB649249249B6DB6DB2492493";
defparam ram_block1a82.mem_init0 = "6DB6D924924DB6DB24924DB6DB24926DB6C9249B6DB24936DB64926DB64926DB64926DB24936DB249B6C924DB64936D924DB64936D926DB249B64936D926DB24DB649B64936C936C936D926D926D926D926D926D926D926C936C93649B649B24DB26D926C93649B24DB26D93649B24D926C9B64D926C9B64D926C9B24D93649B26C9B64D9364D926C9B26C9B26C9B26C9B26C9B26C9B26C9B26C9B26C9B364D9364D9B26C9B364D9366C9B264D9326C99364C9B264D9B26CD9326CD9326CD9326CD93264D9B364C99366CD93264C9B366CD9B364C993264C993264C993264C99B366CD9B3264C993366CD993266CD993266CD993266CC99B3664CD9933664CD9";

arriav_ram_block ram_block1a98(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a98_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a98.clk0_core_clock_enable = "ena0";
defparam ram_block1a98.clk0_input_clock_enable = "ena0";
defparam ram_block1a98.clk0_output_clock_enable = "ena0";
defparam ram_block1a98.data_interleave_offset_in_bits = 1;
defparam ram_block1a98.data_interleave_width_in_bits = 1;
defparam ram_block1a98.init_file = "DDS_48_v1_nco_ii_0_cos.hex";
defparam ram_block1a98.init_file_layout = "port_a";
defparam ram_block1a98.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0121|altsyncram:altsyncram_component0|altsyncram_78g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a98.operation_mode = "rom";
defparam ram_block1a98.port_a_address_clear = "none";
defparam ram_block1a98.port_a_address_width = 13;
defparam ram_block1a98.port_a_data_out_clear = "none";
defparam ram_block1a98.port_a_data_out_clock = "clock0";
defparam ram_block1a98.port_a_data_width = 1;
defparam ram_block1a98.port_a_first_address = 49152;
defparam ram_block1a98.port_a_first_bit_number = 2;
defparam ram_block1a98.port_a_last_address = 57343;
defparam ram_block1a98.port_a_logical_ram_depth = 65536;
defparam ram_block1a98.port_a_logical_ram_width = 16;
defparam ram_block1a98.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a98.ram_block_type = "auto";
defparam ram_block1a98.mem_init3 = "4CD993266CC99B3266CD993366CC993366CC993366CC993266CD9B3664C993264C993366CD9B366CD9B264C993264C99366CD9B264C99366CD93264D9B264C9B364C9B364C9B364C9B264D9B26CD9366C9B364D9B26C99364D9B26C9B364D9364D9B26C9B26C9B26CD9364D9364D9364D93649B26C9B26C9B26C9364D93649B26C9B64D936C9B26D93649B26D93649B24D936C9B64DB26D936C93649B24DB26D926C936C9B649B649B24DB24DB24DB24DB24DB24DB24DB649B649B6C936C926D926DB24DB64936C926DB249B64936D924DB64926DB249B6C924DB64926DB64936DB24936DB64926DB64924DB6D924936DB64924DB6DB24924DB6DB249249B6DB";
defparam ram_block1a98.mem_init2 = "6D9249249B6DB6DB24924924DB6DB6DB6C924924924936DB6DB6DB6DB6DB6D92492492492492492492492492492492492492492496DB6DB6DB6DB6DB6DA492492492496DB6DB6DB6924924925B6DB6DA4924925B6DB6D24924B6DB6D24924B6DB692492DB6DA4924B6DB4924B6DB4924B6DB4924B6DA4925B6D2496DB4925B6D2496DB4925B6D24B6DA496DB492DB6925B6924B6D24B6D24B6D24B6D24B6D24B6D24B6925B6925B492DA496DA4B6D25B692DB496DA4B6925B492DA4B6925B496D24B692DA4B6D25B496D25B496D25B496D25B496D25B496D25B496D25A4B692DA4B496D25B4B692DA5B496D2DA4B496D2DA4B496D2DA4B496D2DA5B49692D25A";
defparam ram_block1a98.mem_init1 = "4B496D2DA5B4B696D2DA5B4B49692D25A4B49696D2DA5A4B49696D2D25A4B4B69692D2DA5A4B4B69696D2D25A5B4B4B69696D2D2DA5A5B4B4B4969692D2D2DA5A5A4B4B4B496969692D2D2D2DA5A5A5A4B4B4B4B4969696969692D2D2D2D2D2D2DA5A5A5A5A5A5A5A5A5B4B4B4B4B4B4B4B4B4B4B4B4B4B4B4B4B4B4B4B4B4B4B4B4B4B4A5A5A5A5A5A5A5A5A5A5AD2D2D2D2D2D2D69696969696B4B4B4B4B5A5A5A5A5AD2D2D2D296969694B4B4B5A5A5A5AD2D2D2969694B4B4B5A5A5AD2D2D69696B4B4B5A5A5AD2D29696B4B4B5A5A52D2D69694B4B5A5A52D29696B4B4A5A52D2D696B4B4A5A52D29696B4B5A5AD2D696B4B5A5AD2D696B4B5A5AD2D696";
defparam ram_block1a98.mem_init0 = "B4B5A52D29694B4A5AD2D696B4A5A52D696B4B5A52D296B4B5A52D696B4A5A52D694B4A5AD29694B5A52D296B4A5AD2D694B5A52D694B4A5AD296B4A5AD296B4A5A52D694B5A52D694B5A52D694B5A52D694B5A5296B4A5AD296B4A5AD296B4A52D694B5A52D6B4A5AD296B4A52D694B5A5296B4A5AD694B5A52D6B4A5AD694B5A5296B4A5AD694B5AD296B5A52D6B4A5AD694B5AD296B5A52D6B4A5AD694B5AD294B5A5296B4A52D6B4A5AD694A5AD294B5AD296B5A5296B5A52D6B4A52D6B4A5AD694A5AD694B5AD294B5AD294B5AD296B5A5296B5A5296B5A5296B4A52D6B4A52D6B4A52D6B4A52D6B4A52D694A5AD694A5AD694A5AD694A5AD694A5AD694";

arriav_ram_block ram_block1a114(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a114_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a114.clk0_core_clock_enable = "ena0";
defparam ram_block1a114.clk0_input_clock_enable = "ena0";
defparam ram_block1a114.clk0_output_clock_enable = "ena0";
defparam ram_block1a114.data_interleave_offset_in_bits = 1;
defparam ram_block1a114.data_interleave_width_in_bits = 1;
defparam ram_block1a114.init_file = "DDS_48_v1_nco_ii_0_cos.hex";
defparam ram_block1a114.init_file_layout = "port_a";
defparam ram_block1a114.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0121|altsyncram:altsyncram_component0|altsyncram_78g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a114.operation_mode = "rom";
defparam ram_block1a114.port_a_address_clear = "none";
defparam ram_block1a114.port_a_address_width = 13;
defparam ram_block1a114.port_a_data_out_clear = "none";
defparam ram_block1a114.port_a_data_out_clock = "clock0";
defparam ram_block1a114.port_a_data_width = 1;
defparam ram_block1a114.port_a_first_address = 57344;
defparam ram_block1a114.port_a_first_bit_number = 2;
defparam ram_block1a114.port_a_last_address = 65535;
defparam ram_block1a114.port_a_logical_ram_depth = 65536;
defparam ram_block1a114.port_a_logical_ram_width = 16;
defparam ram_block1a114.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a114.ram_block_type = "auto";
defparam ram_block1a114.mem_init3 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000001FFFFFFFFFFFFF00000000000FFFFFFFFFE000000001FFFFFFFE00000007FFFFFF8000000FFFFFF8000007FFFFF000001FFFFF000007FFFF800007FFFF00003FFFF00003FFFE0000FFFF80007FFF8000FFFF0001FFF8000FFFC000FFFC000FFFC001FFF0007FFC001FFE000FFF000FFF000FFE001FFE003FF800FFE003FF800FFE007FF003FF801FF801FF801FF801FF803FF007FE00FFC01FF007FC01FF007FC01FF007F803FE01FF00FF007F807FC03FC03FC03FC03FC03FC03FC07F807F00FF01FE03FC07F00FE03FC07F01FC03F80FE03F80FE03F80FC07F01FC0FE03F01FC0FE03F0";
defparam ram_block1a114.mem_init2 = "1F80FC0FE07F03F01F81FC0FC0FE07E07E07E03F03F03F03F03F07E07E07E07E0FC0FC1F81F83F03E07E0FC1F81F03E07C0F81F07E0FC1F83E07C1F83E0FC1F07E0F83F07C1F07C0F83E0F83E0F83E0F83E0F83E0F83E0F87C1F07C1E0F83E1F07C3E0F87C1E0F83C1F0F87C1E0F87C3E1F0783C1E0F0783C1E0F0F87C3E1E0F0787C3C1E1F0F0787C3C3E1E1F0F0F878783C3C3E1E1E1F0F0F0F0F878787878787878783C3C3C3C3C787878787878787870F0F0F0E1E1E1E3C3C3C787870F0F1E1E3C3C7878F0F1E1C3C3878F0E1E3C3878F1E1C3C78F0E1C3C78F1E1C3870E1C3C78F1E3C78F1E3C70E1C3870E3C78F1E3870E3C78E1C78F1C38F1E3871E38";
defparam ram_block1a114.mem_init1 = "71E38F1C38F1C78E1C70E3871C38E1C70E3871C78E3871C78E38F1C71E38E3C71C70E38E38F1C71C70E38E38E3871C71C71C71C71C38E38E38E38E38E38E38E38E39C71C71C71C71C718E38E38E39C71C71CE38E38C71C718E38E71C718E38C71C638E71C738E31C738E31C638E71CE39C718E31C638C738E71CE31C639C738C718E718E718E31CE31CE31CE318E718E718C738C639C631CE318E738C639CE718C739CE318C739CE718C6318E739CE739C6318C6318C6318C6318C6318C6318C6739CE739CE6318C6339CE7318C6739CC6319CE6318CE7318CE7318CE7319CE6319CC63398CE7319CC67398CE63398CE63398CE63398CE67319CC663398CC673";
defparam ram_block1a114.mem_init0 = "198CE673198CC673399CC6633198CC6633198CC6633199CCE6733198CCE6633199CCC66733199CCC667333998CCE667333999CCCE6673339998CCC666733319998CCCE666733339999CCCCC666673333399999CCCCCE6666673333339999999CCCCCCCC666666667333333333399999999999999CCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCC9999999999999933333333332666666666CCCCCCCD99999993333336666664CCCCC99999B3333266664CCCC99999333366664CCCD999B3336666CCCD999B3336664CCD9993336664CCD999332666CCD99B332664CC999332664CD99B33664CC99B33664CD99B3266CC9993366";

arriav_ram_block ram_block1a34(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a34_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a34.clk0_core_clock_enable = "ena0";
defparam ram_block1a34.clk0_input_clock_enable = "ena0";
defparam ram_block1a34.clk0_output_clock_enable = "ena0";
defparam ram_block1a34.data_interleave_offset_in_bits = 1;
defparam ram_block1a34.data_interleave_width_in_bits = 1;
defparam ram_block1a34.init_file = "DDS_48_v1_nco_ii_0_cos.hex";
defparam ram_block1a34.init_file_layout = "port_a";
defparam ram_block1a34.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0121|altsyncram:altsyncram_component0|altsyncram_78g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a34.operation_mode = "rom";
defparam ram_block1a34.port_a_address_clear = "none";
defparam ram_block1a34.port_a_address_width = 13;
defparam ram_block1a34.port_a_data_out_clear = "none";
defparam ram_block1a34.port_a_data_out_clock = "clock0";
defparam ram_block1a34.port_a_data_width = 1;
defparam ram_block1a34.port_a_first_address = 16384;
defparam ram_block1a34.port_a_first_bit_number = 2;
defparam ram_block1a34.port_a_last_address = 24575;
defparam ram_block1a34.port_a_logical_ram_depth = 65536;
defparam ram_block1a34.port_a_logical_ram_width = 16;
defparam ram_block1a34.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a34.ram_block_type = "auto";
defparam ram_block1a34.mem_init3 = "3664CD9933664CD9B3266CC993366CC993366CC993366CD993264C99B366CD9B3264C993264C993264C993264D9B366CD9B264C99366CD93264D9B364C99366C99366C99366C99366C9B364C9B264D9326C99364C9B26CD9364D9B26C9B364D9364D9B26C9B26C9B26C9B26C9B26C9B26C9B26C9B26C9B26C9364D9364DB26C9B24D93649B26C9364DB26C9364DB26C93649B24D936C9B649B24D926C936C9B649B24DB24D926D926C936C936C936C936C936C936C936D926D926D924DB24DB649B6C936D924DB249B6C936D924DB64936D924DB64926DB249B6D9249B6C924DB6C924DB6C924DB6D9249B6DB24926DB6C9249B6DB649249B6DB64924936DB6D";
defparam ram_block1a34.mem_init2 = "9249249B6DB6DB24924924DB6DB6DB649249249249B6DB6DB6DB6DB6C924924924924924924924924924924924924924924924924924925B6DB6DB6DB6DB6D24924924924B6DB6DB6D24924924B6DB6DB4924924B6DB6D2492496DB6DA4924B6DB6D24925B6DA4924B6DB4924B6DB4924B6DB4924B6DA4925B6D2496DB4925B6D2496DB4925B6924B6DA496DA492DB4925B6925B6925B6D24B6D24B6D24B6925B6925B692DB492DB496DA496D24B6925B492DA496D25B692DB496D24B692DA496D25B496DA4B692DA4B692DA496D25B496D25B496D2DA4B692DA4B692DA5B496D25B4B692DA4B496D25A4B692D25B4B692D25B4B692D25A4B696D2DA4B49692D";
defparam ram_block1a34.mem_init1 = "25B4B696D2DA5B4B696D2DA5B4B69692D25A4B4B696D2DA5A4B4B696D2D25A5B4B49696D2D25A5B4B4969692D2DA5A5B4B4B69696D2D2DA5A5B4B4B4969696D2D2D25A5A5A4B4B4B496969692D2D2D2D25A5A5A5A4B4B4B4B4B496969696969692D2D2D2D2D2D2D2D2D2DA5A5A5A5A5A5A5A5A5A5A5A5A5A5A5A5A5A5A5A5A5A5A5A5A5A52D2D2D2D2D2D2D2D2D296969696969696B4B4B4B4B4B5A5A5A5A5AD2D2D2D2D6969696B4B4B4B5A5A5A5AD2D2D2969696B4B4B4A5A5A5AD2D2D69696B4B4B5A5A5AD2D2969694B4B5A5A52D2D29696B4B4A5A5AD2D69694B4B5A5AD2D29696B4B5A5AD2D29694B4A5A5AD2D696B4B5A5AD2D696B4B5A5AD2D696B4B";
defparam ram_block1a34.mem_init0 = "5A52D29694B4A5AD2D696B4A5A52D296B4B5A52D296B4B5A52D296B4B5A52D696B4A5A52D694B5A5AD296B4B5A52D694B5A5AD296B4A5AD29694B5A52D694B5A52D694B5A52D694B4A5AD296B4A52D694B5A52D694B5A52D694B5A52D6B4A5AD296B4A5AD294B5A52D694B5AD296B4A5AD694B5A5296B4A5AD294B5A52D6B4A5AD694B5A5296B4A52D694A5AD296B5A52D6B4A5AD694B5AD296B5A5296B4A52D694A5AD694B5AD296B5A5296B4A52D6B4A5AD694A5AD694B5AD294B5A5296B5A5296B5A52D6B4A52D6B4A52D694A5AD694A5AD694A5AD294B5AD294B5AD294B5AD294B5A5296B5A5296B5A5296B5A5296B5A5296B5A5296B5A52D6B4A52D6B4A";

arriav_ram_block ram_block1a50(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a50_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a50.clk0_core_clock_enable = "ena0";
defparam ram_block1a50.clk0_input_clock_enable = "ena0";
defparam ram_block1a50.clk0_output_clock_enable = "ena0";
defparam ram_block1a50.data_interleave_offset_in_bits = 1;
defparam ram_block1a50.data_interleave_width_in_bits = 1;
defparam ram_block1a50.init_file = "DDS_48_v1_nco_ii_0_cos.hex";
defparam ram_block1a50.init_file_layout = "port_a";
defparam ram_block1a50.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0121|altsyncram:altsyncram_component0|altsyncram_78g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a50.operation_mode = "rom";
defparam ram_block1a50.port_a_address_clear = "none";
defparam ram_block1a50.port_a_address_width = 13;
defparam ram_block1a50.port_a_data_out_clear = "none";
defparam ram_block1a50.port_a_data_out_clock = "clock0";
defparam ram_block1a50.port_a_data_width = 1;
defparam ram_block1a50.port_a_first_address = 24576;
defparam ram_block1a50.port_a_first_bit_number = 2;
defparam ram_block1a50.port_a_last_address = 32767;
defparam ram_block1a50.port_a_logical_ram_depth = 65536;
defparam ram_block1a50.port_a_logical_ram_width = 16;
defparam ram_block1a50.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a50.ram_block_type = "auto";
defparam ram_block1a50.mem_init3 = "00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFE00000000000000FFFFFFFFFFFC0000000003FFFFFFFFC00000001FFFFFFFC0000003FFFFFF8000001FFFFFE000001FFFFF800001FFFFF00000FFFFF00001FFFFC0000FFFFC0001FFFF0000FFFF80007FFF0000FFFE0003FFF0001FFF8001FFF8003FFF0007FFC001FFE000FFF0007FF8007FF8007FF000FFE003FFC007FF001FF800FFE007FF003FF001FF801FF801FF003FF007FE00FFC01FF803FE00FF803FE00FF803FC01FF00FF803FC03FE01FE00FF00FF00FF00FF00FF00FF00FE01FE03FC03F807F00FE01FC07F80FE03F807F01FC07F01FC07F01FC07F03F80FE07F01F80FE07F03F";
defparam ram_block1a50.mem_init2 = "81FC0FE07F03F01F81FC0FC07E07E07F03F03F03F03F03F03F03F03F03F07E07E07C0FC0F81F81F03F07E0FC0F81F03E07C0F81F03E0FC1F83E07C1F83E0FC1F07E0F83E07C1F07C1F83E0F83E0F83E0F83E0F83E0F83C1F07C1F0783E0F87C1F0F83E1F07C3E0F07C3E0F07C3E1F0783C1E0F07C3E1F0F8783C1E0F0787C3E1E0F0787C3C1E1F0F0F8783C3C1E1E0F0F0F878783C3C3C1E1E1E1E1F0F0F0F0F0F0F0F0F87878787870F0F0F0F0F0F0F0F1E1E1E1E1C3C3C38787870F0F1E1E1C3C387870F0E1E1C3C7878F0E1E3C3878F0E1E3C7870E1E3C7870E1E3C78F1E1C3870E1C3870E1C3870E1C78F1E3C78E1C38F1E3C70E1C78E1C38F1C38F1C38F";
defparam ram_block1a50.mem_init1 = "1C38F1C38E1C78E3C70E3871C38E1C70E38F1C78E3871C78E38F1C70E38E3C71C70E38E3871C71C78E38E38E1C71C71C71C71E38E38E38E38E38E38E38E38E38E38E38E39C71C71C71C718E38E38E39C71C718E38E39C71C738E38C71C638E39C718E38C71CE38C71CE38C71CE39C718E31C638C718E31C639C738E718E31CE31C639C639C638C738C738C739C639C639C631CE318E718C739C631CE718C739C6318E739C6318E739CE318C631CE739CE739C6318C6318C6318C6318C6318CE739CE739CE6318C6339CE7318C6339CE6318CE7318C67398C67398C67398CE7318CE6319CC63398CE6319CC67319CC67319CC67319CC673198CE63399CC673398";
defparam ram_block1a50.mem_init0 = "CE673198CE673398CC663319CCE673399CCE6733998CC6633199CCE6633199CCC66733998CCE66733199CCC666333199CCCE667333999CCCC66633339998CCCE666733319998CCCC66667333319999CCCCCE66667333331999998CCCCCCE6666667333333339999999998CCCCCCCCCCCE666666666666666663333333333333333333333333333333333333333332666666666666666666CCCCCCCCCCCD999999999B3333333266666664CCCCCC999999B33333666666CCCCC999993333266664CCCC9999B33366664CCC9999B3336664CCC999B3336664CCD9993336664CC999B33666CCC999332664CC99933266CCD99B32664CD99B3266CCD9933664CD993";

arriav_ram_block ram_block1a2(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a2_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.clk0_input_clock_enable = "ena0";
defparam ram_block1a2.clk0_output_clock_enable = "ena0";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.init_file = "DDS_48_v1_nco_ii_0_cos.hex";
defparam ram_block1a2.init_file_layout = "port_a";
defparam ram_block1a2.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0121|altsyncram:altsyncram_component0|altsyncram_78g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.operation_mode = "rom";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 13;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "clock0";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 8191;
defparam ram_block1a2.port_a_logical_ram_depth = 65536;
defparam ram_block1a2.port_a_logical_ram_width = 16;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.ram_block_type = "auto";
defparam ram_block1a2.mem_init3 = "CD9933266CC99B33664CD99B32664CD99B33664CC999332664CC999B33666CCC9993336664CCD9993336664CCD999B3336666CCCD999B33366664CCCD99993333266664CCCC99999B33332666664CCCCCD999999333333366666666CCCCCCCCC9999999999933333333333332666666666666666666666666666666666666666666666666666666666666667333333333333339999999999CCCCCCCCC666666673333333999999CCCCCCE666673333399999CCCCC6666733339999CCCCE66633331999CCCC6663333999CCCE667333999CCCE66333999CCC66733199CCC66733198CCE6633199CCE6733198CC6633198CC6633198CC673399CC663319CCE6331";
defparam ram_block1a2.mem_init2 = "9CC663398CC67319CCE63398CE63398CE63398CE6339CC67319CE63398C67318CE7319CE6319CE6319CE6318CE7318C6739CC6319CE7398C6318CE739CE739CC6318C6318C6318C6318C6318C6318C739CE739CE318C631CE739C6318E739C631CE738C639CE318E718C738C639C631CE31CE318E718E718E718E31CE31CE31C639C738C718E71CE39C638C718E31C738E71CE38C718E39C718E39C71CE38C71C638E31C71CE38E31C71C638E38E71C71C738E38E38E31C71C71C71C71C738E38E38E38E38E38E38E38E3871C71C71C71C71C38E38E38E1C71C71E38E38E1C71C78E38F1C71E38E3C71C38E3C71C38E1C70E3871C38E1C70E3C71E3871E38F1C";
defparam ram_block1a2.mem_init1 = "38F1C38F1E3871E3C70E3C78E1C38F1E3C78E1C3870E1C78F1E3C78F1E3C7870E1C3870F1E3C7870E1E3C7870F1E3C3878F0E1E3C387870F1E1E3C3C7878F0F1E1E1C3C3C787878F0F0F0E1E1E1E1C3C3C3C3C3C3C3C3C78787878783C3C3C3C3C3C3C3C3E1E1E1E1F0F0F0F878783C3C3E1E1F0F0F8787C3C1E1F0F0787C3C1E0F0F87C3E1E0F0783C1E0F0783C1F0F87C3E0F07C3E1F0783E0F07C3E0F87C1F0F83E0F07C1F07C3E0F83E0F83E0F83E0F83E0F83E0F83E07C1F07C1F83E0FC1F07E0F83F07C0F83F07E0FC1F03E07C0F81F03F07E0FC0F81F83F03F07E07E0FC0FC0FC0FC1F81F81F81F81F80FC0FC0FC0FE07E07F03F01F81FC0FE07E03F0";
defparam ram_block1a2.mem_init0 = "1F80FE07F01F80FE07F01FC07E03F80FE03F80FE03F807F01FC07F80FE01FC07F80FF01FE01FC03FC07F807F807F807F807F807F807FC03FC01FE01FF00FF803FC01FF007FC01FF007FC01FF007FE00FFC01FF803FF003FF003FF003FF003FF801FFC00FFE003FF800FFE003FF800FFF000FFE001FFE001FFE000FFF0007FFC001FFF0007FFE0007FFE0007FFE0003FFF0001FFFE0003FFFC0003FFFE0000FFFF80001FFFF80001FFFFC00003FFFFC00001FFFFF000001FFFFFC000003FFFFFE0000003FFFFFFC0000000FFFFFFFF000000000FFFFFFFFFE00000000001FFFFFFFFFFFFF000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

arriav_ram_block ram_block1a18(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a18_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a18.clk0_core_clock_enable = "ena0";
defparam ram_block1a18.clk0_input_clock_enable = "ena0";
defparam ram_block1a18.clk0_output_clock_enable = "ena0";
defparam ram_block1a18.data_interleave_offset_in_bits = 1;
defparam ram_block1a18.data_interleave_width_in_bits = 1;
defparam ram_block1a18.init_file = "DDS_48_v1_nco_ii_0_cos.hex";
defparam ram_block1a18.init_file_layout = "port_a";
defparam ram_block1a18.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0121|altsyncram:altsyncram_component0|altsyncram_78g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a18.operation_mode = "rom";
defparam ram_block1a18.port_a_address_clear = "none";
defparam ram_block1a18.port_a_address_width = 13;
defparam ram_block1a18.port_a_data_out_clear = "none";
defparam ram_block1a18.port_a_data_out_clock = "clock0";
defparam ram_block1a18.port_a_data_width = 1;
defparam ram_block1a18.port_a_first_address = 8192;
defparam ram_block1a18.port_a_first_bit_number = 2;
defparam ram_block1a18.port_a_last_address = 16383;
defparam ram_block1a18.port_a_logical_ram_depth = 65536;
defparam ram_block1a18.port_a_logical_ram_width = 16;
defparam ram_block1a18.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a18.ram_block_type = "auto";
defparam ram_block1a18.mem_init3 = "52D6B4A52D6B4A52D6B4A52D6B4A52D6B4A52D694A5AD694A5AD694A5AD694A5AD694A5AD294B5AD294B5AD294B5AD296B5A5296B5A5296B5A52D6B4A52D6B4A5AD694A5AD694B5AD294B5AD296B5A5296B4A52D6B4A5AD694A5AD294B5A5296B5A52D6B4A5AD694B5AD296B5A52D6B4A5AD694B5AD296B5A52D6B4A5AD294B5A52D6B4A5AD694B5A52D6B4A5AD294B5A52D694A5AD296B4A5AD694B5A52D694A5AD296B4A5AD296B4A5AD294B5A52D694B5A52D694B5A52D694B5A52D694B4A5AD296B4A5AD296B4A5A52D694B5A52D696B4A5AD29694B5A52D296B4A5A52D694B4A5AD2D694B5A5AD29694B5A5AD2D694B4A5AD2D696B4A5A52D29694B5A5A";
defparam ram_block1a18.mem_init2 = "D2D696B4B5A5AD2D696B4B5A5AD2D696B4B5A5AD2D29694B4A5A5AD2D69694B4A5A5AD2D29694B4B5A5A52D2D69694B4B5A5A5AD2D29696B4B4B5A5A5AD2D2D69696B4B4B5A5A5A52D2D2969696B4B4B4B5A5A5A52D2D2D296969696B4B4B4B4B5A5A5A5A5AD2D2D2D2D2D6969696969696B4B4B4B4B4B4B4B4B4B4A5A5A5A5A5A5A5A5A5A5A5A5A5A5A5A5A5A5A5A5A5A5A5A5A5A5B4B4B4B4B4B4B4B4B4B696969696969692D2D2D2D2D25A5A5A5A4B4B4B4B696969692D2D2D25A5A5A4B4B4B6969692D2D25A5A5B4B4B69696D2D2DA5A5B4B49696D2D2DA5A4B4B69692D2DA5A4B49696D2D25A4B4B696D2D25A4B49692D25A5B4B696D2DA5B4B696D25A4";
defparam ram_block1a18.mem_init1 = "B49692D25B4B696D25A4B696D25A4B696D25A4B696D25B4B692DA5B496D25A4B692DA4B496D25B496D25B496D25B496D25B496D25B496D25B496DA4B692DA496D25B492DA4B6925B492DA4B6D25B692DB496DA4B6D24B6925B492DB492DA496DA496DA496DA496DA496DA496DA492DB492DB6925B6D24B6DA496DB4925B6D2496DB4925B6D2496DB4924B6DA4925B6DA4925B6DA4925B6DA4924B6DB692492DB6DA492496DB6DA492496DB6DB4924924B6DB6DB492492492DB6DB6DB6D24924924924B6DB6DB6DB6DB6DB6D24924924924924924924924924924924924924924936DB6DB6DB6DB6DB6D924924924926DB6DB6DB649249249B6DB6DB24924936D";
defparam ram_block1a18.mem_init0 = "B6DB249249B6DB649249B6DB64924DB6D924936DB64924DB6C924DB6D9249B6D924DB6C924DB64926DB249B6C924DB64936D924DB249B6C926D924DB649B6C936C926D926DB24DB24DB649B649B649B649B649B649B649B24DB24DB26D926C936C9B649B24D926D936C9B64DB26D93649B24D936C9B24D936C9B26D9364DB26C9B24D9364D926C9B26C9B26C9B24D9364D9364D9364D9366C9B26C9B26C9B364D9364D9B26C9B364D9326C9B364D9B26CD9366C9B364C9B264D9B264D9B264D9B264C9B364C99366CD93264C9B366CD93264C993264C9B366CD9B366CD993264C993264CD9B366CC993266CD993266CD993266CD993366CC99B3266CC9933664";

arriav_ram_block ram_block1a67(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a67_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a67.clk0_core_clock_enable = "ena0";
defparam ram_block1a67.clk0_input_clock_enable = "ena0";
defparam ram_block1a67.clk0_output_clock_enable = "ena0";
defparam ram_block1a67.data_interleave_offset_in_bits = 1;
defparam ram_block1a67.data_interleave_width_in_bits = 1;
defparam ram_block1a67.init_file = "DDS_48_v1_nco_ii_0_cos.hex";
defparam ram_block1a67.init_file_layout = "port_a";
defparam ram_block1a67.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0121|altsyncram:altsyncram_component0|altsyncram_78g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a67.operation_mode = "rom";
defparam ram_block1a67.port_a_address_clear = "none";
defparam ram_block1a67.port_a_address_width = 13;
defparam ram_block1a67.port_a_data_out_clear = "none";
defparam ram_block1a67.port_a_data_out_clock = "clock0";
defparam ram_block1a67.port_a_data_width = 1;
defparam ram_block1a67.port_a_first_address = 32768;
defparam ram_block1a67.port_a_first_bit_number = 3;
defparam ram_block1a67.port_a_last_address = 40959;
defparam ram_block1a67.port_a_logical_ram_depth = 65536;
defparam ram_block1a67.port_a_logical_ram_width = 16;
defparam ram_block1a67.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a67.ram_block_type = "auto";
defparam ram_block1a67.mem_init3 = "E3C7870E1E3C7870F1E3C3878F0E1C3C7870F1E1C3C7870F1E1C3C7870F1E1C3C3878F0E1E1C3C7878F0E1E1C3C387870F1E1E3C3C387870F0E1E1C3C3C787870F0F1E1E1C3C3C787870F0F0E1E1E1C3C3C3C78787870F0F0F0E1E1E1E1C3C3C3C3C38787878787870F0F0F0F0F0F0F0F0F1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E0F0F0F0F0F0F0F0F0F078787878787C3C3C3C3C3E1E1E1E1F0F0F0F07878783C3C3C1E1E1E0F0F0F878783C3C1E1E1F0F0F8787C3C3E1E1F0F0F8783C3C1E1F0F078783C3E1E0F0F8783C1E1F0F0787C3E1E0F0F87C3C1E0F0787C3E1F0F0783C1E0F0783C3E1F0F87C3E1F0F87C1E0F0783C1E0F07C3E1F0F8";
defparam ram_block1a67.mem_init2 = "3C1E0F87C3E0F07C3E1F0783E1F0783E1F0783E1F0783E0F07C3E0F87C1F0F83E1F07C3E0F83C1F07C3E0F83E1F07C1F0F83E0F83E1F07C1F07C1F0F83E0F83E0F83E0F83E0F83E0F83E0F83E0F83E0F83E0F81F07C1F07C1F03E0F83E0FC1F07C1F83E0F81F07C1F83E0FC1F07E0F83F07C0F83E07C1F83E07C0F83F07C0F81F07E0FC1F03E07C0F81F03E07C0F81F03E07C0F81F83F07E07C0F81F83F03E07C0FC0F81F83F03E07E07C0FC0FC1F81F83F03F03F03E07E07E07E07C0FC0FC0FC0FC0FC0FC0FC0FC0FC0FC0FC0FE07E07E07E07F03F03F03F81F81FC0FC0FE07E07F03F01F81FC0FC07E03F03F81FC0FE07F03F81FC0FE07F03F80FC07E03F81";
defparam ram_block1a67.mem_init1 = "FC07E03F81FC07F03F80FE07F01FC07F03F80FE03F80FE03F80FE03F80FE03F80FE03F80FF01FC07F00FE03F80FF01FC03F80FF01FC03F807F00FE01FC03F807F00FE01FE03FC03F807F80FF00FF01FE01FE01FE01FE01FC03FC03FC01FE01FE01FE01FE00FF00FF007F807FC03FC01FE00FF007F803FC01FE00FF807FC01FF00FF803FE00FF803FC01FF007FE00FF803FE00FF801FF007FE00FF801FF003FE007FC00FFC01FF801FF803FF003FF003FF003FF003FF003FF801FF800FFC00FFE007FF003FF800FFC007FF001FFC007FF001FFC007FF001FFE003FFC007FF800FFF001FFE001FFE001FFE001FFE001FFE000FFF0007FF8003FFE001FFF0007FFC";
defparam ram_block1a67.mem_init0 = "001FFF0003FFE000FFFC001FFF8001FFF8001FFF8001FFFC000FFFC0007FFF0001FFFC0007FFF0000FFFE0001FFFE0001FFFE0001FFFF0000FFFF80003FFFE00007FFFC0000FFFFC0000FFFFC00007FFFF00001FFFFE00003FFFFC00001FFFFE00000FFFFFC00001FFFFF800000FFFFFE000003FFFFFC000001FFFFFF0000007FFFFFE0000003FFFFFFC0000001FFFFFFF00000001FFFFFFFC00000001FFFFFFFF8000000007FFFFFFFFE0000000001FFFFFFFFFFC00000000000FFFFFFFFFFFFC00000000000007FFFFFFFFFFFFFFF80000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000000000000000000000000000";

arriav_ram_block ram_block1a83(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a83_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a83.clk0_core_clock_enable = "ena0";
defparam ram_block1a83.clk0_input_clock_enable = "ena0";
defparam ram_block1a83.clk0_output_clock_enable = "ena0";
defparam ram_block1a83.data_interleave_offset_in_bits = 1;
defparam ram_block1a83.data_interleave_width_in_bits = 1;
defparam ram_block1a83.init_file = "DDS_48_v1_nco_ii_0_cos.hex";
defparam ram_block1a83.init_file_layout = "port_a";
defparam ram_block1a83.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0121|altsyncram:altsyncram_component0|altsyncram_78g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a83.operation_mode = "rom";
defparam ram_block1a83.port_a_address_clear = "none";
defparam ram_block1a83.port_a_address_width = 13;
defparam ram_block1a83.port_a_data_out_clear = "none";
defparam ram_block1a83.port_a_data_out_clock = "clock0";
defparam ram_block1a83.port_a_data_width = 1;
defparam ram_block1a83.port_a_first_address = 40960;
defparam ram_block1a83.port_a_first_bit_number = 3;
defparam ram_block1a83.port_a_last_address = 49151;
defparam ram_block1a83.port_a_logical_ram_depth = 65536;
defparam ram_block1a83.port_a_logical_ram_width = 16;
defparam ram_block1a83.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a83.ram_block_type = "auto";
defparam ram_block1a83.mem_init3 = "C6318E739CE718C631CE739CE318C631CE739CE318C631CE739CE318C639CE739C6318C639CE739C6318C739CE738C6318C739CE718C6318E739CE718C631CE739CE318C639CE739C6318C739CE738C6318E739CE318C631CE739C6318C739CE718C631CE739CE318C639CE738C6318E739CE318C739CE718C631CE739C6318C739CE718C639CE738C631CE739C6318C739CE318C639CE718C639CE738C631CE738C6318E739C6318E739C6318E739C6318E739CE318C739C6318E739C6318E739C6318E739C631CE738C631CE738C639CE718C639CE318C739C6318E738C631CE718C639CE318E739C631CE718C639CE318E738C631CE718C739C631CE718C6";
defparam ram_block1a83.mem_init2 = "39CE318E738C639CE318E738C639CE318E738C739C631CE718C739C631CE318E738C639C631CE718C738C639CE31CE718E738C639C631CE318E738C739C639CE31CE718E738C738C639C631CE31CE718E738C738C639C639CE31CE318E718E718C738C738C639C639C639CE31CE31CE31CE318E718E718E718E718E738C738C738C738C738C738C738C738C738C738C738C738C738C718E718E718E718E718E31CE31CE31CE39C639C639C738C738C718E718E71CE31CE39C639C738C738E718E71CE31C639C638C738E718E31CE39C638C738E71CE31C639C738E718E31C639C738E718E31C638C738E71CE39C738E71CE31C638C718E31C638C718E31C638E";
defparam ram_block1a83.mem_init1 = "71CE39C738E71CE38C718E31C638E71CE39C718E31C738E71C638C71CE39C718E39C738E31C738E31C738E71C638E71C638E71C738E31C738E31C738E39C718E38C71CE38E71C638E31C718E38C71C638E31C718E38C71C638E39C71CE38E31C71CE38E71C718E38E71C71CE38E31C71C638E38C71C738E38E31C71C638E38E71C71C638E38E71C71C738E38E39C71C71C638E38E39C71C71C738E38E38E71C71C71C738E38E38E38E71C71C71C71C638E38E38E38E38E71C71C71C71C71C71C718E38E38E38E38E38E38E38E38E38E38E38E38E38E38E38E38E38E38E38E38E38E38E38E38E38E38E38E3C71C71C71C71C71C71C78E38E38E38E38E3C71C71C";
defparam ram_block1a83.mem_init0 = "71C71E38E38E38E3C71C71C71C38E38E38F1C71C71C38E38E3871C71C78E38E3871C71C38E38E3C71C70E38E3871C71E38E3871C71E38E3C71C78E38E1C71C38E3871C78E38F1C70E38E1C71E38E1C71E38E1C71E38E1C70E38F1C78E3871C38E3C71E38F1C78E3C71C38E1C78E3C71E38F1C78E1C70E3871E38F1C38E1C78E3C70E3871E3871E38F1C38F1C38F1C38F1C38F1C38F1C38F1C38F1C38F1C3871E3871E3C70E3C78E1C78F1C3871E3C70E1C78F1C3871E3C70E1C38F1E3C70E1C38F1E3C78E1C3870E1C78F1E3C78F1C3870E1C3870E1C3870E1C3870E1C3870E1C3870E1C3C78F1E3C78F1E1C3870E1E3C78F1E1C3870F1E3C7870E1E3C7870E1";

arriav_ram_block ram_block1a99(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a99_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a99.clk0_core_clock_enable = "ena0";
defparam ram_block1a99.clk0_input_clock_enable = "ena0";
defparam ram_block1a99.clk0_output_clock_enable = "ena0";
defparam ram_block1a99.data_interleave_offset_in_bits = 1;
defparam ram_block1a99.data_interleave_width_in_bits = 1;
defparam ram_block1a99.init_file = "DDS_48_v1_nco_ii_0_cos.hex";
defparam ram_block1a99.init_file_layout = "port_a";
defparam ram_block1a99.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0121|altsyncram:altsyncram_component0|altsyncram_78g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a99.operation_mode = "rom";
defparam ram_block1a99.port_a_address_clear = "none";
defparam ram_block1a99.port_a_address_width = 13;
defparam ram_block1a99.port_a_data_out_clear = "none";
defparam ram_block1a99.port_a_data_out_clock = "clock0";
defparam ram_block1a99.port_a_data_width = 1;
defparam ram_block1a99.port_a_first_address = 49152;
defparam ram_block1a99.port_a_first_bit_number = 3;
defparam ram_block1a99.port_a_last_address = 57343;
defparam ram_block1a99.port_a_logical_ram_depth = 65536;
defparam ram_block1a99.port_a_logical_ram_width = 16;
defparam ram_block1a99.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a99.ram_block_type = "auto";
defparam ram_block1a99.mem_init3 = "70E1E3C78F0E1C3C78F1E1C3870F1E3C78F0E1C3870F1E3C78F1E3C7870E1C3870E1C3870E1C3870E1C3870E1C3870E1C78F1E3C78F1E3870E1C3871E3C78F1C3870E3C78F1C3870E3C78E1C38F1E3870E3C78E1C38F1E3871E3C70E3C78E1C78E1C38F1C38F1C38F1E3871E3871E3871E3871C38F1C38F1C38F1C78E1C78E3C70E3871E38F1C38E1C78E3C71E3871C38E1C70E3871C38E1C70E3871C38E3C71E38F1C70E3871C78E3C71C38E3C71C38E3C71C38E3C71C78E3871C70E38F1C71E38E3C71C78E38F1C71C38E3871C71E38E3871C71C38E38F1C71C78E38E3871C71C38E38E3871C71C78E38E38E1C71C71C78E38E38E3C71C71C71C38E38E38E3";
defparam ram_block1a99.mem_init2 = "8E1C71C71C71C71C38E38E38E38E38E38F1C71C71C71C71C71C71C71C71C71E38E38E38E38E38E38E38E38E38E38E38E38E38E38E71C71C71C71C71C71C71C71C71C718E38E38E38E38E38E39C71C71C71C71C638E38E38E38C71C71C71C738E38E38E31C71C71C738E38E38C71C71C738E38E38C71C71C638E38E71C71C638E38E71C71C638E38C71C718E38E31C71C638E38C71C738E38C71C738E38C71C738E38C71C638E39C71CE38E71C738E39C71CE38E71C738E39C71CE38C71C638E71C738E31C738E39C718E39C718E39C718E39C718E39C718E39C718E39C738E31C738E71C638C71CE39C718E31C738E71CE38C718E31C738E71CE39C718E31C63";
defparam ram_block1a99.mem_init1 = "8C718E31C638C718E31C638C718E31C638C718E71CE39C738E718E31C638C738E71CE31C638C738E718E31C639C738C718E71CE31C639C738C718E71CE31CE39C638C738C718E718E31CE31CE39C639C738C738C718E718E718E31CE31CE31CE31C639C639C639C639C638C738C738C738C738C738C738C738C738C738C738C738C738C739C639C639C639C639C631CE31CE31CE318E718E718E738C738C739C639C639CE31CE31CE718E718C738C639C639CE31CE318E718C738C639C631CE318E718C738C639C631CE318E738C739C639CE318E718C739C639CE318E738C739C631CE718C738C639CE318E738C639CE318E738C639CE318E738C639CE318E7";
defparam ram_block1a99.mem_init0 = "38C639CE318E738C631CE718C739C6318E738C639CE318C739C6318E738C639CE718C739CE318E739C631CE738C631CE718C639CE718C739CE318C739CE318C739C6318E739C6318E739C6318E739C6318E739C6318C739CE318C739CE318C739CE718C639CE738C631CE738C6318E739C6318C739CE718C639CE738C6318E739C6318C739CE718C631CE739C6318C739CE718C631CE739C6318C739CE718C631CE739C6318C739CE738C6318E739CE318C631CE739C6318C639CE738C6318C739CE718C6318E739CE318C631CE739CE318C639CE739C6318C639CE738C6318C739CE738C6318C739CE738C6318E739CE718C6318E739CE718C6318E739CE718";

arriav_ram_block ram_block1a115(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a115_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a115.clk0_core_clock_enable = "ena0";
defparam ram_block1a115.clk0_input_clock_enable = "ena0";
defparam ram_block1a115.clk0_output_clock_enable = "ena0";
defparam ram_block1a115.data_interleave_offset_in_bits = 1;
defparam ram_block1a115.data_interleave_width_in_bits = 1;
defparam ram_block1a115.init_file = "DDS_48_v1_nco_ii_0_cos.hex";
defparam ram_block1a115.init_file_layout = "port_a";
defparam ram_block1a115.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0121|altsyncram:altsyncram_component0|altsyncram_78g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a115.operation_mode = "rom";
defparam ram_block1a115.port_a_address_clear = "none";
defparam ram_block1a115.port_a_address_width = 13;
defparam ram_block1a115.port_a_data_out_clear = "none";
defparam ram_block1a115.port_a_data_out_clock = "clock0";
defparam ram_block1a115.port_a_data_width = 1;
defparam ram_block1a115.port_a_first_address = 57344;
defparam ram_block1a115.port_a_first_bit_number = 3;
defparam ram_block1a115.port_a_last_address = 65535;
defparam ram_block1a115.port_a_logical_ram_depth = 65536;
defparam ram_block1a115.port_a_logical_ram_width = 16;
defparam ram_block1a115.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a115.ram_block_type = "auto";
defparam ram_block1a115.mem_init3 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000FFFFFFFFFFFFFFFFFFE0000000000000007FFFFFFFFFFFFF0000000000007FFFFFFFFFFE00000000007FFFFFFFFF8000000003FFFFFFFFC00000000FFFFFFFF80000000FFFFFFFE0000000FFFFFFF0000000FFFFFFE0000007FFFFFE000000FFFFFF000000FFFFFE000003FFFFF000003FFFFF000007FFFFC00001FFFFE00001FFFFE00003FFFF80000FFFFE00007FFFE00007FFFE00007FFFC0001FFFF00007FFF80003FFFC0003FFFC0003FFFC0007FFF8000FFFE0003FFF8000FFFC0007FFE0003FFF0003FFF0003FFF0007FFE000FFFC001FFF0003FF";
defparam ram_block1a115.mem_init2 = "E000FFF0007FFC001FFE000FFF0007FF8007FFC003FFC003FFC007FF8007FF800FFF001FFE003FFC007FF001FFE003FF800FFE007FF001FFC007FE003FF001FF800FFC007FE007FF003FF003FF003FF003FF003FF003FF007FE007FE00FFC01FF803FF007FE00FFC01FF007FE00FF803FE007FC01FF007FC01FF00FF803FE00FF807FC01FE00FF807FC03FE01FF00FF807FC03FC01FE01FF00FF00FF807F807F807F807FC03FC03FC07F807F807F807F807F00FF00FE01FE03FC03F807F80FF01FE03FC07F80FF01FE03FC07F00FE03FC07F01FE03F80FF01FC07F01FE03F80FE03F80FE03F80FE03F80FE03F80FC07F01FC07F03F80FE07F01FC0FE03F81FC0";
defparam ram_block1a115.mem_init1 = "7E03F01FC0FE07F01F80FC07E03F01F80FC07E07F03F81F80FC0FE07E03F03F81F80FC0FC0FE07E07F03F03F03F81F81F81F81F81FC0FC0FC0FC0FC0FC0FC0FC0FC1F81F81F81F81F81F03F03F03E07E07E0FC0FC0F81F81F03F07E07E0FC0F81F83F07E07C0FC1F83F03E07C0F81F03E07E0FC1F83F07C0F81F03E07C1F83F07E0F81F07E0FC1F03E0FC1F03E0F81F07E0F83F07C1F83E0FC1F07C0F83E0F81F07C1F03E0F83E0F81F07C1F07C1F07C1F83E0F83E0F83E0F83E0F83E0F83E0F87C1F07C1F07C1F07C3E0F83E0F87C1F07C1E0F83E0F07C1F0F83E0F07C1E0F83E1F07C3E0F07C1E0F87C1F0F83C1F0F83C1F0F83C1F0F87C1E0F87C3E0F0783";
defparam ram_block1a115.mem_init0 = "E1F0F87C1E0F0783C1E0F87C3E1F0F87C3E1F0F87C3E1E0F0783C1E0F0F87C3E1E0F0787C3E1E0F0787C3C1E0F0F8783C3E1E0F0F8783C3E1E0F0F8787C3C1E1E0F0F078783C3C1E1E0F0F078787C3C3C1E1E1F0F0F07878783C3C3C1E1E1E1F0F0F0F0787878787C3C3C3C3C3E1E1E1E1E1E1E1F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F1E1E1E1E1E1E1E3C3C3C3C3C3878787878F0F0F0F1E1E1E1E3C3C3C78787870F0F0E1E1E3C3C3C787870F0F1E1E1C3C387878F0F1E1E3C3C7878F0F1E1E3C3C7878F0E1E1C3C7878F0E1E1C3C7870F1E1C3C3878F0E1E3C3878F1E1C3C7870F1E3C3878F1E1C3C78F0E1E3C78";

arriav_ram_block ram_block1a35(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a35_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a35.clk0_core_clock_enable = "ena0";
defparam ram_block1a35.clk0_input_clock_enable = "ena0";
defparam ram_block1a35.clk0_output_clock_enable = "ena0";
defparam ram_block1a35.data_interleave_offset_in_bits = 1;
defparam ram_block1a35.data_interleave_width_in_bits = 1;
defparam ram_block1a35.init_file = "DDS_48_v1_nco_ii_0_cos.hex";
defparam ram_block1a35.init_file_layout = "port_a";
defparam ram_block1a35.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0121|altsyncram:altsyncram_component0|altsyncram_78g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a35.operation_mode = "rom";
defparam ram_block1a35.port_a_address_clear = "none";
defparam ram_block1a35.port_a_address_width = 13;
defparam ram_block1a35.port_a_data_out_clear = "none";
defparam ram_block1a35.port_a_data_out_clock = "clock0";
defparam ram_block1a35.port_a_data_width = 1;
defparam ram_block1a35.port_a_first_address = 16384;
defparam ram_block1a35.port_a_first_bit_number = 3;
defparam ram_block1a35.port_a_last_address = 24575;
defparam ram_block1a35.port_a_logical_ram_depth = 65536;
defparam ram_block1a35.port_a_logical_ram_width = 16;
defparam ram_block1a35.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a35.ram_block_type = "auto";
defparam ram_block1a35.mem_init3 = "0E1C3C78F0E1C3C78F1E1C3870F1E3C78F0E1C3870F1E3C78F1E3C7870E1C3870E1C3870E1C3870E1C3870E1C3870E1C3871E3C78F1E3C70E1C3870E3C78F1E3870E1C78F1E3870E1C78F1C3871E3C70E1C78F1C3871E3C70E3C78E1C78F1C38F1C3871E3871E3871E3871E3871E3871E3871E3871E3871E38F1C38F1C38E1C78E3C70E3871E38F1C38E1C70E3C71E38F1C78E3C70E3871C78E3C71E38F1C78E3871C38E3C71E38E1C70E38F1C70E38F1C70E38F1C70E38E1C71E38E3C71C38E3871C70E38E3C71C78E38F1C71C38E38F1C71C38E38E1C71C78E38E3871C71C38E38E3C71C71C38E38E3871C71C71E38E38E3871C71C71C78E38E38E38F1C71C";
defparam ram_block1a35.mem_init2 = "71C71C78E38E38E38E38E3C71C71C71C71C71C71C78E38E38E38E38E38E38E38E38E38E38E38E38E38E38E38E38E38E38E38E38E38E38E38E38E38E38E38E31C71C71C71C71C71C71CE38E38E38E38E38C71C71C71C71CE38E38E38E39C71C71C71CE38E38E39C71C71C738E38E38C71C71C738E38E39C71C71CE38E38C71C71CE38E38C71C718E38E39C71C638E38C71C718E38E71C71CE38E31C71CE38E71C718E38E71C738E38C71C638E31C718E38C71C638E31C718E38C71CE38E71C638E31C738E39C718E39C718E39C71CE38C71CE38C71CE39C718E39C718E39C738E31C738E71C638C71CE39C718E31C738E71CE38C718E31C638E71CE39C738E71C";
defparam ram_block1a35.mem_init1 = "E38C718E31C638C718E31C638C718E71CE39C738E71CE39C638C718E31CE39C738C718E31CE39C738C718E71CE39C638C738E718E31CE39C638C738C718E71CE31CE39C639C738C738E718E71CE31CE31C639C639C738C738C738E718E718E718E31CE31CE31CE31CE31C639C639C639C639C639C639C639C639C639C639C639C639C639CE31CE31CE31CE31CE318E718E718E718E738C738C738C639C639C631CE31CE318E718E738C738C639C639CE31CE718E718C738C639C639CE31CE718E738C739C639CE318E718C738C639CE31CE718E738C639C631CE718C738C639CE318E718C739C631CE718C739C639CE318E738C639CE318E738C639CE318E738";
defparam ram_block1a35.mem_init0 = "C631CE718C739C631CE718C639CE318E738C631CE718C739CE318E738C631CE718C639CE318C739C6318E738C631CE738C639CE718C639CE718C739CE318C739CE318C739CE318C739C6318E739CE318C739CE318C739CE318C739CE318C639CE718C639CE738C631CE738C6318E739C6318C739CE718C639CE738C631CE739C6318C739CE718C631CE739C6318E739CE318C639CE738C6318E739CE718C631CE739C6318C739CE718C6318E739CE318C639CE739C6318C739CE738C6318E739CE718C631CE739CE318C631CE739C6318C639CE739C6318C739CE738C6318C739CE738C6318E739CE718C6318E739CE718C6318E739CE718C631CE739CE318C6";

arriav_ram_block ram_block1a51(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a51_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a51.clk0_core_clock_enable = "ena0";
defparam ram_block1a51.clk0_input_clock_enable = "ena0";
defparam ram_block1a51.clk0_output_clock_enable = "ena0";
defparam ram_block1a51.data_interleave_offset_in_bits = 1;
defparam ram_block1a51.data_interleave_width_in_bits = 1;
defparam ram_block1a51.init_file = "DDS_48_v1_nco_ii_0_cos.hex";
defparam ram_block1a51.init_file_layout = "port_a";
defparam ram_block1a51.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0121|altsyncram:altsyncram_component0|altsyncram_78g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a51.operation_mode = "rom";
defparam ram_block1a51.port_a_address_clear = "none";
defparam ram_block1a51.port_a_address_width = 13;
defparam ram_block1a51.port_a_data_out_clear = "none";
defparam ram_block1a51.port_a_data_out_clock = "clock0";
defparam ram_block1a51.port_a_data_width = 1;
defparam ram_block1a51.port_a_first_address = 24576;
defparam ram_block1a51.port_a_first_bit_number = 3;
defparam ram_block1a51.port_a_last_address = 32767;
defparam ram_block1a51.port_a_logical_ram_depth = 65536;
defparam ram_block1a51.port_a_logical_ram_width = 16;
defparam ram_block1a51.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a51.ram_block_type = "auto";
defparam ram_block1a51.mem_init3 = "0000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000003FFFFFFFFFFFFFFFC00000000000007FFFFFFFFFFFE000000000007FFFFFFFFFF0000000000FFFFFFFFFC000000003FFFFFFFF000000007FFFFFFF00000001FFFFFFF00000007FFFFFF8000000FFFFFFC000001FFFFFF0000007FFFFF800000FFFFFE000003FFFFF000007FFFFE00000FFFFF000007FFFF80000FFFFF00001FFFFC00007FFFE00007FFFE00007FFFC0000FFFF80003FFFE0001FFFF0000FFFF0000FFFF0000FFFE0001FFFC0007FFF0001FFFC0007FFE0007FFF0003FFF0003FFF0003FFF0007FFE000FFF8001FFF000";
defparam ram_block1a51.mem_init2 = "7FFC001FFF000FFF8003FFC001FFE000FFF000FFF000FFF000FFF000FFF001FFE003FFC007FF800FFF001FFC007FF001FFC007FF001FFC007FE003FF801FFC00FFE007FE003FF003FF801FF801FF801FF801FF801FF803FF003FF007FE007FC00FF801FF003FE00FFC01FF003FE00FF803FE00FFC01FF007F803FE00FF803FE01FF007FC03FE00FF007F803FC01FE00FF007F807FC03FC01FE01FE00FF00FF00FF00FF007F807F807F00FF00FF00FF00FF01FE01FE03FC03F807F80FF00FE01FC03F807F00FE01FC03F807F01FE03F807F01FE03F80FE01FC07F01FE03F80FE03F80FE03F80FE03F80FE03F80FE03F81FC07F01FC0FE03F81FC07F03F80FC07F";
defparam ram_block1a51.mem_init1 = "03F80FC07E03F81FC0FE07F03F81FC0FE07F03F81F80FC07E07F03F01F81FC0FC0FE07E07F03F03F81F81F81FC0FC0FC0FC0FE07E07E07E07E07E07E07E07E07E07E07E07C0FC0FC0FC0F81F81F81F83F03F07E07E07C0FC0F81F83F03E07E07C0F81F83F03E07C0FC1F83F03E07C0F81F03E07C0F81F03E07C0F81F07E0FC1F03E07C1F83E07C0F83F07C0F83E07C1F83E0FC1F07E0F83F07C1F03E0F83F07C1F07E0F83E0F81F07C1F07C1F03E0F83E0F83E0F83E0F83E0F83E0F83E0F83E0F83E0F83E1F07C1F07C1F0F83E0F83E1F07C1F0F83E0F87C1F0783E0F87C1F0F83E1F07C3E0F87C1E0F83C1F0F83C1F0F83C1F0F83C1F0F87C1E0F87C3E0F078";
defparam ram_block1a51.mem_init0 = "3E1F0F87C1E0F0783C1E0F07C3E1F0F87C3E1F0F8783C1E0F0783C1E1F0F87C3C1E0F0787C3E1E0F0F87C3C1E1F0F0783C3E1E0F0F8783C3C1E1F0F078783C3E1E1F0F0F8787C3C3E1E1F0F0F078783C3C3E1E1E0F0F0F07878783C3C3C1E1E1E1F0F0F0F0F8787878787C3C3C3C3C3C1E1E1E1E1E1E1E1E1E0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F1E1E1E1E1E1E1E1E1E1C3C3C3C3C3C387878787870F0F0F0E1E1E1E1C3C3C3C78787870F0F0E1E1E1C3C3C787870F0F1E1E1C3C3C787870F0E1E1C3C387878F0F1E1C3C387870F0E1E3C3C7870F0E1E3C387870F1E1C3C7870F1E1C3C7870F1E1C3C7870E1E3C3878F1E1C3C78F0E1C3C78F";

arriav_ram_block ram_block1a3(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a3_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.clk0_input_clock_enable = "ena0";
defparam ram_block1a3.clk0_output_clock_enable = "ena0";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.init_file = "DDS_48_v1_nco_ii_0_cos.hex";
defparam ram_block1a3.init_file_layout = "port_a";
defparam ram_block1a3.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0121|altsyncram:altsyncram_component0|altsyncram_78g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.operation_mode = "rom";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 13;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "clock0";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 8191;
defparam ram_block1a3.port_a_logical_ram_depth = 65536;
defparam ram_block1a3.port_a_logical_ram_width = 16;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.ram_block_type = "auto";
defparam ram_block1a3.mem_init3 = "3C78F0E1E3C7870F1E3C3878F1E1C3C7870F1E3C3878F0E1E3C387870F1E1C3C7870F0E1E3C3C7870F0E1E3C3C7878F0F1E1E3C3C7878F0F1E1E3C3C387870F0F1E1E1C3C3C787878F0F0E1E1E1C3C3C3C787878F0F0F0F1E1E1E1E3C3C3C3C387878787878F0F0F0F0F0F0F1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1F0F0F0F0F0F0F0F8787878787C3C3C3C3C1E1E1E1F0F0F0F07878783C3C3C1E1E1F0F0F078787C3C3C1E1E0F0F078783C3C1E1E0F0F0787C3C3E1E0F0F8783C3E1E0F0F8783C3E1E0F0787C3C1E0F0F87C3C1E0F0F87C3E1E0F0783C1E0F0F87C3E1F0F87C3E1F0F87C3E0F0783C1E0F07C3E1F0F";
defparam ram_block1a3.mem_init2 = "83C1E0F87C3E0F07C3E1F0783E1F0783E1F0783E1F07C3E0F07C1E0F87C1F0F83E0F07C1E0F83E1F07C1E0F83E0F07C1F07C3E0F83E0F87C1F07C1F07C1F07C3E0F83E0F83E0F83E0F83E0F83E0F83F07C1F07C1F07C1F03E0F83E0F81F07C1F03E0F83E07C1F07E0F83F07C1F83E0FC1F03E0F81F07E0F81F07E0FC1F03E0FC1F83F07C0F81F03E07C1F83F07E0FC0F81F03E07C0F81F83F07E07C0FC1F83F03E07E0FC0FC1F81F03F03E07E07E0FC0FC0F81F81F81F03F03F03F03F03F07E07E07E07E07E07E07E07E07F03F03F03F03F03F81F81F81FC0FC0FE07E07E03F03F81F80FC0FE07E03F03F81FC0FC07E03F01F80FC07E03F01FC0FE07F01F80FC";
defparam ram_block1a3.mem_init1 = "07F03F80FE07F01FC0FE03F81FC07F01FC07E03F80FE03F80FE03F80FE03F80FE03F80FF01FC07F01FE03F80FF01FC07F80FE01FC07F80FF01FE03FC07F80FF01FE03FC03F807F80FF00FE01FE01FC03FC03FC03FC03FC07F807F807FC03FC03FC03FC03FE01FE01FF00FF007F807FC03FE01FF00FF807FC03FE00FF007FC03FE00FF803FE01FF007FC01FF007FC00FF803FE00FFC01FF007FE00FFC01FF803FF007FE00FFC00FFC01FF801FF801FF801FF801FF801FF801FFC00FFC007FE003FF001FF800FFC007FF001FFC00FFE003FF800FFF001FFC007FF800FFF001FFE003FFC003FFC007FF8007FF8007FFC003FFC001FFE000FFF0007FFC001FFE000F";
defparam ram_block1a3.mem_init0 = "FF8001FFF0007FFE000FFFC001FFF8001FFF8001FFF8000FFFC0007FFE0003FFF8000FFFE0003FFFC0007FFF80007FFF80007FFF80003FFFC0001FFFF00007FFFC0000FFFFC0000FFFFC0000FFFFE00003FFFF80000FFFFF00000FFFFF000007FFFFC00001FFFFF800001FFFFF800000FFFFFE000001FFFFFE000000FFFFFFC000000FFFFFFE0000001FFFFFFE0000000FFFFFFFE00000003FFFFFFFE000000007FFFFFFFF8000000003FFFFFFFFFC0000000000FFFFFFFFFFFC000000000001FFFFFFFFFFFFFC000000000000000FFFFFFFFFFFFFFFFFFE000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

arriav_ram_block ram_block1a19(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a19_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a19.clk0_core_clock_enable = "ena0";
defparam ram_block1a19.clk0_input_clock_enable = "ena0";
defparam ram_block1a19.clk0_output_clock_enable = "ena0";
defparam ram_block1a19.data_interleave_offset_in_bits = 1;
defparam ram_block1a19.data_interleave_width_in_bits = 1;
defparam ram_block1a19.init_file = "DDS_48_v1_nco_ii_0_cos.hex";
defparam ram_block1a19.init_file_layout = "port_a";
defparam ram_block1a19.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0121|altsyncram:altsyncram_component0|altsyncram_78g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a19.operation_mode = "rom";
defparam ram_block1a19.port_a_address_clear = "none";
defparam ram_block1a19.port_a_address_width = 13;
defparam ram_block1a19.port_a_data_out_clear = "none";
defparam ram_block1a19.port_a_data_out_clock = "clock0";
defparam ram_block1a19.port_a_data_width = 1;
defparam ram_block1a19.port_a_first_address = 8192;
defparam ram_block1a19.port_a_first_bit_number = 3;
defparam ram_block1a19.port_a_last_address = 16383;
defparam ram_block1a19.port_a_logical_ram_depth = 65536;
defparam ram_block1a19.port_a_logical_ram_width = 16;
defparam ram_block1a19.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a19.ram_block_type = "auto";
defparam ram_block1a19.mem_init3 = "31CE739CE318C631CE739CE318C631CE739CE318C639CE739C6318C639CE739C6318C639CE738C6318C739CE738C6318E739CE718C6318E739CE318C631CE739C6318C639CE738C6318C739CE718C6318E739CE318C639CE739C6318C739CE718C631CE739C6318C739CE718C631CE739C6318C739CE718C631CE739C6318C739CE318C639CE738C631CE739C6318C739CE318C639CE718C639CE738C631CE739C6318E739C6318E739C6318C739CE318C739CE318C739CE318C739CE318C739C6318E739C6318E739C631CE738C631CE718C639CE718C739CE318E739C631CE738C639CE318C739C6318E738C639CE318C739C631CE718C639CE318E738C639";
defparam ram_block1a19.mem_init2 = "CE318E738C639CE318E738C639CE318E738C639CE318E738C639C631CE718C739C639CE318E738C739C631CE318E738C739C639CE318E718C738C639C631CE318E718C738C639C631CE318E718E738C738C639C631CE31CE718E718E738C738C739C639C639CE31CE31CE318E718E718E718C738C738C738C738C739C639C639C639C639C639C639C639C639C639C639C639C639C638C738C738C738C738C718E718E718E718E31CE31CE31C639C639C738C738E718E718E31CE31C639C638C738E718E71CE31C639C738C718E71CE31C639C738C718E31CE39C638C718E71CE39C638C718E31CE39C738E71CE31C638C718E31C638C718E31C638C718E31C63";
defparam ram_block1a19.mem_init1 = "8C718E31C738E71CE39C718E31C638E71CE39C718E31C738E71C638C71CE39C718E39C738E31C738E31C738E31C738E31C738E31C738E31C738E39C718E39C71CE38C71C638E71C738E39C71CE38E71C738E39C71CE38E71C738E38C71C638E39C71C638E39C71C638E39C71C638E38C71C718E38E31C71C638E38C71C71CE38E38C71C71CE38E38C71C71C638E38E39C71C71C638E38E39C71C71C718E38E38E39C71C71C71C638E38E38E38C71C71C71C71C738E38E38E38E38E38E31C71C71C71C71C71C71C71C71C71CE38E38E38E38E38E38E38E38E38E38E38E38E38E38F1C71C71C71C71C71C71C71C71C71E38E38E38E38E38E3871C71C71C71C70E3";
defparam ram_block1a19.mem_init0 = "8E38E38E3871C71C71C78E38E38E3C71C71C70E38E38E3C71C71C38E38E3871C71C38E38E3C71C71E38E3871C71C38E38F1C71C38E3871C71E38E3C71C78E38F1C71E38E1C71C38E3C71C78E3871C78E3871C78E3871C78E3C71C38E1C71E38F1C78E3871C38E1C70E3871C38E1C70E3871C38F1C78E3C70E3871E38F1C38E1C78E3C70E3C71E3871E3871E3871C38F1C38F1C38F1C38F1E3871E3871E3870E3C70E3C78E1C78F1C38F1E3870E3C78E1C38F1E3870E3C78E1C3871E3C78E1C3871E3C78F1C3870E1C38F1E3C78F1E3C70E1C3870E1C3870E1C3870E1C3870E1C3870E1C3C78F1E3C78F1E1C3870E1E3C78F1E1C3870F1E3C7870E1E3C78F0E1C";

arriav_ram_block ram_block1a68(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a68_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a68.clk0_core_clock_enable = "ena0";
defparam ram_block1a68.clk0_input_clock_enable = "ena0";
defparam ram_block1a68.clk0_output_clock_enable = "ena0";
defparam ram_block1a68.data_interleave_offset_in_bits = 1;
defparam ram_block1a68.data_interleave_width_in_bits = 1;
defparam ram_block1a68.init_file = "DDS_48_v1_nco_ii_0_cos.hex";
defparam ram_block1a68.init_file_layout = "port_a";
defparam ram_block1a68.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0121|altsyncram:altsyncram_component0|altsyncram_78g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a68.operation_mode = "rom";
defparam ram_block1a68.port_a_address_clear = "none";
defparam ram_block1a68.port_a_address_width = 13;
defparam ram_block1a68.port_a_data_out_clear = "none";
defparam ram_block1a68.port_a_data_out_clock = "clock0";
defparam ram_block1a68.port_a_data_width = 1;
defparam ram_block1a68.port_a_first_address = 32768;
defparam ram_block1a68.port_a_first_bit_number = 4;
defparam ram_block1a68.port_a_last_address = 40959;
defparam ram_block1a68.port_a_logical_ram_depth = 65536;
defparam ram_block1a68.port_a_logical_ram_width = 16;
defparam ram_block1a68.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a68.ram_block_type = "auto";
defparam ram_block1a68.mem_init3 = "FC07F80FE03F807F01FC03F80FF01FC07F80FE01FC07F80FE01FC07F80FE01FC03F80FF01FE03F807F00FE01FC03F807F01FE03FC03F807F00FE01FC03F807F80FF01FE01FC03F807F80FF00FE01FE03FC03F807F807F00FF00FE01FE01FC03FC03FC07F807F807F80FF00FF00FF00FF00FE01FE01FE01FE01FE01FE01FE01FE01FE01FE01FE00FF00FF00FF00FF00FF807F807F807FC03FC03FC01FE01FE00FF00FF807F803FC03FE01FE00FF00FF807FC03FE01FE00FF007F803FC01FE00FF007FC03FE01FF007F803FC01FF00FF803FE01FF007F803FE00FF007FC01FF007F803FE00FF803FE00FF803FC01FF007FC01FF007FE00FF803FE00FF803FE00FF";
defparam ram_block1a68.mem_init2 = "C01FF007FC00FF803FE007FC01FF803FE007FC01FF803FF007FC00FF801FF003FE007FC00FFC01FF803FF003FE007FE00FFC00FFC01FF801FF801FF003FF003FF003FF003FF003FF003FF003FF003FF003FF001FF801FF801FFC00FFC00FFE007FE003FF001FF801FFC00FFE007FF003FF800FFC007FE003FF800FFC007FF001FF800FFE003FF800FFE003FF800FFE003FF800FFE003FF8007FF001FFC003FF800FFF001FFC003FF8007FF000FFE001FFC003FFC003FF8007FF8007FF000FFF000FFF000FFF000FFF000FFF000FFF8007FF8007FFC003FFC001FFE000FFF0007FF8003FFE001FFF0007FFC003FFE000FFF8003FFE000FFF8003FFF0007FFC001";
defparam ram_block1a68.mem_init1 = "FFF8003FFE0007FFC000FFF8001FFF8003FFF0003FFF0003FFF0003FFF0003FFF0003FFF0001FFF8000FFFC000FFFE0003FFF0001FFFC0007FFF0001FFFC0007FFF0001FFFC0003FFF8000FFFF0001FFFE0001FFFE0001FFFC0003FFFE0001FFFE0001FFFF0000FFFF80007FFFC0001FFFF00007FFFC0001FFFF00007FFFE0000FFFFC0000FFFFC0001FFFF80000FFFFC0000FFFFE00007FFFF00001FFFFC00007FFFF00001FFFFE00003FFFFC00003FFFFC00003FFFFC00001FFFFF00000FFFFF800003FFFFF000007FFFFE000007FFFFE000007FFFFE000003FFFFF800000FFFFFE000001FFFFFE000001FFFFFE000000FFFFFF8000003FFFFFE0000007FFF";
defparam ram_block1a68.mem_init0 = "FFE0000003FFFFFF0000001FFFFFFE0000001FFFFFFE0000000FFFFFFF80000001FFFFFFF80000000FFFFFFFE00000001FFFFFFFE00000000FFFFFFFFC000000007FFFFFFFF000000000FFFFFFFFF8000000001FFFFFFFFFC0000000001FFFFFFFFFF00000000001FFFFFFFFFFF000000000003FFFFFFFFFFFE0000000000007FFFFFFFFFFFFC00000000000001FFFFFFFFFFFFFFE0000000000000001FFFFFFFFFFFFFFFFF80000000000000000001FFFFFFFFFFFFFFFFFFFFFF000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000000000000000000000000000000000000000000000000000";

arriav_ram_block ram_block1a84(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a84_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a84.clk0_core_clock_enable = "ena0";
defparam ram_block1a84.clk0_input_clock_enable = "ena0";
defparam ram_block1a84.clk0_output_clock_enable = "ena0";
defparam ram_block1a84.data_interleave_offset_in_bits = 1;
defparam ram_block1a84.data_interleave_width_in_bits = 1;
defparam ram_block1a84.init_file = "DDS_48_v1_nco_ii_0_cos.hex";
defparam ram_block1a84.init_file_layout = "port_a";
defparam ram_block1a84.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0121|altsyncram:altsyncram_component0|altsyncram_78g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a84.operation_mode = "rom";
defparam ram_block1a84.port_a_address_clear = "none";
defparam ram_block1a84.port_a_address_width = 13;
defparam ram_block1a84.port_a_data_out_clear = "none";
defparam ram_block1a84.port_a_data_out_clock = "clock0";
defparam ram_block1a84.port_a_data_width = 1;
defparam ram_block1a84.port_a_first_address = 40960;
defparam ram_block1a84.port_a_first_bit_number = 4;
defparam ram_block1a84.port_a_last_address = 49151;
defparam ram_block1a84.port_a_logical_ram_depth = 65536;
defparam ram_block1a84.port_a_logical_ram_width = 16;
defparam ram_block1a84.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a84.ram_block_type = "auto";
defparam ram_block1a84.mem_init3 = "F83E0F83E0F81F07C1F07C1F03E0F83E0F83E0FC1F07C1F07C1F03E0F83E0F83E07C1F07C1F07C1F83E0F83E0F83F07C1F07C1F07E0F83E0F83E0F81F07C1F07C1F03E0F83E0F83E07C1F07C1F07C0F83E0F83E0FC1F07C1F07C1F83E0F83E0F81F07C1F07C1F03E0F83E0F83F07C1F07C1F03E0F83E0F81F07C1F07C1F83E0F83E0F81F07C1F07C0F83E0F83E07C1F07C1F03E0F83E0F81F07C1F07C0F83E0F83F07C1F07C1F83E0F83E07C1F07C1F83E0F83E0FC1F07C1F83E0F83E07C1F07C1F83E0F83E07C1F07C0F83E0F83F07C1F07E0F83E0FC1F07C1F83E0F83F07C1F07E0F83E0FC1F07C1F83E0F81F07C1F03E0F83F07C1F07E0F83E07C1F07E0F8";
defparam ram_block1a84.mem_init2 = "3E0FC1F07C0F83E0FC1F07C0F83E0FC1F07C0F83E07C1F07E0F83E07C1F03E0F83F07C1F83E0F81F07C0F83E0FC1F07E0F83F07C1F83E0FC1F07C0F83E07C1F03E0F81F07C0F83F07C1F83E0FC1F07E0F83F07C0F83E07C1F03E0FC1F07E0F81F07C0F83F07C1F83E07C1F03E0FC1F03E0FC1F07E0F81F07E0F81F07C0F83F07C0F83F07C0F83F07C0F83F07C0F83F07C0F83F07C0F81F07E0F81F07E0F81F03E0FC1F03E0FC1F83E07C1F83F07C0F81F07E0F81F03E0FC1F83E07C0F83F07E0F81F03E07C1F83F07C0F81F03E0FC1F83F07C0F81F03E07C1F83F07E0FC1F83E07C0F81F03E07C0F83F07E0FC1F83F07E0FC1F83F07E0FC1F83F07E0FC1F83F0";
defparam ram_block1a84.mem_init1 = "7E0FC1F83F07E0FC0F81F03E07C0F81F03E07E0FC1F83F07E07C0F81F03E07E0FC1F83F03E07C0FC1F83F07E07C0F81F83F07E07C0FC1F83F03E07C0FC1F81F03F07E0FC0F81F83F03E07E0FC0F81F83F03E07E0FC0F81F83F03E07E0FC0FC1F81F03F07E07E0FC0F81F81F03F03E07E07C0FC0F81F83F03F03E07E07C0FC0F81F81F83F03F07E07E07C0FC0FC1F81F81F83F03F03E07E07E07C0FC0FC0F81F81F81F83F03F03F03F07E07E07E07E07C0FC0FC0FC0FC0F81F81F81F81F81F81F81F03F03F03F03F03F03F03F03F03F03F03F03F03F03F03F03F03F03F03F03F03F03F03F03F03F03F03F03F81F81F81F81F81F81F80FC0FC0FC0FC0FC07E07E0";
defparam ram_block1a84.mem_init0 = "7E07E03F03F03F03F81F81F81FC0FC0FC0FE07E07E03F03F03F81F81F80FC0FC07E07E03F03F03F81F80FC0FC07E07E03F03F81F81FC0FC07E07F03F01F81FC0FC07E07F03F01F80FC0FE07E03F01F81FC0FE07E03F01F80FC0FE07F03F81FC0FC07E03F01F80FC07E03F01F80FC07E03F01F80FE07F03F81FC0FE03F01F80FC07F03F81FC07E03F01FC0FE03F01FC0FE03F01FC0FE03F01FC0FE03F01FC07E03F81FC07F03F80FE07F01FC07E03F80FE07F01FC07E03F80FE03F01FC07F01FC0FE03F80FE03F80FE07F01FC07F01FC07F01FC07F01FC07F01FC07F01FC07F01FC07F01FC07F01FC07F01FE03F80FE03F80FE01FC07F01FC07F80FE03F807F01";

arriav_ram_block ram_block1a100(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a100_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a100.clk0_core_clock_enable = "ena0";
defparam ram_block1a100.clk0_input_clock_enable = "ena0";
defparam ram_block1a100.clk0_output_clock_enable = "ena0";
defparam ram_block1a100.data_interleave_offset_in_bits = 1;
defparam ram_block1a100.data_interleave_width_in_bits = 1;
defparam ram_block1a100.init_file = "DDS_48_v1_nco_ii_0_cos.hex";
defparam ram_block1a100.init_file_layout = "port_a";
defparam ram_block1a100.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0121|altsyncram:altsyncram_component0|altsyncram_78g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a100.operation_mode = "rom";
defparam ram_block1a100.port_a_address_clear = "none";
defparam ram_block1a100.port_a_address_width = 13;
defparam ram_block1a100.port_a_data_out_clear = "none";
defparam ram_block1a100.port_a_data_out_clock = "clock0";
defparam ram_block1a100.port_a_data_width = 1;
defparam ram_block1a100.port_a_first_address = 49152;
defparam ram_block1a100.port_a_first_bit_number = 4;
defparam ram_block1a100.port_a_last_address = 57343;
defparam ram_block1a100.port_a_logical_ram_depth = 65536;
defparam ram_block1a100.port_a_logical_ram_width = 16;
defparam ram_block1a100.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a100.ram_block_type = "auto";
defparam ram_block1a100.mem_init3 = "7F01FC07F00FE03F80FE01FC07F01FC07F00FE03F80FE03F80FE03F807F01FC07F01FC07F01FC07F01FC07F01FC07F01F80FE03F80FE03F80FE03F81FC07F01FC07F03F80FE03F80FC07F01FC0FE03F80FC07F01FC0FE03F81FC07F03F80FE07F01FC0FE03F01FC0FE03F81FC07E03F81FC07E03F01FC0FE03F01F80FE07F03F80FC07E03F01FC0FE07F03F81FC07E03F01F80FC07E03F01F80FC07E03F03F81FC0FE07F03F81F80FC07E03F03F81FC0FC07E03F03F81F80FC07E07F03F01F81FC0FC07E07F03F01F81FC0FC07E07E03F03F81F81FC0FC0FE07E07F03F03F81F81FC0FC0FC07E07E07F03F03F01F81F81F80FC0FC0FC07E07E07E03F03F03F03";
defparam ram_block1a100.mem_init2 = "F01F81F81F81F81FC0FC0FC0FC0FC0FC0FE07E07E07E07E07E07E07E07E07E03F03F03F03F03F03F03F03F03F03F03F03F03F03F07E07E07E07E07E07E07E07E07E07E0FC0FC0FC0FC0FC0FC1F81F81F81F81F83F03F03F03F07E07E07E07C0FC0FC0FC1F81F81F83F03F03F07E07E07C0FC0FC0F81F81F83F03F07E07E07C0FC0F81F81F83F03F07E07E0FC0FC1F81F83F03F07E07C0FC0F81F83F03F07E07C0FC0F81F83F03E07E0FC0F81F83F03E07E0FC0F81F83F03E07E0FC0F81F83F07E07C0FC1F83F03E07E0FC1F81F03E07E0FC1F81F03E07E0FC1F81F03E07C0FC1F83F07E07C0F81F03E07E0FC1F83F07E0FC0F81F03E07C0F81F03E07E0FC1F83";
defparam ram_block1a100.mem_init1 = "F07E0FC1F83F07E0FC1F83F07E0FC1F83F07E0F81F03E07C0F81F03E07C0F83F07E0FC1F83F07C0F81F03E07C1F83F07E0F81F03E07C1F83F07E0F81F03E0FC1F83F07C0F81F07E0FC1F03E0FC1F83E07C0F83F07E0F81F07E0FC1F03E0FC1F03E07C1F83E07C1F83E07C0F83F07C0F83F07C0F83F07C0F83F07C0F83F07C0F83F07C0F83E07C1F83E07C1F83E07C1F03E0FC1F03E0F81F07E0F83F07C0F83E07C1F83E0FC1F03E0F81F07E0F83F07C1F83E0FC1F03E0F81F07C0F83E07C1F03E0F81F07C0F83E07C1F03E0F83F07C1F83E0FC1F07E0F83E07C1F03E0F83F07C1F83E0F81F07C0F83E0FC1F07C0F83E0FC1F07C0F83E0FC1F07C0F83E0FC1F07";
defparam ram_block1a100.mem_init0 = "C0F83E0FC1F07C0F83E0F81F07C1F83E0F83F07C1F03E0F83E07C1F07C0F83E0F81F07C1F03E0F83E07C1F07C0F83E0F81F07C1F07E0F83E0FC1F07C1F03E0F83E07C1F07C1F83E0F83E07C1F07C1F83E0F83E07C1F07C1F03E0F83E0FC1F07C1F07E0F83E0F83F07C1F07C0F83E0F83E07C1F07C1F07E0F83E0F83F07C1F07C1F83E0F83E0F81F07C1F07C1F83E0F83E0F81F07C1F07C1F83E0F83E0F81F07C1F07C1F83E0F83E0F83F07C1F07C1F03E0F83E0F83E07C1F07C1F07C0F83E0F83E0F81F07C1F07C1F03E0F83E0F83E0FC1F07C1F07C1F83E0F83E0F83F07C1F07C1F07C0F83E0F83E0F83F07C1F07C1F07E0F83E0F83E0F81F07C1F07C1F07E0";

arriav_ram_block ram_block1a116(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a116_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a116.clk0_core_clock_enable = "ena0";
defparam ram_block1a116.clk0_input_clock_enable = "ena0";
defparam ram_block1a116.clk0_output_clock_enable = "ena0";
defparam ram_block1a116.data_interleave_offset_in_bits = 1;
defparam ram_block1a116.data_interleave_width_in_bits = 1;
defparam ram_block1a116.init_file = "DDS_48_v1_nco_ii_0_cos.hex";
defparam ram_block1a116.init_file_layout = "port_a";
defparam ram_block1a116.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0121|altsyncram:altsyncram_component0|altsyncram_78g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a116.operation_mode = "rom";
defparam ram_block1a116.port_a_address_clear = "none";
defparam ram_block1a116.port_a_address_width = 13;
defparam ram_block1a116.port_a_data_out_clear = "none";
defparam ram_block1a116.port_a_data_out_clock = "clock0";
defparam ram_block1a116.port_a_data_width = 1;
defparam ram_block1a116.port_a_first_address = 57344;
defparam ram_block1a116.port_a_first_bit_number = 4;
defparam ram_block1a116.port_a_last_address = 65535;
defparam ram_block1a116.port_a_logical_ram_depth = 65536;
defparam ram_block1a116.port_a_logical_ram_width = 16;
defparam ram_block1a116.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a116.ram_block_type = "auto";
defparam ram_block1a116.mem_init3 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000007FFFFFFFFFFFFFFFFFFC00000000000000000FFFFFFFFFFFFFFFF000000000000000FFFFFFFFFFFFFF00000000000007FFFFFFFFFFFF000000000000FFFFFFFFFFFC00000000003FFFFFFFFFF80000000001FFFFFFFFFE0000000003FFFFFFFFF0000000007FFFFFFFF8000000007FFFFFFFE000000007FFFFFFFC00000003FFFFFFFC00000007FFFFFFF00000003FFFFFFF00000007FFFFFFC0000003FFFFFFC0000007FFFFFF0000001FFFFFFC00";
defparam ram_block1a116.mem_init2 = "0000FFFFFF8000001FFFFFF0000007FFFFF8000003FFFFFC000007FFFFF800000FFFFFE000003FFFFF800001FFFFFC00000FFFFF800001FFFFF800003FFFFE00000FFFFF800007FFFFC00003FFFFC00003FFFFC00003FFFF800007FFFF00001FFFFC00007FFFF00001FFFF80000FFFFC00007FFFE00007FFFE0000FFFFC0000FFFF80001FFFF00007FFFC0001FFFF00007FFFC0001FFFE0000FFFF00007FFF80007FFF80003FFFC0007FFF80007FFF80007FFF0000FFFE0003FFFC0007FFF0001FFFC0007FFF0001FFFC0007FFF0003FFF8001FFFC000FFFE0007FFE0003FFF0003FFF0003FFF0003FFF0003FFF0007FFE0007FFC000FFF8001FFF0003FFE000";
defparam ram_block1a116.mem_init1 = "7FFC001FFF0007FFE000FFF8003FFE000FFF8007FFC001FFF000FFF8003FFC001FFF000FFF0007FF8003FFC003FFE001FFE001FFE000FFF000FFF000FFF000FFF001FFE001FFE001FFE003FFC003FF8007FF000FFF001FFE003FF8007FF000FFE003FF8007FF001FFC003FF800FFE003FF800FFE003FF800FFE003FF801FFC007FF001FF800FFE003FF001FFC00FFE007FF003FF801FFC00FFE007FF003FF001FF801FFC00FFC00FFE007FE007FE007FE003FF003FF003FF003FF003FF003FF007FE007FE007FE007FC00FFC00FF801FF801FF003FF007FE00FFC00FF801FF003FE007FC00FF801FF007FE00FFC01FF003FE00FFC01FF007FE00FF803FF007FC";
defparam ram_block1a116.mem_init0 = "01FF007FE00FF803FE00FF803FE00FF803FE00FF803FE00FF803FE00FF007FC01FF007F803FE00FF807FC01FF00FF803FC01FF00FF803FC01FF00FF807FC01FE00FF007F803FC01FE00FF007F807FC03FE01FE00FF007F807FC03FC01FE01FE00FF00FF807F807F803FC03FC03FE01FE01FE01FE00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FE01FE01FE01FE03FC03FC03FC07F807F80FF00FF01FE01FE03FC03F807F807F00FF01FE03FC03F807F80FF01FE01FC03F807F00FE01FC03F807F00FE01FC03F807F00FE01FC07F80FF01FE03F807F01FE03FC07F00FE03FC07F01FE03F807F01FC03F80FE01FC07F00FE03F80";

arriav_ram_block ram_block1a36(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a36_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a36.clk0_core_clock_enable = "ena0";
defparam ram_block1a36.clk0_input_clock_enable = "ena0";
defparam ram_block1a36.clk0_output_clock_enable = "ena0";
defparam ram_block1a36.data_interleave_offset_in_bits = 1;
defparam ram_block1a36.data_interleave_width_in_bits = 1;
defparam ram_block1a36.init_file = "DDS_48_v1_nco_ii_0_cos.hex";
defparam ram_block1a36.init_file_layout = "port_a";
defparam ram_block1a36.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0121|altsyncram:altsyncram_component0|altsyncram_78g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a36.operation_mode = "rom";
defparam ram_block1a36.port_a_address_clear = "none";
defparam ram_block1a36.port_a_address_width = 13;
defparam ram_block1a36.port_a_data_out_clear = "none";
defparam ram_block1a36.port_a_data_out_clock = "clock0";
defparam ram_block1a36.port_a_data_width = 1;
defparam ram_block1a36.port_a_first_address = 16384;
defparam ram_block1a36.port_a_first_bit_number = 4;
defparam ram_block1a36.port_a_last_address = 24575;
defparam ram_block1a36.port_a_logical_ram_depth = 65536;
defparam ram_block1a36.port_a_logical_ram_width = 16;
defparam ram_block1a36.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a36.ram_block_type = "auto";
defparam ram_block1a36.mem_init3 = "01FC03F80FE03FC07F01FC07F00FE03F80FE03F80FF01FC07F01FC07F01FC07F01FC07F01FC07F01FC07F01FC07F01FC07F01FC07F01FC0FE03F80FE03F80FE07F01FC07F01F80FE03F80FC07F01FC0FE03F80FC07F01FC0FE03F81FC07F03F80FC07F01F80FE07F01F80FE07F01F80FE07F01F80FE07F01F80FC07F03F81FC07E03F01F80FE07F03F81FC0FE03F01F80FC07E03F01F80FC07E03F01F80FC07E07F03F81FC0FE07E03F01F80FC0FE07F03F01F80FC0FE07E03F01F81FC0FC07E07F03F01F81FC0FC07E07F03F03F81F80FC0FC07E07E03F03F81F81F80FC0FC07E07E03F03F03F81F81F80FC0FC0FE07E07E07F03F03F03F81F81F81F80FC0FC";
defparam ram_block1a36.mem_init2 = "0FC0FC07E07E07E07E07E03F03F03F03F03F03F03F81F81F81F81F81F81F81F81F81F81F81F81F81F81F81F81F81F81F81F81F81F81F81F81F81F81F81F81F03F03F03F03F03F03F03E07E07E07E07E07C0FC0FC0FC0FC1F81F81F81F83F03F03F03E07E07E07C0FC0FC0F81F81F83F03F03F07E07E07C0FC0FC1F81F83F03F03E07E07C0FC0F81F81F83F03E07E07C0FC0F81F81F03F03E07E0FC0FC1F81F03F07E07E0FC0F81F83F03E07E0FC0F81F83F03E07E0FC0F81F83F03E07E0FC1F81F03F07E07C0F81F83F07E07C0FC1F83F03E07C0FC1F83F07E07C0F81F83F07E0FC0F81F03E07C0FC1F83F07E0FC0F81F03E07C0F81F03E07E0FC1F83F07E0FC";
defparam ram_block1a36.mem_init1 = "1F83F07E0FC1F83F07E0FC1F83F07E0FC1F83F07E0FC1F83E07C0F81F03E07C0F83F07E0FC1F83F07C0F81F03E07C1F83F07E0F81F03E07C1F83F07C0F81F03E0FC1F83E07C0F83F07E0F81F03E0FC1F03E07C1F83F07C0F83F07E0F81F07E0F81F03E0FC1F03E0FC1F03E07C1F83E07C1F83E07C1F83E07C1F83E07C1F83E07C1F83E07C1F03E0FC1F03E0FC1F07E0F81F07E0F81F07C0F83F07C1F83E07C1F03E0FC1F07E0F81F07C0F83E07C1F83E0FC1F07E0F83F07C1F83E07C1F03E0F81F07C0F83E07C1F07E0F83F07C1F83E0FC1F07E0F83E07C1F03E0F83F07C1F83E0F81F07C0F83E0FC1F07C0F83E07C1F07E0F83E07C1F07E0F83E07C1F07E0F8";
defparam ram_block1a36.mem_init0 = "3E0FC1F07C0F83E0FC1F07C1F83E0F81F07C1F03E0F83F07C1F07E0F83E0FC1F07C1F83E0F83F07C1F07E0F83E0FC1F07C1F83E0F83E07C1F07C0F83E0F83F07C1F07C0F83E0F83F07C1F07E0F83E0F83F07C1F07C0F83E0F83F07C1F07C1F83E0F83E07C1F07C1F03E0F83E0F81F07C1F07C0F83E0F83E07C1F07C1F03E0F83E0F83F07C1F07C1F03E0F83E0F81F07C1F07C1F83E0F83E0F81F07C1F07C1F03E0F83E0F83F07C1F07C1F07E0F83E0F83E07C1F07C1F07C0F83E0F83E0F81F07C1F07C1F03E0F83E0F83E0FC1F07C1F07C1F83E0F83E0F83F07C1F07C1F07C0F83E0F83E0F81F07C1F07C1F07E0F83E0F83E0F81F07C1F07C1F03E0F83E0F83E";

arriav_ram_block ram_block1a52(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a52_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a52.clk0_core_clock_enable = "ena0";
defparam ram_block1a52.clk0_input_clock_enable = "ena0";
defparam ram_block1a52.clk0_output_clock_enable = "ena0";
defparam ram_block1a52.data_interleave_offset_in_bits = 1;
defparam ram_block1a52.data_interleave_width_in_bits = 1;
defparam ram_block1a52.init_file = "DDS_48_v1_nco_ii_0_cos.hex";
defparam ram_block1a52.init_file_layout = "port_a";
defparam ram_block1a52.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0121|altsyncram:altsyncram_component0|altsyncram_78g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a52.operation_mode = "rom";
defparam ram_block1a52.port_a_address_clear = "none";
defparam ram_block1a52.port_a_address_width = 13;
defparam ram_block1a52.port_a_data_out_clear = "none";
defparam ram_block1a52.port_a_data_out_clock = "clock0";
defparam ram_block1a52.port_a_data_width = 1;
defparam ram_block1a52.port_a_first_address = 24576;
defparam ram_block1a52.port_a_first_bit_number = 4;
defparam ram_block1a52.port_a_last_address = 32767;
defparam ram_block1a52.port_a_logical_ram_depth = 65536;
defparam ram_block1a52.port_a_logical_ram_width = 16;
defparam ram_block1a52.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a52.ram_block_type = "auto";
defparam ram_block1a52.mem_init3 = "000000000000000000000000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000001FFFFFFFFFFFFFFFFFFFFFF00000000000000000003FFFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFF000000000000007FFFFFFFFFFFFC000000000000FFFFFFFFFFFF800000000001FFFFFFFFFFF00000000001FFFFFFFFFF00000000007FFFFFFFFF0000000003FFFFFFFFE000000001FFFFFFFFC000000007FFFFFFFE00000000FFFFFFFF00000000FFFFFFFE00000003FFFFFFF00000003FFFFFFE0000000FFFFFFF0000000FFFFFFF0000001FFFFFF8000000FFF";
defparam ram_block1a52.mem_init2 = "FFFC000000FFFFFF8000003FFFFFE000000FFFFFF000000FFFFFF000000FFFFFE000003FFFFF800000FFFFFC00000FFFFFC00000FFFFFC00001FFFFF800003FFFFE00001FFFFF000007FFFF800007FFFF800007FFFF80000FFFFF00001FFFFC00007FFFF00001FFFFC0000FFFFE00007FFFE00003FFFF00007FFFE00007FFFE0000FFFFC0001FFFF00007FFFC0001FFFF00007FFFC0003FFFE0001FFFF0000FFFF0000FFFF80007FFF0000FFFF0000FFFF0001FFFE0003FFF80007FFF0001FFFC0007FFF0001FFFC0007FFF0001FFF8000FFFE0007FFE0003FFF0001FFF8001FFF8001FFF8001FFF8001FFF8001FFF8003FFF0003FFE0007FFC000FFF8003FFF";
defparam ram_block1a52.mem_init1 = "0007FFC001FFF8003FFE000FFF8003FFE000FFF8007FFC001FFF000FFF8003FFC001FFE000FFF0007FF8007FFC003FFC003FFE001FFE001FFE001FFE001FFE001FFE001FFC003FFC003FF8007FF8007FF000FFE001FFC003FF8007FF001FFE003FF8007FF001FFC003FF800FFE003FF800FFE003FF800FFE003FF800FFE003FF001FFC007FE003FF800FFC007FE003FF801FFC00FFE007FF003FF001FF800FFC00FFE007FE007FF003FF003FF001FF801FF801FF801FF801FF801FF801FF801FF801FF801FF003FF003FF007FE007FE00FFC00FF801FF803FF007FE007FC00FF801FF003FE007FC01FF803FF007FC00FF803FF007FC00FF803FE007FC01FF007";
defparam ram_block1a52.mem_init0 = "FE00FF803FE00FF803FE00FFC01FF007FC01FF007F803FE00FF803FE00FF803FC01FF007FC01FE00FF803FC01FF00FF803FE01FF007F803FC01FF00FF807FC01FE00FF007F803FC01FE00FF00FF807FC03FE01FE00FF00FF807F803FC03FE01FE00FF00FF007F807F807FC03FC03FC03FE01FE01FE01FE01FE00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FE01FE01FE01FE01FE03FC03FC03FC07F807F807F00FF00FE01FE01FC03FC03F807F80FF00FE01FE03FC03F807F00FF01FE03FC03F807F00FE01FC03F807F80FF01FC03F807F00FE01FC03F80FF01FE03F807F00FE03FC07F00FE03FC07F00FE03FC07F01FE03F807F01FC03F80FE03FC07F";

arriav_ram_block ram_block1a4(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a4_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.clk0_input_clock_enable = "ena0";
defparam ram_block1a4.clk0_output_clock_enable = "ena0";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.init_file = "DDS_48_v1_nco_ii_0_cos.hex";
defparam ram_block1a4.init_file_layout = "port_a";
defparam ram_block1a4.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0121|altsyncram:altsyncram_component0|altsyncram_78g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.operation_mode = "rom";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 13;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "clock0";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 8191;
defparam ram_block1a4.port_a_logical_ram_depth = 65536;
defparam ram_block1a4.port_a_logical_ram_width = 16;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.ram_block_type = "auto";
defparam ram_block1a4.mem_init3 = "03F80FE01FC07F00FE03F807F01FC03F80FF01FC07F80FE01FC07F80FF01FC03F80FF01FE03FC07F00FE01FC03F807F00FE01FC03F807F00FE01FC03F807F00FF01FE03FC03F807F80FF01FE01FC03FC03F807F80FF00FF01FE01FE03FC03FC07F807F807F80FF00FF00FF00FE01FE01FE01FE01FE01FE01FE01FE01FE01FE01FE01FE01FE01FE01FE01FE00FF00FF00FF00FF807F807F803FC03FC03FE01FE00FF00FF007F807FC03FC01FE00FF00FF807FC03FC01FE00FF007F803FC01FE00FF007FC03FE01FF007F803FE01FF007F803FE01FF007FC03FE00FF803FC01FF007FC01FE00FF803FE00FF803FE00FF803FE00FF803FE00FF803FE00FFC01FF00";
defparam ram_block1a4.mem_init2 = "7FC01FF803FE00FFC01FF007FE00FF801FF007FE00FFC01FF003FE007FC00FF801FF003FE007FE00FFC01FF801FF003FF003FE007FE007FC00FFC00FFC00FFC01FF801FF801FF801FF801FF801FF800FFC00FFC00FFC00FFE007FE007FF003FF001FF801FFC00FFE007FF003FF801FFC00FFE007FF001FF800FFE003FF001FFC007FF003FF800FFE003FF800FFE003FF800FFE003FF8007FF001FFC003FF800FFE001FFC003FF800FFF001FFE001FFC003FF8007FF800FFF000FFF000FFF001FFE001FFE001FFE001FFE000FFF000FFF000FFF8007FF8003FFC001FFE001FFF0007FF8003FFE001FFF0007FFC003FFE000FFF8003FFE000FFFC001FFF0007FFC";
defparam ram_block1a4.mem_init1 = "000FFF8001FFF0003FFE0007FFC000FFFC001FFF8001FFF8001FFF8001FFF8001FFF8000FFFC000FFFE0007FFF0003FFF8001FFFC0007FFF0001FFFC0007FFF0001FFFC0007FFF8000FFFE0001FFFC0003FFFC0003FFFC0007FFF80003FFFC0003FFFC0001FFFE0000FFFF00007FFFC0001FFFF00007FFFC0001FFFF00003FFFE00007FFFE0000FFFFC0000FFFFC00007FFFE00003FFFF00001FFFFC00007FFFF00001FFFFC00003FFFF800007FFFF800007FFFF800007FFFFC00003FFFFE00000FFFFF800003FFFFF000003FFFFE000007FFFFF000003FFFFF800000FFFFFE000003FFFFFC000007FFFFF8000003FFFFFC000001FFFFFF0000003FFFFFE0000";
defparam ram_block1a4.mem_init0 = "007FFFFFF0000001FFFFFFC0000007FFFFFF80000007FFFFFFC0000001FFFFFFF80000001FFFFFFFC00000007FFFFFFF800000007FFFFFFFC00000000FFFFFFFFC000000003FFFFFFFFC000000001FFFFFFFFF8000000000FFFFFFFFFF00000000003FFFFFFFFFF800000000007FFFFFFFFFFE000000000001FFFFFFFFFFFFC0000000000001FFFFFFFFFFFFFE000000000000001FFFFFFFFFFFFFFFE000000000000000007FFFFFFFFFFFFFFFFFFC0000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

arriav_ram_block ram_block1a20(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a20_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a20.clk0_core_clock_enable = "ena0";
defparam ram_block1a20.clk0_input_clock_enable = "ena0";
defparam ram_block1a20.clk0_output_clock_enable = "ena0";
defparam ram_block1a20.data_interleave_offset_in_bits = 1;
defparam ram_block1a20.data_interleave_width_in_bits = 1;
defparam ram_block1a20.init_file = "DDS_48_v1_nco_ii_0_cos.hex";
defparam ram_block1a20.init_file_layout = "port_a";
defparam ram_block1a20.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0121|altsyncram:altsyncram_component0|altsyncram_78g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a20.operation_mode = "rom";
defparam ram_block1a20.port_a_address_clear = "none";
defparam ram_block1a20.port_a_address_width = 13;
defparam ram_block1a20.port_a_data_out_clear = "none";
defparam ram_block1a20.port_a_data_out_clock = "clock0";
defparam ram_block1a20.port_a_data_width = 1;
defparam ram_block1a20.port_a_first_address = 8192;
defparam ram_block1a20.port_a_first_bit_number = 4;
defparam ram_block1a20.port_a_last_address = 16383;
defparam ram_block1a20.port_a_logical_ram_depth = 65536;
defparam ram_block1a20.port_a_logical_ram_width = 16;
defparam ram_block1a20.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a20.ram_block_type = "auto";
defparam ram_block1a20.mem_init3 = "0FC1F07C1F07C1F03E0F83E0F83E0FC1F07C1F07C1F83E0F83E0F83E07C1F07C1F07C1F83E0F83E0F83F07C1F07C1F07E0F83E0F83E0F81F07C1F07C1F03E0F83E0F83E07C1F07C1F07C0F83E0F83E0F81F07C1F07C1F83E0F83E0F83F07C1F07C1F03E0F83E0F83F07C1F07C1F03E0F83E0F83F07C1F07C1F03E0F83E0F83F07C1F07C1F83E0F83E0FC1F07C1F07C0F83E0F83E07C1F07C1F83E0F83E0FC1F07C1F07E0F83E0F81F07C1F07C0F83E0F83F07C1F07C0F83E0F83F07C1F07C0F83E0F81F07C1F07E0F83E0FC1F07C1F03E0F83E07C1F07C0F83E0F81F07C1F03E0F83E07C1F07C0F83E0F81F07C1F83E0F83F07C1F03E0F83E07C1F07E0F83E07";
defparam ram_block1a20.mem_init2 = "C1F07E0F83E07C1F07E0F83E07C1F07E0F83E07C1F07E0F83E07C1F03E0F83F07C1F83E0F81F07C0F83E0FC1F07E0F83F07C1F83E0F81F07C0F83E07C1F03E0F81F07C0F83E07C1F03E0F81F07E0F83F07C1F83E0FC1F03E0F81F07E0F83F07C0F83E07C1F83E0FC1F03E0F81F07E0F81F07C0F83F07C0F83F07C0F83E07C1F83E07C1F83E07C1F83E07C1F83E07C1F83E07C1F83E07C0F83F07C0F83F07C0F81F07E0F81F07E0FC1F03E0FC1F83E07C0F83F07E0F81F07E0FC1F03E07C1F83F07E0F81F03E0FC1F83F07C0F81F03E0FC1F83F07C0F81F03E07C1F83F07E0FC1F83E07C0F81F03E07C0F81F03E0FC1F83F07E0FC1F83F07E0FC1F83F07E0FC1F";
defparam ram_block1a20.mem_init1 = "83F07E0FC0F81F03E07C0F81F03E07E0FC1F83F07E0FC0F81F03E07C0FC1F83F07E07C0F81F03F07E0FC0F81F03F07E0FC0F81F03F07E0FC0F81F83F07E07C0FC1F83F03E07E0FC0F81F83F03E07E0FC0F81F83F03E07E0FC0F81F83F03E07E07C0FC1F81F83F03E07E07C0FC1F81F83F03F07E07E0FC0FC1F81F83F03F03E07E07C0FC0FC1F81F83F03F03E07E07E07C0FC0FC1F81F81F83F03F03F07E07E07E07C0FC0FC0FC1F81F81F81F83F03F03F03F03F07E07E07E07E07E07E0FC0FC0FC0FC0FC0FC0FC0FC0FC0FC1F81F81F81F81F81F81F81F81F81F81F81F81F81F80FC0FC0FC0FC0FC0FC0FC0FC0FC0FE07E07E07E07E07E07F03F03F03F03F01F";
defparam ram_block1a20.mem_init0 = "81F81F81F80FC0FC0FC07E07E07E03F03F03F01F81F81FC0FC0FC07E07E07F03F03F81F81FC0FC0FE07E07F03F03F81F80FC0FC07E07F03F01F81FC0FC07E07F03F01F81FC0FC07E03F03F81F80FC07E07F03F81F80FC07E03F03F81FC0FE07F03F81F80FC07E03F01F80FC07E03F01F80FC07F03F81FC0FE07F01F80FC07E03F81FC0FE03F01F80FE07F01F80FC07F03F80FC07F03F80FE07F01F80FE07F01FC0FE03F81FC07F03F80FE07F01FC07E03F80FE07F01FC07E03F80FE03F81FC07F01FC07F03F80FE03F80FE03F80FE03F01FC07F01FC07F01FC07F01FC07F01FC07F01FC03F80FE03F80FE03F80FE01FC07F01FC07F00FE03F80FE01FC07F01FC";

arriav_ram_block ram_block1a69(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a69_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a69.clk0_core_clock_enable = "ena0";
defparam ram_block1a69.clk0_input_clock_enable = "ena0";
defparam ram_block1a69.clk0_output_clock_enable = "ena0";
defparam ram_block1a69.data_interleave_offset_in_bits = 1;
defparam ram_block1a69.data_interleave_width_in_bits = 1;
defparam ram_block1a69.init_file = "DDS_48_v1_nco_ii_0_cos.hex";
defparam ram_block1a69.init_file_layout = "port_a";
defparam ram_block1a69.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0121|altsyncram:altsyncram_component0|altsyncram_78g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a69.operation_mode = "rom";
defparam ram_block1a69.port_a_address_clear = "none";
defparam ram_block1a69.port_a_address_width = 13;
defparam ram_block1a69.port_a_data_out_clear = "none";
defparam ram_block1a69.port_a_data_out_clock = "clock0";
defparam ram_block1a69.port_a_data_width = 1;
defparam ram_block1a69.port_a_first_address = 32768;
defparam ram_block1a69.port_a_first_bit_number = 5;
defparam ram_block1a69.port_a_last_address = 40959;
defparam ram_block1a69.port_a_logical_ram_depth = 65536;
defparam ram_block1a69.port_a_logical_ram_width = 16;
defparam ram_block1a69.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a69.ram_block_type = "auto";
defparam ram_block1a69.mem_init3 = "FFF8000FFFC0007FFE0003FFF0001FFF8000FFFE0007FFF0001FFF8000FFFE0003FFF0001FFFC0007FFF0001FFFC0007FFE0003FFFC0007FFF0001FFFC0007FFF0001FFFE0003FFF8000FFFF0001FFFC0003FFF80007FFF0000FFFE0001FFFC0003FFF80007FFF8000FFFF0000FFFF0000FFFE0001FFFE0001FFFE0001FFFE0001FFFE0001FFFF0000FFFF0000FFFF00007FFF80007FFFC0003FFFE0001FFFF0000FFFF80003FFFC0001FFFF0000FFFF80003FFFE0000FFFF80003FFFE0000FFFF80003FFFE00007FFFC0001FFFF00003FFFE00007FFFC0000FFFF80001FFFF80003FFFF00003FFFF00003FFFE00007FFFE00007FFFF00003FFFF00003FFFF00";
defparam ram_block1a69.mem_init2 = "001FFFF80000FFFFC00007FFFE00003FFFF80001FFFFC00007FFFF00001FFFFC00007FFFF00001FFFFC00003FFFF80000FFFFF00001FFFFE00001FFFFC00003FFFFC00003FFFFC00003FFFFC00003FFFFC00001FFFFE00001FFFFF00000FFFFF800003FFFFE00001FFFFF000007FFFFC00000FFFFF800003FFFFF000007FFFFE00000FFFFFC00000FFFFFC00000FFFFFC00000FFFFFC000007FFFFE000003FFFFF000001FFFFFC000007FFFFF000001FFFFFC000003FFFFF8000007FFFFF000000FFFFFF000000FFFFFF000000FFFFFF8000007FFFFFC000001FFFFFF0000007FFFFFC000001FFFFFF8000003FFFFFF0000003FFFFFF0000003FFFFFF8000001";
defparam ram_block1a69.mem_init1 = "FFFFFFC0000007FFFFFF0000001FFFFFFC0000003FFFFFFC0000003FFFFFFC0000003FFFFFFE0000000FFFFFFF00000003FFFFFFE00000007FFFFFFE00000007FFFFFFE00000003FFFFFFF00000001FFFFFFFE00000001FFFFFFFC00000001FFFFFFFE00000000FFFFFFFF800000001FFFFFFFF800000001FFFFFFFF800000000FFFFFFFFF000000001FFFFFFFFF000000000FFFFFFFFF8000000001FFFFFFFFF8000000001FFFFFFFFFC0000000003FFFFFFFFFC0000000001FFFFFFFFFF00000000003FFFFFFFFFF800000000007FFFFFFFFFF800000000003FFFFFFFFFFF000000000001FFFFFFFFFFFE000000000000FFFFFFFFFFFFC0000000000007FFF";
defparam ram_block1a69.mem_init0 = "FFFFFFFFFC0000000000001FFFFFFFFFFFFFE00000000000000FFFFFFFFFFFFFFE000000000000000FFFFFFFFFFFFFFFE0000000000000000FFFFFFFFFFFFFFFFF800000000000000000FFFFFFFFFFFFFFFFFFE00000000000000000001FFFFFFFFFFFFFFFFFFFFE00000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

arriav_ram_block ram_block1a85(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a85_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a85.clk0_core_clock_enable = "ena0";
defparam ram_block1a85.clk0_input_clock_enable = "ena0";
defparam ram_block1a85.clk0_output_clock_enable = "ena0";
defparam ram_block1a85.data_interleave_offset_in_bits = 1;
defparam ram_block1a85.data_interleave_width_in_bits = 1;
defparam ram_block1a85.init_file = "DDS_48_v1_nco_ii_0_cos.hex";
defparam ram_block1a85.init_file_layout = "port_a";
defparam ram_block1a85.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0121|altsyncram:altsyncram_component0|altsyncram_78g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a85.operation_mode = "rom";
defparam ram_block1a85.port_a_address_clear = "none";
defparam ram_block1a85.port_a_address_width = 13;
defparam ram_block1a85.port_a_data_out_clear = "none";
defparam ram_block1a85.port_a_data_out_clock = "clock0";
defparam ram_block1a85.port_a_data_width = 1;
defparam ram_block1a85.port_a_first_address = 40960;
defparam ram_block1a85.port_a_first_bit_number = 5;
defparam ram_block1a85.port_a_last_address = 49151;
defparam ram_block1a85.port_a_logical_ram_depth = 65536;
defparam ram_block1a85.port_a_logical_ram_width = 16;
defparam ram_block1a85.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a85.ram_block_type = "auto";
defparam ram_block1a85.mem_init3 = "FFC00FFC00FFE007FE007FE003FF003FF003FF001FF801FF801FFC00FFC00FFC007FE007FE007FE003FF003FF003FF801FF801FF800FFC00FFC00FFE007FE007FE003FF003FF003FF801FF801FF800FFC00FFC00FFE007FE007FE003FF003FF001FF801FF801FFC00FFC00FFC007FE007FE003FF003FF001FF801FF801FFC00FFC00FFE007FE007FF003FF003FF801FF801FFC00FFC00FFE007FE007FF003FF003FF801FF801FFC00FFC007FE007FE003FF003FF001FF801FFC00FFC007FE007FE003FF003FF801FF800FFC00FFC007FE007FF003FF001FF801FFC00FFC007FE007FF003FF001FF801FFC00FFE007FE003FF003FF801FF800FFC007FE007FF00";
defparam ram_block1a85.mem_init2 = "3FF001FF800FFC00FFE007FF003FF001FF800FFC007FE007FF003FF801FFC00FFC007FE003FF001FF800FFC00FFE007FF003FF801FFC00FFE007FF003FF801FFC00FFE007FF003FF801FFC00FFE007FF003FF800FFC007FE003FF001FF800FFE007FF003FF801FFC007FE003FF001FFC00FFE007FF001FF800FFE007FF003FF800FFC007FF003FF800FFC007FF003FF800FFC007FF001FF800FFE007FF001FFC00FFE003FF001FFC007FE003FF800FFE007FF001FFC00FFE003FF800FFC007FF001FFC007FE003FF800FFE003FF001FFC007FF001FFC007FE003FF800FFE003FF800FFE003FF800FFC007FF001FFC007FF001FFC007FF001FFC007FF001FFC00";
defparam ram_block1a85.mem_init1 = "7FF001FFC007FF000FFE003FF800FFE003FF800FFE003FF8007FF001FFC007FF001FFC003FF800FFE003FF8007FF001FFC007FF800FFE003FFC007FF001FFE003FF800FFF001FFC003FF800FFF001FFC003FF800FFF001FFC003FF800FFF001FFE003FF8007FF000FFE001FFC003FF8007FF000FFE003FFC003FF8007FF000FFE001FFC003FF8007FF800FFF001FFE001FFC003FFC007FF8007FF000FFF001FFE001FFC003FFC003FF8007FF8007FF800FFF000FFF000FFE001FFE001FFE001FFE003FFC003FFC003FFC003FFC003FFC003FFC003FFC003FFC003FFC003FFC003FFC003FFC003FFC003FFC001FFE001FFE001FFE000FFF000FFF000FFF8007FF";
defparam ram_block1a85.mem_init0 = "8007FFC003FFC003FFE001FFE000FFF000FFF8007FFC003FFC001FFE000FFF0007FF8003FFC003FFE000FFF0007FF8003FFC001FFE000FFF8007FFC001FFE000FFF8007FFC001FFF000FFF8003FFE001FFF0007FFC001FFF000FFF8003FFE000FFF8003FFE000FFF8003FFE000FFF8003FFE000FFF8003FFE000FFFC001FFF0007FFC001FFF8003FFE000FFFC001FFF0003FFE000FFFC001FFF0003FFE0007FFC001FFF8003FFF0007FFE0007FFC000FFF8001FFF8003FFF0003FFE0007FFE000FFFC000FFFC000FFF8001FFF8001FFF8001FFF8001FFF8001FFF8001FFF8001FFF8001FFF8001FFF8001FFFC000FFFC000FFFE0007FFE0007FFF0003FFF8001";

arriav_ram_block ram_block1a101(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a101_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a101.clk0_core_clock_enable = "ena0";
defparam ram_block1a101.clk0_input_clock_enable = "ena0";
defparam ram_block1a101.clk0_output_clock_enable = "ena0";
defparam ram_block1a101.data_interleave_offset_in_bits = 1;
defparam ram_block1a101.data_interleave_width_in_bits = 1;
defparam ram_block1a101.init_file = "DDS_48_v1_nco_ii_0_cos.hex";
defparam ram_block1a101.init_file_layout = "port_a";
defparam ram_block1a101.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0121|altsyncram:altsyncram_component0|altsyncram_78g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a101.operation_mode = "rom";
defparam ram_block1a101.port_a_address_clear = "none";
defparam ram_block1a101.port_a_address_width = 13;
defparam ram_block1a101.port_a_data_out_clear = "none";
defparam ram_block1a101.port_a_data_out_clock = "clock0";
defparam ram_block1a101.port_a_data_width = 1;
defparam ram_block1a101.port_a_first_address = 49152;
defparam ram_block1a101.port_a_first_bit_number = 5;
defparam ram_block1a101.port_a_last_address = 57343;
defparam ram_block1a101.port_a_logical_ram_depth = 65536;
defparam ram_block1a101.port_a_logical_ram_width = 16;
defparam ram_block1a101.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a101.ram_block_type = "auto";
defparam ram_block1a101.mem_init3 = "7FFE0007FFF0003FFF0001FFF8001FFF8000FFFC000FFFC000FFFC0007FFE0007FFE0007FFE0007FFE0007FFE0007FFE000FFFC000FFFC000FFFC001FFF8001FFF8003FFF0003FFF0007FFE000FFFC000FFF8001FFF0003FFE0007FFC000FFF8001FFF0003FFE000FFFC001FFF8003FFE0007FFC001FFF0003FFE000FFF8003FFF0007FFC001FFF0007FFC001FFF8003FFE000FFF8003FFE000FFF8003FFC001FFF0007FFC001FFF0007FFC003FFE000FFF8003FFC001FFF0007FF8003FFE001FFF0007FF8003FFE001FFF0007FF8003FFC001FFE000FFF0007FF8003FFC001FFE000FFF0007FF8007FFC003FFE001FFE000FFF000FFF8007FF8003FFC003FFC";
defparam ram_block1a101.mem_init2 = "001FFE001FFE001FFF000FFF000FFF000FFF8007FF8007FF8007FF8007FF8003FFC003FFC003FFC003FFC003FFC003FFC003FFC007FF8007FF8007FF8007FF8007FF800FFF000FFF000FFF001FFE001FFE001FFC003FFC003FF8007FF8007FF000FFF001FFE001FFC003FFC007FF8007FF000FFF001FFE003FFC007FF8007FF000FFE001FFC003FF8007FF000FFE001FFC003FF8007FF000FFE003FFC007FF800FFF001FFC003FF800FFF001FFC003FF800FFF001FFC003FF800FFF001FFC007FF800FFE003FFC007FF001FFE003FF800FFE001FFC007FF001FFE003FF800FFE003FF8007FF001FFC007FF001FFC007FF000FFE003FF800FFE003FF800FFE003";
defparam ram_block1a101.mem_init1 = "FF800FFE003FF800FFE003FF800FFE003FF800FFE003FF800FFE003FF800FFC007FF001FFC007FF001FFC007FE003FF800FFE003FF801FFC007FF001FFC00FFE003FF800FFE007FF001FFC00FFE003FF800FFC007FF001FF800FFE003FF001FFC007FE003FF801FFC007FF003FF800FFC007FF003FF800FFC007FF003FF800FFC007FF003FF801FFC007FE003FF801FFC00FFE003FF001FF800FFC007FF003FF801FFC00FFE003FF001FF800FFC007FE003FF001FFC00FFE007FF003FF801FFC00FFE007FF003FF801FFC00FFC007FE003FF001FF800FFC007FE003FF003FF801FFC00FFE007FF003FF001FF800FFC00FFE007FF003FF001FF800FFC00FFE007";
defparam ram_block1a101.mem_init0 = "FF003FF001FF800FFC00FFE007FE003FF003FF801FFC00FFC007FE007FF003FF001FF801FFC00FFC007FE007FF003FF001FF801FF800FFC00FFE007FE003FF003FF801FF801FFC00FFC007FE007FE003FF003FF801FF801FFC00FFC00FFE007FE007FF003FF003FF801FF800FFC00FFC007FE007FE007FF003FF003FF801FF801FFC00FFC00FFE007FE007FE003FF003FF001FF801FF801FFC00FFC00FFE007FE007FE003FF003FF003FF801FF801FFC00FFC00FFC007FE007FE007FF003FF003FF001FF801FF801FFC00FFC00FFC00FFE007FE007FE003FF003FF003FF801FF801FF800FFC00FFC00FFC007FE007FE007FF003FF003FF001FF801FF801FF800";

arriav_ram_block ram_block1a117(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a117_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a117.clk0_core_clock_enable = "ena0";
defparam ram_block1a117.clk0_input_clock_enable = "ena0";
defparam ram_block1a117.clk0_output_clock_enable = "ena0";
defparam ram_block1a117.data_interleave_offset_in_bits = 1;
defparam ram_block1a117.data_interleave_width_in_bits = 1;
defparam ram_block1a117.init_file = "DDS_48_v1_nco_ii_0_cos.hex";
defparam ram_block1a117.init_file_layout = "port_a";
defparam ram_block1a117.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0121|altsyncram:altsyncram_component0|altsyncram_78g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a117.operation_mode = "rom";
defparam ram_block1a117.port_a_address_clear = "none";
defparam ram_block1a117.port_a_address_width = 13;
defparam ram_block1a117.port_a_data_out_clear = "none";
defparam ram_block1a117.port_a_data_out_clock = "clock0";
defparam ram_block1a117.port_a_data_width = 1;
defparam ram_block1a117.port_a_first_address = 57344;
defparam ram_block1a117.port_a_first_bit_number = 5;
defparam ram_block1a117.port_a_last_address = 65535;
defparam ram_block1a117.port_a_logical_ram_depth = 65536;
defparam ram_block1a117.port_a_logical_ram_width = 16;
defparam ram_block1a117.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a117.ram_block_type = "auto";
defparam ram_block1a117.mem_init3 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFC000000000000000000001FFFFFFFFFFFFFFFFFFFC0000000000000000007FFFFFFFFFFFFFFFFF800000000000000007FFFFFFFFFFFFFFFC0000000000000007FFFFFFFFFFFFFFC000000000000007FFFFFFFFFFFFFC00000000000007FFFFFFFFFFFFE000000000";
defparam ram_block1a117.mem_init2 = "0000FFFFFFFFFFFFE0000000000007FFFFFFFFFFFC000000000007FFFFFFFFFFF000000000003FFFFFFFFFFE00000000000FFFFFFFFFFE00000000003FFFFFFFFFF00000000007FFFFFFFFFC0000000003FFFFFFFFFC0000000007FFFFFFFFE0000000007FFFFFFFFE000000000FFFFFFFFF8000000007FFFFFFFF000000000FFFFFFFFE000000007FFFFFFFE000000007FFFFFFFE00000000FFFFFFFF800000007FFFFFFFC00000007FFFFFFF800000007FFFFFFF00000003FFFFFFF80000001FFFFFFF80000001FFFFFFF80000003FFFFFFE0000000FFFFFFF80000003FFFFFFC0000003FFFFFFC0000003FFFFFF80000007FFFFFF0000001FFFFFFC000000";
defparam ram_block1a117.mem_init1 = "7FFFFFE0000007FFFFFF0000003FFFFFF0000007FFFFFE000000FFFFFFC000001FFFFFF0000007FFFFFC000003FFFFFE000001FFFFFF000000FFFFFF000000FFFFFE000001FFFFFE000003FFFFFC000007FFFFF000001FFFFFC000007FFFFF000003FFFFF800001FFFFFC00000FFFFFC00000FFFFFC00000FFFFFC00001FFFFF800001FFFFF000003FFFFE00000FFFFF800003FFFFE00000FFFFF800003FFFFE00001FFFFF00000FFFFF800007FFFF800003FFFFC00003FFFFC00003FFFFC00007FFFF800007FFFF80000FFFFF00001FFFFE00003FFFF80000FFFFF00001FFFFC00007FFFF00001FFFF80000FFFFE00003FFFF00001FFFF80000FFFFC00007FF";
defparam ram_block1a117.mem_init0 = "FE00007FFFF00003FFFF00003FFFF00003FFFF00003FFFF00003FFFF00007FFFE00007FFFC0000FFFF80001FFFF00003FFFE0000FFFFC0001FFFF00007FFFE0000FFFF80003FFFE0000FFFF80007FFFC0001FFFF00007FFF80003FFFE0001FFFF0000FFFF80007FFFC0003FFFC0001FFFE0001FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFE0001FFFE0003FFFC0003FFF80007FFF0000FFFE0001FFFC0003FFF80007FFF0001FFFC0003FFF8000FFFE0001FFFC0007FFF0001FFFC0007FFF0001FFFC0007FFF0001FFF8000FFFE0003FFF8001FFFC0007FFF0003FFF8001FFFC0007FFE0003FFF0001FFF8000FFFC000";

arriav_ram_block ram_block1a37(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a37_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a37.clk0_core_clock_enable = "ena0";
defparam ram_block1a37.clk0_input_clock_enable = "ena0";
defparam ram_block1a37.clk0_output_clock_enable = "ena0";
defparam ram_block1a37.data_interleave_offset_in_bits = 1;
defparam ram_block1a37.data_interleave_width_in_bits = 1;
defparam ram_block1a37.init_file = "DDS_48_v1_nco_ii_0_cos.hex";
defparam ram_block1a37.init_file_layout = "port_a";
defparam ram_block1a37.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0121|altsyncram:altsyncram_component0|altsyncram_78g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a37.operation_mode = "rom";
defparam ram_block1a37.port_a_address_clear = "none";
defparam ram_block1a37.port_a_address_width = 13;
defparam ram_block1a37.port_a_data_out_clear = "none";
defparam ram_block1a37.port_a_data_out_clock = "clock0";
defparam ram_block1a37.port_a_data_width = 1;
defparam ram_block1a37.port_a_first_address = 16384;
defparam ram_block1a37.port_a_first_bit_number = 5;
defparam ram_block1a37.port_a_last_address = 24575;
defparam ram_block1a37.port_a_logical_ram_depth = 65536;
defparam ram_block1a37.port_a_logical_ram_width = 16;
defparam ram_block1a37.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a37.ram_block_type = "auto";
defparam ram_block1a37.mem_init3 = "0003FFF8001FFFC000FFFC000FFFE0007FFE0007FFF0003FFF0003FFF0003FFF0003FFF0003FFF0003FFF0003FFF0003FFF0003FFF0003FFE0007FFE0007FFE000FFFC000FFF8001FFF8003FFF0003FFE0007FFC000FFFC001FFF8003FFF0007FFC000FFF8001FFF0007FFE000FFF8001FFF0007FFE000FFF8003FFF0007FFC001FFF0007FFE000FFF8003FFE000FFF8003FFE000FFF8003FFE000FFF8003FFE000FFF8003FFE001FFF0007FFC001FFF000FFF8003FFE001FFF0007FFC003FFE000FFF0007FFC003FFE000FFF0007FF8003FFC001FFE000FFF8007FF8003FFC001FFE000FFF0007FF8007FFC003FFE001FFE000FFF000FFF8007FF8007FFC003";
defparam ram_block1a37.mem_init2 = "FFC003FFE001FFE001FFE000FFF000FFF000FFF0007FF8007FF8007FF8007FF8007FF8007FF8007FF8007FF8007FF8007FF8007FF8007FF8007FF8007FF800FFF000FFF000FFF000FFE001FFE001FFE003FFC003FFC003FF8007FF8007FF000FFF001FFE001FFC003FFC007FF8007FF000FFF001FFE003FFC003FF8007FF000FFE001FFC003FF8007FF800FFE001FFC003FF8007FF000FFE001FFC003FF800FFF001FFE003FF8007FF001FFE003FF8007FF001FFE003FF8007FF001FFE003FF800FFF001FFC007FF800FFE003FFC007FF001FFC003FF800FFE003FF8007FF001FFC007FF001FFC003FF800FFE003FF800FFE003FF800FFE001FFC007FF001FFC";
defparam ram_block1a37.mem_init1 = "007FF001FFC007FF001FFC007FF001FFC007FF001FFC007FE003FF800FFE003FF800FFE003FF800FFC007FF001FFC007FF001FF800FFE003FF800FFC007FF001FFC007FE003FF800FFE007FF001FFC00FFE003FF800FFC007FF001FF800FFE007FF001FFC00FFE003FF001FFC007FE003FF801FFC007FE003FF801FFC007FE003FF801FFC00FFE003FF001FFC00FFE007FF001FF800FFC007FF003FF801FFC00FFE003FF001FF800FFC007FE003FF801FFC00FFE007FF003FF801FFC00FFE007FF003FF801FFC00FFE007FF003FF801FFC00FFE007FE003FF001FF800FFC007FE007FF003FF801FFC00FFC007FE003FF001FF801FFC00FFE007FE003FF001FF8";
defparam ram_block1a37.mem_init0 = "01FFC00FFC007FE003FF003FF801FF800FFC00FFE007FF003FF001FF801FFC00FFC007FE007FF003FF001FF801FFC00FFC007FE007FE003FF003FF801FF800FFC00FFC007FE007FF003FF001FF801FF800FFC00FFC007FE007FF003FF003FF801FF801FFC00FFC00FFE007FE007FF003FF003FF801FF801FFC00FFC00FFE007FE007FF003FF003FF001FF801FF800FFC00FFC007FE007FE007FF003FF003FF001FF801FF800FFC00FFC00FFE007FE007FE003FF003FF003FF801FF801FF800FFC00FFC00FFE007FE007FE003FF003FF003FF801FF801FF800FFC00FFC00FFC007FE007FE007FF003FF003FF001FF801FF801FF800FFC00FFC00FFE007FE007FE";

arriav_ram_block ram_block1a53(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a53_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a53.clk0_core_clock_enable = "ena0";
defparam ram_block1a53.clk0_input_clock_enable = "ena0";
defparam ram_block1a53.clk0_output_clock_enable = "ena0";
defparam ram_block1a53.data_interleave_offset_in_bits = 1;
defparam ram_block1a53.data_interleave_width_in_bits = 1;
defparam ram_block1a53.init_file = "DDS_48_v1_nco_ii_0_cos.hex";
defparam ram_block1a53.init_file_layout = "port_a";
defparam ram_block1a53.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0121|altsyncram:altsyncram_component0|altsyncram_78g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a53.operation_mode = "rom";
defparam ram_block1a53.port_a_address_clear = "none";
defparam ram_block1a53.port_a_address_width = 13;
defparam ram_block1a53.port_a_data_out_clear = "none";
defparam ram_block1a53.port_a_data_out_clock = "clock0";
defparam ram_block1a53.port_a_data_width = 1;
defparam ram_block1a53.port_a_first_address = 24576;
defparam ram_block1a53.port_a_first_bit_number = 5;
defparam ram_block1a53.port_a_last_address = 32767;
defparam ram_block1a53.port_a_logical_ram_depth = 65536;
defparam ram_block1a53.port_a_logical_ram_width = 16;
defparam ram_block1a53.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a53.ram_block_type = "auto";
defparam ram_block1a53.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000FFFFFFFFFFFFFFFFFFFFF00000000000000000000FFFFFFFFFFFFFFFFFFE000000000000000003FFFFFFFFFFFFFFFFE0000000000000000FFFFFFFFFFFFFFFE000000000000000FFFFFFFFFFFFFFE00000000000000FFFFFFFFFFFFFF00000000000007FFFFFFFFF";
defparam ram_block1a53.mem_init2 = "FFFC0000000000007FFFFFFFFFFFE000000000000FFFFFFFFFFFF000000000001FFFFFFFFFFF800000000003FFFFFFFFFFC00000000003FFFFFFFFFF80000000001FFFFFFFFFF00000000007FFFFFFFFF80000000007FFFFFFFFF0000000003FFFFFFFFF0000000003FFFFFFFFE000000001FFFFFFFFF000000001FFFFFFFFE000000003FFFFFFFF000000003FFFFFFFF000000003FFFFFFFE00000000FFFFFFFF000000007FFFFFFF00000000FFFFFFFF00000001FFFFFFF80000000FFFFFFFC0000000FFFFFFFC0000000FFFFFFF80000001FFFFFFE0000000FFFFFFF80000007FFFFFF80000007FFFFFF80000007FFFFFF0000001FFFFFFC0000007FFFFFF";
defparam ram_block1a53.mem_init1 = "0000003FFFFFF8000001FFFFFF8000001FFFFFF8000003FFFFFF0000007FFFFFC000001FFFFFF0000007FFFFFC000003FFFFFE000001FFFFFE000001FFFFFE000001FFFFFC000003FFFFF8000007FFFFF000001FFFFFC000007FFFFF000001FFFFF800000FFFFFC000007FFFFE000007FFFFE000007FFFFE000007FFFFE00000FFFFFC00001FFFFF800003FFFFE000007FFFFC00001FFFFF00000FFFFF800003FFFFE00001FFFFF00000FFFFF000007FFFF800007FFFF800007FFFF800007FFFF800007FFFF00000FFFFF00001FFFFE00003FFFF800007FFFF00001FFFFC00007FFFF00001FFFFC00007FFFF00003FFFF80000FFFFC00007FFFE00003FFFF000";
defparam ram_block1a53.mem_init0 = "01FFFF80001FFFF80001FFFFC0000FFFFC0000FFFF80001FFFF80001FFFF80003FFFF00003FFFE00007FFFC0000FFFF80001FFFF00007FFFC0000FFFF80003FFFE0000FFFF80003FFFE0000FFFF80003FFFE0001FFFF00007FFF80003FFFE0001FFFF0000FFFF80007FFFC0003FFFC0001FFFE0001FFFE0001FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFE0001FFFE0001FFFE0003FFFC0003FFF80007FFF0000FFFE0001FFFC0003FFF80007FFF0001FFFE0003FFF8000FFFF0001FFFC0007FFF0001FFFC0007FFF8000FFFC0007FFF0001FFFC0007FFF0001FFF8000FFFE0003FFF0001FFFC000FFFE0003FFF0001FFF8000FFFC0007FFE0003FFF";

arriav_ram_block ram_block1a5(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a5_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.clk0_input_clock_enable = "ena0";
defparam ram_block1a5.clk0_output_clock_enable = "ena0";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.init_file = "DDS_48_v1_nco_ii_0_cos.hex";
defparam ram_block1a5.init_file_layout = "port_a";
defparam ram_block1a5.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0121|altsyncram:altsyncram_component0|altsyncram_78g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.operation_mode = "rom";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 13;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "clock0";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 8191;
defparam ram_block1a5.port_a_logical_ram_depth = 65536;
defparam ram_block1a5.port_a_logical_ram_width = 16;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.ram_block_type = "auto";
defparam ram_block1a5.mem_init3 = "0007FFE0003FFF0001FFF8000FFFC0007FFF0003FFF8001FFFC0007FFF0003FFF8000FFFE0003FFF0001FFFC0007FFF0001FFFC0007FFF0001FFFC0007FFF0000FFFE0003FFF80007FFF0001FFFC0003FFF80007FFF0000FFFE0001FFFC0003FFF80007FFF8000FFFF0000FFFE0001FFFE0001FFFE0001FFFE0001FFFE0001FFFE0001FFFE0001FFFE0001FFFF0000FFFF00007FFF80007FFFC0003FFFE0001FFFF0000FFFF80003FFFC0001FFFF00007FFFC0003FFFE0000FFFF80003FFFE0000FFFFC0001FFFF00007FFFE0000FFFF80001FFFF00003FFFE00007FFFC0000FFFFC0001FFFF80001FFFF80001FFFF80001FFFF80001FFFF80001FFFFC0000FF";
defparam ram_block1a5.mem_init2 = "FFC00007FFFE00003FFFF00001FFFF80000FFFFE00003FFFF00001FFFFC00007FFFF00001FFFFE00003FFFF80000FFFFF00001FFFFE00003FFFFC00003FFFFC00007FFFF800007FFFF800007FFFF800003FFFFC00003FFFFE00001FFFFF00000FFFFF800003FFFFE00000FFFFF800003FFFFE00000FFFFF800001FFFFF000003FFFFF000007FFFFE000007FFFFE000007FFFFE000007FFFFF000003FFFFF800001FFFFFC000007FFFFF000001FFFFFC000007FFFFF800000FFFFFF000000FFFFFE000001FFFFFE000001FFFFFF000000FFFFFF8000007FFFFFC000001FFFFFF0000007FFFFFE000000FFFFFFC000001FFFFFF8000001FFFFFFC000000FFFFFFC";
defparam ram_block1a5.mem_init1 = "0000007FFFFFF0000001FFFFFFC0000003FFFFFF80000007FFFFFF80000007FFFFFF80000003FFFFFFE0000000FFFFFFF80000003FFFFFFF00000003FFFFFFF00000003FFFFFFF80000001FFFFFFFC00000003FFFFFFFC00000007FFFFFFFC00000003FFFFFFFE00000000FFFFFFFFC00000000FFFFFFFFC00000000FFFFFFFFE000000001FFFFFFFFC000000003FFFFFFFFE000000000FFFFFFFFFC000000000FFFFFFFFFC0000000007FFFFFFFFF80000000007FFFFFFFFFC0000000001FFFFFFFFFF80000000000FFFFFFFFFFE00000000000FFFFFFFFFFF800000000001FFFFFFFFFFFC000000000007FFFFFFFFFFFC000000000000FFFFFFFFFFFFE0000";
defparam ram_block1a5.mem_init0 = "000000000FFFFFFFFFFFFFC00000000000007FFFFFFFFFFFFFC000000000000007FFFFFFFFFFFFFFC0000000000000007FFFFFFFFFFFFFFFC00000000000000003FFFFFFFFFFFFFFFFFC0000000000000000007FFFFFFFFFFFFFFFFFFF0000000000000000000007FFFFFFFFFFFFFFFFFFFFFE0000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

arriav_ram_block ram_block1a21(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a21_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a21.clk0_core_clock_enable = "ena0";
defparam ram_block1a21.clk0_input_clock_enable = "ena0";
defparam ram_block1a21.clk0_output_clock_enable = "ena0";
defparam ram_block1a21.data_interleave_offset_in_bits = 1;
defparam ram_block1a21.data_interleave_width_in_bits = 1;
defparam ram_block1a21.init_file = "DDS_48_v1_nco_ii_0_cos.hex";
defparam ram_block1a21.init_file_layout = "port_a";
defparam ram_block1a21.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0121|altsyncram:altsyncram_component0|altsyncram_78g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a21.operation_mode = "rom";
defparam ram_block1a21.port_a_address_clear = "none";
defparam ram_block1a21.port_a_address_width = 13;
defparam ram_block1a21.port_a_data_out_clear = "none";
defparam ram_block1a21.port_a_data_out_clock = "clock0";
defparam ram_block1a21.port_a_data_width = 1;
defparam ram_block1a21.port_a_first_address = 8192;
defparam ram_block1a21.port_a_first_bit_number = 5;
defparam ram_block1a21.port_a_last_address = 16383;
defparam ram_block1a21.port_a_logical_ram_depth = 65536;
defparam ram_block1a21.port_a_logical_ram_width = 16;
defparam ram_block1a21.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a21.ram_block_type = "auto";
defparam ram_block1a21.mem_init3 = "003FF003FF003FF001FF801FF801FFC00FFC00FFC007FE007FE007FE003FF003FF003FF801FF801FF800FFC00FFC00FFE007FE007FE007FF003FF003FF001FF801FF801FFC00FFC00FFC007FE007FE007FF003FF003FF801FF801FF800FFC00FFC00FFE007FE007FF003FF003FF001FF801FF800FFC00FFC00FFE007FE007FF003FF003FF801FF801FFC00FFC00FFC007FE007FE003FF003FF801FF801FFC00FFC00FFE007FE007FF003FF003FF801FF800FFC00FFC007FE007FF003FF003FF801FF800FFC00FFE007FE003FF003FF001FF801FFC00FFC007FE007FF003FF001FF801FFC00FFC007FE007FF003FF801FF800FFC00FFE007FE003FF001FF801FF";
defparam ram_block1a21.mem_init2 = "C00FFE007FE003FF001FF801FFC00FFE007FE003FF001FF801FFC00FFE007FF003FF801FF800FFC007FE003FF001FF800FFC007FE007FF003FF801FFC00FFE007FF003FF801FFC00FFE007FF001FF800FFC007FE003FF001FF800FFE007FF003FF801FFC007FE003FF001FF800FFE007FF003FF800FFC007FF003FF801FFC007FE003FF801FFC007FE003FF801FFC007FE003FF801FFC007FF003FF800FFC007FF001FF800FFE003FF001FFC007FE003FF800FFE007FF001FFC00FFE003FF800FFE007FF001FFC007FF003FF800FFE003FF800FFC007FF001FFC007FF001FFC007FE003FF800FFE003FF800FFE003FF800FFE003FF800FFE003FF800FFE003FF";
defparam ram_block1a21.mem_init1 = "800FFE003FF800FFE003FF800FFE001FFC007FF001FFC007FF001FFC003FF800FFE003FF800FFF001FFC007FF000FFE003FF800FFF001FFC007FF800FFE003FFC007FF001FFE003FF8007FF001FFE003FF8007FF001FFE003FF8007FF001FFE003FFC007FF800FFE001FFC003FF8007FF000FFE001FFC003FF8007FF000FFE001FFC003FFC007FF800FFF001FFE001FFC003FFC007FF8007FF000FFF001FFE001FFC003FFC003FF8007FF8007FF000FFF000FFF001FFE001FFE001FFE003FFC003FFC003FFC003FFC003FFC007FF8007FF8007FF8007FF8007FF8007FF8007FF8003FFC003FFC003FFC003FFC003FFE001FFE001FFE001FFF000FFF000FFF000";
defparam ram_block1a21.mem_init0 = "7FF8007FF8003FFC003FFE001FFE000FFF000FFF8007FFC003FFC001FFE000FFF0007FF8003FFC001FFE000FFF0007FF8003FFC001FFF000FFF8003FFC001FFF000FFF8003FFC001FFF0007FF8003FFE000FFF8007FFC001FFF0007FFC001FFF0007FF8003FFE000FFF8003FFE000FFF8003FFF0007FFC001FFF0007FFC001FFF8003FFE000FFF8001FFF0007FFC000FFF8003FFF0007FFE000FFF8001FFF0003FFE0007FFC000FFF8001FFF0003FFE0007FFE000FFFC001FFF8001FFF8003FFF0003FFF0007FFE0007FFE0007FFE000FFFC000FFFC000FFFC000FFFC000FFFC000FFFC0007FFE0007FFE0007FFE0003FFF0003FFF0001FFF8001FFFC000FFFC";

arriav_ram_block ram_block1a70(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a70_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a70.clk0_core_clock_enable = "ena0";
defparam ram_block1a70.clk0_input_clock_enable = "ena0";
defparam ram_block1a70.clk0_output_clock_enable = "ena0";
defparam ram_block1a70.data_interleave_offset_in_bits = 1;
defparam ram_block1a70.data_interleave_width_in_bits = 1;
defparam ram_block1a70.init_file = "DDS_48_v1_nco_ii_0_cos.hex";
defparam ram_block1a70.init_file_layout = "port_a";
defparam ram_block1a70.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0121|altsyncram:altsyncram_component0|altsyncram_78g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a70.operation_mode = "rom";
defparam ram_block1a70.port_a_address_clear = "none";
defparam ram_block1a70.port_a_address_width = 13;
defparam ram_block1a70.port_a_data_out_clear = "none";
defparam ram_block1a70.port_a_data_out_clock = "clock0";
defparam ram_block1a70.port_a_data_width = 1;
defparam ram_block1a70.port_a_first_address = 32768;
defparam ram_block1a70.port_a_first_bit_number = 6;
defparam ram_block1a70.port_a_last_address = 40959;
defparam ram_block1a70.port_a_logical_ram_depth = 65536;
defparam ram_block1a70.port_a_logical_ram_width = 16;
defparam ram_block1a70.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a70.ram_block_type = "auto";
defparam ram_block1a70.mem_init3 = "FFFFFFF00000007FFFFFFC0000001FFFFFFF00000007FFFFFFE0000000FFFFFFFC0000001FFFFFFF80000001FFFFFFF80000003FFFFFFF80000001FFFFFFF80000001FFFFFFFC0000000FFFFFFFE00000003FFFFFFF80000000FFFFFFFE00000003FFFFFFF80000000FFFFFFFF00000000FFFFFFFE00000001FFFFFFFE00000001FFFFFFFE00000000FFFFFFFF000000007FFFFFFF800000003FFFFFFFE00000000FFFFFFFFC00000001FFFFFFFF000000003FFFFFFFF000000003FFFFFFFF000000003FFFFFFFF800000001FFFFFFFFC000000007FFFFFFFF000000001FFFFFFFFC000000003FFFFFFFFC000000007FFFFFFFF8000000003FFFFFFFFC000000";
defparam ram_block1a70.mem_init2 = "001FFFFFFFFF0000000007FFFFFFFFC000000001FFFFFFFFF8000000001FFFFFFFFF8000000001FFFFFFFFFC000000000FFFFFFFFFE0000000001FFFFFFFFFC0000000003FFFFFFFFFC0000000003FFFFFFFFFE0000000001FFFFFFFFFF00000000003FFFFFFFFFE00000000007FFFFFFFFFF00000000003FFFFFFFFFF80000000000FFFFFFFFFFF00000000000FFFFFFFFFFF000000000007FFFFFFFFFFC00000000001FFFFFFFFFFF800000000001FFFFFFFFFFFC000000000007FFFFFFFFFFF000000000000FFFFFFFFFFFF0000000000007FFFFFFFFFFFE0000000000007FFFFFFFFFFFE0000000000003FFFFFFFFFFFFC0000000000003FFFFFFFFFFFFE";
defparam ram_block1a70.mem_init1 = "00000000000007FFFFFFFFFFFFE00000000000003FFFFFFFFFFFFFC00000000000003FFFFFFFFFFFFFF000000000000003FFFFFFFFFFFFFF8000000000000007FFFFFFFFFFFFFFC000000000000001FFFFFFFFFFFFFFFE0000000000000001FFFFFFFFFFFFFFFF00000000000000001FFFFFFFFFFFFFFFFE00000000000000000FFFFFFFFFFFFFFFFFE000000000000000000FFFFFFFFFFFFFFFFFFE0000000000000000001FFFFFFFFFFFFFFFFFFFC00000000000000000001FFFFFFFFFFFFFFFFFFFFC0000000000000000000007FFFFFFFFFFFFFFFFFFFFFC00000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000007FFF";
defparam ram_block1a70.mem_init0 = "FFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

arriav_ram_block ram_block1a86(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a86_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a86.clk0_core_clock_enable = "ena0";
defparam ram_block1a86.clk0_input_clock_enable = "ena0";
defparam ram_block1a86.clk0_output_clock_enable = "ena0";
defparam ram_block1a86.data_interleave_offset_in_bits = 1;
defparam ram_block1a86.data_interleave_width_in_bits = 1;
defparam ram_block1a86.init_file = "DDS_48_v1_nco_ii_0_cos.hex";
defparam ram_block1a86.init_file_layout = "port_a";
defparam ram_block1a86.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0121|altsyncram:altsyncram_component0|altsyncram_78g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a86.operation_mode = "rom";
defparam ram_block1a86.port_a_address_clear = "none";
defparam ram_block1a86.port_a_address_width = 13;
defparam ram_block1a86.port_a_data_out_clear = "none";
defparam ram_block1a86.port_a_data_out_clock = "clock0";
defparam ram_block1a86.port_a_data_width = 1;
defparam ram_block1a86.port_a_first_address = 40960;
defparam ram_block1a86.port_a_first_bit_number = 6;
defparam ram_block1a86.port_a_last_address = 49151;
defparam ram_block1a86.port_a_logical_ram_depth = 65536;
defparam ram_block1a86.port_a_logical_ram_width = 16;
defparam ram_block1a86.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a86.ram_block_type = "auto";
defparam ram_block1a86.mem_init3 = "FFFFF00000FFFFF800007FFFFC00003FFFFC00001FFFFE00001FFFFF00000FFFFF800007FFFF800003FFFFC00003FFFFE00001FFFFF00000FFFFF000007FFFF800003FFFFC00003FFFFE00001FFFFF00000FFFFF000007FFFF800003FFFFC00001FFFFE00001FFFFF00000FFFFF800007FFFFC00003FFFFE00001FFFFE00000FFFFF000007FFFF800003FFFFC00001FFFFE00000FFFFF000007FFFF800003FFFFC00001FFFFE00000FFFFF800007FFFFC00003FFFFE00001FFFFF000007FFFF800003FFFFC00001FFFFF00000FFFFF800007FFFFC00001FFFFE00000FFFFF800007FFFFC00001FFFFE00000FFFFF800003FFFFC00001FFFFF000007FFFF80000";
defparam ram_block1a86.mem_init2 = "3FFFFE00000FFFFF000007FFFFC00001FFFFF000007FFFF800003FFFFE00000FFFFF800003FFFFE00000FFFFF000007FFFFC00001FFFFF000007FFFFC00001FFFFF000007FFFFC00001FFFFF000007FFFFC00000FFFFF800003FFFFE00000FFFFF800003FFFFE000007FFFFC00001FFFFF000007FFFFE00000FFFFF800003FFFFF000007FFFFC00000FFFFF800003FFFFF000007FFFFE00000FFFFF800001FFFFF000003FFFFE000007FFFFC00000FFFFF800001FFFFF000003FFFFF000007FFFFE000007FFFFC00000FFFFFC00001FFFFF800001FFFFF800003FFFFF000003FFFFF000003FFFFF000007FFFFE000007FFFFE000007FFFFE000007FFFFE00000";
defparam ram_block1a86.mem_init1 = "7FFFFE000007FFFFF000003FFFFF000003FFFFF000003FFFFF800001FFFFF800001FFFFFC00000FFFFFC000007FFFFE000007FFFFF000003FFFFF800001FFFFFC00000FFFFFE000003FFFFF000001FFFFFC00000FFFFFE000003FFFFF000001FFFFFC000007FFFFF000001FFFFFC000007FFFFF000003FFFFFC000007FFFFF000001FFFFFC000007FFFFF000001FFFFFE000003FFFFF8000007FFFFF000001FFFFFE000003FFFFFC000007FFFFF800000FFFFFF000000FFFFFE000001FFFFFE000003FFFFFC000003FFFFFC000003FFFFFC000003FFFFFC000003FFFFFC000003FFFFFC000003FFFFFC000001FFFFFE000001FFFFFF000000FFFFFF0000007FF";
defparam ram_block1a86.mem_init0 = "FFF8000003FFFFFC000001FFFFFF000000FFFFFF8000003FFFFFE000000FFFFFF8000003FFFFFC000000FFFFFF8000003FFFFFE000000FFFFFF8000001FFFFFF0000007FFFFFE000000FFFFFFC000001FFFFFF8000001FFFFFF0000003FFFFFF0000003FFFFFF0000003FFFFFF0000003FFFFFF0000003FFFFFF0000001FFFFFF8000001FFFFFFC000000FFFFFFE0000003FFFFFF0000001FFFFFFC0000007FFFFFE0000003FFFFFF80000007FFFFFF0000001FFFFFFC0000003FFFFFF8000000FFFFFFF0000000FFFFFFE0000001FFFFFFE0000001FFFFFFE0000001FFFFFFE0000001FFFFFFE0000001FFFFFFF0000000FFFFFFF80000007FFFFFFC0000001";

arriav_ram_block ram_block1a102(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a102_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a102.clk0_core_clock_enable = "ena0";
defparam ram_block1a102.clk0_input_clock_enable = "ena0";
defparam ram_block1a102.clk0_output_clock_enable = "ena0";
defparam ram_block1a102.data_interleave_offset_in_bits = 1;
defparam ram_block1a102.data_interleave_width_in_bits = 1;
defparam ram_block1a102.init_file = "DDS_48_v1_nco_ii_0_cos.hex";
defparam ram_block1a102.init_file_layout = "port_a";
defparam ram_block1a102.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0121|altsyncram:altsyncram_component0|altsyncram_78g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a102.operation_mode = "rom";
defparam ram_block1a102.port_a_address_clear = "none";
defparam ram_block1a102.port_a_address_width = 13;
defparam ram_block1a102.port_a_data_out_clear = "none";
defparam ram_block1a102.port_a_data_out_clock = "clock0";
defparam ram_block1a102.port_a_data_width = 1;
defparam ram_block1a102.port_a_first_address = 49152;
defparam ram_block1a102.port_a_first_bit_number = 6;
defparam ram_block1a102.port_a_last_address = 57343;
defparam ram_block1a102.port_a_logical_ram_depth = 65536;
defparam ram_block1a102.port_a_logical_ram_width = 16;
defparam ram_block1a102.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a102.ram_block_type = "auto";
defparam ram_block1a102.mem_init3 = "7FFFFFF80000003FFFFFFE0000001FFFFFFF0000000FFFFFFF00000007FFFFFF80000007FFFFFF80000007FFFFFF8000000FFFFFFF0000000FFFFFFE0000001FFFFFFC0000003FFFFFF8000000FFFFFFF0000001FFFFFFC0000007FFFFFF0000001FFFFFFC000000FFFFFFE0000003FFFFFF8000001FFFFFFC000000FFFFFFC0000007FFFFFE0000007FFFFFE0000003FFFFFF0000003FFFFFF0000003FFFFFE0000007FFFFFE0000007FFFFFC000000FFFFFFC000001FFFFFF8000003FFFFFE0000007FFFFFC000001FFFFFF8000003FFFFFE000000FFFFFF8000003FFFFFE000000FFFFFF8000007FFFFFC000001FFFFFF000000FFFFFF8000003FFFFFC000";
defparam ram_block1a102.mem_init2 = "001FFFFFE000001FFFFFF000000FFFFFF0000007FFFFF8000007FFFFF8000003FFFFFC000003FFFFFC000003FFFFFC000003FFFFF8000007FFFFF8000007FFFFF800000FFFFFF000000FFFFFE000001FFFFFE000003FFFFFC000007FFFFF800000FFFFFE000001FFFFFC000007FFFFF800000FFFFFE000003FFFFF8000007FFFFF000001FFFFFC000007FFFFF000001FFFFFC000007FFFFF000003FFFFF800000FFFFFE000003FFFFF000001FFFFFC00000FFFFFE000003FFFFF000001FFFFF800000FFFFFC000007FFFFE000003FFFFF000001FFFFF800001FFFFFC00000FFFFFC000007FFFFE000007FFFFE000007FFFFF000003FFFFF000003FFFFF000003";
defparam ram_block1a102.mem_init1 = "FFFFF000003FFFFF000003FFFFF000003FFFFF000003FFFFF000003FFFFF000007FFFFE000007FFFFE000007FFFFC00000FFFFFC00001FFFFF800001FFFFF000003FFFFF000007FFFFE00000FFFFFC00000FFFFF800001FFFFF000003FFFFE000007FFFFC00001FFFFF800003FFFFF000007FFFFC00000FFFFF800003FFFFF000007FFFFC00001FFFFF800003FFFFE00000FFFFFC00001FFFFF000007FFFFC00001FFFFF000003FFFFE00000FFFFF800003FFFFE00000FFFFF800003FFFFE00000FFFFF800003FFFFE00000FFFFF800003FFFFE00000FFFFF800003FFFFC00001FFFFF000007FFFFC00001FFFFF00000FFFFF800003FFFFE00000FFFFF000007";
defparam ram_block1a102.mem_init0 = "FFFFC00001FFFFF00000FFFFF800003FFFFC00001FFFFF000007FFFF800003FFFFE00001FFFFF000007FFFF800003FFFFE00001FFFFF00000FFFFF800003FFFFC00001FFFFE00000FFFFF800007FFFFC00003FFFFE00001FFFFF00000FFFFF800007FFFFC00003FFFFE00000FFFFF000007FFFF800007FFFFC00003FFFFE00001FFFFF00000FFFFF800007FFFFC00003FFFFE00001FFFFE00000FFFFF000007FFFF800003FFFFC00003FFFFE00001FFFFF00000FFFFF800007FFFF800003FFFFC00001FFFFE00001FFFFF00000FFFFF000007FFFF800003FFFFC00003FFFFE00001FFFFF00000FFFFF000007FFFF800007FFFFC00003FFFFE00001FFFFE00000";

arriav_ram_block ram_block1a118(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a118_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a118.clk0_core_clock_enable = "ena0";
defparam ram_block1a118.clk0_input_clock_enable = "ena0";
defparam ram_block1a118.clk0_output_clock_enable = "ena0";
defparam ram_block1a118.data_interleave_offset_in_bits = 1;
defparam ram_block1a118.data_interleave_width_in_bits = 1;
defparam ram_block1a118.init_file = "DDS_48_v1_nco_ii_0_cos.hex";
defparam ram_block1a118.init_file_layout = "port_a";
defparam ram_block1a118.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0121|altsyncram:altsyncram_component0|altsyncram_78g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a118.operation_mode = "rom";
defparam ram_block1a118.port_a_address_clear = "none";
defparam ram_block1a118.port_a_address_width = 13;
defparam ram_block1a118.port_a_data_out_clear = "none";
defparam ram_block1a118.port_a_data_out_clock = "clock0";
defparam ram_block1a118.port_a_data_width = 1;
defparam ram_block1a118.port_a_first_address = 57344;
defparam ram_block1a118.port_a_first_bit_number = 6;
defparam ram_block1a118.port_a_last_address = 65535;
defparam ram_block1a118.port_a_logical_ram_depth = 65536;
defparam ram_block1a118.port_a_logical_ram_width = 16;
defparam ram_block1a118.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a118.ram_block_type = "auto";
defparam ram_block1a118.mem_init3 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000";
defparam ram_block1a118.mem_init2 = "0000FFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000FFFFFFFFFFFFFFFFFFFFFC000000000000000000007FFFFFFFFFFFFFFFFFFFC00000000000000000007FFFFFFFFFFFFFFFFFF8000000000000000000FFFFFFFFFFFFFFFFFF800000000000000000FFFFFFFFFFFFFFFFF800000000000000007FFFFFFFFFFFFFFFF00000000000000007FFFFFFFFFFFFFFF80000000000000007FFFFFFFFFFFFFFC000000000000001FFFFFFFFFFFFFFE000000000000003FFFFFFFFFFFFFF000000000000003FFFFFFFFFFFFFC00000000000003FFFFFFFFFFFFF80000000000001FFFFFFFFFFFFF";
defparam ram_block1a118.mem_init1 = "80000000000007FFFFFFFFFFFFC0000000000007FFFFFFFFFFFF0000000000001FFFFFFFFFFFF8000000000003FFFFFFFFFFFE000000000000FFFFFFFFFFFF000000000001FFFFFFFFFFFC000000000007FFFFFFFFFFE000000000007FFFFFFFFFFC00000000001FFFFFFFFFFF00000000000FFFFFFFFFFF00000000001FFFFFFFFFFE00000000003FFFFFFFFFF00000000003FFFFFFFFFF00000000003FFFFFFFFFE0000000000FFFFFFFFFF80000000003FFFFFFFFFC0000000003FFFFFFFFF80000000007FFFFFFFFF0000000001FFFFFFFFFC000000000FFFFFFFFFE0000000007FFFFFFFFE000000000FFFFFFFFFC000000001FFFFFFFFF0000000007FF";
defparam ram_block1a118.mem_init0 = "FFFFFF8000000003FFFFFFFFC000000003FFFFFFFFC000000003FFFFFFFF8000000007FFFFFFFF000000001FFFFFFFFC00000000FFFFFFFFE000000007FFFFFFFF000000003FFFFFFFF000000007FFFFFFFE000000007FFFFFFFC00000001FFFFFFFF000000007FFFFFFFC00000001FFFFFFFE00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000001FFFFFFFC00000003FFFFFFF80000000FFFFFFFE00000003FFFFFFF80000001FFFFFFFC0000000FFFFFFFE00000007FFFFFFE00000007FFFFFFE00000007FFFFFFE0000000FFFFFFFC0000001FFFFFFF80000003FFFFFFE00000007FFFFFFC0000001FFFFFFF0000000";

arriav_ram_block ram_block1a38(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a38_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a38.clk0_core_clock_enable = "ena0";
defparam ram_block1a38.clk0_input_clock_enable = "ena0";
defparam ram_block1a38.clk0_output_clock_enable = "ena0";
defparam ram_block1a38.data_interleave_offset_in_bits = 1;
defparam ram_block1a38.data_interleave_width_in_bits = 1;
defparam ram_block1a38.init_file = "DDS_48_v1_nco_ii_0_cos.hex";
defparam ram_block1a38.init_file_layout = "port_a";
defparam ram_block1a38.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0121|altsyncram:altsyncram_component0|altsyncram_78g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a38.operation_mode = "rom";
defparam ram_block1a38.port_a_address_clear = "none";
defparam ram_block1a38.port_a_address_width = 13;
defparam ram_block1a38.port_a_data_out_clear = "none";
defparam ram_block1a38.port_a_data_out_clock = "clock0";
defparam ram_block1a38.port_a_data_width = 1;
defparam ram_block1a38.port_a_first_address = 16384;
defparam ram_block1a38.port_a_first_bit_number = 6;
defparam ram_block1a38.port_a_last_address = 24575;
defparam ram_block1a38.port_a_logical_ram_depth = 65536;
defparam ram_block1a38.port_a_logical_ram_width = 16;
defparam ram_block1a38.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a38.ram_block_type = "auto";
defparam ram_block1a38.mem_init3 = "00000007FFFFFFC0000003FFFFFFE0000001FFFFFFF0000000FFFFFFF0000000FFFFFFF0000000FFFFFFF0000000FFFFFFF0000000FFFFFFE0000001FFFFFFE0000003FFFFFF80000007FFFFFF0000001FFFFFFC0000003FFFFFF8000000FFFFFFC0000007FFFFFF0000001FFFFFF8000000FFFFFFE0000007FFFFFF0000003FFFFFF0000001FFFFFF8000001FFFFFF8000001FFFFFF8000001FFFFFF8000001FFFFFF8000001FFFFFF0000003FFFFFF0000007FFFFFE000000FFFFFFC000001FFFFFF0000003FFFFFE000000FFFFFF8000003FFFFFE0000007FFFFF8000003FFFFFE000000FFFFFF8000003FFFFFE000001FFFFFF0000007FFFFF8000003FFF";
defparam ram_block1a38.mem_init2 = "FFC000001FFFFFE000001FFFFFF000000FFFFFF0000007FFFFF8000007FFFFF8000007FFFFF8000007FFFFF8000007FFFFF8000007FFFFF8000007FFFFF800000FFFFFF000000FFFFFE000001FFFFFE000003FFFFFC000007FFFFF800000FFFFFF000001FFFFFC000003FFFFF800000FFFFFF000001FFFFFC000007FFFFF000001FFFFFC000007FFFFF800001FFFFFC000007FFFFF000001FFFFFC000007FFFFF000001FFFFF800000FFFFFE000007FFFFF000001FFFFF800000FFFFFE000007FFFFF000003FFFFF800001FFFFFC00000FFFFFC000007FFFFE000007FFFFF000003FFFFF000003FFFFF800001FFFFF800001FFFFF800001FFFFFC00000FFFFFC";
defparam ram_block1a38.mem_init1 = "00000FFFFFC00000FFFFFC00000FFFFFC00000FFFFFC00001FFFFF800001FFFFF800001FFFFF800003FFFFF000003FFFFF000007FFFFE000007FFFFC00000FFFFFC00001FFFFF800001FFFFF000003FFFFE000007FFFFC00000FFFFF800001FFFFF000003FFFFE00000FFFFFC00001FFFFF800003FFFFE000007FFFFC00001FFFFF800003FFFFE00000FFFFFC00001FFFFF000007FFFFC00000FFFFF800003FFFFE00000FFFFF800003FFFFE000007FFFFC00001FFFFF000007FFFFC00001FFFFF000007FFFFC00001FFFFF000007FFFFC00001FFFFE00000FFFFF800003FFFFE00000FFFFF800003FFFFC00001FFFFF000007FFFFC00001FFFFE00000FFFFF8";
defparam ram_block1a38.mem_init0 = "00003FFFFC00001FFFFF000007FFFF800003FFFFE00000FFFFF000007FFFFC00003FFFFE00000FFFFF000007FFFFC00003FFFFE00001FFFFF000007FFFF800003FFFFC00001FFFFF00000FFFFF800007FFFFC00003FFFFE00000FFFFF000007FFFF800003FFFFC00001FFFFE00000FFFFF000007FFFF800003FFFFC00001FFFFE00000FFFFF00000FFFFF800007FFFFC00003FFFFE00001FFFFF00000FFFFF000007FFFF800003FFFFC00001FFFFE00001FFFFF00000FFFFF800007FFFF800003FFFFC00001FFFFE00001FFFFF00000FFFFF800007FFFF800003FFFFC00003FFFFE00001FFFFF00000FFFFF000007FFFF800007FFFFC00003FFFFE00001FFFFE";

arriav_ram_block ram_block1a54(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a54_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a54.clk0_core_clock_enable = "ena0";
defparam ram_block1a54.clk0_input_clock_enable = "ena0";
defparam ram_block1a54.clk0_output_clock_enable = "ena0";
defparam ram_block1a54.data_interleave_offset_in_bits = 1;
defparam ram_block1a54.data_interleave_width_in_bits = 1;
defparam ram_block1a54.init_file = "DDS_48_v1_nco_ii_0_cos.hex";
defparam ram_block1a54.init_file_layout = "port_a";
defparam ram_block1a54.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0121|altsyncram:altsyncram_component0|altsyncram_78g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a54.operation_mode = "rom";
defparam ram_block1a54.port_a_address_clear = "none";
defparam ram_block1a54.port_a_address_width = 13;
defparam ram_block1a54.port_a_data_out_clear = "none";
defparam ram_block1a54.port_a_data_out_clock = "clock0";
defparam ram_block1a54.port_a_data_width = 1;
defparam ram_block1a54.port_a_first_address = 24576;
defparam ram_block1a54.port_a_first_bit_number = 6;
defparam ram_block1a54.port_a_last_address = 32767;
defparam ram_block1a54.port_a_logical_ram_depth = 65536;
defparam ram_block1a54.port_a_logical_ram_width = 16;
defparam ram_block1a54.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a54.ram_block_type = "auto";
defparam ram_block1a54.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a54.mem_init2 = "FFFC0000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000007FFFFFFFFFFFFFFFFFFFFFC0000000000000000000007FFFFFFFFFFFFFFFFFFFF000000000000000000007FFFFFFFFFFFFFFFFFFF0000000000000000000FFFFFFFFFFFFFFFFFFE000000000000000000FFFFFFFFFFFFFFFFFE00000000000000000FFFFFFFFFFFFFFFFF00000000000000001FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF0000000000000007FFFFFFFFFFFFFFC000000000000003FFFFFFFFFFFFFF800000000000001FFFFFFFFFFFFFF800000000000007FFFFFFFFFFFFF80000000000000FFFFFFFFFFFFFC0000000000000";
defparam ram_block1a54.mem_init1 = "FFFFFFFFFFFFF80000000000007FFFFFFFFFFFF8000000000000FFFFFFFFFFFFC000000000000FFFFFFFFFFFFC000000000001FFFFFFFFFFFE000000000001FFFFFFFFFFFC000000000007FFFFFFFFFFF000000000003FFFFFFFFFFF000000000007FFFFFFFFFFC00000000001FFFFFFFFFFE00000000001FFFFFFFFFFE00000000003FFFFFFFFFF80000000001FFFFFFFFFFC0000000000FFFFFFFFFF80000000001FFFFFFFFFF0000000000FFFFFFFFFF80000000007FFFFFFFFF80000000007FFFFFFFFF0000000000FFFFFFFFFE0000000007FFFFFFFFF0000000003FFFFFFFFF0000000003FFFFFFFFF0000000007FFFFFFFFC000000001FFFFFFFFF000";
defparam ram_block1a54.mem_init0 = "0000007FFFFFFFF8000000003FFFFFFFFC000000007FFFFFFFF8000000007FFFFFFFF000000001FFFFFFFFC000000007FFFFFFFF000000003FFFFFFFF800000001FFFFFFFF800000001FFFFFFFF800000001FFFFFFFF000000007FFFFFFFE00000000FFFFFFFF800000003FFFFFFFC00000001FFFFFFFE00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFE00000001FFFFFFFE00000003FFFFFFF80000000FFFFFFFE00000003FFFFFFF80000000FFFFFFFE00000007FFFFFFF00000003FFFFFFF00000003FFFFFFF80000003FFFFFFF00000003FFFFFFF00000007FFFFFFE0000000FFFFFFFC0000001FFFFFFF00000007FFFFFFC0000001FFFFFFF";

arriav_ram_block ram_block1a6(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a6_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.clk0_input_clock_enable = "ena0";
defparam ram_block1a6.clk0_output_clock_enable = "ena0";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.init_file = "DDS_48_v1_nco_ii_0_cos.hex";
defparam ram_block1a6.init_file_layout = "port_a";
defparam ram_block1a6.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0121|altsyncram:altsyncram_component0|altsyncram_78g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.operation_mode = "rom";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 13;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "clock0";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 8191;
defparam ram_block1a6.port_a_logical_ram_depth = 65536;
defparam ram_block1a6.port_a_logical_ram_width = 16;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.ram_block_type = "auto";
defparam ram_block1a6.mem_init3 = "0000001FFFFFFF00000007FFFFFFC0000000FFFFFFF80000003FFFFFFF00000007FFFFFFE0000000FFFFFFFC0000000FFFFFFFC0000000FFFFFFFC0000000FFFFFFFE00000007FFFFFFF00000003FFFFFFF80000000FFFFFFFE00000003FFFFFFF800000007FFFFFFF00000001FFFFFFFE00000001FFFFFFFE00000001FFFFFFFE00000001FFFFFFFE00000000FFFFFFFF000000007FFFFFFFC00000001FFFFFFFF000000007FFFFFFFC00000000FFFFFFFFC00000001FFFFFFFF800000001FFFFFFFFC00000000FFFFFFFFE000000007FFFFFFFF000000001FFFFFFFFC000000003FFFFFFFF8000000007FFFFFFFF8000000007FFFFFFFF8000000003FFFFFF";
defparam ram_block1a6.mem_init2 = "FFC000000001FFFFFFFFF0000000007FFFFFFFFE000000000FFFFFFFFFC000000000FFFFFFFFFE0000000007FFFFFFFFF0000000001FFFFFFFFFC0000000003FFFFFFFFF80000000007FFFFFFFFF80000000003FFFFFFFFFE0000000000FFFFFFFFFF80000000001FFFFFFFFFF80000000001FFFFFFFFFF80000000000FFFFFFFFFFF00000000001FFFFFFFFFFE00000000001FFFFFFFFFFF000000000007FFFFFFFFFFC00000000000FFFFFFFFFFFC000000000007FFFFFFFFFFF000000000001FFFFFFFFFFFE000000000000FFFFFFFFFFFF8000000000003FFFFFFFFFFFF0000000000001FFFFFFFFFFFFC0000000000007FFFFFFFFFFFFC0000000000003";
defparam ram_block1a6.mem_init1 = "FFFFFFFFFFFFF00000000000003FFFFFFFFFFFFF800000000000007FFFFFFFFFFFFF800000000000001FFFFFFFFFFFFFF800000000000000FFFFFFFFFFFFFFF0000000000000007FFFFFFFFFFFFFFC0000000000000003FFFFFFFFFFFFFFFC0000000000000001FFFFFFFFFFFFFFFFC00000000000000003FFFFFFFFFFFFFFFFE000000000000000003FFFFFFFFFFFFFFFFFE0000000000000000003FFFFFFFFFFFFFFFFFFC00000000000000000007FFFFFFFFFFFFFFFFFFFC000000000000000000007FFFFFFFFFFFFFFFFFFFFE00000000000000000000007FFFFFFFFFFFFFFFFFFFFFFC000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFE0000";
defparam ram_block1a6.mem_init0 = "00000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

arriav_ram_block ram_block1a22(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a22_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a22.clk0_core_clock_enable = "ena0";
defparam ram_block1a22.clk0_input_clock_enable = "ena0";
defparam ram_block1a22.clk0_output_clock_enable = "ena0";
defparam ram_block1a22.data_interleave_offset_in_bits = 1;
defparam ram_block1a22.data_interleave_width_in_bits = 1;
defparam ram_block1a22.init_file = "DDS_48_v1_nco_ii_0_cos.hex";
defparam ram_block1a22.init_file_layout = "port_a";
defparam ram_block1a22.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0121|altsyncram:altsyncram_component0|altsyncram_78g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a22.operation_mode = "rom";
defparam ram_block1a22.port_a_address_clear = "none";
defparam ram_block1a22.port_a_address_width = 13;
defparam ram_block1a22.port_a_data_out_clear = "none";
defparam ram_block1a22.port_a_data_out_clock = "clock0";
defparam ram_block1a22.port_a_data_width = 1;
defparam ram_block1a22.port_a_first_address = 8192;
defparam ram_block1a22.port_a_first_bit_number = 6;
defparam ram_block1a22.port_a_last_address = 16383;
defparam ram_block1a22.port_a_logical_ram_depth = 65536;
defparam ram_block1a22.port_a_logical_ram_width = 16;
defparam ram_block1a22.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a22.ram_block_type = "auto";
defparam ram_block1a22.mem_init3 = "00000FFFFF00000FFFFF800007FFFFC00003FFFFC00001FFFFE00001FFFFF00000FFFFF800007FFFF800003FFFFC00001FFFFE00001FFFFF00000FFFFF000007FFFF800003FFFFC00003FFFFE00001FFFFF00000FFFFF800007FFFF800003FFFFC00001FFFFE00000FFFFF00000FFFFF800007FFFFC00003FFFFE00001FFFFF00000FFFFF800007FFFFC00003FFFFC00001FFFFE00000FFFFF800007FFFFC00003FFFFE00001FFFFF00000FFFFF800007FFFFC00003FFFFE00000FFFFF000007FFFF800003FFFFE00001FFFFF00000FFFFF800003FFFFC00001FFFFF00000FFFFF800003FFFFC00001FFFFF000007FFFF800003FFFFE00001FFFFF000007FFFF";
defparam ram_block1a22.mem_init2 = "C00001FFFFE00000FFFFF800003FFFFE00001FFFFF000007FFFFC00001FFFFF000007FFFF800003FFFFE00000FFFFF800003FFFFE00000FFFFF800003FFFFE00000FFFFF800003FFFFE00000FFFFF800003FFFFE00000FFFFF800001FFFFF000007FFFFC00001FFFFF000007FFFFE00000FFFFF800003FFFFF000007FFFFC00001FFFFF800003FFFFE000007FFFFC00001FFFFF800003FFFFF000007FFFFC00000FFFFF800001FFFFF000003FFFFE000007FFFFE00000FFFFFC00001FFFFF800001FFFFF000003FFFFF000007FFFFE000007FFFFC00000FFFFFC00000FFFFFC00001FFFFF800001FFFFF800001FFFFF800001FFFFF800001FFFFF800001FFFFF";
defparam ram_block1a22.mem_init1 = "800001FFFFF800001FFFFF800001FFFFFC00000FFFFFC00000FFFFFC000007FFFFE000007FFFFF000003FFFFF000001FFFFF800000FFFFFC000007FFFFE000003FFFFF000001FFFFF800000FFFFFE000007FFFFF000001FFFFF800000FFFFFE000003FFFFF800001FFFFFC000007FFFFF000001FFFFFC000007FFFFF000001FFFFFC000003FFFFF800000FFFFFE000003FFFFFC000007FFFFF000000FFFFFE000003FFFFFC000007FFFFF800000FFFFFF000000FFFFFE000001FFFFFE000003FFFFFC000003FFFFFC000003FFFFF8000007FFFFF8000007FFFFF8000007FFFFF8000003FFFFFC000003FFFFFC000001FFFFFE000001FFFFFF000000FFFFFF000";
defparam ram_block1a22.mem_init0 = "0007FFFFF8000003FFFFFE000001FFFFFF0000007FFFFFC000003FFFFFE000000FFFFFF8000003FFFFFE000000FFFFFF8000003FFFFFF0000007FFFFFC000000FFFFFF8000003FFFFFF0000007FFFFFE0000007FFFFFC000000FFFFFFC000000FFFFFF8000001FFFFFF8000001FFFFFF8000000FFFFFFC000000FFFFFFC0000007FFFFFE0000007FFFFFF0000003FFFFFF8000000FFFFFFE0000007FFFFFF0000001FFFFFFC0000007FFFFFF0000001FFFFFFE0000003FFFFFF80000007FFFFFF0000000FFFFFFE0000001FFFFFFE0000003FFFFFFC0000003FFFFFFC0000003FFFFFFC0000001FFFFFFE0000001FFFFFFF0000000FFFFFFF80000003FFFFFFC";

arriav_ram_block ram_block1a71(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a71_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a71.clk0_core_clock_enable = "ena0";
defparam ram_block1a71.clk0_input_clock_enable = "ena0";
defparam ram_block1a71.clk0_output_clock_enable = "ena0";
defparam ram_block1a71.data_interleave_offset_in_bits = 1;
defparam ram_block1a71.data_interleave_width_in_bits = 1;
defparam ram_block1a71.init_file = "DDS_48_v1_nco_ii_0_cos.hex";
defparam ram_block1a71.init_file_layout = "port_a";
defparam ram_block1a71.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0121|altsyncram:altsyncram_component0|altsyncram_78g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a71.operation_mode = "rom";
defparam ram_block1a71.port_a_address_clear = "none";
defparam ram_block1a71.port_a_address_width = 13;
defparam ram_block1a71.port_a_data_out_clear = "none";
defparam ram_block1a71.port_a_data_out_clock = "clock0";
defparam ram_block1a71.port_a_data_width = 1;
defparam ram_block1a71.port_a_first_address = 32768;
defparam ram_block1a71.port_a_first_bit_number = 7;
defparam ram_block1a71.port_a_last_address = 40959;
defparam ram_block1a71.port_a_logical_ram_depth = 65536;
defparam ram_block1a71.port_a_logical_ram_width = 16;
defparam ram_block1a71.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a71.ram_block_type = "auto";
defparam ram_block1a71.mem_init3 = "000000000000007FFFFFFFFFFFFFE000000000000007FFFFFFFFFFFFFF000000000000001FFFFFFFFFFFFFFE000000000000003FFFFFFFFFFFFFFE000000000000001FFFFFFFFFFFFFFF0000000000000003FFFFFFFFFFFFFFF0000000000000003FFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFE0000000000000001FFFFFFFFFFFFFFFF00000000000000007FFFFFFFFFFFFFFFC0000000000000000FFFFFFFFFFFFFFFFE00000000000000003FFFFFFFFFFFFFFFFC00000000000000003FFFFFFFFFFFFFFFFE000000000000000007FFFFFFFFFFFFFFFFE000000000000000003FFFFFFFFFFFFFFFFF8000000000000000003FFFFFFFFFFFFFFF";
defparam ram_block1a71.mem_init2 = "FFE0000000000000000007FFFFFFFFFFFFFFFFFE0000000000000000001FFFFFFFFFFFFFFFFFFE0000000000000000000FFFFFFFFFFFFFFFFFFFE00000000000000000003FFFFFFFFFFFFFFFFFFFC00000000000000000001FFFFFFFFFFFFFFFFFFFFC000000000000000000007FFFFFFFFFFFFFFFFFFFFC000000000000000000000FFFFFFFFFFFFFFFFFFFFFF00000000000000000000007FFFFFFFFFFFFFFFFFFFFFE00000000000000000000001FFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000003FFFFFFFFFFFFF";
defparam ram_block1a71.mem_init1 = "FFFFFFFFFFFFF8000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000";
defparam ram_block1a71.mem_init0 = "000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

arriav_ram_block ram_block1a87(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a87_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a87.clk0_core_clock_enable = "ena0";
defparam ram_block1a87.clk0_input_clock_enable = "ena0";
defparam ram_block1a87.clk0_output_clock_enable = "ena0";
defparam ram_block1a87.data_interleave_offset_in_bits = 1;
defparam ram_block1a87.data_interleave_width_in_bits = 1;
defparam ram_block1a87.init_file = "DDS_48_v1_nco_ii_0_cos.hex";
defparam ram_block1a87.init_file_layout = "port_a";
defparam ram_block1a87.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0121|altsyncram:altsyncram_component0|altsyncram_78g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a87.operation_mode = "rom";
defparam ram_block1a87.port_a_address_clear = "none";
defparam ram_block1a87.port_a_address_width = 13;
defparam ram_block1a87.port_a_data_out_clear = "none";
defparam ram_block1a87.port_a_data_out_clock = "clock0";
defparam ram_block1a87.port_a_data_width = 1;
defparam ram_block1a87.port_a_first_address = 40960;
defparam ram_block1a87.port_a_first_bit_number = 7;
defparam ram_block1a87.port_a_last_address = 49151;
defparam ram_block1a87.port_a_logical_ram_depth = 65536;
defparam ram_block1a87.port_a_logical_ram_width = 16;
defparam ram_block1a87.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a87.ram_block_type = "auto";
defparam ram_block1a87.mem_init3 = "FFFFFFFFFF00000000007FFFFFFFFFC0000000001FFFFFFFFFE0000000000FFFFFFFFFF80000000003FFFFFFFFFC0000000001FFFFFFFFFF00000000007FFFFFFFFFC0000000003FFFFFFFFFE0000000000FFFFFFFFFF80000000003FFFFFFFFFE0000000001FFFFFFFFFF00000000007FFFFFFFFFC0000000001FFFFFFFFFF00000000007FFFFFFFFFC0000000001FFFFFFFFFF00000000007FFFFFFFFFC0000000001FFFFFFFFFF00000000007FFFFFFFFFC0000000001FFFFFFFFFF80000000003FFFFFFFFFE0000000000FFFFFFFFFF80000000001FFFFFFFFFF00000000007FFFFFFFFFE0000000000FFFFFFFFFFC0000000001FFFFFFFFFF8000000000";
defparam ram_block1a87.mem_init2 = "3FFFFFFFFFF00000000007FFFFFFFFFE00000000007FFFFFFFFFC0000000000FFFFFFFFFFC0000000000FFFFFFFFFF80000000001FFFFFFFFFF80000000001FFFFFFFFFF80000000001FFFFFFFFFF80000000000FFFFFFFFFFC0000000000FFFFFFFFFFC00000000007FFFFFFFFFE00000000007FFFFFFFFFF00000000003FFFFFFFFFF80000000000FFFFFFFFFFC00000000007FFFFFFFFFF00000000001FFFFFFFFFFC00000000007FFFFFFFFFF00000000001FFFFFFFFFFC00000000007FFFFFFFFFF80000000000FFFFFFFFFFE00000000001FFFFFFFFFFC00000000003FFFFFFFFFFC00000000007FFFFFFFFFF800000000007FFFFFFFFFF80000000000";
defparam ram_block1a87.mem_init1 = "7FFFFFFFFFF800000000003FFFFFFFFFFC00000000003FFFFFFFFFFE00000000001FFFFFFFFFFF000000000007FFFFFFFFFF800000000003FFFFFFFFFFE00000000000FFFFFFFFFFFC00000000001FFFFFFFFFFF000000000003FFFFFFFFFFE000000000007FFFFFFFFFFE000000000007FFFFFFFFFFC000000000007FFFFFFFFFFE000000000007FFFFFFFFFFE000000000003FFFFFFFFFFF800000000001FFFFFFFFFFFC000000000007FFFFFFFFFFF000000000000FFFFFFFFFFFE000000000003FFFFFFFFFFFC000000000003FFFFFFFFFFFC000000000003FFFFFFFFFFFC000000000003FFFFFFFFFFFE000000000001FFFFFFFFFFFF0000000000007FF";
defparam ram_block1a87.mem_init0 = "FFFFFFFFFC000000000001FFFFFFFFFFFF0000000000003FFFFFFFFFFFF0000000000003FFFFFFFFFFFF0000000000003FFFFFFFFFFFF0000000000001FFFFFFFFFFFF8000000000000FFFFFFFFFFFFE0000000000001FFFFFFFFFFFFC0000000000003FFFFFFFFFFFFC0000000000003FFFFFFFFFFFFC0000000000001FFFFFFFFFFFFE0000000000000FFFFFFFFFFFFFC0000000000001FFFFFFFFFFFFF80000000000003FFFFFFFFFFFFF80000000000001FFFFFFFFFFFFFC0000000000000FFFFFFFFFFFFFF00000000000001FFFFFFFFFFFFFE00000000000001FFFFFFFFFFFFFE00000000000001FFFFFFFFFFFFFF000000000000007FFFFFFFFFFFFFE";

arriav_ram_block ram_block1a103(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a103_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a103.clk0_core_clock_enable = "ena0";
defparam ram_block1a103.clk0_input_clock_enable = "ena0";
defparam ram_block1a103.clk0_output_clock_enable = "ena0";
defparam ram_block1a103.data_interleave_offset_in_bits = 1;
defparam ram_block1a103.data_interleave_width_in_bits = 1;
defparam ram_block1a103.init_file = "DDS_48_v1_nco_ii_0_cos.hex";
defparam ram_block1a103.init_file_layout = "port_a";
defparam ram_block1a103.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0121|altsyncram:altsyncram_component0|altsyncram_78g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a103.operation_mode = "rom";
defparam ram_block1a103.port_a_address_clear = "none";
defparam ram_block1a103.port_a_address_width = 13;
defparam ram_block1a103.port_a_data_out_clear = "none";
defparam ram_block1a103.port_a_data_out_clock = "clock0";
defparam ram_block1a103.port_a_data_width = 1;
defparam ram_block1a103.port_a_first_address = 49152;
defparam ram_block1a103.port_a_first_bit_number = 7;
defparam ram_block1a103.port_a_last_address = 57343;
defparam ram_block1a103.port_a_logical_ram_depth = 65536;
defparam ram_block1a103.port_a_logical_ram_width = 16;
defparam ram_block1a103.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a103.ram_block_type = "auto";
defparam ram_block1a103.mem_init3 = "800000000000003FFFFFFFFFFFFFE00000000000000FFFFFFFFFFFFFF800000000000007FFFFFFFFFFFFF80000000000000FFFFFFFFFFFFFF00000000000001FFFFFFFFFFFFFC0000000000000FFFFFFFFFFFFFE00000000000007FFFFFFFFFFFFE0000000000000FFFFFFFFFFFFFC0000000000001FFFFFFFFFFFFF00000000000007FFFFFFFFFFFF80000000000003FFFFFFFFFFFFC0000000000003FFFFFFFFFFFF80000000000007FFFFFFFFFFFF0000000000001FFFFFFFFFFFFC0000000000007FFFFFFFFFFFE0000000000003FFFFFFFFFFFF0000000000003FFFFFFFFFFFF0000000000007FFFFFFFFFFFE000000000000FFFFFFFFFFFFC000000000";
defparam ram_block1a103.mem_init2 = "001FFFFFFFFFFFE000000000000FFFFFFFFFFFF8000000000007FFFFFFFFFFFC000000000003FFFFFFFFFFFC000000000003FFFFFFFFFFF8000000000007FFFFFFFFFFF000000000000FFFFFFFFFFFE000000000003FFFFFFFFFFF800000000000FFFFFFFFFFFE000000000007FFFFFFFFFFF000000000003FFFFFFFFFFF800000000001FFFFFFFFFFF800000000001FFFFFFFFFFF800000000003FFFFFFFFFFF000000000003FFFFFFFFFFE00000000000FFFFFFFFFFFC00000000001FFFFFFFFFFF000000000007FFFFFFFFFFC00000000001FFFFFFFFFFE00000000000FFFFFFFFFFF800000000007FFFFFFFFFF800000000003FFFFFFFFFFC00000000003";
defparam ram_block1a103.mem_init1 = "FFFFFFFFFFC00000000003FFFFFFFFFFC00000000003FFFFFFFFFFC00000000007FFFFFFFFFF800000000007FFFFFFFFFF00000000001FFFFFFFFFFE00000000003FFFFFFFFFF80000000000FFFFFFFFFFF00000000001FFFFFFFFFFC00000000007FFFFFFFFFE00000000003FFFFFFFFFF80000000000FFFFFFFFFFC00000000007FFFFFFFFFE00000000003FFFFFFFFFF00000000001FFFFFFFFFF80000000001FFFFFFFFFFC0000000000FFFFFFFFFFC0000000000FFFFFFFFFFC0000000000FFFFFFFFFFC0000000000FFFFFFFFFFC0000000000FFFFFFFFFFC0000000001FFFFFFFFFF80000000001FFFFFFFFFF00000000003FFFFFFFFFF00000000007";
defparam ram_block1a103.mem_init0 = "FFFFFFFFFE0000000000FFFFFFFFFFC0000000001FFFFFFFFFF80000000003FFFFFFFFFE00000000007FFFFFFFFFC0000000001FFFFFFFFFF00000000003FFFFFFFFFE0000000000FFFFFFFFFF80000000003FFFFFFFFFE0000000000FFFFFFFFFF80000000003FFFFFFFFFF00000000007FFFFFFFFF80000000003FFFFFFFFFE0000000000FFFFFFFFFF80000000003FFFFFFFFFE0000000000FFFFFFFFFF80000000003FFFFFFFFFC0000000001FFFFFFFFFF00000000007FFFFFFFFFC0000000001FFFFFFFFFE0000000000FFFFFFFFFF80000000003FFFFFFFFFC0000000001FFFFFFFFFF00000000007FFFFFFFFF80000000003FFFFFFFFFE0000000000";

arriav_ram_block ram_block1a119(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a119_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a119.clk0_core_clock_enable = "ena0";
defparam ram_block1a119.clk0_input_clock_enable = "ena0";
defparam ram_block1a119.clk0_output_clock_enable = "ena0";
defparam ram_block1a119.data_interleave_offset_in_bits = 1;
defparam ram_block1a119.data_interleave_width_in_bits = 1;
defparam ram_block1a119.init_file = "DDS_48_v1_nco_ii_0_cos.hex";
defparam ram_block1a119.init_file_layout = "port_a";
defparam ram_block1a119.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0121|altsyncram:altsyncram_component0|altsyncram_78g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a119.operation_mode = "rom";
defparam ram_block1a119.port_a_address_clear = "none";
defparam ram_block1a119.port_a_address_width = 13;
defparam ram_block1a119.port_a_data_out_clear = "none";
defparam ram_block1a119.port_a_data_out_clock = "clock0";
defparam ram_block1a119.port_a_data_width = 1;
defparam ram_block1a119.port_a_first_address = 57344;
defparam ram_block1a119.port_a_first_bit_number = 7;
defparam ram_block1a119.port_a_last_address = 65535;
defparam ram_block1a119.port_a_logical_ram_depth = 65536;
defparam ram_block1a119.port_a_logical_ram_width = 16;
defparam ram_block1a119.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a119.ram_block_type = "auto";
defparam ram_block1a119.mem_init3 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a119.mem_init2 = "FFFF00000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000";
defparam ram_block1a119.mem_init1 = "00000000000007FFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000007FFFFFFFFFFFFFFFFFFFFFF80000000000000000000001FFFFFFFFFFFFFFFFFFFFFF0000000000000000000001FFFFFFFFFFFFFFFFFFFFFC000000000000000000003FFFFFFFFFFFFFFFFFFFFC00000000000000000000FFFFFFFFFFFFFFFFFFFFC00000000000000000003FFFFFFFFFFFFFFFFFFF80000000000000000001FFFFFFFFFFFFFFFFFFF00000000000000000007FFFFFFFFFFFFFFFFFF0000000000000000001FFFFFFFFFFFFFFFFFF800";
defparam ram_block1a119.mem_init0 = "0000000000000003FFFFFFFFFFFFFFFFFC000000000000000003FFFFFFFFFFFFFFFFF800000000000000001FFFFFFFFFFFFFFFFF000000000000000007FFFFFFFFFFFFFFFFC00000000000000007FFFFFFFFFFFFFFFF80000000000000001FFFFFFFFFFFFFFFF80000000000000001FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFE0000000000000003FFFFFFFFFFFFFFF0000000000000003FFFFFFFFFFFFFFE000000000000000FFFFFFFFFFFFFFF8000000000000007FFFFFFFFFFFFFF800000000000000FFFFFFFFFFFFFFE000000000000003FFFFFFFFFFFFFF800000000000001FFFFFFFFFFFFFF";

arriav_ram_block ram_block1a39(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a39_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a39.clk0_core_clock_enable = "ena0";
defparam ram_block1a39.clk0_input_clock_enable = "ena0";
defparam ram_block1a39.clk0_output_clock_enable = "ena0";
defparam ram_block1a39.data_interleave_offset_in_bits = 1;
defparam ram_block1a39.data_interleave_width_in_bits = 1;
defparam ram_block1a39.init_file = "DDS_48_v1_nco_ii_0_cos.hex";
defparam ram_block1a39.init_file_layout = "port_a";
defparam ram_block1a39.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0121|altsyncram:altsyncram_component0|altsyncram_78g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a39.operation_mode = "rom";
defparam ram_block1a39.port_a_address_clear = "none";
defparam ram_block1a39.port_a_address_width = 13;
defparam ram_block1a39.port_a_data_out_clear = "none";
defparam ram_block1a39.port_a_data_out_clock = "clock0";
defparam ram_block1a39.port_a_data_width = 1;
defparam ram_block1a39.port_a_first_address = 16384;
defparam ram_block1a39.port_a_first_bit_number = 7;
defparam ram_block1a39.port_a_last_address = 24575;
defparam ram_block1a39.port_a_logical_ram_depth = 65536;
defparam ram_block1a39.port_a_logical_ram_width = 16;
defparam ram_block1a39.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a39.ram_block_type = "auto";
defparam ram_block1a39.mem_init3 = "FFFFFFFFFFFFFFC00000000000001FFFFFFFFFFFFFF00000000000000FFFFFFFFFFFFFF00000000000000FFFFFFFFFFFFFF00000000000001FFFFFFFFFFFFFE00000000000007FFFFFFFFFFFFF00000000000003FFFFFFFFFFFFF80000000000003FFFFFFFFFFFFF00000000000007FFFFFFFFFFFFE0000000000000FFFFFFFFFFFFF00000000000007FFFFFFFFFFFF80000000000007FFFFFFFFFFFF80000000000007FFFFFFFFFFFF0000000000000FFFFFFFFFFFFE0000000000003FFFFFFFFFFFF0000000000001FFFFFFFFFFFF8000000000001FFFFFFFFFFFF8000000000001FFFFFFFFFFFF8000000000001FFFFFFFFFFFF0000000000007FFFFFFFFF";
defparam ram_block1a39.mem_init2 = "FFC000000000001FFFFFFFFFFFF000000000000FFFFFFFFFFFF8000000000007FFFFFFFFFFF8000000000007FFFFFFFFFFF8000000000007FFFFFFFFFFF800000000000FFFFFFFFFFFE000000000001FFFFFFFFFFFC000000000007FFFFFFFFFFF000000000003FFFFFFFFFFF800000000000FFFFFFFFFFFC00000000000FFFFFFFFFFFC000000000007FFFFFFFFFFC00000000000FFFFFFFFFFFC00000000000FFFFFFFFFFF800000000001FFFFFFFFFFF000000000007FFFFFFFFFFE00000000000FFFFFFFFFFF800000000003FFFFFFFFFFC00000000001FFFFFFFFFFF00000000000FFFFFFFFFFF800000000007FFFFFFFFFF800000000003FFFFFFFFFFC";
defparam ram_block1a39.mem_init1 = "00000000003FFFFFFFFFFC00000000003FFFFFFFFFFC00000000007FFFFFFFFFF800000000007FFFFFFFFFF00000000000FFFFFFFFFFE00000000003FFFFFFFFFFC00000000007FFFFFFFFFF00000000001FFFFFFFFFFC00000000007FFFFFFFFFF00000000001FFFFFFFFFFC00000000007FFFFFFFFFE00000000003FFFFFFFFFF80000000001FFFFFFFFFFC0000000000FFFFFFFFFFC00000000007FFFFFFFFFE00000000007FFFFFFFFFE00000000003FFFFFFFFFF00000000003FFFFFFFFFF00000000003FFFFFFFFFF00000000003FFFFFFFFFE00000000007FFFFFFFFFE00000000007FFFFFFFFFC0000000000FFFFFFFFFFC0000000001FFFFFFFFFF8";
defparam ram_block1a39.mem_init0 = "0000000003FFFFFFFFFF00000000007FFFFFFFFFE0000000000FFFFFFFFFFC0000000001FFFFFFFFFF00000000003FFFFFFFFFE0000000000FFFFFFFFFF80000000003FFFFFFFFFF00000000007FFFFFFFFFC0000000001FFFFFFFFFF00000000007FFFFFFFFFC0000000001FFFFFFFFFF00000000007FFFFFFFFFC0000000001FFFFFFFFFF00000000007FFFFFFFFFC0000000001FFFFFFFFFF0000000000FFFFFFFFFF80000000003FFFFFFFFFE0000000000FFFFFFFFFF80000000007FFFFFFFFFC0000000001FFFFFFFFFF00000000007FFFFFFFFF80000000003FFFFFFFFFE0000000000FFFFFFFFFF00000000007FFFFFFFFFC0000000001FFFFFFFFFE";

arriav_ram_block ram_block1a55(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a55_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a55.clk0_core_clock_enable = "ena0";
defparam ram_block1a55.clk0_input_clock_enable = "ena0";
defparam ram_block1a55.clk0_output_clock_enable = "ena0";
defparam ram_block1a55.data_interleave_offset_in_bits = 1;
defparam ram_block1a55.data_interleave_width_in_bits = 1;
defparam ram_block1a55.init_file = "DDS_48_v1_nco_ii_0_cos.hex";
defparam ram_block1a55.init_file_layout = "port_a";
defparam ram_block1a55.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0121|altsyncram:altsyncram_component0|altsyncram_78g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a55.operation_mode = "rom";
defparam ram_block1a55.port_a_address_clear = "none";
defparam ram_block1a55.port_a_address_width = 13;
defparam ram_block1a55.port_a_data_out_clear = "none";
defparam ram_block1a55.port_a_data_out_clock = "clock0";
defparam ram_block1a55.port_a_data_width = 1;
defparam ram_block1a55.port_a_first_address = 24576;
defparam ram_block1a55.port_a_first_bit_number = 7;
defparam ram_block1a55.port_a_last_address = 32767;
defparam ram_block1a55.port_a_logical_ram_depth = 65536;
defparam ram_block1a55.port_a_logical_ram_width = 16;
defparam ram_block1a55.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a55.ram_block_type = "auto";
defparam ram_block1a55.mem_init3 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000000000000000000000000000000";
defparam ram_block1a55.mem_init2 = "0003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000003FFFFFFFFFFFFF";
defparam ram_block1a55.mem_init1 = "FFFFFFFFFFFFF800000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000FFFFFFFFFFFFFFFFFFFFFFC0000000000000000000001FFFFFFFFFFFFFFFFFFFFFE0000000000000000000007FFFFFFFFFFFFFFFFFFFFC000000000000000000007FFFFFFFFFFFFFFFFFFFF000000000000000000007FFFFFFFFFFFFFFFFFFF80000000000000000000FFFFFFFFFFFFFFFFFFFE0000000000000000000FFFFFFFFFFFFFFFFFFF0000000000000000000FFFFFFFFFFFFFFFFFFC000000000000000000FFF";
defparam ram_block1a55.mem_init0 = "FFFFFFFFFFFFFFF8000000000000000003FFFFFFFFFFFFFFFFF800000000000000000FFFFFFFFFFFFFFFFFC00000000000000000FFFFFFFFFFFFFFFFF800000000000000007FFFFFFFFFFFFFFFF80000000000000000FFFFFFFFFFFFFFFFE00000000000000007FFFFFFFFFFFFFFFC0000000000000001FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFE0000000000000001FFFFFFFFFFFFFFF8000000000000001FFFFFFFFFFFFFFF8000000000000001FFFFFFFFFFFFFFF000000000000000FFFFFFFFFFFFFFF800000000000000FFFFFFFFFFFFFFF000000000000001FFFFFFFFFFFFFFC00000000000000FFFFFFFFFFFFFFC00000000000000";

arriav_ram_block ram_block1a7(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a7_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.clk0_input_clock_enable = "ena0";
defparam ram_block1a7.clk0_output_clock_enable = "ena0";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.init_file = "DDS_48_v1_nco_ii_0_cos.hex";
defparam ram_block1a7.init_file_layout = "port_a";
defparam ram_block1a7.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0121|altsyncram:altsyncram_component0|altsyncram_78g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.operation_mode = "rom";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 13;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "clock0";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 8191;
defparam ram_block1a7.port_a_logical_ram_depth = 65536;
defparam ram_block1a7.port_a_logical_ram_width = 16;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.ram_block_type = "auto";
defparam ram_block1a7.mem_init3 = "FFFFFFFFFFFFFF000000000000003FFFFFFFFFFFFFF800000000000000FFFFFFFFFFFFFFE000000000000003FFFFFFFFFFFFFFC000000000000003FFFFFFFFFFFFFFE000000000000000FFFFFFFFFFFFFFF8000000000000001FFFFFFFFFFFFFFF8000000000000000FFFFFFFFFFFFFFFE0000000000000001FFFFFFFFFFFFFFFE0000000000000001FFFFFFFFFFFFFFFF00000000000000003FFFFFFFFFFFFFFFF00000000000000003FFFFFFFFFFFFFFFFC00000000000000007FFFFFFFFFFFFFFFFC00000000000000001FFFFFFFFFFFFFFFFF000000000000000003FFFFFFFFFFFFFFFFF8000000000000000007FFFFFFFFFFFFFFFFF8000000000000000";
defparam ram_block1a7.mem_init2 = "003FFFFFFFFFFFFFFFFFF0000000000000000001FFFFFFFFFFFFFFFFFFC0000000000000000001FFFFFFFFFFFFFFFFFFF00000000000000000003FFFFFFFFFFFFFFFFFFF800000000000000000007FFFFFFFFFFFFFFFFFFFE000000000000000000007FFFFFFFFFFFFFFFFFFFF8000000000000000000007FFFFFFFFFFFFFFFFFFFFF0000000000000000000001FFFFFFFFFFFFFFFFFFFFFF00000000000000000000003FFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000";
defparam ram_block1a7.mem_init1 = "0000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000000000000000000000000001FFFF";
defparam ram_block1a7.mem_init0 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

arriav_ram_block ram_block1a23(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a23_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a23.clk0_core_clock_enable = "ena0";
defparam ram_block1a23.clk0_input_clock_enable = "ena0";
defparam ram_block1a23.clk0_output_clock_enable = "ena0";
defparam ram_block1a23.data_interleave_offset_in_bits = 1;
defparam ram_block1a23.data_interleave_width_in_bits = 1;
defparam ram_block1a23.init_file = "DDS_48_v1_nco_ii_0_cos.hex";
defparam ram_block1a23.init_file_layout = "port_a";
defparam ram_block1a23.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0121|altsyncram:altsyncram_component0|altsyncram_78g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a23.operation_mode = "rom";
defparam ram_block1a23.port_a_address_clear = "none";
defparam ram_block1a23.port_a_address_width = 13;
defparam ram_block1a23.port_a_data_out_clear = "none";
defparam ram_block1a23.port_a_data_out_clock = "clock0";
defparam ram_block1a23.port_a_data_width = 1;
defparam ram_block1a23.port_a_first_address = 8192;
defparam ram_block1a23.port_a_first_bit_number = 7;
defparam ram_block1a23.port_a_last_address = 16383;
defparam ram_block1a23.port_a_logical_ram_depth = 65536;
defparam ram_block1a23.port_a_logical_ram_width = 16;
defparam ram_block1a23.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a23.ram_block_type = "auto";
defparam ram_block1a23.mem_init3 = "0000000000FFFFFFFFFF80000000003FFFFFFFFFC0000000001FFFFFFFFFF00000000007FFFFFFFFF80000000003FFFFFFFFFE0000000000FFFFFFFFFF00000000007FFFFFFFFFC0000000001FFFFFFFFFF00000000007FFFFFFFFF80000000003FFFFFFFFFE0000000000FFFFFFFFFF80000000003FFFFFFFFFE0000000000FFFFFFFFFF80000000003FFFFFFFFFC0000000001FFFFFFFFFF80000000003FFFFFFFFFE0000000000FFFFFFFFFF80000000003FFFFFFFFFE0000000000FFFFFFFFFF80000000001FFFFFFFFFF00000000007FFFFFFFFFC0000000000FFFFFFFFFF80000000003FFFFFFFFFF00000000007FFFFFFFFFE0000000000FFFFFFFFFF";
defparam ram_block1a23.mem_init2 = "C0000000001FFFFFFFFFF80000000001FFFFFFFFFF00000000003FFFFFFFFFF00000000007FFFFFFFFFE00000000007FFFFFFFFFE00000000007FFFFFFFFFE00000000007FFFFFFFFFE00000000007FFFFFFFFFE00000000007FFFFFFFFFF00000000003FFFFFFFFFF00000000001FFFFFFFFFF80000000000FFFFFFFFFFC00000000007FFFFFFFFFE00000000003FFFFFFFFFF80000000000FFFFFFFFFFC00000000007FFFFFFFFFF00000000001FFFFFFFFFFE00000000003FFFFFFFFFF80000000000FFFFFFFFFFF00000000001FFFFFFFFFFC00000000003FFFFFFFFFFC00000000007FFFFFFFFFF800000000007FFFFFFFFFF800000000007FFFFFFFFFF";
defparam ram_block1a23.mem_init1 = "800000000007FFFFFFFFFF800000000003FFFFFFFFFFC00000000003FFFFFFFFFFE00000000000FFFFFFFFFFF000000000007FFFFFFFFFFC00000000001FFFFFFFFFFF000000000007FFFFFFFFFFE00000000000FFFFFFFFFFF800000000001FFFFFFFFFFF800000000003FFFFFFFFFFF000000000003FFFFFFFFFFF000000000003FFFFFFFFFFF800000000001FFFFFFFFFFFC00000000000FFFFFFFFFFFE000000000003FFFFFFFFFFF800000000000FFFFFFFFFFFE000000000001FFFFFFFFFFFC000000000003FFFFFFFFFFF8000000000007FFFFFFFFFFF8000000000007FFFFFFFFFFFC000000000003FFFFFFFFFFFE000000000000FFFFFFFFFFFF000";
defparam ram_block1a23.mem_init0 = "0000000007FFFFFFFFFFFE000000000000FFFFFFFFFFFFC000000000001FFFFFFFFFFFF8000000000001FFFFFFFFFFFF8000000000000FFFFFFFFFFFFC0000000000007FFFFFFFFFFFF0000000000001FFFFFFFFFFFFC0000000000003FFFFFFFFFFFF80000000000007FFFFFFFFFFFF80000000000003FFFFFFFFFFFFC0000000000001FFFFFFFFFFFFF00000000000007FFFFFFFFFFFFE0000000000000FFFFFFFFFFFFFC0000000000000FFFFFFFFFFFFFE00000000000007FFFFFFFFFFFFF00000000000001FFFFFFFFFFFFFE00000000000003FFFFFFFFFFFFFC00000000000003FFFFFFFFFFFFFE00000000000000FFFFFFFFFFFFFF800000000000003";

arriav_ram_block ram_block1a72(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a72_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a72.clk0_core_clock_enable = "ena0";
defparam ram_block1a72.clk0_input_clock_enable = "ena0";
defparam ram_block1a72.clk0_output_clock_enable = "ena0";
defparam ram_block1a72.data_interleave_offset_in_bits = 1;
defparam ram_block1a72.data_interleave_width_in_bits = 1;
defparam ram_block1a72.init_file = "DDS_48_v1_nco_ii_0_cos.hex";
defparam ram_block1a72.init_file_layout = "port_a";
defparam ram_block1a72.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0121|altsyncram:altsyncram_component0|altsyncram_78g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a72.operation_mode = "rom";
defparam ram_block1a72.port_a_address_clear = "none";
defparam ram_block1a72.port_a_address_width = 13;
defparam ram_block1a72.port_a_data_out_clear = "none";
defparam ram_block1a72.port_a_data_out_clock = "clock0";
defparam ram_block1a72.port_a_data_width = 1;
defparam ram_block1a72.port_a_first_address = 32768;
defparam ram_block1a72.port_a_first_bit_number = 8;
defparam ram_block1a72.port_a_last_address = 40959;
defparam ram_block1a72.port_a_logical_ram_depth = 65536;
defparam ram_block1a72.port_a_logical_ram_width = 16;
defparam ram_block1a72.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a72.ram_block_type = "auto";
defparam ram_block1a72.mem_init3 = "FFFFFFFFFFFFFF800000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000000000003FFFFFFFFFFFFFFF";
defparam ram_block1a72.mem_init2 = "FFFFFFFFFFFFFFFFFFFFF80000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000000003FFFFFFFFFFFFF";
defparam ram_block1a72.mem_init1 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000000000000000000000";
defparam ram_block1a72.mem_init0 = "000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

arriav_ram_block ram_block1a88(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a88_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a88.clk0_core_clock_enable = "ena0";
defparam ram_block1a88.clk0_input_clock_enable = "ena0";
defparam ram_block1a88.clk0_output_clock_enable = "ena0";
defparam ram_block1a88.data_interleave_offset_in_bits = 1;
defparam ram_block1a88.data_interleave_width_in_bits = 1;
defparam ram_block1a88.init_file = "DDS_48_v1_nco_ii_0_cos.hex";
defparam ram_block1a88.init_file_layout = "port_a";
defparam ram_block1a88.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0121|altsyncram:altsyncram_component0|altsyncram_78g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a88.operation_mode = "rom";
defparam ram_block1a88.port_a_address_clear = "none";
defparam ram_block1a88.port_a_address_width = 13;
defparam ram_block1a88.port_a_data_out_clear = "none";
defparam ram_block1a88.port_a_data_out_clock = "clock0";
defparam ram_block1a88.port_a_data_width = 1;
defparam ram_block1a88.port_a_first_address = 40960;
defparam ram_block1a88.port_a_first_bit_number = 8;
defparam ram_block1a88.port_a_last_address = 49151;
defparam ram_block1a88.port_a_logical_ram_depth = 65536;
defparam ram_block1a88.port_a_logical_ram_width = 16;
defparam ram_block1a88.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a88.ram_block_type = "auto";
defparam ram_block1a88.mem_init3 = "FFFFFFFFFFFFFFFFFFFF800000000000000000001FFFFFFFFFFFFFFFFFFFF000000000000000000003FFFFFFFFFFFFFFFFFFFE000000000000000000007FFFFFFFFFFFFFFFFFFFC00000000000000000000FFFFFFFFFFFFFFFFFFFFC00000000000000000001FFFFFFFFFFFFFFFFFFFF800000000000000000001FFFFFFFFFFFFFFFFFFFF800000000000000000001FFFFFFFFFFFFFFFFFFFF800000000000000000001FFFFFFFFFFFFFFFFFFFF800000000000000000001FFFFFFFFFFFFFFFFFFFFC00000000000000000000FFFFFFFFFFFFFFFFFFFFE000000000000000000007FFFFFFFFFFFFFFFFFFFF000000000000000000001FFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a88.mem_init2 = "C000000000000000000007FFFFFFFFFFFFFFFFFFFF800000000000000000000FFFFFFFFFFFFFFFFFFFFF000000000000000000001FFFFFFFFFFFFFFFFFFFFE000000000000000000001FFFFFFFFFFFFFFFFFFFFF000000000000000000000FFFFFFFFFFFFFFFFFFFFF8000000000000000000007FFFFFFFFFFFFFFFFFFFFC000000000000000000000FFFFFFFFFFFFFFFFFFFFF8000000000000000000001FFFFFFFFFFFFFFFFFFFFF8000000000000000000001FFFFFFFFFFFFFFFFFFFFF8000000000000000000000FFFFFFFFFFFFFFFFFFFFFE0000000000000000000003FFFFFFFFFFFFFFFFFFFFF80000000000000000000007FFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a88.mem_init1 = "80000000000000000000003FFFFFFFFFFFFFFFFFFFFFC0000000000000000000001FFFFFFFFFFFFFFFFFFFFFF80000000000000000000003FFFFFFFFFFFFFFFFFFFFFF00000000000000000000001FFFFFFFFFFFFFFFFFFFFFFC00000000000000000000007FFFFFFFFFFFFFFFFFFFFFF800000000000000000000007FFFFFFFFFFFFFFFFFFFFFF800000000000000000000003FFFFFFFFFFFFFFFFFFFFFFE000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFF000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFF800";
defparam ram_block1a88.mem_init0 = "0000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000007FFFFFFFFFFFFFF";

arriav_ram_block ram_block1a104(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a104_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a104.clk0_core_clock_enable = "ena0";
defparam ram_block1a104.clk0_input_clock_enable = "ena0";
defparam ram_block1a104.clk0_output_clock_enable = "ena0";
defparam ram_block1a104.data_interleave_offset_in_bits = 1;
defparam ram_block1a104.data_interleave_width_in_bits = 1;
defparam ram_block1a104.init_file = "DDS_48_v1_nco_ii_0_cos.hex";
defparam ram_block1a104.init_file_layout = "port_a";
defparam ram_block1a104.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0121|altsyncram:altsyncram_component0|altsyncram_78g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a104.operation_mode = "rom";
defparam ram_block1a104.port_a_address_clear = "none";
defparam ram_block1a104.port_a_address_width = 13;
defparam ram_block1a104.port_a_data_out_clear = "none";
defparam ram_block1a104.port_a_data_out_clock = "clock0";
defparam ram_block1a104.port_a_data_width = 1;
defparam ram_block1a104.port_a_first_address = 49152;
defparam ram_block1a104.port_a_first_bit_number = 8;
defparam ram_block1a104.port_a_last_address = 57343;
defparam ram_block1a104.port_a_logical_ram_depth = 65536;
defparam ram_block1a104.port_a_logical_ram_width = 16;
defparam ram_block1a104.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a104.ram_block_type = "auto";
defparam ram_block1a104.mem_init3 = "000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000FFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a104.mem_init2 = "FFE000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFF000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFF000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFC00000000000000000000001FFFFFFFFFFFFFFFFFFFFFFE00000000000000000000003FFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000FFFFFFFFFFFFFFFFFFFFFFE00000000000000000000007FFFFFFFFFFFFFFFFFFFFFE0000000000000000000000FFFFFFFFFFFFFFFFFFFFFF80000000000000000000003FFFFFFFFFFFFFFFFFFFFFC";
defparam ram_block1a104.mem_init1 = "0000000000000000000003FFFFFFFFFFFFFFFFFFFFFC0000000000000000000007FFFFFFFFFFFFFFFFFFFFF8000000000000000000001FFFFFFFFFFFFFFFFFFFFFC000000000000000000000FFFFFFFFFFFFFFFFFFFFFE0000000000000000000007FFFFFFFFFFFFFFFFFFFFC000000000000000000000FFFFFFFFFFFFFFFFFFFFF8000000000000000000003FFFFFFFFFFFFFFFFFFFFE000000000000000000001FFFFFFFFFFFFFFFFFFFFF000000000000000000000FFFFFFFFFFFFFFFFFFFFF000000000000000000000FFFFFFFFFFFFFFFFFFFFF000000000000000000001FFFFFFFFFFFFFFFFFFFFE000000000000000000003FFFFFFFFFFFFFFFFFFFF8";
defparam ram_block1a104.mem_init0 = "00000000000000000000FFFFFFFFFFFFFFFFFFFFE000000000000000000003FFFFFFFFFFFFFFFFFFFF800000000000000000001FFFFFFFFFFFFFFFFFFFFC00000000000000000000FFFFFFFFFFFFFFFFFFFFC00000000000000000000FFFFFFFFFFFFFFFFFFFFC000000000000000000007FFFFFFFFFFFFFFFFFFFC00000000000000000000FFFFFFFFFFFFFFFFFFFFC00000000000000000000FFFFFFFFFFFFFFFFFFFFC00000000000000000001FFFFFFFFFFFFFFFFFFFF800000000000000000001FFFFFFFFFFFFFFFFFFFF000000000000000000003FFFFFFFFFFFFFFFFFFFE000000000000000000007FFFFFFFFFFFFFFFFFFFC00000000000000000000";

arriav_ram_block ram_block1a120(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a120_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a120.clk0_core_clock_enable = "ena0";
defparam ram_block1a120.clk0_input_clock_enable = "ena0";
defparam ram_block1a120.clk0_output_clock_enable = "ena0";
defparam ram_block1a120.data_interleave_offset_in_bits = 1;
defparam ram_block1a120.data_interleave_width_in_bits = 1;
defparam ram_block1a120.init_file = "DDS_48_v1_nco_ii_0_cos.hex";
defparam ram_block1a120.init_file_layout = "port_a";
defparam ram_block1a120.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0121|altsyncram:altsyncram_component0|altsyncram_78g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a120.operation_mode = "rom";
defparam ram_block1a120.port_a_address_clear = "none";
defparam ram_block1a120.port_a_address_width = 13;
defparam ram_block1a120.port_a_data_out_clear = "none";
defparam ram_block1a120.port_a_data_out_clock = "clock0";
defparam ram_block1a120.port_a_data_width = 1;
defparam ram_block1a120.port_a_first_address = 57344;
defparam ram_block1a120.port_a_first_bit_number = 8;
defparam ram_block1a120.port_a_last_address = 65535;
defparam ram_block1a120.port_a_logical_ram_depth = 65536;
defparam ram_block1a120.port_a_logical_ram_width = 16;
defparam ram_block1a120.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a120.ram_block_type = "auto";
defparam ram_block1a120.mem_init3 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a120.mem_init2 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000000000000000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000000000000000000";
defparam ram_block1a120.mem_init1 = "00000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000";
defparam ram_block1a120.mem_init0 = "0000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000";

arriav_ram_block ram_block1a40(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a40_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a40.clk0_core_clock_enable = "ena0";
defparam ram_block1a40.clk0_input_clock_enable = "ena0";
defparam ram_block1a40.clk0_output_clock_enable = "ena0";
defparam ram_block1a40.data_interleave_offset_in_bits = 1;
defparam ram_block1a40.data_interleave_width_in_bits = 1;
defparam ram_block1a40.init_file = "DDS_48_v1_nco_ii_0_cos.hex";
defparam ram_block1a40.init_file_layout = "port_a";
defparam ram_block1a40.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0121|altsyncram:altsyncram_component0|altsyncram_78g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a40.operation_mode = "rom";
defparam ram_block1a40.port_a_address_clear = "none";
defparam ram_block1a40.port_a_address_width = 13;
defparam ram_block1a40.port_a_data_out_clear = "none";
defparam ram_block1a40.port_a_data_out_clock = "clock0";
defparam ram_block1a40.port_a_data_width = 1;
defparam ram_block1a40.port_a_first_address = 16384;
defparam ram_block1a40.port_a_first_bit_number = 8;
defparam ram_block1a40.port_a_last_address = 24575;
defparam ram_block1a40.port_a_logical_ram_depth = 65536;
defparam ram_block1a40.port_a_logical_ram_width = 16;
defparam ram_block1a40.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a40.ram_block_type = "auto";
defparam ram_block1a40.mem_init3 = "FFFFFFFFFFFFFFC0000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000";
defparam ram_block1a40.mem_init2 = "003FFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFF800000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000FFFFFFFFFFFFFFFFFFFFFFF800000000000000000000003FFFFFFFFFFFFFFFFFFFFFFC00000000000000000000003FFFFFFFFFFFFFFFFFFFFFFC00000000000000000000007FFFFFFFFFFFFFFFFFFFFFF00000000000000000000001FFFFFFFFFFFFFFFFFFFFFF80000000000000000000003FFFFFFFFFFFFFFFFFFFFFF00000000000000000000007FFFFFFFFFFFFFFFFFFFFF80000000000000000000003";
defparam ram_block1a40.mem_init1 = "FFFFFFFFFFFFFFFFFFFFFC0000000000000000000003FFFFFFFFFFFFFFFFFFFFF8000000000000000000000FFFFFFFFFFFFFFFFFFFFFE0000000000000000000003FFFFFFFFFFFFFFFFFFFFF0000000000000000000003FFFFFFFFFFFFFFFFFFFFF0000000000000000000003FFFFFFFFFFFFFFFFFFFFE0000000000000000000007FFFFFFFFFFFFFFFFFFFFC000000000000000000003FFFFFFFFFFFFFFFFFFFFE000000000000000000001FFFFFFFFFFFFFFFFFFFFF000000000000000000000FFFFFFFFFFFFFFFFFFFFF000000000000000000001FFFFFFFFFFFFFFFFFFFFE000000000000000000003FFFFFFFFFFFFFFFFFFFFC000000000000000000007";
defparam ram_block1a40.mem_init0 = "FFFFFFFFFFFFFFFFFFFF000000000000000000001FFFFFFFFFFFFFFFFFFFFC00000000000000000000FFFFFFFFFFFFFFFFFFFFE000000000000000000007FFFFFFFFFFFFFFFFFFFF000000000000000000003FFFFFFFFFFFFFFFFFFFF000000000000000000003FFFFFFFFFFFFFFFFFFFF000000000000000000003FFFFFFFFFFFFFFFFFFFF000000000000000000003FFFFFFFFFFFFFFFFFFFF000000000000000000007FFFFFFFFFFFFFFFFFFFE000000000000000000007FFFFFFFFFFFFFFFFFFFC00000000000000000000FFFFFFFFFFFFFFFFFFFF800000000000000000001FFFFFFFFFFFFFFFFFFFF000000000000000000003FFFFFFFFFFFFFFFFFFFE";

arriav_ram_block ram_block1a56(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a56_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a56.clk0_core_clock_enable = "ena0";
defparam ram_block1a56.clk0_input_clock_enable = "ena0";
defparam ram_block1a56.clk0_output_clock_enable = "ena0";
defparam ram_block1a56.data_interleave_offset_in_bits = 1;
defparam ram_block1a56.data_interleave_width_in_bits = 1;
defparam ram_block1a56.init_file = "DDS_48_v1_nco_ii_0_cos.hex";
defparam ram_block1a56.init_file_layout = "port_a";
defparam ram_block1a56.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0121|altsyncram:altsyncram_component0|altsyncram_78g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a56.operation_mode = "rom";
defparam ram_block1a56.port_a_address_clear = "none";
defparam ram_block1a56.port_a_address_width = 13;
defparam ram_block1a56.port_a_data_out_clear = "none";
defparam ram_block1a56.port_a_data_out_clock = "clock0";
defparam ram_block1a56.port_a_data_width = 1;
defparam ram_block1a56.port_a_first_address = 24576;
defparam ram_block1a56.port_a_first_bit_number = 8;
defparam ram_block1a56.port_a_last_address = 32767;
defparam ram_block1a56.port_a_logical_ram_depth = 65536;
defparam ram_block1a56.port_a_logical_ram_width = 16;
defparam ram_block1a56.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a56.ram_block_type = "auto";
defparam ram_block1a56.mem_init3 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000000000000000000000000000000";
defparam ram_block1a56.mem_init2 = "00000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a56.mem_init1 = "FFFFFFFFFFFFF8000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a56.mem_init0 = "FFFFFFFFFFFFFFF8000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000003FFFFFFFFFFFFFF";

arriav_ram_block ram_block1a8(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a8_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a8.clk0_core_clock_enable = "ena0";
defparam ram_block1a8.clk0_input_clock_enable = "ena0";
defparam ram_block1a8.clk0_output_clock_enable = "ena0";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.init_file = "DDS_48_v1_nco_ii_0_cos.hex";
defparam ram_block1a8.init_file_layout = "port_a";
defparam ram_block1a8.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0121|altsyncram:altsyncram_component0|altsyncram_78g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a8.operation_mode = "rom";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 13;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "clock0";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 8191;
defparam ram_block1a8.port_a_logical_ram_depth = 65536;
defparam ram_block1a8.port_a_logical_ram_width = 16;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a8.ram_block_type = "auto";
defparam ram_block1a8.mem_init3 = "00000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000";
defparam ram_block1a8.mem_init2 = "000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000";
defparam ram_block1a8.mem_init1 = "00000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000000000000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a8.mem_init0 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

arriav_ram_block ram_block1a24(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a24_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a24.clk0_core_clock_enable = "ena0";
defparam ram_block1a24.clk0_input_clock_enable = "ena0";
defparam ram_block1a24.clk0_output_clock_enable = "ena0";
defparam ram_block1a24.data_interleave_offset_in_bits = 1;
defparam ram_block1a24.data_interleave_width_in_bits = 1;
defparam ram_block1a24.init_file = "DDS_48_v1_nco_ii_0_cos.hex";
defparam ram_block1a24.init_file_layout = "port_a";
defparam ram_block1a24.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0121|altsyncram:altsyncram_component0|altsyncram_78g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a24.operation_mode = "rom";
defparam ram_block1a24.port_a_address_clear = "none";
defparam ram_block1a24.port_a_address_width = 13;
defparam ram_block1a24.port_a_data_out_clear = "none";
defparam ram_block1a24.port_a_data_out_clock = "clock0";
defparam ram_block1a24.port_a_data_width = 1;
defparam ram_block1a24.port_a_first_address = 8192;
defparam ram_block1a24.port_a_first_bit_number = 8;
defparam ram_block1a24.port_a_last_address = 16383;
defparam ram_block1a24.port_a_logical_ram_depth = 65536;
defparam ram_block1a24.port_a_logical_ram_width = 16;
defparam ram_block1a24.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a24.ram_block_type = "auto";
defparam ram_block1a24.mem_init3 = "000000000000000000007FFFFFFFFFFFFFFFFFFFC00000000000000000000FFFFFFFFFFFFFFFFFFFF800000000000000000001FFFFFFFFFFFFFFFFFFFF000000000000000000003FFFFFFFFFFFFFFFFFFFF000000000000000000007FFFFFFFFFFFFFFFFFFFE000000000000000000007FFFFFFFFFFFFFFFFFFFE000000000000000000007FFFFFFFFFFFFFFFFFFFC000000000000000000007FFFFFFFFFFFFFFFFFFFE000000000000000000007FFFFFFFFFFFFFFFFFFFE000000000000000000007FFFFFFFFFFFFFFFFFFFF000000000000000000003FFFFFFFFFFFFFFFFFFFF800000000000000000000FFFFFFFFFFFFFFFFFFFFE00000000000000000000";
defparam ram_block1a24.mem_init2 = "3FFFFFFFFFFFFFFFFFFFF800000000000000000000FFFFFFFFFFFFFFFFFFFFF000000000000000000001FFFFFFFFFFFFFFFFFFFFE000000000000000000001FFFFFFFFFFFFFFFFFFFFE000000000000000000001FFFFFFFFFFFFFFFFFFFFF000000000000000000000FFFFFFFFFFFFFFFFFFFFF8000000000000000000003FFFFFFFFFFFFFFFFFFFFE0000000000000000000007FFFFFFFFFFFFFFFFFFFFC000000000000000000000FFFFFFFFFFFFFFFFFFFFFE0000000000000000000007FFFFFFFFFFFFFFFFFFFFF0000000000000000000003FFFFFFFFFFFFFFFFFFFFFC0000000000000000000007FFFFFFFFFFFFFFFFFFFFF8000000000000000000000";
defparam ram_block1a24.mem_init1 = "7FFFFFFFFFFFFFFFFFFFFF80000000000000000000003FFFFFFFFFFFFFFFFFFFFFE0000000000000000000000FFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000FFFFFFFFFFFFFFFFFFFFFFE00000000000000000000007FFFFFFFFFFFFFFFFFFFFFF80000000000000000000000FFFFFFFFFFFFFFFFFFFFFFF000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFC00000000000000000000001FFFFFFFFFFFFFFFFFFFFFFF800000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000FFF";
defparam ram_block1a24.mem_init0 = "FFFFFFFFFFFFFFFFFFFFFE0000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000";

arriav_ram_block ram_block1a73(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a73_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a73.clk0_core_clock_enable = "ena0";
defparam ram_block1a73.clk0_input_clock_enable = "ena0";
defparam ram_block1a73.clk0_output_clock_enable = "ena0";
defparam ram_block1a73.data_interleave_offset_in_bits = 1;
defparam ram_block1a73.data_interleave_width_in_bits = 1;
defparam ram_block1a73.init_file = "DDS_48_v1_nco_ii_0_cos.hex";
defparam ram_block1a73.init_file_layout = "port_a";
defparam ram_block1a73.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0121|altsyncram:altsyncram_component0|altsyncram_78g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a73.operation_mode = "rom";
defparam ram_block1a73.port_a_address_clear = "none";
defparam ram_block1a73.port_a_address_width = 13;
defparam ram_block1a73.port_a_data_out_clear = "none";
defparam ram_block1a73.port_a_data_out_clock = "clock0";
defparam ram_block1a73.port_a_data_width = 1;
defparam ram_block1a73.port_a_first_address = 32768;
defparam ram_block1a73.port_a_first_bit_number = 9;
defparam ram_block1a73.port_a_last_address = 40959;
defparam ram_block1a73.port_a_logical_ram_depth = 65536;
defparam ram_block1a73.port_a_logical_ram_width = 16;
defparam ram_block1a73.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a73.ram_block_type = "auto";
defparam ram_block1a73.mem_init3 = "00000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000";
defparam ram_block1a73.mem_init2 = "00000000000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000000000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000";
defparam ram_block1a73.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a73.mem_init0 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

arriav_ram_block ram_block1a89(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a89_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a89.clk0_core_clock_enable = "ena0";
defparam ram_block1a89.clk0_input_clock_enable = "ena0";
defparam ram_block1a89.clk0_output_clock_enable = "ena0";
defparam ram_block1a89.data_interleave_offset_in_bits = 1;
defparam ram_block1a89.data_interleave_width_in_bits = 1;
defparam ram_block1a89.init_file = "DDS_48_v1_nco_ii_0_cos.hex";
defparam ram_block1a89.init_file_layout = "port_a";
defparam ram_block1a89.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0121|altsyncram:altsyncram_component0|altsyncram_78g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a89.operation_mode = "rom";
defparam ram_block1a89.port_a_address_clear = "none";
defparam ram_block1a89.port_a_address_width = 13;
defparam ram_block1a89.port_a_data_out_clear = "none";
defparam ram_block1a89.port_a_data_out_clock = "clock0";
defparam ram_block1a89.port_a_data_width = 1;
defparam ram_block1a89.port_a_first_address = 40960;
defparam ram_block1a89.port_a_first_bit_number = 9;
defparam ram_block1a89.port_a_last_address = 49151;
defparam ram_block1a89.port_a_logical_ram_depth = 65536;
defparam ram_block1a89.port_a_logical_ram_width = 16;
defparam ram_block1a89.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a89.ram_block_type = "auto";
defparam ram_block1a89.mem_init3 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a89.mem_init2 = "FFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a89.mem_init1 = "FFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000000";
defparam ram_block1a89.mem_init0 = "0000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000";

arriav_ram_block ram_block1a105(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a105_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a105.clk0_core_clock_enable = "ena0";
defparam ram_block1a105.clk0_input_clock_enable = "ena0";
defparam ram_block1a105.clk0_output_clock_enable = "ena0";
defparam ram_block1a105.data_interleave_offset_in_bits = 1;
defparam ram_block1a105.data_interleave_width_in_bits = 1;
defparam ram_block1a105.init_file = "DDS_48_v1_nco_ii_0_cos.hex";
defparam ram_block1a105.init_file_layout = "port_a";
defparam ram_block1a105.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0121|altsyncram:altsyncram_component0|altsyncram_78g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a105.operation_mode = "rom";
defparam ram_block1a105.port_a_address_clear = "none";
defparam ram_block1a105.port_a_address_width = 13;
defparam ram_block1a105.port_a_data_out_clear = "none";
defparam ram_block1a105.port_a_data_out_clock = "clock0";
defparam ram_block1a105.port_a_data_width = 1;
defparam ram_block1a105.port_a_first_address = 49152;
defparam ram_block1a105.port_a_first_bit_number = 9;
defparam ram_block1a105.port_a_last_address = 57343;
defparam ram_block1a105.port_a_logical_ram_depth = 65536;
defparam ram_block1a105.port_a_logical_ram_width = 16;
defparam ram_block1a105.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a105.ram_block_type = "auto";
defparam ram_block1a105.mem_init3 = "FFFFFFFFFFFFFFC000000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a105.mem_init2 = "FFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000";
defparam ram_block1a105.mem_init1 = "0000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000";
defparam ram_block1a105.mem_init0 = "00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000000000000000000";

arriav_ram_block ram_block1a121(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a121_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a121.clk0_core_clock_enable = "ena0";
defparam ram_block1a121.clk0_input_clock_enable = "ena0";
defparam ram_block1a121.clk0_output_clock_enable = "ena0";
defparam ram_block1a121.data_interleave_offset_in_bits = 1;
defparam ram_block1a121.data_interleave_width_in_bits = 1;
defparam ram_block1a121.init_file = "DDS_48_v1_nco_ii_0_cos.hex";
defparam ram_block1a121.init_file_layout = "port_a";
defparam ram_block1a121.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0121|altsyncram:altsyncram_component0|altsyncram_78g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a121.operation_mode = "rom";
defparam ram_block1a121.port_a_address_clear = "none";
defparam ram_block1a121.port_a_address_width = 13;
defparam ram_block1a121.port_a_data_out_clear = "none";
defparam ram_block1a121.port_a_data_out_clock = "clock0";
defparam ram_block1a121.port_a_data_width = 1;
defparam ram_block1a121.port_a_first_address = 57344;
defparam ram_block1a121.port_a_first_bit_number = 9;
defparam ram_block1a121.port_a_last_address = 65535;
defparam ram_block1a121.port_a_logical_ram_depth = 65536;
defparam ram_block1a121.port_a_logical_ram_width = 16;
defparam ram_block1a121.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a121.ram_block_type = "auto";
defparam ram_block1a121.mem_init3 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000000000000000000000000";
defparam ram_block1a121.mem_init2 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a121.mem_init1 = "FFFFFFFFFFFFF80000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000000000000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a121.mem_init0 = "FFFFFFFFFFFFFFFC00000000000000000000000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

arriav_ram_block ram_block1a41(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a41_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a41.clk0_core_clock_enable = "ena0";
defparam ram_block1a41.clk0_input_clock_enable = "ena0";
defparam ram_block1a41.clk0_output_clock_enable = "ena0";
defparam ram_block1a41.data_interleave_offset_in_bits = 1;
defparam ram_block1a41.data_interleave_width_in_bits = 1;
defparam ram_block1a41.init_file = "DDS_48_v1_nco_ii_0_cos.hex";
defparam ram_block1a41.init_file_layout = "port_a";
defparam ram_block1a41.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0121|altsyncram:altsyncram_component0|altsyncram_78g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a41.operation_mode = "rom";
defparam ram_block1a41.port_a_address_clear = "none";
defparam ram_block1a41.port_a_address_width = 13;
defparam ram_block1a41.port_a_data_out_clear = "none";
defparam ram_block1a41.port_a_data_out_clock = "clock0";
defparam ram_block1a41.port_a_data_width = 1;
defparam ram_block1a41.port_a_first_address = 16384;
defparam ram_block1a41.port_a_first_bit_number = 9;
defparam ram_block1a41.port_a_last_address = 24575;
defparam ram_block1a41.port_a_logical_ram_depth = 65536;
defparam ram_block1a41.port_a_logical_ram_width = 16;
defparam ram_block1a41.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a41.ram_block_type = "auto";
defparam ram_block1a41.mem_init3 = "000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000";
defparam ram_block1a41.mem_init2 = "000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a41.mem_init1 = "FFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a41.mem_init0 = "FFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE";

arriav_ram_block ram_block1a57(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a57_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a57.clk0_core_clock_enable = "ena0";
defparam ram_block1a57.clk0_input_clock_enable = "ena0";
defparam ram_block1a57.clk0_output_clock_enable = "ena0";
defparam ram_block1a57.data_interleave_offset_in_bits = 1;
defparam ram_block1a57.data_interleave_width_in_bits = 1;
defparam ram_block1a57.init_file = "DDS_48_v1_nco_ii_0_cos.hex";
defparam ram_block1a57.init_file_layout = "port_a";
defparam ram_block1a57.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0121|altsyncram:altsyncram_component0|altsyncram_78g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a57.operation_mode = "rom";
defparam ram_block1a57.port_a_address_clear = "none";
defparam ram_block1a57.port_a_address_width = 13;
defparam ram_block1a57.port_a_data_out_clear = "none";
defparam ram_block1a57.port_a_data_out_clock = "clock0";
defparam ram_block1a57.port_a_data_width = 1;
defparam ram_block1a57.port_a_first_address = 24576;
defparam ram_block1a57.port_a_first_bit_number = 9;
defparam ram_block1a57.port_a_last_address = 32767;
defparam ram_block1a57.port_a_logical_ram_depth = 65536;
defparam ram_block1a57.port_a_logical_ram_width = 16;
defparam ram_block1a57.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a57.ram_block_type = "auto";
defparam ram_block1a57.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a57.mem_init2 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a57.mem_init1 = "00000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000000000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a57.mem_init0 = "0000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000000000000000000000";

arriav_ram_block ram_block1a9(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a9_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a9.clk0_core_clock_enable = "ena0";
defparam ram_block1a9.clk0_input_clock_enable = "ena0";
defparam ram_block1a9.clk0_output_clock_enable = "ena0";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.init_file = "DDS_48_v1_nco_ii_0_cos.hex";
defparam ram_block1a9.init_file_layout = "port_a";
defparam ram_block1a9.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0121|altsyncram:altsyncram_component0|altsyncram_78g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a9.operation_mode = "rom";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 13;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "clock0";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 8191;
defparam ram_block1a9.port_a_logical_ram_depth = 65536;
defparam ram_block1a9.port_a_logical_ram_width = 16;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a9.ram_block_type = "auto";
defparam ram_block1a9.mem_init3 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFF";
defparam ram_block1a9.mem_init2 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFF";
defparam ram_block1a9.mem_init1 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a9.mem_init0 = "000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

arriav_ram_block ram_block1a25(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a25_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a25.clk0_core_clock_enable = "ena0";
defparam ram_block1a25.clk0_input_clock_enable = "ena0";
defparam ram_block1a25.clk0_output_clock_enable = "ena0";
defparam ram_block1a25.data_interleave_offset_in_bits = 1;
defparam ram_block1a25.data_interleave_width_in_bits = 1;
defparam ram_block1a25.init_file = "DDS_48_v1_nco_ii_0_cos.hex";
defparam ram_block1a25.init_file_layout = "port_a";
defparam ram_block1a25.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0121|altsyncram:altsyncram_component0|altsyncram_78g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a25.operation_mode = "rom";
defparam ram_block1a25.port_a_address_clear = "none";
defparam ram_block1a25.port_a_address_width = 13;
defparam ram_block1a25.port_a_data_out_clear = "none";
defparam ram_block1a25.port_a_data_out_clock = "clock0";
defparam ram_block1a25.port_a_data_width = 1;
defparam ram_block1a25.port_a_first_address = 8192;
defparam ram_block1a25.port_a_first_bit_number = 9;
defparam ram_block1a25.port_a_last_address = 16383;
defparam ram_block1a25.port_a_logical_ram_depth = 65536;
defparam ram_block1a25.port_a_logical_ram_width = 16;
defparam ram_block1a25.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a25.ram_block_type = "auto";
defparam ram_block1a25.mem_init3 = "00000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000";
defparam ram_block1a25.mem_init2 = "0000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000";
defparam ram_block1a25.mem_init1 = "00000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a25.mem_init0 = "FFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFF";

arriav_ram_block ram_block1a74(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a74_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a74.clk0_core_clock_enable = "ena0";
defparam ram_block1a74.clk0_input_clock_enable = "ena0";
defparam ram_block1a74.clk0_output_clock_enable = "ena0";
defparam ram_block1a74.data_interleave_offset_in_bits = 1;
defparam ram_block1a74.data_interleave_width_in_bits = 1;
defparam ram_block1a74.init_file = "DDS_48_v1_nco_ii_0_cos.hex";
defparam ram_block1a74.init_file_layout = "port_a";
defparam ram_block1a74.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0121|altsyncram:altsyncram_component0|altsyncram_78g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a74.operation_mode = "rom";
defparam ram_block1a74.port_a_address_clear = "none";
defparam ram_block1a74.port_a_address_width = 13;
defparam ram_block1a74.port_a_data_out_clear = "none";
defparam ram_block1a74.port_a_data_out_clock = "clock0";
defparam ram_block1a74.port_a_data_width = 1;
defparam ram_block1a74.port_a_first_address = 32768;
defparam ram_block1a74.port_a_first_bit_number = 10;
defparam ram_block1a74.port_a_last_address = 40959;
defparam ram_block1a74.port_a_logical_ram_depth = 65536;
defparam ram_block1a74.port_a_logical_ram_width = 16;
defparam ram_block1a74.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a74.ram_block_type = "auto";
defparam ram_block1a74.mem_init3 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a74.mem_init2 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a74.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a74.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

arriav_ram_block ram_block1a90(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a90_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a90.clk0_core_clock_enable = "ena0";
defparam ram_block1a90.clk0_input_clock_enable = "ena0";
defparam ram_block1a90.clk0_output_clock_enable = "ena0";
defparam ram_block1a90.data_interleave_offset_in_bits = 1;
defparam ram_block1a90.data_interleave_width_in_bits = 1;
defparam ram_block1a90.init_file = "DDS_48_v1_nco_ii_0_cos.hex";
defparam ram_block1a90.init_file_layout = "port_a";
defparam ram_block1a90.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0121|altsyncram:altsyncram_component0|altsyncram_78g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a90.operation_mode = "rom";
defparam ram_block1a90.port_a_address_clear = "none";
defparam ram_block1a90.port_a_address_width = 13;
defparam ram_block1a90.port_a_data_out_clear = "none";
defparam ram_block1a90.port_a_data_out_clock = "clock0";
defparam ram_block1a90.port_a_data_width = 1;
defparam ram_block1a90.port_a_first_address = 40960;
defparam ram_block1a90.port_a_first_bit_number = 10;
defparam ram_block1a90.port_a_last_address = 49151;
defparam ram_block1a90.port_a_logical_ram_depth = 65536;
defparam ram_block1a90.port_a_logical_ram_width = 16;
defparam ram_block1a90.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a90.ram_block_type = "auto";
defparam ram_block1a90.mem_init3 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000000000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a90.mem_init2 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000000000000000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000000000000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a90.mem_init1 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a90.mem_init0 = "0000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

arriav_ram_block ram_block1a106(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a106_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a106.clk0_core_clock_enable = "ena0";
defparam ram_block1a106.clk0_input_clock_enable = "ena0";
defparam ram_block1a106.clk0_output_clock_enable = "ena0";
defparam ram_block1a106.data_interleave_offset_in_bits = 1;
defparam ram_block1a106.data_interleave_width_in_bits = 1;
defparam ram_block1a106.init_file = "DDS_48_v1_nco_ii_0_cos.hex";
defparam ram_block1a106.init_file_layout = "port_a";
defparam ram_block1a106.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0121|altsyncram:altsyncram_component0|altsyncram_78g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a106.operation_mode = "rom";
defparam ram_block1a106.port_a_address_clear = "none";
defparam ram_block1a106.port_a_address_width = 13;
defparam ram_block1a106.port_a_data_out_clear = "none";
defparam ram_block1a106.port_a_data_out_clock = "clock0";
defparam ram_block1a106.port_a_data_width = 1;
defparam ram_block1a106.port_a_first_address = 49152;
defparam ram_block1a106.port_a_first_bit_number = 10;
defparam ram_block1a106.port_a_last_address = 57343;
defparam ram_block1a106.port_a_logical_ram_depth = 65536;
defparam ram_block1a106.port_a_logical_ram_width = 16;
defparam ram_block1a106.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a106.ram_block_type = "auto";
defparam ram_block1a106.mem_init3 = "000000000000000000000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a106.mem_init2 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a106.mem_init1 = "0000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000000000000000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a106.mem_init0 = "00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000000000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000000000000000000000000000000000000000000000000000000000";

arriav_ram_block ram_block1a122(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a122_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a122.clk0_core_clock_enable = "ena0";
defparam ram_block1a122.clk0_input_clock_enable = "ena0";
defparam ram_block1a122.clk0_output_clock_enable = "ena0";
defparam ram_block1a122.data_interleave_offset_in_bits = 1;
defparam ram_block1a122.data_interleave_width_in_bits = 1;
defparam ram_block1a122.init_file = "DDS_48_v1_nco_ii_0_cos.hex";
defparam ram_block1a122.init_file_layout = "port_a";
defparam ram_block1a122.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0121|altsyncram:altsyncram_component0|altsyncram_78g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a122.operation_mode = "rom";
defparam ram_block1a122.port_a_address_clear = "none";
defparam ram_block1a122.port_a_address_width = 13;
defparam ram_block1a122.port_a_data_out_clear = "none";
defparam ram_block1a122.port_a_data_out_clock = "clock0";
defparam ram_block1a122.port_a_data_width = 1;
defparam ram_block1a122.port_a_first_address = 57344;
defparam ram_block1a122.port_a_first_bit_number = 10;
defparam ram_block1a122.port_a_last_address = 65535;
defparam ram_block1a122.port_a_logical_ram_depth = 65536;
defparam ram_block1a122.port_a_logical_ram_width = 16;
defparam ram_block1a122.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a122.ram_block_type = "auto";
defparam ram_block1a122.mem_init3 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a122.mem_init2 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a122.mem_init1 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a122.mem_init0 = "000000000000000000000000000000000000000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000000000000000000000";

arriav_ram_block ram_block1a42(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a42_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a42.clk0_core_clock_enable = "ena0";
defparam ram_block1a42.clk0_input_clock_enable = "ena0";
defparam ram_block1a42.clk0_output_clock_enable = "ena0";
defparam ram_block1a42.data_interleave_offset_in_bits = 1;
defparam ram_block1a42.data_interleave_width_in_bits = 1;
defparam ram_block1a42.init_file = "DDS_48_v1_nco_ii_0_cos.hex";
defparam ram_block1a42.init_file_layout = "port_a";
defparam ram_block1a42.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0121|altsyncram:altsyncram_component0|altsyncram_78g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a42.operation_mode = "rom";
defparam ram_block1a42.port_a_address_clear = "none";
defparam ram_block1a42.port_a_address_width = 13;
defparam ram_block1a42.port_a_data_out_clear = "none";
defparam ram_block1a42.port_a_data_out_clock = "clock0";
defparam ram_block1a42.port_a_data_width = 1;
defparam ram_block1a42.port_a_first_address = 16384;
defparam ram_block1a42.port_a_first_bit_number = 10;
defparam ram_block1a42.port_a_last_address = 24575;
defparam ram_block1a42.port_a_logical_ram_depth = 65536;
defparam ram_block1a42.port_a_logical_ram_width = 16;
defparam ram_block1a42.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a42.ram_block_type = "auto";
defparam ram_block1a42.mem_init3 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000";
defparam ram_block1a42.mem_init2 = "0000000000000000000000000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a42.mem_init1 = "FFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000000000000000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a42.mem_init0 = "FFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE";

arriav_ram_block ram_block1a58(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a58_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a58.clk0_core_clock_enable = "ena0";
defparam ram_block1a58.clk0_input_clock_enable = "ena0";
defparam ram_block1a58.clk0_output_clock_enable = "ena0";
defparam ram_block1a58.data_interleave_offset_in_bits = 1;
defparam ram_block1a58.data_interleave_width_in_bits = 1;
defparam ram_block1a58.init_file = "DDS_48_v1_nco_ii_0_cos.hex";
defparam ram_block1a58.init_file_layout = "port_a";
defparam ram_block1a58.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0121|altsyncram:altsyncram_component0|altsyncram_78g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a58.operation_mode = "rom";
defparam ram_block1a58.port_a_address_clear = "none";
defparam ram_block1a58.port_a_address_width = 13;
defparam ram_block1a58.port_a_data_out_clear = "none";
defparam ram_block1a58.port_a_data_out_clock = "clock0";
defparam ram_block1a58.port_a_data_width = 1;
defparam ram_block1a58.port_a_first_address = 24576;
defparam ram_block1a58.port_a_first_bit_number = 10;
defparam ram_block1a58.port_a_last_address = 32767;
defparam ram_block1a58.port_a_logical_ram_depth = 65536;
defparam ram_block1a58.port_a_logical_ram_width = 16;
defparam ram_block1a58.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a58.ram_block_type = "auto";
defparam ram_block1a58.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a58.mem_init2 = "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a58.mem_init1 = "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a58.mem_init0 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

arriav_ram_block ram_block1a10(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a10_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a10.clk0_core_clock_enable = "ena0";
defparam ram_block1a10.clk0_input_clock_enable = "ena0";
defparam ram_block1a10.clk0_output_clock_enable = "ena0";
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.init_file = "DDS_48_v1_nco_ii_0_cos.hex";
defparam ram_block1a10.init_file_layout = "port_a";
defparam ram_block1a10.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0121|altsyncram:altsyncram_component0|altsyncram_78g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a10.operation_mode = "rom";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 13;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "clock0";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 8191;
defparam ram_block1a10.port_a_logical_ram_depth = 65536;
defparam ram_block1a10.port_a_logical_ram_width = 16;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a10.ram_block_type = "auto";
defparam ram_block1a10.mem_init3 = "00000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a10.mem_init2 = "00000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a10.mem_init1 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a10.mem_init0 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

arriav_ram_block ram_block1a26(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a26_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a26.clk0_core_clock_enable = "ena0";
defparam ram_block1a26.clk0_input_clock_enable = "ena0";
defparam ram_block1a26.clk0_output_clock_enable = "ena0";
defparam ram_block1a26.data_interleave_offset_in_bits = 1;
defparam ram_block1a26.data_interleave_width_in_bits = 1;
defparam ram_block1a26.init_file = "DDS_48_v1_nco_ii_0_cos.hex";
defparam ram_block1a26.init_file_layout = "port_a";
defparam ram_block1a26.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0121|altsyncram:altsyncram_component0|altsyncram_78g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a26.operation_mode = "rom";
defparam ram_block1a26.port_a_address_clear = "none";
defparam ram_block1a26.port_a_address_width = 13;
defparam ram_block1a26.port_a_data_out_clear = "none";
defparam ram_block1a26.port_a_data_out_clock = "clock0";
defparam ram_block1a26.port_a_data_width = 1;
defparam ram_block1a26.port_a_first_address = 8192;
defparam ram_block1a26.port_a_first_bit_number = 10;
defparam ram_block1a26.port_a_last_address = 16383;
defparam ram_block1a26.port_a_logical_ram_depth = 65536;
defparam ram_block1a26.port_a_logical_ram_width = 16;
defparam ram_block1a26.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a26.ram_block_type = "auto";
defparam ram_block1a26.mem_init3 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000000000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000";
defparam ram_block1a26.mem_init2 = "000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000000000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000";
defparam ram_block1a26.mem_init1 = "0000000000000000000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a26.mem_init0 = "FFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000000000000000000000000000000000000000000000";

arriav_ram_block ram_block1a75(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a75_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a75.clk0_core_clock_enable = "ena0";
defparam ram_block1a75.clk0_input_clock_enable = "ena0";
defparam ram_block1a75.clk0_output_clock_enable = "ena0";
defparam ram_block1a75.data_interleave_offset_in_bits = 1;
defparam ram_block1a75.data_interleave_width_in_bits = 1;
defparam ram_block1a75.init_file = "DDS_48_v1_nco_ii_0_cos.hex";
defparam ram_block1a75.init_file_layout = "port_a";
defparam ram_block1a75.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0121|altsyncram:altsyncram_component0|altsyncram_78g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a75.operation_mode = "rom";
defparam ram_block1a75.port_a_address_clear = "none";
defparam ram_block1a75.port_a_address_width = 13;
defparam ram_block1a75.port_a_data_out_clear = "none";
defparam ram_block1a75.port_a_data_out_clock = "clock0";
defparam ram_block1a75.port_a_data_width = 1;
defparam ram_block1a75.port_a_first_address = 32768;
defparam ram_block1a75.port_a_first_bit_number = 11;
defparam ram_block1a75.port_a_last_address = 40959;
defparam ram_block1a75.port_a_logical_ram_depth = 65536;
defparam ram_block1a75.port_a_logical_ram_width = 16;
defparam ram_block1a75.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a75.ram_block_type = "auto";
defparam ram_block1a75.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a75.mem_init2 = "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a75.mem_init1 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a75.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

arriav_ram_block ram_block1a91(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a91_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a91.clk0_core_clock_enable = "ena0";
defparam ram_block1a91.clk0_input_clock_enable = "ena0";
defparam ram_block1a91.clk0_output_clock_enable = "ena0";
defparam ram_block1a91.data_interleave_offset_in_bits = 1;
defparam ram_block1a91.data_interleave_width_in_bits = 1;
defparam ram_block1a91.init_file = "DDS_48_v1_nco_ii_0_cos.hex";
defparam ram_block1a91.init_file_layout = "port_a";
defparam ram_block1a91.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0121|altsyncram:altsyncram_component0|altsyncram_78g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a91.operation_mode = "rom";
defparam ram_block1a91.port_a_address_clear = "none";
defparam ram_block1a91.port_a_address_width = 13;
defparam ram_block1a91.port_a_data_out_clear = "none";
defparam ram_block1a91.port_a_data_out_clock = "clock0";
defparam ram_block1a91.port_a_data_width = 1;
defparam ram_block1a91.port_a_first_address = 40960;
defparam ram_block1a91.port_a_first_bit_number = 11;
defparam ram_block1a91.port_a_last_address = 49151;
defparam ram_block1a91.port_a_logical_ram_depth = 65536;
defparam ram_block1a91.port_a_logical_ram_width = 16;
defparam ram_block1a91.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a91.ram_block_type = "auto";
defparam ram_block1a91.mem_init3 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000";
defparam ram_block1a91.mem_init2 = "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a91.mem_init1 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a91.mem_init0 = "FFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000000000000000000000000000000000000000";

arriav_ram_block ram_block1a107(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a107_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a107.clk0_core_clock_enable = "ena0";
defparam ram_block1a107.clk0_input_clock_enable = "ena0";
defparam ram_block1a107.clk0_output_clock_enable = "ena0";
defparam ram_block1a107.data_interleave_offset_in_bits = 1;
defparam ram_block1a107.data_interleave_width_in_bits = 1;
defparam ram_block1a107.init_file = "DDS_48_v1_nco_ii_0_cos.hex";
defparam ram_block1a107.init_file_layout = "port_a";
defparam ram_block1a107.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0121|altsyncram:altsyncram_component0|altsyncram_78g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a107.operation_mode = "rom";
defparam ram_block1a107.port_a_address_clear = "none";
defparam ram_block1a107.port_a_address_width = 13;
defparam ram_block1a107.port_a_data_out_clear = "none";
defparam ram_block1a107.port_a_data_out_clock = "clock0";
defparam ram_block1a107.port_a_data_width = 1;
defparam ram_block1a107.port_a_first_address = 49152;
defparam ram_block1a107.port_a_first_bit_number = 11;
defparam ram_block1a107.port_a_last_address = 57343;
defparam ram_block1a107.port_a_logical_ram_depth = 65536;
defparam ram_block1a107.port_a_logical_ram_width = 16;
defparam ram_block1a107.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a107.ram_block_type = "auto";
defparam ram_block1a107.mem_init3 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000";
defparam ram_block1a107.mem_init2 = "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a107.mem_init1 = "0000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a107.mem_init0 = "FFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

arriav_ram_block ram_block1a123(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a123_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a123.clk0_core_clock_enable = "ena0";
defparam ram_block1a123.clk0_input_clock_enable = "ena0";
defparam ram_block1a123.clk0_output_clock_enable = "ena0";
defparam ram_block1a123.data_interleave_offset_in_bits = 1;
defparam ram_block1a123.data_interleave_width_in_bits = 1;
defparam ram_block1a123.init_file = "DDS_48_v1_nco_ii_0_cos.hex";
defparam ram_block1a123.init_file_layout = "port_a";
defparam ram_block1a123.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0121|altsyncram:altsyncram_component0|altsyncram_78g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a123.operation_mode = "rom";
defparam ram_block1a123.port_a_address_clear = "none";
defparam ram_block1a123.port_a_address_width = 13;
defparam ram_block1a123.port_a_data_out_clear = "none";
defparam ram_block1a123.port_a_data_out_clock = "clock0";
defparam ram_block1a123.port_a_data_width = 1;
defparam ram_block1a123.port_a_first_address = 57344;
defparam ram_block1a123.port_a_first_bit_number = 11;
defparam ram_block1a123.port_a_last_address = 65535;
defparam ram_block1a123.port_a_logical_ram_depth = 65536;
defparam ram_block1a123.port_a_logical_ram_width = 16;
defparam ram_block1a123.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a123.ram_block_type = "auto";
defparam ram_block1a123.mem_init3 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a123.mem_init2 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a123.mem_init1 = "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a123.mem_init0 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

arriav_ram_block ram_block1a43(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a43_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a43.clk0_core_clock_enable = "ena0";
defparam ram_block1a43.clk0_input_clock_enable = "ena0";
defparam ram_block1a43.clk0_output_clock_enable = "ena0";
defparam ram_block1a43.data_interleave_offset_in_bits = 1;
defparam ram_block1a43.data_interleave_width_in_bits = 1;
defparam ram_block1a43.init_file = "DDS_48_v1_nco_ii_0_cos.hex";
defparam ram_block1a43.init_file_layout = "port_a";
defparam ram_block1a43.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0121|altsyncram:altsyncram_component0|altsyncram_78g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a43.operation_mode = "rom";
defparam ram_block1a43.port_a_address_clear = "none";
defparam ram_block1a43.port_a_address_width = 13;
defparam ram_block1a43.port_a_data_out_clear = "none";
defparam ram_block1a43.port_a_data_out_clock = "clock0";
defparam ram_block1a43.port_a_data_width = 1;
defparam ram_block1a43.port_a_first_address = 16384;
defparam ram_block1a43.port_a_first_bit_number = 11;
defparam ram_block1a43.port_a_last_address = 24575;
defparam ram_block1a43.port_a_logical_ram_depth = 65536;
defparam ram_block1a43.port_a_logical_ram_width = 16;
defparam ram_block1a43.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a43.ram_block_type = "auto";
defparam ram_block1a43.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a43.mem_init2 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a43.mem_init1 = "FFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a43.mem_init0 = "00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE";

arriav_ram_block ram_block1a59(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a59_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a59.clk0_core_clock_enable = "ena0";
defparam ram_block1a59.clk0_input_clock_enable = "ena0";
defparam ram_block1a59.clk0_output_clock_enable = "ena0";
defparam ram_block1a59.data_interleave_offset_in_bits = 1;
defparam ram_block1a59.data_interleave_width_in_bits = 1;
defparam ram_block1a59.init_file = "DDS_48_v1_nco_ii_0_cos.hex";
defparam ram_block1a59.init_file_layout = "port_a";
defparam ram_block1a59.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0121|altsyncram:altsyncram_component0|altsyncram_78g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a59.operation_mode = "rom";
defparam ram_block1a59.port_a_address_clear = "none";
defparam ram_block1a59.port_a_address_width = 13;
defparam ram_block1a59.port_a_data_out_clear = "none";
defparam ram_block1a59.port_a_data_out_clock = "clock0";
defparam ram_block1a59.port_a_data_width = 1;
defparam ram_block1a59.port_a_first_address = 24576;
defparam ram_block1a59.port_a_first_bit_number = 11;
defparam ram_block1a59.port_a_last_address = 32767;
defparam ram_block1a59.port_a_logical_ram_depth = 65536;
defparam ram_block1a59.port_a_logical_ram_width = 16;
defparam ram_block1a59.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a59.ram_block_type = "auto";
defparam ram_block1a59.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a59.mem_init2 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a59.mem_init1 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a59.mem_init0 = "000000000000000000000000000000000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

arriav_ram_block ram_block1a11(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a11_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a11.clk0_core_clock_enable = "ena0";
defparam ram_block1a11.clk0_input_clock_enable = "ena0";
defparam ram_block1a11.clk0_output_clock_enable = "ena0";
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.init_file = "DDS_48_v1_nco_ii_0_cos.hex";
defparam ram_block1a11.init_file_layout = "port_a";
defparam ram_block1a11.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0121|altsyncram:altsyncram_component0|altsyncram_78g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a11.operation_mode = "rom";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 13;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "clock0";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 8191;
defparam ram_block1a11.port_a_logical_ram_depth = 65536;
defparam ram_block1a11.port_a_logical_ram_width = 16;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a11.ram_block_type = "auto";
defparam ram_block1a11.mem_init3 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a11.mem_init2 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a11.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a11.mem_init0 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

arriav_ram_block ram_block1a27(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a27_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a27.clk0_core_clock_enable = "ena0";
defparam ram_block1a27.clk0_input_clock_enable = "ena0";
defparam ram_block1a27.clk0_output_clock_enable = "ena0";
defparam ram_block1a27.data_interleave_offset_in_bits = 1;
defparam ram_block1a27.data_interleave_width_in_bits = 1;
defparam ram_block1a27.init_file = "DDS_48_v1_nco_ii_0_cos.hex";
defparam ram_block1a27.init_file_layout = "port_a";
defparam ram_block1a27.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0121|altsyncram:altsyncram_component0|altsyncram_78g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a27.operation_mode = "rom";
defparam ram_block1a27.port_a_address_clear = "none";
defparam ram_block1a27.port_a_address_width = 13;
defparam ram_block1a27.port_a_data_out_clear = "none";
defparam ram_block1a27.port_a_data_out_clock = "clock0";
defparam ram_block1a27.port_a_data_width = 1;
defparam ram_block1a27.port_a_first_address = 8192;
defparam ram_block1a27.port_a_first_bit_number = 11;
defparam ram_block1a27.port_a_last_address = 16383;
defparam ram_block1a27.port_a_logical_ram_depth = 65536;
defparam ram_block1a27.port_a_logical_ram_width = 16;
defparam ram_block1a27.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a27.ram_block_type = "auto";
defparam ram_block1a27.mem_init3 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a27.mem_init2 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000";
defparam ram_block1a27.mem_init1 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a27.mem_init0 = "0000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

arriav_ram_block ram_block1a76(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a76_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a76.clk0_core_clock_enable = "ena0";
defparam ram_block1a76.clk0_input_clock_enable = "ena0";
defparam ram_block1a76.clk0_output_clock_enable = "ena0";
defparam ram_block1a76.data_interleave_offset_in_bits = 1;
defparam ram_block1a76.data_interleave_width_in_bits = 1;
defparam ram_block1a76.init_file = "DDS_48_v1_nco_ii_0_cos.hex";
defparam ram_block1a76.init_file_layout = "port_a";
defparam ram_block1a76.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0121|altsyncram:altsyncram_component0|altsyncram_78g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a76.operation_mode = "rom";
defparam ram_block1a76.port_a_address_clear = "none";
defparam ram_block1a76.port_a_address_width = 13;
defparam ram_block1a76.port_a_data_out_clear = "none";
defparam ram_block1a76.port_a_data_out_clock = "clock0";
defparam ram_block1a76.port_a_data_width = 1;
defparam ram_block1a76.port_a_first_address = 32768;
defparam ram_block1a76.port_a_first_bit_number = 12;
defparam ram_block1a76.port_a_last_address = 40959;
defparam ram_block1a76.port_a_logical_ram_depth = 65536;
defparam ram_block1a76.port_a_logical_ram_width = 16;
defparam ram_block1a76.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a76.ram_block_type = "auto";
defparam ram_block1a76.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a76.mem_init2 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a76.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a76.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

arriav_ram_block ram_block1a92(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a92_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a92.clk0_core_clock_enable = "ena0";
defparam ram_block1a92.clk0_input_clock_enable = "ena0";
defparam ram_block1a92.clk0_output_clock_enable = "ena0";
defparam ram_block1a92.data_interleave_offset_in_bits = 1;
defparam ram_block1a92.data_interleave_width_in_bits = 1;
defparam ram_block1a92.init_file = "DDS_48_v1_nco_ii_0_cos.hex";
defparam ram_block1a92.init_file_layout = "port_a";
defparam ram_block1a92.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0121|altsyncram:altsyncram_component0|altsyncram_78g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a92.operation_mode = "rom";
defparam ram_block1a92.port_a_address_clear = "none";
defparam ram_block1a92.port_a_address_width = 13;
defparam ram_block1a92.port_a_data_out_clear = "none";
defparam ram_block1a92.port_a_data_out_clock = "clock0";
defparam ram_block1a92.port_a_data_width = 1;
defparam ram_block1a92.port_a_first_address = 40960;
defparam ram_block1a92.port_a_first_bit_number = 12;
defparam ram_block1a92.port_a_last_address = 49151;
defparam ram_block1a92.port_a_logical_ram_depth = 65536;
defparam ram_block1a92.port_a_logical_ram_width = 16;
defparam ram_block1a92.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a92.ram_block_type = "auto";
defparam ram_block1a92.mem_init3 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a92.mem_init2 = "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000";
defparam ram_block1a92.mem_init1 = "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a92.mem_init0 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

arriav_ram_block ram_block1a108(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a108_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a108.clk0_core_clock_enable = "ena0";
defparam ram_block1a108.clk0_input_clock_enable = "ena0";
defparam ram_block1a108.clk0_output_clock_enable = "ena0";
defparam ram_block1a108.data_interleave_offset_in_bits = 1;
defparam ram_block1a108.data_interleave_width_in_bits = 1;
defparam ram_block1a108.init_file = "DDS_48_v1_nco_ii_0_cos.hex";
defparam ram_block1a108.init_file_layout = "port_a";
defparam ram_block1a108.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0121|altsyncram:altsyncram_component0|altsyncram_78g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a108.operation_mode = "rom";
defparam ram_block1a108.port_a_address_clear = "none";
defparam ram_block1a108.port_a_address_width = 13;
defparam ram_block1a108.port_a_data_out_clear = "none";
defparam ram_block1a108.port_a_data_out_clock = "clock0";
defparam ram_block1a108.port_a_data_width = 1;
defparam ram_block1a108.port_a_first_address = 49152;
defparam ram_block1a108.port_a_first_bit_number = 12;
defparam ram_block1a108.port_a_last_address = 57343;
defparam ram_block1a108.port_a_logical_ram_depth = 65536;
defparam ram_block1a108.port_a_logical_ram_width = 16;
defparam ram_block1a108.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a108.ram_block_type = "auto";
defparam ram_block1a108.mem_init3 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a108.mem_init2 = "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a108.mem_init1 = "FFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a108.mem_init0 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

arriav_ram_block ram_block1a124(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a124_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a124.clk0_core_clock_enable = "ena0";
defparam ram_block1a124.clk0_input_clock_enable = "ena0";
defparam ram_block1a124.clk0_output_clock_enable = "ena0";
defparam ram_block1a124.data_interleave_offset_in_bits = 1;
defparam ram_block1a124.data_interleave_width_in_bits = 1;
defparam ram_block1a124.init_file = "DDS_48_v1_nco_ii_0_cos.hex";
defparam ram_block1a124.init_file_layout = "port_a";
defparam ram_block1a124.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0121|altsyncram:altsyncram_component0|altsyncram_78g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a124.operation_mode = "rom";
defparam ram_block1a124.port_a_address_clear = "none";
defparam ram_block1a124.port_a_address_width = 13;
defparam ram_block1a124.port_a_data_out_clear = "none";
defparam ram_block1a124.port_a_data_out_clock = "clock0";
defparam ram_block1a124.port_a_data_width = 1;
defparam ram_block1a124.port_a_first_address = 57344;
defparam ram_block1a124.port_a_first_bit_number = 12;
defparam ram_block1a124.port_a_last_address = 65535;
defparam ram_block1a124.port_a_logical_ram_depth = 65536;
defparam ram_block1a124.port_a_logical_ram_width = 16;
defparam ram_block1a124.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a124.ram_block_type = "auto";
defparam ram_block1a124.mem_init3 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a124.mem_init2 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a124.mem_init1 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a124.mem_init0 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

arriav_ram_block ram_block1a44(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a44_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a44.clk0_core_clock_enable = "ena0";
defparam ram_block1a44.clk0_input_clock_enable = "ena0";
defparam ram_block1a44.clk0_output_clock_enable = "ena0";
defparam ram_block1a44.data_interleave_offset_in_bits = 1;
defparam ram_block1a44.data_interleave_width_in_bits = 1;
defparam ram_block1a44.init_file = "DDS_48_v1_nco_ii_0_cos.hex";
defparam ram_block1a44.init_file_layout = "port_a";
defparam ram_block1a44.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0121|altsyncram:altsyncram_component0|altsyncram_78g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a44.operation_mode = "rom";
defparam ram_block1a44.port_a_address_clear = "none";
defparam ram_block1a44.port_a_address_width = 13;
defparam ram_block1a44.port_a_data_out_clear = "none";
defparam ram_block1a44.port_a_data_out_clock = "clock0";
defparam ram_block1a44.port_a_data_width = 1;
defparam ram_block1a44.port_a_first_address = 16384;
defparam ram_block1a44.port_a_first_bit_number = 12;
defparam ram_block1a44.port_a_last_address = 24575;
defparam ram_block1a44.port_a_logical_ram_depth = 65536;
defparam ram_block1a44.port_a_logical_ram_width = 16;
defparam ram_block1a44.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a44.ram_block_type = "auto";
defparam ram_block1a44.mem_init3 = "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a44.mem_init2 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a44.mem_init1 = "0000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a44.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE";

arriav_ram_block ram_block1a60(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a60_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a60.clk0_core_clock_enable = "ena0";
defparam ram_block1a60.clk0_input_clock_enable = "ena0";
defparam ram_block1a60.clk0_output_clock_enable = "ena0";
defparam ram_block1a60.data_interleave_offset_in_bits = 1;
defparam ram_block1a60.data_interleave_width_in_bits = 1;
defparam ram_block1a60.init_file = "DDS_48_v1_nco_ii_0_cos.hex";
defparam ram_block1a60.init_file_layout = "port_a";
defparam ram_block1a60.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0121|altsyncram:altsyncram_component0|altsyncram_78g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a60.operation_mode = "rom";
defparam ram_block1a60.port_a_address_clear = "none";
defparam ram_block1a60.port_a_address_width = 13;
defparam ram_block1a60.port_a_data_out_clear = "none";
defparam ram_block1a60.port_a_data_out_clock = "clock0";
defparam ram_block1a60.port_a_data_width = 1;
defparam ram_block1a60.port_a_first_address = 24576;
defparam ram_block1a60.port_a_first_bit_number = 12;
defparam ram_block1a60.port_a_last_address = 32767;
defparam ram_block1a60.port_a_logical_ram_depth = 65536;
defparam ram_block1a60.port_a_logical_ram_width = 16;
defparam ram_block1a60.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a60.ram_block_type = "auto";
defparam ram_block1a60.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a60.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a60.mem_init1 = "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a60.mem_init0 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

arriav_ram_block ram_block1a12(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a12_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a12.clk0_core_clock_enable = "ena0";
defparam ram_block1a12.clk0_input_clock_enable = "ena0";
defparam ram_block1a12.clk0_output_clock_enable = "ena0";
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.init_file = "DDS_48_v1_nco_ii_0_cos.hex";
defparam ram_block1a12.init_file_layout = "port_a";
defparam ram_block1a12.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0121|altsyncram:altsyncram_component0|altsyncram_78g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a12.operation_mode = "rom";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 13;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "clock0";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 8191;
defparam ram_block1a12.port_a_logical_ram_depth = 65536;
defparam ram_block1a12.port_a_logical_ram_width = 16;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a12.ram_block_type = "auto";
defparam ram_block1a12.mem_init3 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a12.mem_init2 = "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a12.mem_init1 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a12.mem_init0 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

arriav_ram_block ram_block1a28(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a28_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a28.clk0_core_clock_enable = "ena0";
defparam ram_block1a28.clk0_input_clock_enable = "ena0";
defparam ram_block1a28.clk0_output_clock_enable = "ena0";
defparam ram_block1a28.data_interleave_offset_in_bits = 1;
defparam ram_block1a28.data_interleave_width_in_bits = 1;
defparam ram_block1a28.init_file = "DDS_48_v1_nco_ii_0_cos.hex";
defparam ram_block1a28.init_file_layout = "port_a";
defparam ram_block1a28.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0121|altsyncram:altsyncram_component0|altsyncram_78g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a28.operation_mode = "rom";
defparam ram_block1a28.port_a_address_clear = "none";
defparam ram_block1a28.port_a_address_width = 13;
defparam ram_block1a28.port_a_data_out_clear = "none";
defparam ram_block1a28.port_a_data_out_clock = "clock0";
defparam ram_block1a28.port_a_data_width = 1;
defparam ram_block1a28.port_a_first_address = 8192;
defparam ram_block1a28.port_a_first_bit_number = 12;
defparam ram_block1a28.port_a_last_address = 16383;
defparam ram_block1a28.port_a_logical_ram_depth = 65536;
defparam ram_block1a28.port_a_logical_ram_width = 16;
defparam ram_block1a28.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a28.ram_block_type = "auto";
defparam ram_block1a28.mem_init3 = "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a28.mem_init2 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a28.mem_init1 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a28.mem_init0 = "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

arriav_ram_block ram_block1a77(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a77_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a77.clk0_core_clock_enable = "ena0";
defparam ram_block1a77.clk0_input_clock_enable = "ena0";
defparam ram_block1a77.clk0_output_clock_enable = "ena0";
defparam ram_block1a77.data_interleave_offset_in_bits = 1;
defparam ram_block1a77.data_interleave_width_in_bits = 1;
defparam ram_block1a77.init_file = "DDS_48_v1_nco_ii_0_cos.hex";
defparam ram_block1a77.init_file_layout = "port_a";
defparam ram_block1a77.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0121|altsyncram:altsyncram_component0|altsyncram_78g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a77.operation_mode = "rom";
defparam ram_block1a77.port_a_address_clear = "none";
defparam ram_block1a77.port_a_address_width = 13;
defparam ram_block1a77.port_a_data_out_clear = "none";
defparam ram_block1a77.port_a_data_out_clock = "clock0";
defparam ram_block1a77.port_a_data_width = 1;
defparam ram_block1a77.port_a_first_address = 32768;
defparam ram_block1a77.port_a_first_bit_number = 13;
defparam ram_block1a77.port_a_last_address = 40959;
defparam ram_block1a77.port_a_logical_ram_depth = 65536;
defparam ram_block1a77.port_a_logical_ram_width = 16;
defparam ram_block1a77.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a77.ram_block_type = "auto";
defparam ram_block1a77.mem_init3 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a77.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a77.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a77.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

arriav_ram_block ram_block1a93(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a93_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a93.clk0_core_clock_enable = "ena0";
defparam ram_block1a93.clk0_input_clock_enable = "ena0";
defparam ram_block1a93.clk0_output_clock_enable = "ena0";
defparam ram_block1a93.data_interleave_offset_in_bits = 1;
defparam ram_block1a93.data_interleave_width_in_bits = 1;
defparam ram_block1a93.init_file = "DDS_48_v1_nco_ii_0_cos.hex";
defparam ram_block1a93.init_file_layout = "port_a";
defparam ram_block1a93.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0121|altsyncram:altsyncram_component0|altsyncram_78g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a93.operation_mode = "rom";
defparam ram_block1a93.port_a_address_clear = "none";
defparam ram_block1a93.port_a_address_width = 13;
defparam ram_block1a93.port_a_data_out_clear = "none";
defparam ram_block1a93.port_a_data_out_clock = "clock0";
defparam ram_block1a93.port_a_data_width = 1;
defparam ram_block1a93.port_a_first_address = 40960;
defparam ram_block1a93.port_a_first_bit_number = 13;
defparam ram_block1a93.port_a_last_address = 49151;
defparam ram_block1a93.port_a_logical_ram_depth = 65536;
defparam ram_block1a93.port_a_logical_ram_width = 16;
defparam ram_block1a93.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a93.ram_block_type = "auto";
defparam ram_block1a93.mem_init3 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a93.mem_init2 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a93.mem_init1 = "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a93.mem_init0 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

arriav_ram_block ram_block1a109(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a109_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a109.clk0_core_clock_enable = "ena0";
defparam ram_block1a109.clk0_input_clock_enable = "ena0";
defparam ram_block1a109.clk0_output_clock_enable = "ena0";
defparam ram_block1a109.data_interleave_offset_in_bits = 1;
defparam ram_block1a109.data_interleave_width_in_bits = 1;
defparam ram_block1a109.init_file = "DDS_48_v1_nco_ii_0_cos.hex";
defparam ram_block1a109.init_file_layout = "port_a";
defparam ram_block1a109.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0121|altsyncram:altsyncram_component0|altsyncram_78g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a109.operation_mode = "rom";
defparam ram_block1a109.port_a_address_clear = "none";
defparam ram_block1a109.port_a_address_width = 13;
defparam ram_block1a109.port_a_data_out_clear = "none";
defparam ram_block1a109.port_a_data_out_clock = "clock0";
defparam ram_block1a109.port_a_data_width = 1;
defparam ram_block1a109.port_a_first_address = 49152;
defparam ram_block1a109.port_a_first_bit_number = 13;
defparam ram_block1a109.port_a_last_address = 57343;
defparam ram_block1a109.port_a_logical_ram_depth = 65536;
defparam ram_block1a109.port_a_logical_ram_width = 16;
defparam ram_block1a109.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a109.ram_block_type = "auto";
defparam ram_block1a109.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a109.mem_init2 = "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a109.mem_init1 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a109.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

arriav_ram_block ram_block1a125(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a125_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a125.clk0_core_clock_enable = "ena0";
defparam ram_block1a125.clk0_input_clock_enable = "ena0";
defparam ram_block1a125.clk0_output_clock_enable = "ena0";
defparam ram_block1a125.data_interleave_offset_in_bits = 1;
defparam ram_block1a125.data_interleave_width_in_bits = 1;
defparam ram_block1a125.init_file = "DDS_48_v1_nco_ii_0_cos.hex";
defparam ram_block1a125.init_file_layout = "port_a";
defparam ram_block1a125.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0121|altsyncram:altsyncram_component0|altsyncram_78g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a125.operation_mode = "rom";
defparam ram_block1a125.port_a_address_clear = "none";
defparam ram_block1a125.port_a_address_width = 13;
defparam ram_block1a125.port_a_data_out_clear = "none";
defparam ram_block1a125.port_a_data_out_clock = "clock0";
defparam ram_block1a125.port_a_data_width = 1;
defparam ram_block1a125.port_a_first_address = 57344;
defparam ram_block1a125.port_a_first_bit_number = 13;
defparam ram_block1a125.port_a_last_address = 65535;
defparam ram_block1a125.port_a_logical_ram_depth = 65536;
defparam ram_block1a125.port_a_logical_ram_width = 16;
defparam ram_block1a125.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a125.ram_block_type = "auto";
defparam ram_block1a125.mem_init3 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a125.mem_init2 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a125.mem_init1 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a125.mem_init0 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

arriav_ram_block ram_block1a45(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a45_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a45.clk0_core_clock_enable = "ena0";
defparam ram_block1a45.clk0_input_clock_enable = "ena0";
defparam ram_block1a45.clk0_output_clock_enable = "ena0";
defparam ram_block1a45.data_interleave_offset_in_bits = 1;
defparam ram_block1a45.data_interleave_width_in_bits = 1;
defparam ram_block1a45.init_file = "DDS_48_v1_nco_ii_0_cos.hex";
defparam ram_block1a45.init_file_layout = "port_a";
defparam ram_block1a45.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0121|altsyncram:altsyncram_component0|altsyncram_78g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a45.operation_mode = "rom";
defparam ram_block1a45.port_a_address_clear = "none";
defparam ram_block1a45.port_a_address_width = 13;
defparam ram_block1a45.port_a_data_out_clear = "none";
defparam ram_block1a45.port_a_data_out_clock = "clock0";
defparam ram_block1a45.port_a_data_width = 1;
defparam ram_block1a45.port_a_first_address = 16384;
defparam ram_block1a45.port_a_first_bit_number = 13;
defparam ram_block1a45.port_a_last_address = 24575;
defparam ram_block1a45.port_a_logical_ram_depth = 65536;
defparam ram_block1a45.port_a_logical_ram_width = 16;
defparam ram_block1a45.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a45.ram_block_type = "auto";
defparam ram_block1a45.mem_init3 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a45.mem_init2 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a45.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a45.mem_init0 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE";

arriav_ram_block ram_block1a61(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a61_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a61.clk0_core_clock_enable = "ena0";
defparam ram_block1a61.clk0_input_clock_enable = "ena0";
defparam ram_block1a61.clk0_output_clock_enable = "ena0";
defparam ram_block1a61.data_interleave_offset_in_bits = 1;
defparam ram_block1a61.data_interleave_width_in_bits = 1;
defparam ram_block1a61.init_file = "DDS_48_v1_nco_ii_0_cos.hex";
defparam ram_block1a61.init_file_layout = "port_a";
defparam ram_block1a61.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0121|altsyncram:altsyncram_component0|altsyncram_78g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a61.operation_mode = "rom";
defparam ram_block1a61.port_a_address_clear = "none";
defparam ram_block1a61.port_a_address_width = 13;
defparam ram_block1a61.port_a_data_out_clear = "none";
defparam ram_block1a61.port_a_data_out_clock = "clock0";
defparam ram_block1a61.port_a_data_width = 1;
defparam ram_block1a61.port_a_first_address = 24576;
defparam ram_block1a61.port_a_first_bit_number = 13;
defparam ram_block1a61.port_a_last_address = 32767;
defparam ram_block1a61.port_a_logical_ram_depth = 65536;
defparam ram_block1a61.port_a_logical_ram_width = 16;
defparam ram_block1a61.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a61.ram_block_type = "auto";
defparam ram_block1a61.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a61.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a61.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a61.mem_init0 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

arriav_ram_block ram_block1a13(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a13_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a13.clk0_core_clock_enable = "ena0";
defparam ram_block1a13.clk0_input_clock_enable = "ena0";
defparam ram_block1a13.clk0_output_clock_enable = "ena0";
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.init_file = "DDS_48_v1_nco_ii_0_cos.hex";
defparam ram_block1a13.init_file_layout = "port_a";
defparam ram_block1a13.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0121|altsyncram:altsyncram_component0|altsyncram_78g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a13.operation_mode = "rom";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 13;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "clock0";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 8191;
defparam ram_block1a13.port_a_logical_ram_depth = 65536;
defparam ram_block1a13.port_a_logical_ram_width = 16;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a13.ram_block_type = "auto";
defparam ram_block1a13.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a13.mem_init2 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a13.mem_init1 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a13.mem_init0 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

arriav_ram_block ram_block1a29(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a29_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a29.clk0_core_clock_enable = "ena0";
defparam ram_block1a29.clk0_input_clock_enable = "ena0";
defparam ram_block1a29.clk0_output_clock_enable = "ena0";
defparam ram_block1a29.data_interleave_offset_in_bits = 1;
defparam ram_block1a29.data_interleave_width_in_bits = 1;
defparam ram_block1a29.init_file = "DDS_48_v1_nco_ii_0_cos.hex";
defparam ram_block1a29.init_file_layout = "port_a";
defparam ram_block1a29.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0121|altsyncram:altsyncram_component0|altsyncram_78g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a29.operation_mode = "rom";
defparam ram_block1a29.port_a_address_clear = "none";
defparam ram_block1a29.port_a_address_width = 13;
defparam ram_block1a29.port_a_data_out_clear = "none";
defparam ram_block1a29.port_a_data_out_clock = "clock0";
defparam ram_block1a29.port_a_data_width = 1;
defparam ram_block1a29.port_a_first_address = 8192;
defparam ram_block1a29.port_a_first_bit_number = 13;
defparam ram_block1a29.port_a_last_address = 16383;
defparam ram_block1a29.port_a_logical_ram_depth = 65536;
defparam ram_block1a29.port_a_logical_ram_width = 16;
defparam ram_block1a29.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a29.ram_block_type = "auto";
defparam ram_block1a29.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a29.mem_init2 = "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a29.mem_init1 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a29.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

arriav_ram_block ram_block1a78(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a78_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a78.clk0_core_clock_enable = "ena0";
defparam ram_block1a78.clk0_input_clock_enable = "ena0";
defparam ram_block1a78.clk0_output_clock_enable = "ena0";
defparam ram_block1a78.data_interleave_offset_in_bits = 1;
defparam ram_block1a78.data_interleave_width_in_bits = 1;
defparam ram_block1a78.init_file = "DDS_48_v1_nco_ii_0_cos.hex";
defparam ram_block1a78.init_file_layout = "port_a";
defparam ram_block1a78.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0121|altsyncram:altsyncram_component0|altsyncram_78g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a78.operation_mode = "rom";
defparam ram_block1a78.port_a_address_clear = "none";
defparam ram_block1a78.port_a_address_width = 13;
defparam ram_block1a78.port_a_data_out_clear = "none";
defparam ram_block1a78.port_a_data_out_clock = "clock0";
defparam ram_block1a78.port_a_data_width = 1;
defparam ram_block1a78.port_a_first_address = 32768;
defparam ram_block1a78.port_a_first_bit_number = 14;
defparam ram_block1a78.port_a_last_address = 40959;
defparam ram_block1a78.port_a_logical_ram_depth = 65536;
defparam ram_block1a78.port_a_logical_ram_width = 16;
defparam ram_block1a78.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a78.ram_block_type = "auto";
defparam ram_block1a78.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a78.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a78.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a78.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

arriav_ram_block ram_block1a94(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a94_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a94.clk0_core_clock_enable = "ena0";
defparam ram_block1a94.clk0_input_clock_enable = "ena0";
defparam ram_block1a94.clk0_output_clock_enable = "ena0";
defparam ram_block1a94.data_interleave_offset_in_bits = 1;
defparam ram_block1a94.data_interleave_width_in_bits = 1;
defparam ram_block1a94.init_file = "DDS_48_v1_nco_ii_0_cos.hex";
defparam ram_block1a94.init_file_layout = "port_a";
defparam ram_block1a94.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0121|altsyncram:altsyncram_component0|altsyncram_78g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a94.operation_mode = "rom";
defparam ram_block1a94.port_a_address_clear = "none";
defparam ram_block1a94.port_a_address_width = 13;
defparam ram_block1a94.port_a_data_out_clear = "none";
defparam ram_block1a94.port_a_data_out_clock = "clock0";
defparam ram_block1a94.port_a_data_width = 1;
defparam ram_block1a94.port_a_first_address = 40960;
defparam ram_block1a94.port_a_first_bit_number = 14;
defparam ram_block1a94.port_a_last_address = 49151;
defparam ram_block1a94.port_a_logical_ram_depth = 65536;
defparam ram_block1a94.port_a_logical_ram_width = 16;
defparam ram_block1a94.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a94.ram_block_type = "auto";
defparam ram_block1a94.mem_init3 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a94.mem_init2 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a94.mem_init1 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a94.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

arriav_ram_block ram_block1a110(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a110_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a110.clk0_core_clock_enable = "ena0";
defparam ram_block1a110.clk0_input_clock_enable = "ena0";
defparam ram_block1a110.clk0_output_clock_enable = "ena0";
defparam ram_block1a110.data_interleave_offset_in_bits = 1;
defparam ram_block1a110.data_interleave_width_in_bits = 1;
defparam ram_block1a110.init_file = "DDS_48_v1_nco_ii_0_cos.hex";
defparam ram_block1a110.init_file_layout = "port_a";
defparam ram_block1a110.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0121|altsyncram:altsyncram_component0|altsyncram_78g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a110.operation_mode = "rom";
defparam ram_block1a110.port_a_address_clear = "none";
defparam ram_block1a110.port_a_address_width = 13;
defparam ram_block1a110.port_a_data_out_clear = "none";
defparam ram_block1a110.port_a_data_out_clock = "clock0";
defparam ram_block1a110.port_a_data_width = 1;
defparam ram_block1a110.port_a_first_address = 49152;
defparam ram_block1a110.port_a_first_bit_number = 14;
defparam ram_block1a110.port_a_last_address = 57343;
defparam ram_block1a110.port_a_logical_ram_depth = 65536;
defparam ram_block1a110.port_a_logical_ram_width = 16;
defparam ram_block1a110.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a110.ram_block_type = "auto";
defparam ram_block1a110.mem_init3 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a110.mem_init2 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a110.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a110.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

arriav_ram_block ram_block1a126(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a126_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a126.clk0_core_clock_enable = "ena0";
defparam ram_block1a126.clk0_input_clock_enable = "ena0";
defparam ram_block1a126.clk0_output_clock_enable = "ena0";
defparam ram_block1a126.data_interleave_offset_in_bits = 1;
defparam ram_block1a126.data_interleave_width_in_bits = 1;
defparam ram_block1a126.init_file = "DDS_48_v1_nco_ii_0_cos.hex";
defparam ram_block1a126.init_file_layout = "port_a";
defparam ram_block1a126.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0121|altsyncram:altsyncram_component0|altsyncram_78g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a126.operation_mode = "rom";
defparam ram_block1a126.port_a_address_clear = "none";
defparam ram_block1a126.port_a_address_width = 13;
defparam ram_block1a126.port_a_data_out_clear = "none";
defparam ram_block1a126.port_a_data_out_clock = "clock0";
defparam ram_block1a126.port_a_data_width = 1;
defparam ram_block1a126.port_a_first_address = 57344;
defparam ram_block1a126.port_a_first_bit_number = 14;
defparam ram_block1a126.port_a_last_address = 65535;
defparam ram_block1a126.port_a_logical_ram_depth = 65536;
defparam ram_block1a126.port_a_logical_ram_width = 16;
defparam ram_block1a126.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a126.ram_block_type = "auto";
defparam ram_block1a126.mem_init3 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a126.mem_init2 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a126.mem_init1 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a126.mem_init0 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

arriav_ram_block ram_block1a46(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a46_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a46.clk0_core_clock_enable = "ena0";
defparam ram_block1a46.clk0_input_clock_enable = "ena0";
defparam ram_block1a46.clk0_output_clock_enable = "ena0";
defparam ram_block1a46.data_interleave_offset_in_bits = 1;
defparam ram_block1a46.data_interleave_width_in_bits = 1;
defparam ram_block1a46.init_file = "DDS_48_v1_nco_ii_0_cos.hex";
defparam ram_block1a46.init_file_layout = "port_a";
defparam ram_block1a46.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0121|altsyncram:altsyncram_component0|altsyncram_78g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a46.operation_mode = "rom";
defparam ram_block1a46.port_a_address_clear = "none";
defparam ram_block1a46.port_a_address_width = 13;
defparam ram_block1a46.port_a_data_out_clear = "none";
defparam ram_block1a46.port_a_data_out_clock = "clock0";
defparam ram_block1a46.port_a_data_width = 1;
defparam ram_block1a46.port_a_first_address = 16384;
defparam ram_block1a46.port_a_first_bit_number = 14;
defparam ram_block1a46.port_a_last_address = 24575;
defparam ram_block1a46.port_a_logical_ram_depth = 65536;
defparam ram_block1a46.port_a_logical_ram_width = 16;
defparam ram_block1a46.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a46.ram_block_type = "auto";
defparam ram_block1a46.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a46.mem_init2 = "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a46.mem_init1 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a46.mem_init0 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE";

arriav_ram_block ram_block1a62(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a62_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a62.clk0_core_clock_enable = "ena0";
defparam ram_block1a62.clk0_input_clock_enable = "ena0";
defparam ram_block1a62.clk0_output_clock_enable = "ena0";
defparam ram_block1a62.data_interleave_offset_in_bits = 1;
defparam ram_block1a62.data_interleave_width_in_bits = 1;
defparam ram_block1a62.init_file = "DDS_48_v1_nco_ii_0_cos.hex";
defparam ram_block1a62.init_file_layout = "port_a";
defparam ram_block1a62.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0121|altsyncram:altsyncram_component0|altsyncram_78g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a62.operation_mode = "rom";
defparam ram_block1a62.port_a_address_clear = "none";
defparam ram_block1a62.port_a_address_width = 13;
defparam ram_block1a62.port_a_data_out_clear = "none";
defparam ram_block1a62.port_a_data_out_clock = "clock0";
defparam ram_block1a62.port_a_data_width = 1;
defparam ram_block1a62.port_a_first_address = 24576;
defparam ram_block1a62.port_a_first_bit_number = 14;
defparam ram_block1a62.port_a_last_address = 32767;
defparam ram_block1a62.port_a_logical_ram_depth = 65536;
defparam ram_block1a62.port_a_logical_ram_width = 16;
defparam ram_block1a62.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a62.ram_block_type = "auto";
defparam ram_block1a62.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a62.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a62.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a62.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

arriav_ram_block ram_block1a14(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a14_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a14.clk0_core_clock_enable = "ena0";
defparam ram_block1a14.clk0_input_clock_enable = "ena0";
defparam ram_block1a14.clk0_output_clock_enable = "ena0";
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.init_file = "DDS_48_v1_nco_ii_0_cos.hex";
defparam ram_block1a14.init_file_layout = "port_a";
defparam ram_block1a14.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0121|altsyncram:altsyncram_component0|altsyncram_78g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a14.operation_mode = "rom";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 13;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "clock0";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 8191;
defparam ram_block1a14.port_a_logical_ram_depth = 65536;
defparam ram_block1a14.port_a_logical_ram_width = 16;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a14.ram_block_type = "auto";
defparam ram_block1a14.mem_init3 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a14.mem_init2 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a14.mem_init1 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a14.mem_init0 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

arriav_ram_block ram_block1a30(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a30_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a30.clk0_core_clock_enable = "ena0";
defparam ram_block1a30.clk0_input_clock_enable = "ena0";
defparam ram_block1a30.clk0_output_clock_enable = "ena0";
defparam ram_block1a30.data_interleave_offset_in_bits = 1;
defparam ram_block1a30.data_interleave_width_in_bits = 1;
defparam ram_block1a30.init_file = "DDS_48_v1_nco_ii_0_cos.hex";
defparam ram_block1a30.init_file_layout = "port_a";
defparam ram_block1a30.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0121|altsyncram:altsyncram_component0|altsyncram_78g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a30.operation_mode = "rom";
defparam ram_block1a30.port_a_address_clear = "none";
defparam ram_block1a30.port_a_address_width = 13;
defparam ram_block1a30.port_a_data_out_clear = "none";
defparam ram_block1a30.port_a_data_out_clock = "clock0";
defparam ram_block1a30.port_a_data_width = 1;
defparam ram_block1a30.port_a_first_address = 8192;
defparam ram_block1a30.port_a_first_bit_number = 14;
defparam ram_block1a30.port_a_last_address = 16383;
defparam ram_block1a30.port_a_logical_ram_depth = 65536;
defparam ram_block1a30.port_a_logical_ram_width = 16;
defparam ram_block1a30.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a30.ram_block_type = "auto";
defparam ram_block1a30.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a30.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a30.mem_init1 = "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a30.mem_init0 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

arriav_ram_block ram_block1a79(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a79_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a79.clk0_core_clock_enable = "ena0";
defparam ram_block1a79.clk0_input_clock_enable = "ena0";
defparam ram_block1a79.clk0_output_clock_enable = "ena0";
defparam ram_block1a79.data_interleave_offset_in_bits = 1;
defparam ram_block1a79.data_interleave_width_in_bits = 1;
defparam ram_block1a79.init_file = "DDS_48_v1_nco_ii_0_cos.hex";
defparam ram_block1a79.init_file_layout = "port_a";
defparam ram_block1a79.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0121|altsyncram:altsyncram_component0|altsyncram_78g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a79.operation_mode = "rom";
defparam ram_block1a79.port_a_address_clear = "none";
defparam ram_block1a79.port_a_address_width = 13;
defparam ram_block1a79.port_a_data_out_clear = "none";
defparam ram_block1a79.port_a_data_out_clock = "clock0";
defparam ram_block1a79.port_a_data_width = 1;
defparam ram_block1a79.port_a_first_address = 32768;
defparam ram_block1a79.port_a_first_bit_number = 15;
defparam ram_block1a79.port_a_last_address = 40959;
defparam ram_block1a79.port_a_logical_ram_depth = 65536;
defparam ram_block1a79.port_a_logical_ram_width = 16;
defparam ram_block1a79.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a79.ram_block_type = "auto";
defparam ram_block1a79.mem_init3 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a79.mem_init2 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a79.mem_init1 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a79.mem_init0 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

arriav_ram_block ram_block1a95(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a95_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a95.clk0_core_clock_enable = "ena0";
defparam ram_block1a95.clk0_input_clock_enable = "ena0";
defparam ram_block1a95.clk0_output_clock_enable = "ena0";
defparam ram_block1a95.data_interleave_offset_in_bits = 1;
defparam ram_block1a95.data_interleave_width_in_bits = 1;
defparam ram_block1a95.init_file = "DDS_48_v1_nco_ii_0_cos.hex";
defparam ram_block1a95.init_file_layout = "port_a";
defparam ram_block1a95.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0121|altsyncram:altsyncram_component0|altsyncram_78g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a95.operation_mode = "rom";
defparam ram_block1a95.port_a_address_clear = "none";
defparam ram_block1a95.port_a_address_width = 13;
defparam ram_block1a95.port_a_data_out_clear = "none";
defparam ram_block1a95.port_a_data_out_clock = "clock0";
defparam ram_block1a95.port_a_data_width = 1;
defparam ram_block1a95.port_a_first_address = 40960;
defparam ram_block1a95.port_a_first_bit_number = 15;
defparam ram_block1a95.port_a_last_address = 49151;
defparam ram_block1a95.port_a_logical_ram_depth = 65536;
defparam ram_block1a95.port_a_logical_ram_width = 16;
defparam ram_block1a95.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a95.ram_block_type = "auto";
defparam ram_block1a95.mem_init3 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a95.mem_init2 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a95.mem_init1 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a95.mem_init0 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

arriav_ram_block ram_block1a111(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a111_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a111.clk0_core_clock_enable = "ena0";
defparam ram_block1a111.clk0_input_clock_enable = "ena0";
defparam ram_block1a111.clk0_output_clock_enable = "ena0";
defparam ram_block1a111.data_interleave_offset_in_bits = 1;
defparam ram_block1a111.data_interleave_width_in_bits = 1;
defparam ram_block1a111.init_file = "DDS_48_v1_nco_ii_0_cos.hex";
defparam ram_block1a111.init_file_layout = "port_a";
defparam ram_block1a111.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0121|altsyncram:altsyncram_component0|altsyncram_78g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a111.operation_mode = "rom";
defparam ram_block1a111.port_a_address_clear = "none";
defparam ram_block1a111.port_a_address_width = 13;
defparam ram_block1a111.port_a_data_out_clear = "none";
defparam ram_block1a111.port_a_data_out_clock = "clock0";
defparam ram_block1a111.port_a_data_width = 1;
defparam ram_block1a111.port_a_first_address = 49152;
defparam ram_block1a111.port_a_first_bit_number = 15;
defparam ram_block1a111.port_a_last_address = 57343;
defparam ram_block1a111.port_a_logical_ram_depth = 65536;
defparam ram_block1a111.port_a_logical_ram_width = 16;
defparam ram_block1a111.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a111.ram_block_type = "auto";
defparam ram_block1a111.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a111.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a111.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a111.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

arriav_ram_block ram_block1a127(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a127_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a127.clk0_core_clock_enable = "ena0";
defparam ram_block1a127.clk0_input_clock_enable = "ena0";
defparam ram_block1a127.clk0_output_clock_enable = "ena0";
defparam ram_block1a127.data_interleave_offset_in_bits = 1;
defparam ram_block1a127.data_interleave_width_in_bits = 1;
defparam ram_block1a127.init_file = "DDS_48_v1_nco_ii_0_cos.hex";
defparam ram_block1a127.init_file_layout = "port_a";
defparam ram_block1a127.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0121|altsyncram:altsyncram_component0|altsyncram_78g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a127.operation_mode = "rom";
defparam ram_block1a127.port_a_address_clear = "none";
defparam ram_block1a127.port_a_address_width = 13;
defparam ram_block1a127.port_a_data_out_clear = "none";
defparam ram_block1a127.port_a_data_out_clock = "clock0";
defparam ram_block1a127.port_a_data_width = 1;
defparam ram_block1a127.port_a_first_address = 57344;
defparam ram_block1a127.port_a_first_bit_number = 15;
defparam ram_block1a127.port_a_last_address = 65535;
defparam ram_block1a127.port_a_logical_ram_depth = 65536;
defparam ram_block1a127.port_a_logical_ram_width = 16;
defparam ram_block1a127.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a127.ram_block_type = "auto";
defparam ram_block1a127.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a127.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a127.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a127.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

arriav_ram_block ram_block1a47(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a47_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a47.clk0_core_clock_enable = "ena0";
defparam ram_block1a47.clk0_input_clock_enable = "ena0";
defparam ram_block1a47.clk0_output_clock_enable = "ena0";
defparam ram_block1a47.data_interleave_offset_in_bits = 1;
defparam ram_block1a47.data_interleave_width_in_bits = 1;
defparam ram_block1a47.init_file = "DDS_48_v1_nco_ii_0_cos.hex";
defparam ram_block1a47.init_file_layout = "port_a";
defparam ram_block1a47.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0121|altsyncram:altsyncram_component0|altsyncram_78g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a47.operation_mode = "rom";
defparam ram_block1a47.port_a_address_clear = "none";
defparam ram_block1a47.port_a_address_width = 13;
defparam ram_block1a47.port_a_data_out_clear = "none";
defparam ram_block1a47.port_a_data_out_clock = "clock0";
defparam ram_block1a47.port_a_data_width = 1;
defparam ram_block1a47.port_a_first_address = 16384;
defparam ram_block1a47.port_a_first_bit_number = 15;
defparam ram_block1a47.port_a_last_address = 24575;
defparam ram_block1a47.port_a_logical_ram_depth = 65536;
defparam ram_block1a47.port_a_logical_ram_width = 16;
defparam ram_block1a47.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a47.ram_block_type = "auto";
defparam ram_block1a47.mem_init3 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a47.mem_init2 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a47.mem_init1 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a47.mem_init0 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE";

arriav_ram_block ram_block1a63(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a63_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a63.clk0_core_clock_enable = "ena0";
defparam ram_block1a63.clk0_input_clock_enable = "ena0";
defparam ram_block1a63.clk0_output_clock_enable = "ena0";
defparam ram_block1a63.data_interleave_offset_in_bits = 1;
defparam ram_block1a63.data_interleave_width_in_bits = 1;
defparam ram_block1a63.init_file = "DDS_48_v1_nco_ii_0_cos.hex";
defparam ram_block1a63.init_file_layout = "port_a";
defparam ram_block1a63.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0121|altsyncram:altsyncram_component0|altsyncram_78g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a63.operation_mode = "rom";
defparam ram_block1a63.port_a_address_clear = "none";
defparam ram_block1a63.port_a_address_width = 13;
defparam ram_block1a63.port_a_data_out_clear = "none";
defparam ram_block1a63.port_a_data_out_clock = "clock0";
defparam ram_block1a63.port_a_data_width = 1;
defparam ram_block1a63.port_a_first_address = 24576;
defparam ram_block1a63.port_a_first_bit_number = 15;
defparam ram_block1a63.port_a_last_address = 32767;
defparam ram_block1a63.port_a_logical_ram_depth = 65536;
defparam ram_block1a63.port_a_logical_ram_width = 16;
defparam ram_block1a63.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a63.ram_block_type = "auto";
defparam ram_block1a63.mem_init3 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a63.mem_init2 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a63.mem_init1 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a63.mem_init0 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

arriav_ram_block ram_block1a15(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a15_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a15.clk0_core_clock_enable = "ena0";
defparam ram_block1a15.clk0_input_clock_enable = "ena0";
defparam ram_block1a15.clk0_output_clock_enable = "ena0";
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.init_file = "DDS_48_v1_nco_ii_0_cos.hex";
defparam ram_block1a15.init_file_layout = "port_a";
defparam ram_block1a15.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0121|altsyncram:altsyncram_component0|altsyncram_78g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a15.operation_mode = "rom";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 13;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "clock0";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 8191;
defparam ram_block1a15.port_a_logical_ram_depth = 65536;
defparam ram_block1a15.port_a_logical_ram_width = 16;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a15.ram_block_type = "auto";
defparam ram_block1a15.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a15.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a15.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a15.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

arriav_ram_block ram_block1a31(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a31_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a31.clk0_core_clock_enable = "ena0";
defparam ram_block1a31.clk0_input_clock_enable = "ena0";
defparam ram_block1a31.clk0_output_clock_enable = "ena0";
defparam ram_block1a31.data_interleave_offset_in_bits = 1;
defparam ram_block1a31.data_interleave_width_in_bits = 1;
defparam ram_block1a31.init_file = "DDS_48_v1_nco_ii_0_cos.hex";
defparam ram_block1a31.init_file_layout = "port_a";
defparam ram_block1a31.logical_ram_name = "DDS_48_v1_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0121|altsyncram:altsyncram_component0|altsyncram_78g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a31.operation_mode = "rom";
defparam ram_block1a31.port_a_address_clear = "none";
defparam ram_block1a31.port_a_address_width = 13;
defparam ram_block1a31.port_a_data_out_clear = "none";
defparam ram_block1a31.port_a_data_out_clock = "clock0";
defparam ram_block1a31.port_a_data_width = 1;
defparam ram_block1a31.port_a_first_address = 8192;
defparam ram_block1a31.port_a_first_bit_number = 15;
defparam ram_block1a31.port_a_last_address = 16383;
defparam ram_block1a31.port_a_logical_ram_depth = 65536;
defparam ram_block1a31.port_a_logical_ram_width = 16;
defparam ram_block1a31.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a31.ram_block_type = "auto";
defparam ram_block1a31.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a31.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a31.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a31.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

endmodule

module DDS_48_v1_asj_nco_fxx (
	pipeline_dffe_32,
	pipeline_dffe_33,
	pipeline_dffe_34,
	pipeline_dffe_35,
	pipeline_dffe_36,
	pipeline_dffe_37,
	pipeline_dffe_38,
	pipeline_dffe_39,
	pipeline_dffe_40,
	pipeline_dffe_41,
	pipeline_dffe_42,
	pipeline_dffe_43,
	pipeline_dffe_44,
	pipeline_dffe_47,
	pipeline_dffe_31,
	pipeline_dffe_45,
	pipeline_dffe_46,
	pipeline_dffe_30,
	pipeline_dffe_29,
	pipeline_dffe_28,
	pipeline_dffe_27,
	pipeline_dffe_26,
	pipeline_dffe_25,
	pipeline_dffe_24,
	pipeline_dffe_23,
	pipeline_dffe_22,
	pipeline_dffe_21,
	pipeline_dffe_20,
	pipeline_dffe_19,
	pipeline_dffe_18,
	pipeline_dffe_17,
	pipeline_dffe_16,
	pipeline_dffe_15,
	pipeline_dffe_14,
	pipeline_dffe_13,
	pipeline_dffe_12,
	pipeline_dffe_11,
	pipeline_dffe_10,
	pipeline_dffe_9,
	pipeline_dffe_8,
	pipeline_dffe_7,
	pipeline_dffe_6,
	pipeline_dffe_5,
	pipeline_dffe_4,
	pipeline_dffe_3,
	pipeline_dffe_2,
	pipeline_dffe_1,
	pipeline_dffe_0,
	clk,
	reset_n,
	clken,
	freq_mod_i_31,
	phi_inc_i_32,
	phi_inc_i_33,
	phi_inc_i_34,
	phi_inc_i_35,
	phi_inc_i_36,
	phi_inc_i_37,
	phi_inc_i_38,
	phi_inc_i_39,
	phi_inc_i_40,
	phi_inc_i_41,
	phi_inc_i_42,
	phi_inc_i_43,
	phi_inc_i_44,
	phi_inc_i_47,
	phi_inc_i_31,
	phi_inc_i_45,
	phi_inc_i_46,
	freq_mod_i_30,
	phi_inc_i_30,
	freq_mod_i_29,
	phi_inc_i_29,
	freq_mod_i_28,
	phi_inc_i_28,
	freq_mod_i_27,
	phi_inc_i_27,
	freq_mod_i_26,
	phi_inc_i_26,
	freq_mod_i_25,
	phi_inc_i_25,
	freq_mod_i_24,
	phi_inc_i_24,
	freq_mod_i_23,
	phi_inc_i_23,
	freq_mod_i_22,
	phi_inc_i_22,
	freq_mod_i_21,
	phi_inc_i_21,
	freq_mod_i_20,
	phi_inc_i_20,
	freq_mod_i_19,
	phi_inc_i_19,
	freq_mod_i_18,
	phi_inc_i_18,
	freq_mod_i_17,
	phi_inc_i_17,
	freq_mod_i_16,
	phi_inc_i_16,
	freq_mod_i_15,
	phi_inc_i_15,
	freq_mod_i_14,
	phi_inc_i_14,
	freq_mod_i_13,
	phi_inc_i_13,
	freq_mod_i_12,
	phi_inc_i_12,
	freq_mod_i_11,
	phi_inc_i_11,
	freq_mod_i_10,
	phi_inc_i_10,
	freq_mod_i_9,
	phi_inc_i_9,
	freq_mod_i_8,
	phi_inc_i_8,
	freq_mod_i_7,
	phi_inc_i_7,
	freq_mod_i_6,
	phi_inc_i_6,
	freq_mod_i_5,
	phi_inc_i_5,
	freq_mod_i_4,
	phi_inc_i_4,
	freq_mod_i_3,
	phi_inc_i_3,
	freq_mod_i_2,
	phi_inc_i_2,
	freq_mod_i_1,
	phi_inc_i_1,
	freq_mod_i_0,
	phi_inc_i_0)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_32;
output 	pipeline_dffe_33;
output 	pipeline_dffe_34;
output 	pipeline_dffe_35;
output 	pipeline_dffe_36;
output 	pipeline_dffe_37;
output 	pipeline_dffe_38;
output 	pipeline_dffe_39;
output 	pipeline_dffe_40;
output 	pipeline_dffe_41;
output 	pipeline_dffe_42;
output 	pipeline_dffe_43;
output 	pipeline_dffe_44;
output 	pipeline_dffe_47;
output 	pipeline_dffe_31;
output 	pipeline_dffe_45;
output 	pipeline_dffe_46;
output 	pipeline_dffe_30;
output 	pipeline_dffe_29;
output 	pipeline_dffe_28;
output 	pipeline_dffe_27;
output 	pipeline_dffe_26;
output 	pipeline_dffe_25;
output 	pipeline_dffe_24;
output 	pipeline_dffe_23;
output 	pipeline_dffe_22;
output 	pipeline_dffe_21;
output 	pipeline_dffe_20;
output 	pipeline_dffe_19;
output 	pipeline_dffe_18;
output 	pipeline_dffe_17;
output 	pipeline_dffe_16;
output 	pipeline_dffe_15;
output 	pipeline_dffe_14;
output 	pipeline_dffe_13;
output 	pipeline_dffe_12;
output 	pipeline_dffe_11;
output 	pipeline_dffe_10;
output 	pipeline_dffe_9;
output 	pipeline_dffe_8;
output 	pipeline_dffe_7;
output 	pipeline_dffe_6;
output 	pipeline_dffe_5;
output 	pipeline_dffe_4;
output 	pipeline_dffe_3;
output 	pipeline_dffe_2;
output 	pipeline_dffe_1;
output 	pipeline_dffe_0;
input 	clk;
input 	reset_n;
input 	clken;
input 	freq_mod_i_31;
input 	phi_inc_i_32;
input 	phi_inc_i_33;
input 	phi_inc_i_34;
input 	phi_inc_i_35;
input 	phi_inc_i_36;
input 	phi_inc_i_37;
input 	phi_inc_i_38;
input 	phi_inc_i_39;
input 	phi_inc_i_40;
input 	phi_inc_i_41;
input 	phi_inc_i_42;
input 	phi_inc_i_43;
input 	phi_inc_i_44;
input 	phi_inc_i_47;
input 	phi_inc_i_31;
input 	phi_inc_i_45;
input 	phi_inc_i_46;
input 	freq_mod_i_30;
input 	phi_inc_i_30;
input 	freq_mod_i_29;
input 	phi_inc_i_29;
input 	freq_mod_i_28;
input 	phi_inc_i_28;
input 	freq_mod_i_27;
input 	phi_inc_i_27;
input 	freq_mod_i_26;
input 	phi_inc_i_26;
input 	freq_mod_i_25;
input 	phi_inc_i_25;
input 	freq_mod_i_24;
input 	phi_inc_i_24;
input 	freq_mod_i_23;
input 	phi_inc_i_23;
input 	freq_mod_i_22;
input 	phi_inc_i_22;
input 	freq_mod_i_21;
input 	phi_inc_i_21;
input 	freq_mod_i_20;
input 	phi_inc_i_20;
input 	freq_mod_i_19;
input 	phi_inc_i_19;
input 	freq_mod_i_18;
input 	phi_inc_i_18;
input 	freq_mod_i_17;
input 	phi_inc_i_17;
input 	freq_mod_i_16;
input 	phi_inc_i_16;
input 	freq_mod_i_15;
input 	phi_inc_i_15;
input 	freq_mod_i_14;
input 	phi_inc_i_14;
input 	freq_mod_i_13;
input 	phi_inc_i_13;
input 	freq_mod_i_12;
input 	phi_inc_i_12;
input 	freq_mod_i_11;
input 	phi_inc_i_11;
input 	freq_mod_i_10;
input 	phi_inc_i_10;
input 	freq_mod_i_9;
input 	phi_inc_i_9;
input 	freq_mod_i_8;
input 	phi_inc_i_8;
input 	freq_mod_i_7;
input 	phi_inc_i_7;
input 	freq_mod_i_6;
input 	phi_inc_i_6;
input 	freq_mod_i_5;
input 	phi_inc_i_5;
input 	freq_mod_i_4;
input 	phi_inc_i_4;
input 	freq_mod_i_3;
input 	phi_inc_i_3;
input 	freq_mod_i_2;
input 	phi_inc_i_2;
input 	freq_mod_i_1;
input 	phi_inc_i_1;
input 	freq_mod_i_0;
input 	phi_inc_i_0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



DDS_48_v1_lpm_add_sub_2 acc(
	.pipeline_dffe_32(pipeline_dffe_32),
	.pipeline_dffe_33(pipeline_dffe_33),
	.pipeline_dffe_34(pipeline_dffe_34),
	.pipeline_dffe_35(pipeline_dffe_35),
	.pipeline_dffe_36(pipeline_dffe_36),
	.pipeline_dffe_37(pipeline_dffe_37),
	.pipeline_dffe_38(pipeline_dffe_38),
	.pipeline_dffe_39(pipeline_dffe_39),
	.pipeline_dffe_40(pipeline_dffe_40),
	.pipeline_dffe_41(pipeline_dffe_41),
	.pipeline_dffe_42(pipeline_dffe_42),
	.pipeline_dffe_43(pipeline_dffe_43),
	.pipeline_dffe_44(pipeline_dffe_44),
	.pipeline_dffe_47(pipeline_dffe_47),
	.pipeline_dffe_31(pipeline_dffe_31),
	.pipeline_dffe_45(pipeline_dffe_45),
	.pipeline_dffe_46(pipeline_dffe_46),
	.pipeline_dffe_30(pipeline_dffe_30),
	.pipeline_dffe_29(pipeline_dffe_29),
	.pipeline_dffe_28(pipeline_dffe_28),
	.pipeline_dffe_27(pipeline_dffe_27),
	.pipeline_dffe_26(pipeline_dffe_26),
	.pipeline_dffe_25(pipeline_dffe_25),
	.pipeline_dffe_24(pipeline_dffe_24),
	.pipeline_dffe_23(pipeline_dffe_23),
	.pipeline_dffe_22(pipeline_dffe_22),
	.pipeline_dffe_21(pipeline_dffe_21),
	.pipeline_dffe_20(pipeline_dffe_20),
	.pipeline_dffe_19(pipeline_dffe_19),
	.pipeline_dffe_18(pipeline_dffe_18),
	.pipeline_dffe_17(pipeline_dffe_17),
	.pipeline_dffe_16(pipeline_dffe_16),
	.pipeline_dffe_15(pipeline_dffe_15),
	.pipeline_dffe_14(pipeline_dffe_14),
	.pipeline_dffe_13(pipeline_dffe_13),
	.pipeline_dffe_12(pipeline_dffe_12),
	.pipeline_dffe_11(pipeline_dffe_11),
	.pipeline_dffe_10(pipeline_dffe_10),
	.pipeline_dffe_9(pipeline_dffe_9),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_1(pipeline_dffe_1),
	.pipeline_dffe_0(pipeline_dffe_0),
	.clock(clk),
	.reset_n(reset_n),
	.clken(clken),
	.freq_mod_i_31(freq_mod_i_31),
	.phi_inc_i_32(phi_inc_i_32),
	.phi_inc_i_33(phi_inc_i_33),
	.phi_inc_i_34(phi_inc_i_34),
	.phi_inc_i_35(phi_inc_i_35),
	.phi_inc_i_36(phi_inc_i_36),
	.phi_inc_i_37(phi_inc_i_37),
	.phi_inc_i_38(phi_inc_i_38),
	.phi_inc_i_39(phi_inc_i_39),
	.phi_inc_i_40(phi_inc_i_40),
	.phi_inc_i_41(phi_inc_i_41),
	.phi_inc_i_42(phi_inc_i_42),
	.phi_inc_i_43(phi_inc_i_43),
	.phi_inc_i_44(phi_inc_i_44),
	.phi_inc_i_47(phi_inc_i_47),
	.phi_inc_i_31(phi_inc_i_31),
	.phi_inc_i_45(phi_inc_i_45),
	.phi_inc_i_46(phi_inc_i_46),
	.freq_mod_i_30(freq_mod_i_30),
	.phi_inc_i_30(phi_inc_i_30),
	.freq_mod_i_29(freq_mod_i_29),
	.phi_inc_i_29(phi_inc_i_29),
	.freq_mod_i_28(freq_mod_i_28),
	.phi_inc_i_28(phi_inc_i_28),
	.freq_mod_i_27(freq_mod_i_27),
	.phi_inc_i_27(phi_inc_i_27),
	.freq_mod_i_26(freq_mod_i_26),
	.phi_inc_i_26(phi_inc_i_26),
	.freq_mod_i_25(freq_mod_i_25),
	.phi_inc_i_25(phi_inc_i_25),
	.freq_mod_i_24(freq_mod_i_24),
	.phi_inc_i_24(phi_inc_i_24),
	.freq_mod_i_23(freq_mod_i_23),
	.phi_inc_i_23(phi_inc_i_23),
	.freq_mod_i_22(freq_mod_i_22),
	.phi_inc_i_22(phi_inc_i_22),
	.freq_mod_i_21(freq_mod_i_21),
	.phi_inc_i_21(phi_inc_i_21),
	.freq_mod_i_20(freq_mod_i_20),
	.phi_inc_i_20(phi_inc_i_20),
	.freq_mod_i_19(freq_mod_i_19),
	.phi_inc_i_19(phi_inc_i_19),
	.freq_mod_i_18(freq_mod_i_18),
	.phi_inc_i_18(phi_inc_i_18),
	.freq_mod_i_17(freq_mod_i_17),
	.phi_inc_i_17(phi_inc_i_17),
	.freq_mod_i_16(freq_mod_i_16),
	.phi_inc_i_16(phi_inc_i_16),
	.freq_mod_i_15(freq_mod_i_15),
	.phi_inc_i_15(phi_inc_i_15),
	.freq_mod_i_14(freq_mod_i_14),
	.phi_inc_i_14(phi_inc_i_14),
	.freq_mod_i_13(freq_mod_i_13),
	.phi_inc_i_13(phi_inc_i_13),
	.freq_mod_i_12(freq_mod_i_12),
	.phi_inc_i_12(phi_inc_i_12),
	.freq_mod_i_11(freq_mod_i_11),
	.phi_inc_i_11(phi_inc_i_11),
	.freq_mod_i_10(freq_mod_i_10),
	.phi_inc_i_10(phi_inc_i_10),
	.freq_mod_i_9(freq_mod_i_9),
	.phi_inc_i_9(phi_inc_i_9),
	.freq_mod_i_8(freq_mod_i_8),
	.phi_inc_i_8(phi_inc_i_8),
	.freq_mod_i_7(freq_mod_i_7),
	.phi_inc_i_7(phi_inc_i_7),
	.freq_mod_i_6(freq_mod_i_6),
	.phi_inc_i_6(phi_inc_i_6),
	.freq_mod_i_5(freq_mod_i_5),
	.phi_inc_i_5(phi_inc_i_5),
	.freq_mod_i_4(freq_mod_i_4),
	.phi_inc_i_4(phi_inc_i_4),
	.freq_mod_i_3(freq_mod_i_3),
	.phi_inc_i_3(phi_inc_i_3),
	.freq_mod_i_2(freq_mod_i_2),
	.phi_inc_i_2(phi_inc_i_2),
	.freq_mod_i_1(freq_mod_i_1),
	.phi_inc_i_1(phi_inc_i_1),
	.freq_mod_i_0(freq_mod_i_0),
	.phi_inc_i_0(phi_inc_i_0));

endmodule

module DDS_48_v1_lpm_add_sub_2 (
	pipeline_dffe_32,
	pipeline_dffe_33,
	pipeline_dffe_34,
	pipeline_dffe_35,
	pipeline_dffe_36,
	pipeline_dffe_37,
	pipeline_dffe_38,
	pipeline_dffe_39,
	pipeline_dffe_40,
	pipeline_dffe_41,
	pipeline_dffe_42,
	pipeline_dffe_43,
	pipeline_dffe_44,
	pipeline_dffe_47,
	pipeline_dffe_31,
	pipeline_dffe_45,
	pipeline_dffe_46,
	pipeline_dffe_30,
	pipeline_dffe_29,
	pipeline_dffe_28,
	pipeline_dffe_27,
	pipeline_dffe_26,
	pipeline_dffe_25,
	pipeline_dffe_24,
	pipeline_dffe_23,
	pipeline_dffe_22,
	pipeline_dffe_21,
	pipeline_dffe_20,
	pipeline_dffe_19,
	pipeline_dffe_18,
	pipeline_dffe_17,
	pipeline_dffe_16,
	pipeline_dffe_15,
	pipeline_dffe_14,
	pipeline_dffe_13,
	pipeline_dffe_12,
	pipeline_dffe_11,
	pipeline_dffe_10,
	pipeline_dffe_9,
	pipeline_dffe_8,
	pipeline_dffe_7,
	pipeline_dffe_6,
	pipeline_dffe_5,
	pipeline_dffe_4,
	pipeline_dffe_3,
	pipeline_dffe_2,
	pipeline_dffe_1,
	pipeline_dffe_0,
	clock,
	reset_n,
	clken,
	freq_mod_i_31,
	phi_inc_i_32,
	phi_inc_i_33,
	phi_inc_i_34,
	phi_inc_i_35,
	phi_inc_i_36,
	phi_inc_i_37,
	phi_inc_i_38,
	phi_inc_i_39,
	phi_inc_i_40,
	phi_inc_i_41,
	phi_inc_i_42,
	phi_inc_i_43,
	phi_inc_i_44,
	phi_inc_i_47,
	phi_inc_i_31,
	phi_inc_i_45,
	phi_inc_i_46,
	freq_mod_i_30,
	phi_inc_i_30,
	freq_mod_i_29,
	phi_inc_i_29,
	freq_mod_i_28,
	phi_inc_i_28,
	freq_mod_i_27,
	phi_inc_i_27,
	freq_mod_i_26,
	phi_inc_i_26,
	freq_mod_i_25,
	phi_inc_i_25,
	freq_mod_i_24,
	phi_inc_i_24,
	freq_mod_i_23,
	phi_inc_i_23,
	freq_mod_i_22,
	phi_inc_i_22,
	freq_mod_i_21,
	phi_inc_i_21,
	freq_mod_i_20,
	phi_inc_i_20,
	freq_mod_i_19,
	phi_inc_i_19,
	freq_mod_i_18,
	phi_inc_i_18,
	freq_mod_i_17,
	phi_inc_i_17,
	freq_mod_i_16,
	phi_inc_i_16,
	freq_mod_i_15,
	phi_inc_i_15,
	freq_mod_i_14,
	phi_inc_i_14,
	freq_mod_i_13,
	phi_inc_i_13,
	freq_mod_i_12,
	phi_inc_i_12,
	freq_mod_i_11,
	phi_inc_i_11,
	freq_mod_i_10,
	phi_inc_i_10,
	freq_mod_i_9,
	phi_inc_i_9,
	freq_mod_i_8,
	phi_inc_i_8,
	freq_mod_i_7,
	phi_inc_i_7,
	freq_mod_i_6,
	phi_inc_i_6,
	freq_mod_i_5,
	phi_inc_i_5,
	freq_mod_i_4,
	phi_inc_i_4,
	freq_mod_i_3,
	phi_inc_i_3,
	freq_mod_i_2,
	phi_inc_i_2,
	freq_mod_i_1,
	phi_inc_i_1,
	freq_mod_i_0,
	phi_inc_i_0)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_32;
output 	pipeline_dffe_33;
output 	pipeline_dffe_34;
output 	pipeline_dffe_35;
output 	pipeline_dffe_36;
output 	pipeline_dffe_37;
output 	pipeline_dffe_38;
output 	pipeline_dffe_39;
output 	pipeline_dffe_40;
output 	pipeline_dffe_41;
output 	pipeline_dffe_42;
output 	pipeline_dffe_43;
output 	pipeline_dffe_44;
output 	pipeline_dffe_47;
output 	pipeline_dffe_31;
output 	pipeline_dffe_45;
output 	pipeline_dffe_46;
output 	pipeline_dffe_30;
output 	pipeline_dffe_29;
output 	pipeline_dffe_28;
output 	pipeline_dffe_27;
output 	pipeline_dffe_26;
output 	pipeline_dffe_25;
output 	pipeline_dffe_24;
output 	pipeline_dffe_23;
output 	pipeline_dffe_22;
output 	pipeline_dffe_21;
output 	pipeline_dffe_20;
output 	pipeline_dffe_19;
output 	pipeline_dffe_18;
output 	pipeline_dffe_17;
output 	pipeline_dffe_16;
output 	pipeline_dffe_15;
output 	pipeline_dffe_14;
output 	pipeline_dffe_13;
output 	pipeline_dffe_12;
output 	pipeline_dffe_11;
output 	pipeline_dffe_10;
output 	pipeline_dffe_9;
output 	pipeline_dffe_8;
output 	pipeline_dffe_7;
output 	pipeline_dffe_6;
output 	pipeline_dffe_5;
output 	pipeline_dffe_4;
output 	pipeline_dffe_3;
output 	pipeline_dffe_2;
output 	pipeline_dffe_1;
output 	pipeline_dffe_0;
input 	clock;
input 	reset_n;
input 	clken;
input 	freq_mod_i_31;
input 	phi_inc_i_32;
input 	phi_inc_i_33;
input 	phi_inc_i_34;
input 	phi_inc_i_35;
input 	phi_inc_i_36;
input 	phi_inc_i_37;
input 	phi_inc_i_38;
input 	phi_inc_i_39;
input 	phi_inc_i_40;
input 	phi_inc_i_41;
input 	phi_inc_i_42;
input 	phi_inc_i_43;
input 	phi_inc_i_44;
input 	phi_inc_i_47;
input 	phi_inc_i_31;
input 	phi_inc_i_45;
input 	phi_inc_i_46;
input 	freq_mod_i_30;
input 	phi_inc_i_30;
input 	freq_mod_i_29;
input 	phi_inc_i_29;
input 	freq_mod_i_28;
input 	phi_inc_i_28;
input 	freq_mod_i_27;
input 	phi_inc_i_27;
input 	freq_mod_i_26;
input 	phi_inc_i_26;
input 	freq_mod_i_25;
input 	phi_inc_i_25;
input 	freq_mod_i_24;
input 	phi_inc_i_24;
input 	freq_mod_i_23;
input 	phi_inc_i_23;
input 	freq_mod_i_22;
input 	phi_inc_i_22;
input 	freq_mod_i_21;
input 	phi_inc_i_21;
input 	freq_mod_i_20;
input 	phi_inc_i_20;
input 	freq_mod_i_19;
input 	phi_inc_i_19;
input 	freq_mod_i_18;
input 	phi_inc_i_18;
input 	freq_mod_i_17;
input 	phi_inc_i_17;
input 	freq_mod_i_16;
input 	phi_inc_i_16;
input 	freq_mod_i_15;
input 	phi_inc_i_15;
input 	freq_mod_i_14;
input 	phi_inc_i_14;
input 	freq_mod_i_13;
input 	phi_inc_i_13;
input 	freq_mod_i_12;
input 	phi_inc_i_12;
input 	freq_mod_i_11;
input 	phi_inc_i_11;
input 	freq_mod_i_10;
input 	phi_inc_i_10;
input 	freq_mod_i_9;
input 	phi_inc_i_9;
input 	freq_mod_i_8;
input 	phi_inc_i_8;
input 	freq_mod_i_7;
input 	phi_inc_i_7;
input 	freq_mod_i_6;
input 	phi_inc_i_6;
input 	freq_mod_i_5;
input 	phi_inc_i_5;
input 	freq_mod_i_4;
input 	phi_inc_i_4;
input 	freq_mod_i_3;
input 	phi_inc_i_3;
input 	freq_mod_i_2;
input 	phi_inc_i_2;
input 	freq_mod_i_1;
input 	phi_inc_i_1;
input 	freq_mod_i_0;
input 	phi_inc_i_0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



DDS_48_v1_add_sub_3qg auto_generated(
	.pipeline_dffe_32(pipeline_dffe_32),
	.pipeline_dffe_33(pipeline_dffe_33),
	.pipeline_dffe_34(pipeline_dffe_34),
	.pipeline_dffe_35(pipeline_dffe_35),
	.pipeline_dffe_36(pipeline_dffe_36),
	.pipeline_dffe_37(pipeline_dffe_37),
	.pipeline_dffe_38(pipeline_dffe_38),
	.pipeline_dffe_39(pipeline_dffe_39),
	.pipeline_dffe_40(pipeline_dffe_40),
	.pipeline_dffe_41(pipeline_dffe_41),
	.pipeline_dffe_42(pipeline_dffe_42),
	.pipeline_dffe_43(pipeline_dffe_43),
	.pipeline_dffe_44(pipeline_dffe_44),
	.pipeline_dffe_47(pipeline_dffe_47),
	.pipeline_dffe_31(pipeline_dffe_31),
	.pipeline_dffe_45(pipeline_dffe_45),
	.pipeline_dffe_46(pipeline_dffe_46),
	.pipeline_dffe_30(pipeline_dffe_30),
	.pipeline_dffe_29(pipeline_dffe_29),
	.pipeline_dffe_28(pipeline_dffe_28),
	.pipeline_dffe_27(pipeline_dffe_27),
	.pipeline_dffe_26(pipeline_dffe_26),
	.pipeline_dffe_25(pipeline_dffe_25),
	.pipeline_dffe_24(pipeline_dffe_24),
	.pipeline_dffe_23(pipeline_dffe_23),
	.pipeline_dffe_22(pipeline_dffe_22),
	.pipeline_dffe_21(pipeline_dffe_21),
	.pipeline_dffe_20(pipeline_dffe_20),
	.pipeline_dffe_19(pipeline_dffe_19),
	.pipeline_dffe_18(pipeline_dffe_18),
	.pipeline_dffe_17(pipeline_dffe_17),
	.pipeline_dffe_16(pipeline_dffe_16),
	.pipeline_dffe_15(pipeline_dffe_15),
	.pipeline_dffe_14(pipeline_dffe_14),
	.pipeline_dffe_13(pipeline_dffe_13),
	.pipeline_dffe_12(pipeline_dffe_12),
	.pipeline_dffe_11(pipeline_dffe_11),
	.pipeline_dffe_10(pipeline_dffe_10),
	.pipeline_dffe_9(pipeline_dffe_9),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_1(pipeline_dffe_1),
	.pipeline_dffe_0(pipeline_dffe_0),
	.clock(clock),
	.reset_n(reset_n),
	.clken(clken),
	.freq_mod_i_31(freq_mod_i_31),
	.phi_inc_i_32(phi_inc_i_32),
	.phi_inc_i_33(phi_inc_i_33),
	.phi_inc_i_34(phi_inc_i_34),
	.phi_inc_i_35(phi_inc_i_35),
	.phi_inc_i_36(phi_inc_i_36),
	.phi_inc_i_37(phi_inc_i_37),
	.phi_inc_i_38(phi_inc_i_38),
	.phi_inc_i_39(phi_inc_i_39),
	.phi_inc_i_40(phi_inc_i_40),
	.phi_inc_i_41(phi_inc_i_41),
	.phi_inc_i_42(phi_inc_i_42),
	.phi_inc_i_43(phi_inc_i_43),
	.phi_inc_i_44(phi_inc_i_44),
	.phi_inc_i_47(phi_inc_i_47),
	.phi_inc_i_31(phi_inc_i_31),
	.phi_inc_i_45(phi_inc_i_45),
	.phi_inc_i_46(phi_inc_i_46),
	.freq_mod_i_30(freq_mod_i_30),
	.phi_inc_i_30(phi_inc_i_30),
	.freq_mod_i_29(freq_mod_i_29),
	.phi_inc_i_29(phi_inc_i_29),
	.freq_mod_i_28(freq_mod_i_28),
	.phi_inc_i_28(phi_inc_i_28),
	.freq_mod_i_27(freq_mod_i_27),
	.phi_inc_i_27(phi_inc_i_27),
	.freq_mod_i_26(freq_mod_i_26),
	.phi_inc_i_26(phi_inc_i_26),
	.freq_mod_i_25(freq_mod_i_25),
	.phi_inc_i_25(phi_inc_i_25),
	.freq_mod_i_24(freq_mod_i_24),
	.phi_inc_i_24(phi_inc_i_24),
	.freq_mod_i_23(freq_mod_i_23),
	.phi_inc_i_23(phi_inc_i_23),
	.freq_mod_i_22(freq_mod_i_22),
	.phi_inc_i_22(phi_inc_i_22),
	.freq_mod_i_21(freq_mod_i_21),
	.phi_inc_i_21(phi_inc_i_21),
	.freq_mod_i_20(freq_mod_i_20),
	.phi_inc_i_20(phi_inc_i_20),
	.freq_mod_i_19(freq_mod_i_19),
	.phi_inc_i_19(phi_inc_i_19),
	.freq_mod_i_18(freq_mod_i_18),
	.phi_inc_i_18(phi_inc_i_18),
	.freq_mod_i_17(freq_mod_i_17),
	.phi_inc_i_17(phi_inc_i_17),
	.freq_mod_i_16(freq_mod_i_16),
	.phi_inc_i_16(phi_inc_i_16),
	.freq_mod_i_15(freq_mod_i_15),
	.phi_inc_i_15(phi_inc_i_15),
	.freq_mod_i_14(freq_mod_i_14),
	.phi_inc_i_14(phi_inc_i_14),
	.freq_mod_i_13(freq_mod_i_13),
	.phi_inc_i_13(phi_inc_i_13),
	.freq_mod_i_12(freq_mod_i_12),
	.phi_inc_i_12(phi_inc_i_12),
	.freq_mod_i_11(freq_mod_i_11),
	.phi_inc_i_11(phi_inc_i_11),
	.freq_mod_i_10(freq_mod_i_10),
	.phi_inc_i_10(phi_inc_i_10),
	.freq_mod_i_9(freq_mod_i_9),
	.phi_inc_i_9(phi_inc_i_9),
	.freq_mod_i_8(freq_mod_i_8),
	.phi_inc_i_8(phi_inc_i_8),
	.freq_mod_i_7(freq_mod_i_7),
	.phi_inc_i_7(phi_inc_i_7),
	.freq_mod_i_6(freq_mod_i_6),
	.phi_inc_i_6(phi_inc_i_6),
	.freq_mod_i_5(freq_mod_i_5),
	.phi_inc_i_5(phi_inc_i_5),
	.freq_mod_i_4(freq_mod_i_4),
	.phi_inc_i_4(phi_inc_i_4),
	.freq_mod_i_3(freq_mod_i_3),
	.phi_inc_i_3(phi_inc_i_3),
	.freq_mod_i_2(freq_mod_i_2),
	.phi_inc_i_2(phi_inc_i_2),
	.freq_mod_i_1(freq_mod_i_1),
	.phi_inc_i_1(phi_inc_i_1),
	.freq_mod_i_0(freq_mod_i_0),
	.phi_inc_i_0(phi_inc_i_0));

endmodule

module DDS_48_v1_add_sub_3qg (
	pipeline_dffe_32,
	pipeline_dffe_33,
	pipeline_dffe_34,
	pipeline_dffe_35,
	pipeline_dffe_36,
	pipeline_dffe_37,
	pipeline_dffe_38,
	pipeline_dffe_39,
	pipeline_dffe_40,
	pipeline_dffe_41,
	pipeline_dffe_42,
	pipeline_dffe_43,
	pipeline_dffe_44,
	pipeline_dffe_47,
	pipeline_dffe_31,
	pipeline_dffe_45,
	pipeline_dffe_46,
	pipeline_dffe_30,
	pipeline_dffe_29,
	pipeline_dffe_28,
	pipeline_dffe_27,
	pipeline_dffe_26,
	pipeline_dffe_25,
	pipeline_dffe_24,
	pipeline_dffe_23,
	pipeline_dffe_22,
	pipeline_dffe_21,
	pipeline_dffe_20,
	pipeline_dffe_19,
	pipeline_dffe_18,
	pipeline_dffe_17,
	pipeline_dffe_16,
	pipeline_dffe_15,
	pipeline_dffe_14,
	pipeline_dffe_13,
	pipeline_dffe_12,
	pipeline_dffe_11,
	pipeline_dffe_10,
	pipeline_dffe_9,
	pipeline_dffe_8,
	pipeline_dffe_7,
	pipeline_dffe_6,
	pipeline_dffe_5,
	pipeline_dffe_4,
	pipeline_dffe_3,
	pipeline_dffe_2,
	pipeline_dffe_1,
	pipeline_dffe_0,
	clock,
	reset_n,
	clken,
	freq_mod_i_31,
	phi_inc_i_32,
	phi_inc_i_33,
	phi_inc_i_34,
	phi_inc_i_35,
	phi_inc_i_36,
	phi_inc_i_37,
	phi_inc_i_38,
	phi_inc_i_39,
	phi_inc_i_40,
	phi_inc_i_41,
	phi_inc_i_42,
	phi_inc_i_43,
	phi_inc_i_44,
	phi_inc_i_47,
	phi_inc_i_31,
	phi_inc_i_45,
	phi_inc_i_46,
	freq_mod_i_30,
	phi_inc_i_30,
	freq_mod_i_29,
	phi_inc_i_29,
	freq_mod_i_28,
	phi_inc_i_28,
	freq_mod_i_27,
	phi_inc_i_27,
	freq_mod_i_26,
	phi_inc_i_26,
	freq_mod_i_25,
	phi_inc_i_25,
	freq_mod_i_24,
	phi_inc_i_24,
	freq_mod_i_23,
	phi_inc_i_23,
	freq_mod_i_22,
	phi_inc_i_22,
	freq_mod_i_21,
	phi_inc_i_21,
	freq_mod_i_20,
	phi_inc_i_20,
	freq_mod_i_19,
	phi_inc_i_19,
	freq_mod_i_18,
	phi_inc_i_18,
	freq_mod_i_17,
	phi_inc_i_17,
	freq_mod_i_16,
	phi_inc_i_16,
	freq_mod_i_15,
	phi_inc_i_15,
	freq_mod_i_14,
	phi_inc_i_14,
	freq_mod_i_13,
	phi_inc_i_13,
	freq_mod_i_12,
	phi_inc_i_12,
	freq_mod_i_11,
	phi_inc_i_11,
	freq_mod_i_10,
	phi_inc_i_10,
	freq_mod_i_9,
	phi_inc_i_9,
	freq_mod_i_8,
	phi_inc_i_8,
	freq_mod_i_7,
	phi_inc_i_7,
	freq_mod_i_6,
	phi_inc_i_6,
	freq_mod_i_5,
	phi_inc_i_5,
	freq_mod_i_4,
	phi_inc_i_4,
	freq_mod_i_3,
	phi_inc_i_3,
	freq_mod_i_2,
	phi_inc_i_2,
	freq_mod_i_1,
	phi_inc_i_1,
	freq_mod_i_0,
	phi_inc_i_0)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_32;
output 	pipeline_dffe_33;
output 	pipeline_dffe_34;
output 	pipeline_dffe_35;
output 	pipeline_dffe_36;
output 	pipeline_dffe_37;
output 	pipeline_dffe_38;
output 	pipeline_dffe_39;
output 	pipeline_dffe_40;
output 	pipeline_dffe_41;
output 	pipeline_dffe_42;
output 	pipeline_dffe_43;
output 	pipeline_dffe_44;
output 	pipeline_dffe_47;
output 	pipeline_dffe_31;
output 	pipeline_dffe_45;
output 	pipeline_dffe_46;
output 	pipeline_dffe_30;
output 	pipeline_dffe_29;
output 	pipeline_dffe_28;
output 	pipeline_dffe_27;
output 	pipeline_dffe_26;
output 	pipeline_dffe_25;
output 	pipeline_dffe_24;
output 	pipeline_dffe_23;
output 	pipeline_dffe_22;
output 	pipeline_dffe_21;
output 	pipeline_dffe_20;
output 	pipeline_dffe_19;
output 	pipeline_dffe_18;
output 	pipeline_dffe_17;
output 	pipeline_dffe_16;
output 	pipeline_dffe_15;
output 	pipeline_dffe_14;
output 	pipeline_dffe_13;
output 	pipeline_dffe_12;
output 	pipeline_dffe_11;
output 	pipeline_dffe_10;
output 	pipeline_dffe_9;
output 	pipeline_dffe_8;
output 	pipeline_dffe_7;
output 	pipeline_dffe_6;
output 	pipeline_dffe_5;
output 	pipeline_dffe_4;
output 	pipeline_dffe_3;
output 	pipeline_dffe_2;
output 	pipeline_dffe_1;
output 	pipeline_dffe_0;
input 	clock;
input 	reset_n;
input 	clken;
input 	freq_mod_i_31;
input 	phi_inc_i_32;
input 	phi_inc_i_33;
input 	phi_inc_i_34;
input 	phi_inc_i_35;
input 	phi_inc_i_36;
input 	phi_inc_i_37;
input 	phi_inc_i_38;
input 	phi_inc_i_39;
input 	phi_inc_i_40;
input 	phi_inc_i_41;
input 	phi_inc_i_42;
input 	phi_inc_i_43;
input 	phi_inc_i_44;
input 	phi_inc_i_47;
input 	phi_inc_i_31;
input 	phi_inc_i_45;
input 	phi_inc_i_46;
input 	freq_mod_i_30;
input 	phi_inc_i_30;
input 	freq_mod_i_29;
input 	phi_inc_i_29;
input 	freq_mod_i_28;
input 	phi_inc_i_28;
input 	freq_mod_i_27;
input 	phi_inc_i_27;
input 	freq_mod_i_26;
input 	phi_inc_i_26;
input 	freq_mod_i_25;
input 	phi_inc_i_25;
input 	freq_mod_i_24;
input 	phi_inc_i_24;
input 	freq_mod_i_23;
input 	phi_inc_i_23;
input 	freq_mod_i_22;
input 	phi_inc_i_22;
input 	freq_mod_i_21;
input 	phi_inc_i_21;
input 	freq_mod_i_20;
input 	phi_inc_i_20;
input 	freq_mod_i_19;
input 	phi_inc_i_19;
input 	freq_mod_i_18;
input 	phi_inc_i_18;
input 	freq_mod_i_17;
input 	phi_inc_i_17;
input 	freq_mod_i_16;
input 	phi_inc_i_16;
input 	freq_mod_i_15;
input 	phi_inc_i_15;
input 	freq_mod_i_14;
input 	phi_inc_i_14;
input 	freq_mod_i_13;
input 	phi_inc_i_13;
input 	freq_mod_i_12;
input 	phi_inc_i_12;
input 	freq_mod_i_11;
input 	phi_inc_i_11;
input 	freq_mod_i_10;
input 	phi_inc_i_10;
input 	freq_mod_i_9;
input 	phi_inc_i_9;
input 	freq_mod_i_8;
input 	phi_inc_i_8;
input 	freq_mod_i_7;
input 	phi_inc_i_7;
input 	freq_mod_i_6;
input 	phi_inc_i_6;
input 	freq_mod_i_5;
input 	phi_inc_i_5;
input 	freq_mod_i_4;
input 	phi_inc_i_4;
input 	freq_mod_i_3;
input 	phi_inc_i_3;
input 	freq_mod_i_2;
input 	phi_inc_i_2;
input 	freq_mod_i_1;
input 	phi_inc_i_1;
input 	freq_mod_i_0;
input 	phi_inc_i_0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \op_1~190 ;
wire \op_1~186 ;
wire \op_1~182 ;
wire \op_1~178 ;
wire \op_1~174 ;
wire \op_1~170 ;
wire \op_1~166 ;
wire \op_1~162 ;
wire \op_1~158 ;
wire \op_1~154 ;
wire \op_1~150 ;
wire \op_1~146 ;
wire \op_1~142 ;
wire \op_1~138 ;
wire \op_1~134 ;
wire \op_1~130 ;
wire \op_1~126 ;
wire \op_1~122 ;
wire \op_1~118 ;
wire \op_1~114 ;
wire \op_1~110 ;
wire \op_1~106 ;
wire \op_1~102 ;
wire \op_1~98 ;
wire \op_1~94 ;
wire \op_1~90 ;
wire \op_1~86 ;
wire \op_1~82 ;
wire \op_1~78 ;
wire \op_1~74 ;
wire \op_1~70 ;
wire \op_1~58 ;
wire \op_1~1_sumout ;
wire \op_1~2 ;
wire \op_1~5_sumout ;
wire \op_1~6 ;
wire \op_1~9_sumout ;
wire \op_1~10 ;
wire \op_1~13_sumout ;
wire \op_1~14 ;
wire \op_1~17_sumout ;
wire \op_1~18 ;
wire \op_1~21_sumout ;
wire \op_1~22 ;
wire \op_1~25_sumout ;
wire \op_1~26 ;
wire \op_1~29_sumout ;
wire \op_1~30 ;
wire \op_1~33_sumout ;
wire \op_1~34 ;
wire \op_1~37_sumout ;
wire \op_1~38 ;
wire \op_1~41_sumout ;
wire \op_1~42 ;
wire \op_1~45_sumout ;
wire \op_1~46 ;
wire \op_1~49_sumout ;
wire \op_1~50 ;
wire \op_1~62 ;
wire \op_1~66 ;
wire \op_1~53_sumout ;
wire \op_1~57_sumout ;
wire \op_1~61_sumout ;
wire \op_1~65_sumout ;
wire \op_1~69_sumout ;
wire \op_1~73_sumout ;
wire \op_1~77_sumout ;
wire \op_1~81_sumout ;
wire \op_1~85_sumout ;
wire \op_1~89_sumout ;
wire \op_1~93_sumout ;
wire \op_1~97_sumout ;
wire \op_1~101_sumout ;
wire \op_1~105_sumout ;
wire \op_1~109_sumout ;
wire \op_1~113_sumout ;
wire \op_1~117_sumout ;
wire \op_1~121_sumout ;
wire \op_1~125_sumout ;
wire \op_1~129_sumout ;
wire \op_1~133_sumout ;
wire \op_1~137_sumout ;
wire \op_1~141_sumout ;
wire \op_1~145_sumout ;
wire \op_1~149_sumout ;
wire \op_1~153_sumout ;
wire \op_1~157_sumout ;
wire \op_1~161_sumout ;
wire \op_1~165_sumout ;
wire \op_1~169_sumout ;
wire \op_1~173_sumout ;
wire \op_1~177_sumout ;
wire \op_1~181_sumout ;
wire \op_1~185_sumout ;
wire \op_1~189_sumout ;


dffeas \pipeline_dffe[32] (
	.clk(clock),
	.d(\op_1~1_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_32),
	.prn(vcc));
defparam \pipeline_dffe[32] .is_wysiwyg = "true";
defparam \pipeline_dffe[32] .power_up = "low";

dffeas \pipeline_dffe[33] (
	.clk(clock),
	.d(\op_1~5_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_33),
	.prn(vcc));
defparam \pipeline_dffe[33] .is_wysiwyg = "true";
defparam \pipeline_dffe[33] .power_up = "low";

dffeas \pipeline_dffe[34] (
	.clk(clock),
	.d(\op_1~9_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_34),
	.prn(vcc));
defparam \pipeline_dffe[34] .is_wysiwyg = "true";
defparam \pipeline_dffe[34] .power_up = "low";

dffeas \pipeline_dffe[35] (
	.clk(clock),
	.d(\op_1~13_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_35),
	.prn(vcc));
defparam \pipeline_dffe[35] .is_wysiwyg = "true";
defparam \pipeline_dffe[35] .power_up = "low";

dffeas \pipeline_dffe[36] (
	.clk(clock),
	.d(\op_1~17_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_36),
	.prn(vcc));
defparam \pipeline_dffe[36] .is_wysiwyg = "true";
defparam \pipeline_dffe[36] .power_up = "low";

dffeas \pipeline_dffe[37] (
	.clk(clock),
	.d(\op_1~21_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_37),
	.prn(vcc));
defparam \pipeline_dffe[37] .is_wysiwyg = "true";
defparam \pipeline_dffe[37] .power_up = "low";

dffeas \pipeline_dffe[38] (
	.clk(clock),
	.d(\op_1~25_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_38),
	.prn(vcc));
defparam \pipeline_dffe[38] .is_wysiwyg = "true";
defparam \pipeline_dffe[38] .power_up = "low";

dffeas \pipeline_dffe[39] (
	.clk(clock),
	.d(\op_1~29_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_39),
	.prn(vcc));
defparam \pipeline_dffe[39] .is_wysiwyg = "true";
defparam \pipeline_dffe[39] .power_up = "low";

dffeas \pipeline_dffe[40] (
	.clk(clock),
	.d(\op_1~33_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_40),
	.prn(vcc));
defparam \pipeline_dffe[40] .is_wysiwyg = "true";
defparam \pipeline_dffe[40] .power_up = "low";

dffeas \pipeline_dffe[41] (
	.clk(clock),
	.d(\op_1~37_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_41),
	.prn(vcc));
defparam \pipeline_dffe[41] .is_wysiwyg = "true";
defparam \pipeline_dffe[41] .power_up = "low";

dffeas \pipeline_dffe[42] (
	.clk(clock),
	.d(\op_1~41_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_42),
	.prn(vcc));
defparam \pipeline_dffe[42] .is_wysiwyg = "true";
defparam \pipeline_dffe[42] .power_up = "low";

dffeas \pipeline_dffe[43] (
	.clk(clock),
	.d(\op_1~45_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_43),
	.prn(vcc));
defparam \pipeline_dffe[43] .is_wysiwyg = "true";
defparam \pipeline_dffe[43] .power_up = "low";

dffeas \pipeline_dffe[44] (
	.clk(clock),
	.d(\op_1~49_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_44),
	.prn(vcc));
defparam \pipeline_dffe[44] .is_wysiwyg = "true";
defparam \pipeline_dffe[44] .power_up = "low";

dffeas \pipeline_dffe[47] (
	.clk(clock),
	.d(\op_1~53_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_47),
	.prn(vcc));
defparam \pipeline_dffe[47] .is_wysiwyg = "true";
defparam \pipeline_dffe[47] .power_up = "low";

dffeas \pipeline_dffe[31] (
	.clk(clock),
	.d(\op_1~57_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_31),
	.prn(vcc));
defparam \pipeline_dffe[31] .is_wysiwyg = "true";
defparam \pipeline_dffe[31] .power_up = "low";

dffeas \pipeline_dffe[45] (
	.clk(clock),
	.d(\op_1~61_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_45),
	.prn(vcc));
defparam \pipeline_dffe[45] .is_wysiwyg = "true";
defparam \pipeline_dffe[45] .power_up = "low";

dffeas \pipeline_dffe[46] (
	.clk(clock),
	.d(\op_1~65_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_46),
	.prn(vcc));
defparam \pipeline_dffe[46] .is_wysiwyg = "true";
defparam \pipeline_dffe[46] .power_up = "low";

dffeas \pipeline_dffe[30] (
	.clk(clock),
	.d(\op_1~69_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_30),
	.prn(vcc));
defparam \pipeline_dffe[30] .is_wysiwyg = "true";
defparam \pipeline_dffe[30] .power_up = "low";

dffeas \pipeline_dffe[29] (
	.clk(clock),
	.d(\op_1~73_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_29),
	.prn(vcc));
defparam \pipeline_dffe[29] .is_wysiwyg = "true";
defparam \pipeline_dffe[29] .power_up = "low";

dffeas \pipeline_dffe[28] (
	.clk(clock),
	.d(\op_1~77_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_28),
	.prn(vcc));
defparam \pipeline_dffe[28] .is_wysiwyg = "true";
defparam \pipeline_dffe[28] .power_up = "low";

dffeas \pipeline_dffe[27] (
	.clk(clock),
	.d(\op_1~81_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_27),
	.prn(vcc));
defparam \pipeline_dffe[27] .is_wysiwyg = "true";
defparam \pipeline_dffe[27] .power_up = "low";

dffeas \pipeline_dffe[26] (
	.clk(clock),
	.d(\op_1~85_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_26),
	.prn(vcc));
defparam \pipeline_dffe[26] .is_wysiwyg = "true";
defparam \pipeline_dffe[26] .power_up = "low";

dffeas \pipeline_dffe[25] (
	.clk(clock),
	.d(\op_1~89_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_25),
	.prn(vcc));
defparam \pipeline_dffe[25] .is_wysiwyg = "true";
defparam \pipeline_dffe[25] .power_up = "low";

dffeas \pipeline_dffe[24] (
	.clk(clock),
	.d(\op_1~93_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_24),
	.prn(vcc));
defparam \pipeline_dffe[24] .is_wysiwyg = "true";
defparam \pipeline_dffe[24] .power_up = "low";

dffeas \pipeline_dffe[23] (
	.clk(clock),
	.d(\op_1~97_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_23),
	.prn(vcc));
defparam \pipeline_dffe[23] .is_wysiwyg = "true";
defparam \pipeline_dffe[23] .power_up = "low";

dffeas \pipeline_dffe[22] (
	.clk(clock),
	.d(\op_1~101_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_22),
	.prn(vcc));
defparam \pipeline_dffe[22] .is_wysiwyg = "true";
defparam \pipeline_dffe[22] .power_up = "low";

dffeas \pipeline_dffe[21] (
	.clk(clock),
	.d(\op_1~105_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_21),
	.prn(vcc));
defparam \pipeline_dffe[21] .is_wysiwyg = "true";
defparam \pipeline_dffe[21] .power_up = "low";

dffeas \pipeline_dffe[20] (
	.clk(clock),
	.d(\op_1~109_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_20),
	.prn(vcc));
defparam \pipeline_dffe[20] .is_wysiwyg = "true";
defparam \pipeline_dffe[20] .power_up = "low";

dffeas \pipeline_dffe[19] (
	.clk(clock),
	.d(\op_1~113_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_19),
	.prn(vcc));
defparam \pipeline_dffe[19] .is_wysiwyg = "true";
defparam \pipeline_dffe[19] .power_up = "low";

dffeas \pipeline_dffe[18] (
	.clk(clock),
	.d(\op_1~117_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_18),
	.prn(vcc));
defparam \pipeline_dffe[18] .is_wysiwyg = "true";
defparam \pipeline_dffe[18] .power_up = "low";

dffeas \pipeline_dffe[17] (
	.clk(clock),
	.d(\op_1~121_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_17),
	.prn(vcc));
defparam \pipeline_dffe[17] .is_wysiwyg = "true";
defparam \pipeline_dffe[17] .power_up = "low";

dffeas \pipeline_dffe[16] (
	.clk(clock),
	.d(\op_1~125_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_16),
	.prn(vcc));
defparam \pipeline_dffe[16] .is_wysiwyg = "true";
defparam \pipeline_dffe[16] .power_up = "low";

dffeas \pipeline_dffe[15] (
	.clk(clock),
	.d(\op_1~129_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_15),
	.prn(vcc));
defparam \pipeline_dffe[15] .is_wysiwyg = "true";
defparam \pipeline_dffe[15] .power_up = "low";

dffeas \pipeline_dffe[14] (
	.clk(clock),
	.d(\op_1~133_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_14),
	.prn(vcc));
defparam \pipeline_dffe[14] .is_wysiwyg = "true";
defparam \pipeline_dffe[14] .power_up = "low";

dffeas \pipeline_dffe[13] (
	.clk(clock),
	.d(\op_1~137_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_13),
	.prn(vcc));
defparam \pipeline_dffe[13] .is_wysiwyg = "true";
defparam \pipeline_dffe[13] .power_up = "low";

dffeas \pipeline_dffe[12] (
	.clk(clock),
	.d(\op_1~141_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_12),
	.prn(vcc));
defparam \pipeline_dffe[12] .is_wysiwyg = "true";
defparam \pipeline_dffe[12] .power_up = "low";

dffeas \pipeline_dffe[11] (
	.clk(clock),
	.d(\op_1~145_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_11),
	.prn(vcc));
defparam \pipeline_dffe[11] .is_wysiwyg = "true";
defparam \pipeline_dffe[11] .power_up = "low";

dffeas \pipeline_dffe[10] (
	.clk(clock),
	.d(\op_1~149_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_10),
	.prn(vcc));
defparam \pipeline_dffe[10] .is_wysiwyg = "true";
defparam \pipeline_dffe[10] .power_up = "low";

dffeas \pipeline_dffe[9] (
	.clk(clock),
	.d(\op_1~153_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_9),
	.prn(vcc));
defparam \pipeline_dffe[9] .is_wysiwyg = "true";
defparam \pipeline_dffe[9] .power_up = "low";

dffeas \pipeline_dffe[8] (
	.clk(clock),
	.d(\op_1~157_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_8),
	.prn(vcc));
defparam \pipeline_dffe[8] .is_wysiwyg = "true";
defparam \pipeline_dffe[8] .power_up = "low";

dffeas \pipeline_dffe[7] (
	.clk(clock),
	.d(\op_1~161_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_7),
	.prn(vcc));
defparam \pipeline_dffe[7] .is_wysiwyg = "true";
defparam \pipeline_dffe[7] .power_up = "low";

dffeas \pipeline_dffe[6] (
	.clk(clock),
	.d(\op_1~165_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_6),
	.prn(vcc));
defparam \pipeline_dffe[6] .is_wysiwyg = "true";
defparam \pipeline_dffe[6] .power_up = "low";

dffeas \pipeline_dffe[5] (
	.clk(clock),
	.d(\op_1~169_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_5),
	.prn(vcc));
defparam \pipeline_dffe[5] .is_wysiwyg = "true";
defparam \pipeline_dffe[5] .power_up = "low";

dffeas \pipeline_dffe[4] (
	.clk(clock),
	.d(\op_1~173_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_4),
	.prn(vcc));
defparam \pipeline_dffe[4] .is_wysiwyg = "true";
defparam \pipeline_dffe[4] .power_up = "low";

dffeas \pipeline_dffe[3] (
	.clk(clock),
	.d(\op_1~177_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_3),
	.prn(vcc));
defparam \pipeline_dffe[3] .is_wysiwyg = "true";
defparam \pipeline_dffe[3] .power_up = "low";

dffeas \pipeline_dffe[2] (
	.clk(clock),
	.d(\op_1~181_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_2),
	.prn(vcc));
defparam \pipeline_dffe[2] .is_wysiwyg = "true";
defparam \pipeline_dffe[2] .power_up = "low";

dffeas \pipeline_dffe[1] (
	.clk(clock),
	.d(\op_1~185_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_1),
	.prn(vcc));
defparam \pipeline_dffe[1] .is_wysiwyg = "true";
defparam \pipeline_dffe[1] .power_up = "low";

dffeas \pipeline_dffe[0] (
	.clk(clock),
	.d(\op_1~189_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_0),
	.prn(vcc));
defparam \pipeline_dffe[0] .is_wysiwyg = "true";
defparam \pipeline_dffe[0] .power_up = "low";

arriav_lcell_comb \op_1~189 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!freq_mod_i_0),
	.datae(gnd),
	.dataf(!phi_inc_i_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~189_sumout ),
	.cout(\op_1~190 ),
	.shareout());
defparam \op_1~189 .extended_lut = "off";
defparam \op_1~189 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~189 .shared_arith = "off";

arriav_lcell_comb \op_1~185 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!freq_mod_i_1),
	.datae(gnd),
	.dataf(!phi_inc_i_1),
	.datag(gnd),
	.cin(\op_1~190 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~185_sumout ),
	.cout(\op_1~186 ),
	.shareout());
defparam \op_1~185 .extended_lut = "off";
defparam \op_1~185 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~185 .shared_arith = "off";

arriav_lcell_comb \op_1~181 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!freq_mod_i_2),
	.datae(gnd),
	.dataf(!phi_inc_i_2),
	.datag(gnd),
	.cin(\op_1~186 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~181_sumout ),
	.cout(\op_1~182 ),
	.shareout());
defparam \op_1~181 .extended_lut = "off";
defparam \op_1~181 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~181 .shared_arith = "off";

arriav_lcell_comb \op_1~177 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!freq_mod_i_3),
	.datae(gnd),
	.dataf(!phi_inc_i_3),
	.datag(gnd),
	.cin(\op_1~182 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~177_sumout ),
	.cout(\op_1~178 ),
	.shareout());
defparam \op_1~177 .extended_lut = "off";
defparam \op_1~177 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~177 .shared_arith = "off";

arriav_lcell_comb \op_1~173 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!freq_mod_i_4),
	.datae(gnd),
	.dataf(!phi_inc_i_4),
	.datag(gnd),
	.cin(\op_1~178 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~173_sumout ),
	.cout(\op_1~174 ),
	.shareout());
defparam \op_1~173 .extended_lut = "off";
defparam \op_1~173 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~173 .shared_arith = "off";

arriav_lcell_comb \op_1~169 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!freq_mod_i_5),
	.datae(gnd),
	.dataf(!phi_inc_i_5),
	.datag(gnd),
	.cin(\op_1~174 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~169_sumout ),
	.cout(\op_1~170 ),
	.shareout());
defparam \op_1~169 .extended_lut = "off";
defparam \op_1~169 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~169 .shared_arith = "off";

arriav_lcell_comb \op_1~165 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!freq_mod_i_6),
	.datae(gnd),
	.dataf(!phi_inc_i_6),
	.datag(gnd),
	.cin(\op_1~170 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~165_sumout ),
	.cout(\op_1~166 ),
	.shareout());
defparam \op_1~165 .extended_lut = "off";
defparam \op_1~165 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~165 .shared_arith = "off";

arriav_lcell_comb \op_1~161 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!freq_mod_i_7),
	.datae(gnd),
	.dataf(!phi_inc_i_7),
	.datag(gnd),
	.cin(\op_1~166 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~161_sumout ),
	.cout(\op_1~162 ),
	.shareout());
defparam \op_1~161 .extended_lut = "off";
defparam \op_1~161 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~161 .shared_arith = "off";

arriav_lcell_comb \op_1~157 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!freq_mod_i_8),
	.datae(gnd),
	.dataf(!phi_inc_i_8),
	.datag(gnd),
	.cin(\op_1~162 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~157_sumout ),
	.cout(\op_1~158 ),
	.shareout());
defparam \op_1~157 .extended_lut = "off";
defparam \op_1~157 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~157 .shared_arith = "off";

arriav_lcell_comb \op_1~153 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!freq_mod_i_9),
	.datae(gnd),
	.dataf(!phi_inc_i_9),
	.datag(gnd),
	.cin(\op_1~158 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~153_sumout ),
	.cout(\op_1~154 ),
	.shareout());
defparam \op_1~153 .extended_lut = "off";
defparam \op_1~153 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~153 .shared_arith = "off";

arriav_lcell_comb \op_1~149 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!freq_mod_i_10),
	.datae(gnd),
	.dataf(!phi_inc_i_10),
	.datag(gnd),
	.cin(\op_1~154 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~149_sumout ),
	.cout(\op_1~150 ),
	.shareout());
defparam \op_1~149 .extended_lut = "off";
defparam \op_1~149 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~149 .shared_arith = "off";

arriav_lcell_comb \op_1~145 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!freq_mod_i_11),
	.datae(gnd),
	.dataf(!phi_inc_i_11),
	.datag(gnd),
	.cin(\op_1~150 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~145_sumout ),
	.cout(\op_1~146 ),
	.shareout());
defparam \op_1~145 .extended_lut = "off";
defparam \op_1~145 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~145 .shared_arith = "off";

arriav_lcell_comb \op_1~141 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!freq_mod_i_12),
	.datae(gnd),
	.dataf(!phi_inc_i_12),
	.datag(gnd),
	.cin(\op_1~146 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~141_sumout ),
	.cout(\op_1~142 ),
	.shareout());
defparam \op_1~141 .extended_lut = "off";
defparam \op_1~141 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~141 .shared_arith = "off";

arriav_lcell_comb \op_1~137 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!freq_mod_i_13),
	.datae(gnd),
	.dataf(!phi_inc_i_13),
	.datag(gnd),
	.cin(\op_1~142 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~137_sumout ),
	.cout(\op_1~138 ),
	.shareout());
defparam \op_1~137 .extended_lut = "off";
defparam \op_1~137 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~137 .shared_arith = "off";

arriav_lcell_comb \op_1~133 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!freq_mod_i_14),
	.datae(gnd),
	.dataf(!phi_inc_i_14),
	.datag(gnd),
	.cin(\op_1~138 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~133_sumout ),
	.cout(\op_1~134 ),
	.shareout());
defparam \op_1~133 .extended_lut = "off";
defparam \op_1~133 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~133 .shared_arith = "off";

arriav_lcell_comb \op_1~129 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!freq_mod_i_15),
	.datae(gnd),
	.dataf(!phi_inc_i_15),
	.datag(gnd),
	.cin(\op_1~134 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~129_sumout ),
	.cout(\op_1~130 ),
	.shareout());
defparam \op_1~129 .extended_lut = "off";
defparam \op_1~129 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~129 .shared_arith = "off";

arriav_lcell_comb \op_1~125 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!freq_mod_i_16),
	.datae(gnd),
	.dataf(!phi_inc_i_16),
	.datag(gnd),
	.cin(\op_1~130 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~125_sumout ),
	.cout(\op_1~126 ),
	.shareout());
defparam \op_1~125 .extended_lut = "off";
defparam \op_1~125 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~125 .shared_arith = "off";

arriav_lcell_comb \op_1~121 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!freq_mod_i_17),
	.datae(gnd),
	.dataf(!phi_inc_i_17),
	.datag(gnd),
	.cin(\op_1~126 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~121_sumout ),
	.cout(\op_1~122 ),
	.shareout());
defparam \op_1~121 .extended_lut = "off";
defparam \op_1~121 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~121 .shared_arith = "off";

arriav_lcell_comb \op_1~117 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!freq_mod_i_18),
	.datae(gnd),
	.dataf(!phi_inc_i_18),
	.datag(gnd),
	.cin(\op_1~122 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~117_sumout ),
	.cout(\op_1~118 ),
	.shareout());
defparam \op_1~117 .extended_lut = "off";
defparam \op_1~117 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~117 .shared_arith = "off";

arriav_lcell_comb \op_1~113 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!freq_mod_i_19),
	.datae(gnd),
	.dataf(!phi_inc_i_19),
	.datag(gnd),
	.cin(\op_1~118 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~113_sumout ),
	.cout(\op_1~114 ),
	.shareout());
defparam \op_1~113 .extended_lut = "off";
defparam \op_1~113 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~113 .shared_arith = "off";

arriav_lcell_comb \op_1~109 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!freq_mod_i_20),
	.datae(gnd),
	.dataf(!phi_inc_i_20),
	.datag(gnd),
	.cin(\op_1~114 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~109_sumout ),
	.cout(\op_1~110 ),
	.shareout());
defparam \op_1~109 .extended_lut = "off";
defparam \op_1~109 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~109 .shared_arith = "off";

arriav_lcell_comb \op_1~105 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!freq_mod_i_21),
	.datae(gnd),
	.dataf(!phi_inc_i_21),
	.datag(gnd),
	.cin(\op_1~110 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~105_sumout ),
	.cout(\op_1~106 ),
	.shareout());
defparam \op_1~105 .extended_lut = "off";
defparam \op_1~105 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~105 .shared_arith = "off";

arriav_lcell_comb \op_1~101 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!freq_mod_i_22),
	.datae(gnd),
	.dataf(!phi_inc_i_22),
	.datag(gnd),
	.cin(\op_1~106 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~101_sumout ),
	.cout(\op_1~102 ),
	.shareout());
defparam \op_1~101 .extended_lut = "off";
defparam \op_1~101 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~101 .shared_arith = "off";

arriav_lcell_comb \op_1~97 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!freq_mod_i_23),
	.datae(gnd),
	.dataf(!phi_inc_i_23),
	.datag(gnd),
	.cin(\op_1~102 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~97_sumout ),
	.cout(\op_1~98 ),
	.shareout());
defparam \op_1~97 .extended_lut = "off";
defparam \op_1~97 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~97 .shared_arith = "off";

arriav_lcell_comb \op_1~93 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!freq_mod_i_24),
	.datae(gnd),
	.dataf(!phi_inc_i_24),
	.datag(gnd),
	.cin(\op_1~98 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~93_sumout ),
	.cout(\op_1~94 ),
	.shareout());
defparam \op_1~93 .extended_lut = "off";
defparam \op_1~93 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~93 .shared_arith = "off";

arriav_lcell_comb \op_1~89 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!freq_mod_i_25),
	.datae(gnd),
	.dataf(!phi_inc_i_25),
	.datag(gnd),
	.cin(\op_1~94 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~89_sumout ),
	.cout(\op_1~90 ),
	.shareout());
defparam \op_1~89 .extended_lut = "off";
defparam \op_1~89 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~89 .shared_arith = "off";

arriav_lcell_comb \op_1~85 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!freq_mod_i_26),
	.datae(gnd),
	.dataf(!phi_inc_i_26),
	.datag(gnd),
	.cin(\op_1~90 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~85_sumout ),
	.cout(\op_1~86 ),
	.shareout());
defparam \op_1~85 .extended_lut = "off";
defparam \op_1~85 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~85 .shared_arith = "off";

arriav_lcell_comb \op_1~81 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!freq_mod_i_27),
	.datae(gnd),
	.dataf(!phi_inc_i_27),
	.datag(gnd),
	.cin(\op_1~86 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~81_sumout ),
	.cout(\op_1~82 ),
	.shareout());
defparam \op_1~81 .extended_lut = "off";
defparam \op_1~81 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~81 .shared_arith = "off";

arriav_lcell_comb \op_1~77 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!freq_mod_i_28),
	.datae(gnd),
	.dataf(!phi_inc_i_28),
	.datag(gnd),
	.cin(\op_1~82 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~77_sumout ),
	.cout(\op_1~78 ),
	.shareout());
defparam \op_1~77 .extended_lut = "off";
defparam \op_1~77 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~77 .shared_arith = "off";

arriav_lcell_comb \op_1~73 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!freq_mod_i_29),
	.datae(gnd),
	.dataf(!phi_inc_i_29),
	.datag(gnd),
	.cin(\op_1~78 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~73_sumout ),
	.cout(\op_1~74 ),
	.shareout());
defparam \op_1~73 .extended_lut = "off";
defparam \op_1~73 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~73 .shared_arith = "off";

arriav_lcell_comb \op_1~69 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!freq_mod_i_30),
	.datae(gnd),
	.dataf(!phi_inc_i_30),
	.datag(gnd),
	.cin(\op_1~74 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~69_sumout ),
	.cout(\op_1~70 ),
	.shareout());
defparam \op_1~69 .extended_lut = "off";
defparam \op_1~69 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~69 .shared_arith = "off";

arriav_lcell_comb \op_1~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!freq_mod_i_31),
	.datae(gnd),
	.dataf(!phi_inc_i_31),
	.datag(gnd),
	.cin(\op_1~70 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~57_sumout ),
	.cout(\op_1~58 ),
	.shareout());
defparam \op_1~57 .extended_lut = "off";
defparam \op_1~57 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~57 .shared_arith = "off";

arriav_lcell_comb \op_1~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!freq_mod_i_31),
	.datae(gnd),
	.dataf(!phi_inc_i_32),
	.datag(gnd),
	.cin(\op_1~58 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~1_sumout ),
	.cout(\op_1~2 ),
	.shareout());
defparam \op_1~1 .extended_lut = "off";
defparam \op_1~1 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~1 .shared_arith = "off";

arriav_lcell_comb \op_1~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!freq_mod_i_31),
	.datae(gnd),
	.dataf(!phi_inc_i_33),
	.datag(gnd),
	.cin(\op_1~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~5_sumout ),
	.cout(\op_1~6 ),
	.shareout());
defparam \op_1~5 .extended_lut = "off";
defparam \op_1~5 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~5 .shared_arith = "off";

arriav_lcell_comb \op_1~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!freq_mod_i_31),
	.datae(gnd),
	.dataf(!phi_inc_i_34),
	.datag(gnd),
	.cin(\op_1~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~9_sumout ),
	.cout(\op_1~10 ),
	.shareout());
defparam \op_1~9 .extended_lut = "off";
defparam \op_1~9 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~9 .shared_arith = "off";

arriav_lcell_comb \op_1~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!freq_mod_i_31),
	.datae(gnd),
	.dataf(!phi_inc_i_35),
	.datag(gnd),
	.cin(\op_1~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~13_sumout ),
	.cout(\op_1~14 ),
	.shareout());
defparam \op_1~13 .extended_lut = "off";
defparam \op_1~13 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~13 .shared_arith = "off";

arriav_lcell_comb \op_1~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!freq_mod_i_31),
	.datae(gnd),
	.dataf(!phi_inc_i_36),
	.datag(gnd),
	.cin(\op_1~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~17_sumout ),
	.cout(\op_1~18 ),
	.shareout());
defparam \op_1~17 .extended_lut = "off";
defparam \op_1~17 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~17 .shared_arith = "off";

arriav_lcell_comb \op_1~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!freq_mod_i_31),
	.datae(gnd),
	.dataf(!phi_inc_i_37),
	.datag(gnd),
	.cin(\op_1~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~21_sumout ),
	.cout(\op_1~22 ),
	.shareout());
defparam \op_1~21 .extended_lut = "off";
defparam \op_1~21 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~21 .shared_arith = "off";

arriav_lcell_comb \op_1~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!freq_mod_i_31),
	.datae(gnd),
	.dataf(!phi_inc_i_38),
	.datag(gnd),
	.cin(\op_1~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~25_sumout ),
	.cout(\op_1~26 ),
	.shareout());
defparam \op_1~25 .extended_lut = "off";
defparam \op_1~25 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~25 .shared_arith = "off";

arriav_lcell_comb \op_1~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!freq_mod_i_31),
	.datae(gnd),
	.dataf(!phi_inc_i_39),
	.datag(gnd),
	.cin(\op_1~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~29_sumout ),
	.cout(\op_1~30 ),
	.shareout());
defparam \op_1~29 .extended_lut = "off";
defparam \op_1~29 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~29 .shared_arith = "off";

arriav_lcell_comb \op_1~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!freq_mod_i_31),
	.datae(gnd),
	.dataf(!phi_inc_i_40),
	.datag(gnd),
	.cin(\op_1~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~33_sumout ),
	.cout(\op_1~34 ),
	.shareout());
defparam \op_1~33 .extended_lut = "off";
defparam \op_1~33 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~33 .shared_arith = "off";

arriav_lcell_comb \op_1~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!freq_mod_i_31),
	.datae(gnd),
	.dataf(!phi_inc_i_41),
	.datag(gnd),
	.cin(\op_1~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~37_sumout ),
	.cout(\op_1~38 ),
	.shareout());
defparam \op_1~37 .extended_lut = "off";
defparam \op_1~37 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~37 .shared_arith = "off";

arriav_lcell_comb \op_1~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!freq_mod_i_31),
	.datae(gnd),
	.dataf(!phi_inc_i_42),
	.datag(gnd),
	.cin(\op_1~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~41_sumout ),
	.cout(\op_1~42 ),
	.shareout());
defparam \op_1~41 .extended_lut = "off";
defparam \op_1~41 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~41 .shared_arith = "off";

arriav_lcell_comb \op_1~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!freq_mod_i_31),
	.datae(gnd),
	.dataf(!phi_inc_i_43),
	.datag(gnd),
	.cin(\op_1~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~45_sumout ),
	.cout(\op_1~46 ),
	.shareout());
defparam \op_1~45 .extended_lut = "off";
defparam \op_1~45 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~45 .shared_arith = "off";

arriav_lcell_comb \op_1~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!freq_mod_i_31),
	.datae(gnd),
	.dataf(!phi_inc_i_44),
	.datag(gnd),
	.cin(\op_1~46 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~49_sumout ),
	.cout(\op_1~50 ),
	.shareout());
defparam \op_1~49 .extended_lut = "off";
defparam \op_1~49 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~49 .shared_arith = "off";

arriav_lcell_comb \op_1~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!freq_mod_i_31),
	.datae(gnd),
	.dataf(!phi_inc_i_45),
	.datag(gnd),
	.cin(\op_1~50 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~61_sumout ),
	.cout(\op_1~62 ),
	.shareout());
defparam \op_1~61 .extended_lut = "off";
defparam \op_1~61 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~61 .shared_arith = "off";

arriav_lcell_comb \op_1~65 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!freq_mod_i_31),
	.datae(gnd),
	.dataf(!phi_inc_i_46),
	.datag(gnd),
	.cin(\op_1~62 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~65_sumout ),
	.cout(\op_1~66 ),
	.shareout());
defparam \op_1~65 .extended_lut = "off";
defparam \op_1~65 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~65 .shared_arith = "off";

arriav_lcell_comb \op_1~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!freq_mod_i_31),
	.datae(gnd),
	.dataf(!phi_inc_i_47),
	.datag(gnd),
	.cin(\op_1~66 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~53_sumout ),
	.cout(),
	.shareout());
defparam \op_1~53 .extended_lut = "off";
defparam \op_1~53 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~53 .shared_arith = "off";

endmodule

module DDS_48_v1_asj_nco_isdr (
	data_ready1,
	clk,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
output 	data_ready1;
input 	clk;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \lpm_counter_component|auto_generated|counter_reg_bit[3]~q ;
wire \lpm_counter_component|auto_generated|counter_reg_bit[2]~q ;
wire \lpm_counter_component|auto_generated|counter_reg_bit[1]~q ;
wire \lpm_counter_component|auto_generated|counter_reg_bit[0]~q ;
wire \data_ready~0_combout ;


DDS_48_v1_lpm_counter_1 lpm_counter_component(
	.counter_reg_bit_3(\lpm_counter_component|auto_generated|counter_reg_bit[3]~q ),
	.counter_reg_bit_2(\lpm_counter_component|auto_generated|counter_reg_bit[2]~q ),
	.counter_reg_bit_1(\lpm_counter_component|auto_generated|counter_reg_bit[1]~q ),
	.counter_reg_bit_0(\lpm_counter_component|auto_generated|counter_reg_bit[0]~q ),
	.clock(clk),
	.sclr(reset_n),
	.clken(clken));

dffeas data_ready(
	.clk(clk),
	.d(\data_ready~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(vcc),
	.q(data_ready1),
	.prn(vcc));
defparam data_ready.is_wysiwyg = "true";
defparam data_ready.power_up = "low";

arriav_lcell_comb \data_ready~0 (
	.dataa(!data_ready1),
	.datab(!clken),
	.datac(!\lpm_counter_component|auto_generated|counter_reg_bit[3]~q ),
	.datad(!\lpm_counter_component|auto_generated|counter_reg_bit[2]~q ),
	.datae(!\lpm_counter_component|auto_generated|counter_reg_bit[1]~q ),
	.dataf(!\lpm_counter_component|auto_generated|counter_reg_bit[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_ready~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_ready~0 .extended_lut = "off";
defparam \data_ready~0 .lut_mask = 64'hFFFFFFFFFFFFFF7F;
defparam \data_ready~0 .shared_arith = "off";

endmodule

module DDS_48_v1_lpm_counter_1 (
	counter_reg_bit_3,
	counter_reg_bit_2,
	counter_reg_bit_1,
	counter_reg_bit_0,
	clock,
	sclr,
	clken)/* synthesis synthesis_greybox=1 */;
output 	counter_reg_bit_3;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
output 	counter_reg_bit_0;
input 	clock;
input 	sclr;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



DDS_48_v1_cntr_udi auto_generated(
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_1(counter_reg_bit_1),
	.counter_reg_bit_0(counter_reg_bit_0),
	.clock(clock),
	.sclr(sclr),
	.clken(clken));

endmodule

module DDS_48_v1_cntr_udi (
	counter_reg_bit_3,
	counter_reg_bit_2,
	counter_reg_bit_1,
	counter_reg_bit_0,
	clock,
	sclr,
	clken)/* synthesis synthesis_greybox=1 */;
output 	counter_reg_bit_3;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
output 	counter_reg_bit_0;
input 	clock;
input 	sclr;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~sumout ;
wire \counter_comb_bita2~sumout ;
wire \counter_comb_bita1~sumout ;
wire \counter_comb_bita0~sumout ;


dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!sclr),
	.sload(gnd),
	.ena(clken),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!sclr),
	.sload(gnd),
	.ena(clken),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!sclr),
	.sload(gnd),
	.ena(clken),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!sclr),
	.sload(gnd),
	.ena(clken),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

arriav_lcell_comb counter_comb_bita0(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita0~sumout ),
	.cout(\counter_comb_bita0~COUT ),
	.shareout());
defparam counter_comb_bita0.extended_lut = "off";
defparam counter_comb_bita0.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita0.shared_arith = "off";

arriav_lcell_comb counter_comb_bita1(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita0~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita1~sumout ),
	.cout(\counter_comb_bita1~COUT ),
	.shareout());
defparam counter_comb_bita1.extended_lut = "off";
defparam counter_comb_bita1.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita1.shared_arith = "off";

arriav_lcell_comb counter_comb_bita2(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita1~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita2~sumout ),
	.cout(\counter_comb_bita2~COUT ),
	.shareout());
defparam counter_comb_bita2.extended_lut = "off";
defparam counter_comb_bita2.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita2.shared_arith = "off";

arriav_lcell_comb counter_comb_bita3(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita2~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita3~sumout ),
	.cout(),
	.shareout());
defparam counter_comb_bita3.extended_lut = "off";
defparam counter_comb_bita3.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita3.shared_arith = "off";

endmodule

module DDS_48_v1_asj_nco_mob_rw (
	data_out_0,
	data_out_1,
	data_out_2,
	data_out_3,
	data_out_4,
	data_out_5,
	data_out_6,
	data_out_7,
	data_out_8,
	data_out_9,
	data_out_10,
	data_out_11,
	data_out_12,
	data_out_13,
	data_out_14,
	data_out_15,
	ram_block1a64,
	ram_block1a80,
	ram_block1a96,
	ram_block1a112,
	ram_block1a32,
	ram_block1a48,
	ram_block1a0,
	ram_block1a16,
	ram_block1a65,
	ram_block1a81,
	ram_block1a97,
	ram_block1a113,
	ram_block1a33,
	ram_block1a49,
	ram_block1a1,
	ram_block1a17,
	ram_block1a66,
	ram_block1a82,
	ram_block1a98,
	ram_block1a114,
	ram_block1a34,
	ram_block1a50,
	ram_block1a2,
	ram_block1a18,
	ram_block1a67,
	ram_block1a83,
	ram_block1a99,
	ram_block1a115,
	ram_block1a35,
	ram_block1a51,
	ram_block1a3,
	ram_block1a19,
	ram_block1a68,
	ram_block1a84,
	ram_block1a100,
	ram_block1a116,
	ram_block1a36,
	ram_block1a52,
	ram_block1a4,
	ram_block1a20,
	ram_block1a69,
	ram_block1a85,
	ram_block1a101,
	ram_block1a117,
	ram_block1a37,
	ram_block1a53,
	ram_block1a5,
	ram_block1a21,
	ram_block1a70,
	ram_block1a86,
	ram_block1a102,
	ram_block1a118,
	ram_block1a38,
	ram_block1a54,
	ram_block1a6,
	ram_block1a22,
	ram_block1a71,
	ram_block1a87,
	ram_block1a103,
	ram_block1a119,
	ram_block1a39,
	ram_block1a55,
	ram_block1a7,
	ram_block1a23,
	ram_block1a72,
	ram_block1a88,
	ram_block1a104,
	ram_block1a120,
	ram_block1a40,
	ram_block1a56,
	ram_block1a8,
	ram_block1a24,
	ram_block1a73,
	ram_block1a89,
	ram_block1a105,
	ram_block1a121,
	ram_block1a41,
	ram_block1a57,
	ram_block1a9,
	ram_block1a25,
	ram_block1a74,
	ram_block1a90,
	ram_block1a106,
	ram_block1a122,
	ram_block1a42,
	ram_block1a58,
	ram_block1a10,
	ram_block1a26,
	ram_block1a75,
	ram_block1a91,
	ram_block1a107,
	ram_block1a123,
	ram_block1a43,
	ram_block1a59,
	ram_block1a11,
	ram_block1a27,
	ram_block1a76,
	ram_block1a92,
	ram_block1a108,
	ram_block1a124,
	ram_block1a44,
	ram_block1a60,
	ram_block1a12,
	ram_block1a28,
	ram_block1a77,
	ram_block1a93,
	ram_block1a109,
	ram_block1a125,
	ram_block1a45,
	ram_block1a61,
	ram_block1a13,
	ram_block1a29,
	ram_block1a78,
	ram_block1a94,
	ram_block1a110,
	ram_block1a126,
	ram_block1a46,
	ram_block1a62,
	ram_block1a14,
	ram_block1a30,
	ram_block1a79,
	ram_block1a95,
	ram_block1a111,
	ram_block1a127,
	ram_block1a47,
	ram_block1a63,
	ram_block1a15,
	ram_block1a31,
	out_address_reg_a_2,
	out_address_reg_a_0,
	out_address_reg_a_1,
	data_out_121,
	clk,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
output 	data_out_0;
output 	data_out_1;
output 	data_out_2;
output 	data_out_3;
output 	data_out_4;
output 	data_out_5;
output 	data_out_6;
output 	data_out_7;
output 	data_out_8;
output 	data_out_9;
output 	data_out_10;
output 	data_out_11;
output 	data_out_12;
output 	data_out_13;
output 	data_out_14;
output 	data_out_15;
input 	ram_block1a64;
input 	ram_block1a80;
input 	ram_block1a96;
input 	ram_block1a112;
input 	ram_block1a32;
input 	ram_block1a48;
input 	ram_block1a0;
input 	ram_block1a16;
input 	ram_block1a65;
input 	ram_block1a81;
input 	ram_block1a97;
input 	ram_block1a113;
input 	ram_block1a33;
input 	ram_block1a49;
input 	ram_block1a1;
input 	ram_block1a17;
input 	ram_block1a66;
input 	ram_block1a82;
input 	ram_block1a98;
input 	ram_block1a114;
input 	ram_block1a34;
input 	ram_block1a50;
input 	ram_block1a2;
input 	ram_block1a18;
input 	ram_block1a67;
input 	ram_block1a83;
input 	ram_block1a99;
input 	ram_block1a115;
input 	ram_block1a35;
input 	ram_block1a51;
input 	ram_block1a3;
input 	ram_block1a19;
input 	ram_block1a68;
input 	ram_block1a84;
input 	ram_block1a100;
input 	ram_block1a116;
input 	ram_block1a36;
input 	ram_block1a52;
input 	ram_block1a4;
input 	ram_block1a20;
input 	ram_block1a69;
input 	ram_block1a85;
input 	ram_block1a101;
input 	ram_block1a117;
input 	ram_block1a37;
input 	ram_block1a53;
input 	ram_block1a5;
input 	ram_block1a21;
input 	ram_block1a70;
input 	ram_block1a86;
input 	ram_block1a102;
input 	ram_block1a118;
input 	ram_block1a38;
input 	ram_block1a54;
input 	ram_block1a6;
input 	ram_block1a22;
input 	ram_block1a71;
input 	ram_block1a87;
input 	ram_block1a103;
input 	ram_block1a119;
input 	ram_block1a39;
input 	ram_block1a55;
input 	ram_block1a7;
input 	ram_block1a23;
input 	ram_block1a72;
input 	ram_block1a88;
input 	ram_block1a104;
input 	ram_block1a120;
input 	ram_block1a40;
input 	ram_block1a56;
input 	ram_block1a8;
input 	ram_block1a24;
input 	ram_block1a73;
input 	ram_block1a89;
input 	ram_block1a105;
input 	ram_block1a121;
input 	ram_block1a41;
input 	ram_block1a57;
input 	ram_block1a9;
input 	ram_block1a25;
input 	ram_block1a74;
input 	ram_block1a90;
input 	ram_block1a106;
input 	ram_block1a122;
input 	ram_block1a42;
input 	ram_block1a58;
input 	ram_block1a10;
input 	ram_block1a26;
input 	ram_block1a75;
input 	ram_block1a91;
input 	ram_block1a107;
input 	ram_block1a123;
input 	ram_block1a43;
input 	ram_block1a59;
input 	ram_block1a11;
input 	ram_block1a27;
input 	ram_block1a76;
input 	ram_block1a92;
input 	ram_block1a108;
input 	ram_block1a124;
input 	ram_block1a44;
input 	ram_block1a60;
input 	ram_block1a12;
input 	ram_block1a28;
input 	ram_block1a77;
input 	ram_block1a93;
input 	ram_block1a109;
input 	ram_block1a125;
input 	ram_block1a45;
input 	ram_block1a61;
input 	ram_block1a13;
input 	ram_block1a29;
input 	ram_block1a78;
input 	ram_block1a94;
input 	ram_block1a110;
input 	ram_block1a126;
input 	ram_block1a46;
input 	ram_block1a62;
input 	ram_block1a14;
input 	ram_block1a30;
input 	ram_block1a79;
input 	ram_block1a95;
input 	ram_block1a111;
input 	ram_block1a127;
input 	ram_block1a47;
input 	ram_block1a63;
input 	ram_block1a15;
input 	ram_block1a31;
input 	out_address_reg_a_2;
input 	out_address_reg_a_0;
input 	out_address_reg_a_1;
output 	data_out_121;
input 	clk;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \data_out~0_combout ;
wire \data_out~1_combout ;
wire \data_out~2_combout ;
wire \data_out~4_combout ;
wire \data_out~5_combout ;
wire \data_out~6_combout ;
wire \data_out~7_combout ;
wire \data_out~8_combout ;
wire \data_out~9_combout ;
wire \data_out~10_combout ;
wire \data_out~11_combout ;
wire \data_out~12_combout ;
wire \data_out~13_combout ;
wire \data_out~14_combout ;
wire \data_out~15_combout ;
wire \data_out~16_combout ;
wire \data_out~17_combout ;
wire \data_out~18_combout ;
wire \data_out~19_combout ;
wire \data_out~20_combout ;
wire \data_out~21_combout ;
wire \data_out~22_combout ;
wire \data_out~23_combout ;
wire \data_out~24_combout ;
wire \data_out~25_combout ;
wire \data_out~26_combout ;
wire \data_out~27_combout ;
wire \data_out~28_combout ;
wire \data_out~29_combout ;
wire \data_out~30_combout ;
wire \data_out~31_combout ;
wire \data_out~32_combout ;
wire \data_out~33_combout ;
wire \data_out~34_combout ;
wire \data_out~35_combout ;
wire \data_out~36_combout ;
wire \data_out~37_combout ;
wire \data_out~38_combout ;
wire \data_out~39_combout ;
wire \data_out~40_combout ;
wire \data_out~41_combout ;
wire \data_out~42_combout ;
wire \data_out~43_combout ;
wire \data_out~44_combout ;
wire \data_out~45_combout ;
wire \data_out~46_combout ;
wire \data_out~47_combout ;
wire \data_out~48_combout ;


dffeas \data_out[0] (
	.clk(clk),
	.d(\data_out~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_121),
	.q(data_out_0),
	.prn(vcc));
defparam \data_out[0] .is_wysiwyg = "true";
defparam \data_out[0] .power_up = "low";

dffeas \data_out[1] (
	.clk(clk),
	.d(\data_out~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_121),
	.q(data_out_1),
	.prn(vcc));
defparam \data_out[1] .is_wysiwyg = "true";
defparam \data_out[1] .power_up = "low";

dffeas \data_out[2] (
	.clk(clk),
	.d(\data_out~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_121),
	.q(data_out_2),
	.prn(vcc));
defparam \data_out[2] .is_wysiwyg = "true";
defparam \data_out[2] .power_up = "low";

dffeas \data_out[3] (
	.clk(clk),
	.d(\data_out~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_121),
	.q(data_out_3),
	.prn(vcc));
defparam \data_out[3] .is_wysiwyg = "true";
defparam \data_out[3] .power_up = "low";

dffeas \data_out[4] (
	.clk(clk),
	.d(\data_out~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_121),
	.q(data_out_4),
	.prn(vcc));
defparam \data_out[4] .is_wysiwyg = "true";
defparam \data_out[4] .power_up = "low";

dffeas \data_out[5] (
	.clk(clk),
	.d(\data_out~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_121),
	.q(data_out_5),
	.prn(vcc));
defparam \data_out[5] .is_wysiwyg = "true";
defparam \data_out[5] .power_up = "low";

dffeas \data_out[6] (
	.clk(clk),
	.d(\data_out~21_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_121),
	.q(data_out_6),
	.prn(vcc));
defparam \data_out[6] .is_wysiwyg = "true";
defparam \data_out[6] .power_up = "low";

dffeas \data_out[7] (
	.clk(clk),
	.d(\data_out~24_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_121),
	.q(data_out_7),
	.prn(vcc));
defparam \data_out[7] .is_wysiwyg = "true";
defparam \data_out[7] .power_up = "low";

dffeas \data_out[8] (
	.clk(clk),
	.d(\data_out~27_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_121),
	.q(data_out_8),
	.prn(vcc));
defparam \data_out[8] .is_wysiwyg = "true";
defparam \data_out[8] .power_up = "low";

dffeas \data_out[9] (
	.clk(clk),
	.d(\data_out~30_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_121),
	.q(data_out_9),
	.prn(vcc));
defparam \data_out[9] .is_wysiwyg = "true";
defparam \data_out[9] .power_up = "low";

dffeas \data_out[10] (
	.clk(clk),
	.d(\data_out~33_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_121),
	.q(data_out_10),
	.prn(vcc));
defparam \data_out[10] .is_wysiwyg = "true";
defparam \data_out[10] .power_up = "low";

dffeas \data_out[11] (
	.clk(clk),
	.d(\data_out~36_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_121),
	.q(data_out_11),
	.prn(vcc));
defparam \data_out[11] .is_wysiwyg = "true";
defparam \data_out[11] .power_up = "low";

dffeas \data_out[12] (
	.clk(clk),
	.d(\data_out~39_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_121),
	.q(data_out_12),
	.prn(vcc));
defparam \data_out[12] .is_wysiwyg = "true";
defparam \data_out[12] .power_up = "low";

dffeas \data_out[13] (
	.clk(clk),
	.d(\data_out~42_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_121),
	.q(data_out_13),
	.prn(vcc));
defparam \data_out[13] .is_wysiwyg = "true";
defparam \data_out[13] .power_up = "low";

dffeas \data_out[14] (
	.clk(clk),
	.d(\data_out~45_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_121),
	.q(data_out_14),
	.prn(vcc));
defparam \data_out[14] .is_wysiwyg = "true";
defparam \data_out[14] .power_up = "low";

dffeas \data_out[15] (
	.clk(clk),
	.d(\data_out~48_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_121),
	.q(data_out_15),
	.prn(vcc));
defparam \data_out[15] .is_wysiwyg = "true";
defparam \data_out[15] .power_up = "low";

arriav_lcell_comb \data_out[12]~3 (
	.dataa(!reset_n),
	.datab(!clken),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(data_out_121),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out[12]~3 .extended_lut = "off";
defparam \data_out[12]~3 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \data_out[12]~3 .shared_arith = "off";

arriav_lcell_comb \data_out~0 (
	.dataa(!ram_block1a64),
	.datab(!ram_block1a80),
	.datac(!ram_block1a96),
	.datad(!ram_block1a112),
	.datae(!out_address_reg_a_0),
	.dataf(!out_address_reg_a_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~0 .extended_lut = "off";
defparam \data_out~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \data_out~0 .shared_arith = "off";

arriav_lcell_comb \data_out~1 (
	.dataa(!out_address_reg_a_0),
	.datab(!out_address_reg_a_1),
	.datac(!ram_block1a32),
	.datad(!ram_block1a48),
	.datae(!ram_block1a0),
	.dataf(!ram_block1a16),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~1 .extended_lut = "off";
defparam \data_out~1 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \data_out~1 .shared_arith = "off";

arriav_lcell_comb \data_out~2 (
	.dataa(!out_address_reg_a_2),
	.datab(!\data_out~0_combout ),
	.datac(!\data_out~1_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~2 .extended_lut = "off";
defparam \data_out~2 .lut_mask = 64'h2727272727272727;
defparam \data_out~2 .shared_arith = "off";

arriav_lcell_comb \data_out~4 (
	.dataa(!ram_block1a65),
	.datab(!ram_block1a81),
	.datac(!ram_block1a97),
	.datad(!ram_block1a113),
	.datae(!out_address_reg_a_0),
	.dataf(!out_address_reg_a_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~4 .extended_lut = "off";
defparam \data_out~4 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \data_out~4 .shared_arith = "off";

arriav_lcell_comb \data_out~5 (
	.dataa(!out_address_reg_a_0),
	.datab(!out_address_reg_a_1),
	.datac(!ram_block1a33),
	.datad(!ram_block1a49),
	.datae(!ram_block1a1),
	.dataf(!ram_block1a17),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~5 .extended_lut = "off";
defparam \data_out~5 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \data_out~5 .shared_arith = "off";

arriav_lcell_comb \data_out~6 (
	.dataa(!out_address_reg_a_2),
	.datab(!\data_out~4_combout ),
	.datac(!\data_out~5_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~6 .extended_lut = "off";
defparam \data_out~6 .lut_mask = 64'h2727272727272727;
defparam \data_out~6 .shared_arith = "off";

arriav_lcell_comb \data_out~7 (
	.dataa(!ram_block1a66),
	.datab(!ram_block1a82),
	.datac(!ram_block1a98),
	.datad(!ram_block1a114),
	.datae(!out_address_reg_a_0),
	.dataf(!out_address_reg_a_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~7 .extended_lut = "off";
defparam \data_out~7 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \data_out~7 .shared_arith = "off";

arriav_lcell_comb \data_out~8 (
	.dataa(!out_address_reg_a_0),
	.datab(!out_address_reg_a_1),
	.datac(!ram_block1a34),
	.datad(!ram_block1a50),
	.datae(!ram_block1a2),
	.dataf(!ram_block1a18),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~8 .extended_lut = "off";
defparam \data_out~8 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \data_out~8 .shared_arith = "off";

arriav_lcell_comb \data_out~9 (
	.dataa(!out_address_reg_a_2),
	.datab(!\data_out~7_combout ),
	.datac(!\data_out~8_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~9 .extended_lut = "off";
defparam \data_out~9 .lut_mask = 64'h2727272727272727;
defparam \data_out~9 .shared_arith = "off";

arriav_lcell_comb \data_out~10 (
	.dataa(!ram_block1a67),
	.datab(!ram_block1a83),
	.datac(!ram_block1a99),
	.datad(!ram_block1a115),
	.datae(!out_address_reg_a_0),
	.dataf(!out_address_reg_a_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~10 .extended_lut = "off";
defparam \data_out~10 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \data_out~10 .shared_arith = "off";

arriav_lcell_comb \data_out~11 (
	.dataa(!out_address_reg_a_0),
	.datab(!out_address_reg_a_1),
	.datac(!ram_block1a35),
	.datad(!ram_block1a51),
	.datae(!ram_block1a3),
	.dataf(!ram_block1a19),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~11 .extended_lut = "off";
defparam \data_out~11 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \data_out~11 .shared_arith = "off";

arriav_lcell_comb \data_out~12 (
	.dataa(!out_address_reg_a_2),
	.datab(!\data_out~10_combout ),
	.datac(!\data_out~11_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~12 .extended_lut = "off";
defparam \data_out~12 .lut_mask = 64'h2727272727272727;
defparam \data_out~12 .shared_arith = "off";

arriav_lcell_comb \data_out~13 (
	.dataa(!ram_block1a68),
	.datab(!ram_block1a84),
	.datac(!ram_block1a100),
	.datad(!ram_block1a116),
	.datae(!out_address_reg_a_0),
	.dataf(!out_address_reg_a_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~13 .extended_lut = "off";
defparam \data_out~13 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \data_out~13 .shared_arith = "off";

arriav_lcell_comb \data_out~14 (
	.dataa(!out_address_reg_a_0),
	.datab(!out_address_reg_a_1),
	.datac(!ram_block1a36),
	.datad(!ram_block1a52),
	.datae(!ram_block1a4),
	.dataf(!ram_block1a20),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~14 .extended_lut = "off";
defparam \data_out~14 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \data_out~14 .shared_arith = "off";

arriav_lcell_comb \data_out~15 (
	.dataa(!out_address_reg_a_2),
	.datab(!\data_out~13_combout ),
	.datac(!\data_out~14_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~15 .extended_lut = "off";
defparam \data_out~15 .lut_mask = 64'h2727272727272727;
defparam \data_out~15 .shared_arith = "off";

arriav_lcell_comb \data_out~16 (
	.dataa(!ram_block1a69),
	.datab(!ram_block1a85),
	.datac(!ram_block1a101),
	.datad(!ram_block1a117),
	.datae(!out_address_reg_a_0),
	.dataf(!out_address_reg_a_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~16 .extended_lut = "off";
defparam \data_out~16 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \data_out~16 .shared_arith = "off";

arriav_lcell_comb \data_out~17 (
	.dataa(!out_address_reg_a_0),
	.datab(!out_address_reg_a_1),
	.datac(!ram_block1a37),
	.datad(!ram_block1a53),
	.datae(!ram_block1a5),
	.dataf(!ram_block1a21),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~17 .extended_lut = "off";
defparam \data_out~17 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \data_out~17 .shared_arith = "off";

arriav_lcell_comb \data_out~18 (
	.dataa(!out_address_reg_a_2),
	.datab(!\data_out~16_combout ),
	.datac(!\data_out~17_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~18 .extended_lut = "off";
defparam \data_out~18 .lut_mask = 64'h2727272727272727;
defparam \data_out~18 .shared_arith = "off";

arriav_lcell_comb \data_out~19 (
	.dataa(!ram_block1a70),
	.datab(!ram_block1a86),
	.datac(!ram_block1a102),
	.datad(!ram_block1a118),
	.datae(!out_address_reg_a_0),
	.dataf(!out_address_reg_a_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~19 .extended_lut = "off";
defparam \data_out~19 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \data_out~19 .shared_arith = "off";

arriav_lcell_comb \data_out~20 (
	.dataa(!out_address_reg_a_0),
	.datab(!out_address_reg_a_1),
	.datac(!ram_block1a38),
	.datad(!ram_block1a54),
	.datae(!ram_block1a6),
	.dataf(!ram_block1a22),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~20 .extended_lut = "off";
defparam \data_out~20 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \data_out~20 .shared_arith = "off";

arriav_lcell_comb \data_out~21 (
	.dataa(!out_address_reg_a_2),
	.datab(!\data_out~19_combout ),
	.datac(!\data_out~20_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~21_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~21 .extended_lut = "off";
defparam \data_out~21 .lut_mask = 64'h2727272727272727;
defparam \data_out~21 .shared_arith = "off";

arriav_lcell_comb \data_out~22 (
	.dataa(!ram_block1a71),
	.datab(!ram_block1a87),
	.datac(!ram_block1a103),
	.datad(!ram_block1a119),
	.datae(!out_address_reg_a_0),
	.dataf(!out_address_reg_a_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~22_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~22 .extended_lut = "off";
defparam \data_out~22 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \data_out~22 .shared_arith = "off";

arriav_lcell_comb \data_out~23 (
	.dataa(!out_address_reg_a_0),
	.datab(!out_address_reg_a_1),
	.datac(!ram_block1a39),
	.datad(!ram_block1a55),
	.datae(!ram_block1a7),
	.dataf(!ram_block1a23),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~23_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~23 .extended_lut = "off";
defparam \data_out~23 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \data_out~23 .shared_arith = "off";

arriav_lcell_comb \data_out~24 (
	.dataa(!out_address_reg_a_2),
	.datab(!\data_out~22_combout ),
	.datac(!\data_out~23_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~24_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~24 .extended_lut = "off";
defparam \data_out~24 .lut_mask = 64'h2727272727272727;
defparam \data_out~24 .shared_arith = "off";

arriav_lcell_comb \data_out~25 (
	.dataa(!ram_block1a72),
	.datab(!ram_block1a88),
	.datac(!ram_block1a104),
	.datad(!ram_block1a120),
	.datae(!out_address_reg_a_0),
	.dataf(!out_address_reg_a_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~25_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~25 .extended_lut = "off";
defparam \data_out~25 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \data_out~25 .shared_arith = "off";

arriav_lcell_comb \data_out~26 (
	.dataa(!out_address_reg_a_0),
	.datab(!out_address_reg_a_1),
	.datac(!ram_block1a40),
	.datad(!ram_block1a56),
	.datae(!ram_block1a8),
	.dataf(!ram_block1a24),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~26_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~26 .extended_lut = "off";
defparam \data_out~26 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \data_out~26 .shared_arith = "off";

arriav_lcell_comb \data_out~27 (
	.dataa(!out_address_reg_a_2),
	.datab(!\data_out~25_combout ),
	.datac(!\data_out~26_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~27_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~27 .extended_lut = "off";
defparam \data_out~27 .lut_mask = 64'h2727272727272727;
defparam \data_out~27 .shared_arith = "off";

arriav_lcell_comb \data_out~28 (
	.dataa(!ram_block1a73),
	.datab(!ram_block1a89),
	.datac(!ram_block1a105),
	.datad(!ram_block1a121),
	.datae(!out_address_reg_a_0),
	.dataf(!out_address_reg_a_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~28_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~28 .extended_lut = "off";
defparam \data_out~28 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \data_out~28 .shared_arith = "off";

arriav_lcell_comb \data_out~29 (
	.dataa(!out_address_reg_a_0),
	.datab(!out_address_reg_a_1),
	.datac(!ram_block1a41),
	.datad(!ram_block1a57),
	.datae(!ram_block1a9),
	.dataf(!ram_block1a25),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~29_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~29 .extended_lut = "off";
defparam \data_out~29 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \data_out~29 .shared_arith = "off";

arriav_lcell_comb \data_out~30 (
	.dataa(!out_address_reg_a_2),
	.datab(!\data_out~28_combout ),
	.datac(!\data_out~29_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~30_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~30 .extended_lut = "off";
defparam \data_out~30 .lut_mask = 64'h2727272727272727;
defparam \data_out~30 .shared_arith = "off";

arriav_lcell_comb \data_out~31 (
	.dataa(!ram_block1a74),
	.datab(!ram_block1a90),
	.datac(!ram_block1a106),
	.datad(!ram_block1a122),
	.datae(!out_address_reg_a_0),
	.dataf(!out_address_reg_a_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~31_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~31 .extended_lut = "off";
defparam \data_out~31 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \data_out~31 .shared_arith = "off";

arriav_lcell_comb \data_out~32 (
	.dataa(!out_address_reg_a_0),
	.datab(!out_address_reg_a_1),
	.datac(!ram_block1a42),
	.datad(!ram_block1a58),
	.datae(!ram_block1a10),
	.dataf(!ram_block1a26),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~32_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~32 .extended_lut = "off";
defparam \data_out~32 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \data_out~32 .shared_arith = "off";

arriav_lcell_comb \data_out~33 (
	.dataa(!out_address_reg_a_2),
	.datab(!\data_out~31_combout ),
	.datac(!\data_out~32_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~33_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~33 .extended_lut = "off";
defparam \data_out~33 .lut_mask = 64'h2727272727272727;
defparam \data_out~33 .shared_arith = "off";

arriav_lcell_comb \data_out~34 (
	.dataa(!ram_block1a75),
	.datab(!ram_block1a91),
	.datac(!ram_block1a107),
	.datad(!ram_block1a123),
	.datae(!out_address_reg_a_0),
	.dataf(!out_address_reg_a_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~34_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~34 .extended_lut = "off";
defparam \data_out~34 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \data_out~34 .shared_arith = "off";

arriav_lcell_comb \data_out~35 (
	.dataa(!out_address_reg_a_0),
	.datab(!out_address_reg_a_1),
	.datac(!ram_block1a43),
	.datad(!ram_block1a59),
	.datae(!ram_block1a11),
	.dataf(!ram_block1a27),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~35_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~35 .extended_lut = "off";
defparam \data_out~35 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \data_out~35 .shared_arith = "off";

arriav_lcell_comb \data_out~36 (
	.dataa(!out_address_reg_a_2),
	.datab(!\data_out~34_combout ),
	.datac(!\data_out~35_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~36_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~36 .extended_lut = "off";
defparam \data_out~36 .lut_mask = 64'h2727272727272727;
defparam \data_out~36 .shared_arith = "off";

arriav_lcell_comb \data_out~37 (
	.dataa(!ram_block1a76),
	.datab(!ram_block1a92),
	.datac(!ram_block1a108),
	.datad(!ram_block1a124),
	.datae(!out_address_reg_a_0),
	.dataf(!out_address_reg_a_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~37_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~37 .extended_lut = "off";
defparam \data_out~37 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \data_out~37 .shared_arith = "off";

arriav_lcell_comb \data_out~38 (
	.dataa(!out_address_reg_a_0),
	.datab(!out_address_reg_a_1),
	.datac(!ram_block1a44),
	.datad(!ram_block1a60),
	.datae(!ram_block1a12),
	.dataf(!ram_block1a28),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~38_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~38 .extended_lut = "off";
defparam \data_out~38 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \data_out~38 .shared_arith = "off";

arriav_lcell_comb \data_out~39 (
	.dataa(!out_address_reg_a_2),
	.datab(!\data_out~37_combout ),
	.datac(!\data_out~38_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~39_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~39 .extended_lut = "off";
defparam \data_out~39 .lut_mask = 64'h2727272727272727;
defparam \data_out~39 .shared_arith = "off";

arriav_lcell_comb \data_out~40 (
	.dataa(!ram_block1a77),
	.datab(!ram_block1a93),
	.datac(!ram_block1a109),
	.datad(!ram_block1a125),
	.datae(!out_address_reg_a_0),
	.dataf(!out_address_reg_a_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~40_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~40 .extended_lut = "off";
defparam \data_out~40 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \data_out~40 .shared_arith = "off";

arriav_lcell_comb \data_out~41 (
	.dataa(!out_address_reg_a_0),
	.datab(!out_address_reg_a_1),
	.datac(!ram_block1a45),
	.datad(!ram_block1a61),
	.datae(!ram_block1a13),
	.dataf(!ram_block1a29),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~41_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~41 .extended_lut = "off";
defparam \data_out~41 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \data_out~41 .shared_arith = "off";

arriav_lcell_comb \data_out~42 (
	.dataa(!out_address_reg_a_2),
	.datab(!\data_out~40_combout ),
	.datac(!\data_out~41_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~42_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~42 .extended_lut = "off";
defparam \data_out~42 .lut_mask = 64'h2727272727272727;
defparam \data_out~42 .shared_arith = "off";

arriav_lcell_comb \data_out~43 (
	.dataa(!ram_block1a78),
	.datab(!ram_block1a94),
	.datac(!ram_block1a110),
	.datad(!ram_block1a126),
	.datae(!out_address_reg_a_0),
	.dataf(!out_address_reg_a_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~43_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~43 .extended_lut = "off";
defparam \data_out~43 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \data_out~43 .shared_arith = "off";

arriav_lcell_comb \data_out~44 (
	.dataa(!out_address_reg_a_0),
	.datab(!out_address_reg_a_1),
	.datac(!ram_block1a46),
	.datad(!ram_block1a62),
	.datae(!ram_block1a14),
	.dataf(!ram_block1a30),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~44_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~44 .extended_lut = "off";
defparam \data_out~44 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \data_out~44 .shared_arith = "off";

arriav_lcell_comb \data_out~45 (
	.dataa(!out_address_reg_a_2),
	.datab(!\data_out~43_combout ),
	.datac(!\data_out~44_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~45_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~45 .extended_lut = "off";
defparam \data_out~45 .lut_mask = 64'h2727272727272727;
defparam \data_out~45 .shared_arith = "off";

arriav_lcell_comb \data_out~46 (
	.dataa(!ram_block1a79),
	.datab(!ram_block1a95),
	.datac(!ram_block1a111),
	.datad(!ram_block1a127),
	.datae(!out_address_reg_a_0),
	.dataf(!out_address_reg_a_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~46_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~46 .extended_lut = "off";
defparam \data_out~46 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \data_out~46 .shared_arith = "off";

arriav_lcell_comb \data_out~47 (
	.dataa(!out_address_reg_a_0),
	.datab(!out_address_reg_a_1),
	.datac(!ram_block1a47),
	.datad(!ram_block1a63),
	.datae(!ram_block1a15),
	.dataf(!ram_block1a31),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~47_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~47 .extended_lut = "off";
defparam \data_out~47 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \data_out~47 .shared_arith = "off";

arriav_lcell_comb \data_out~48 (
	.dataa(!out_address_reg_a_2),
	.datab(!\data_out~46_combout ),
	.datac(!\data_out~47_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~48_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~48 .extended_lut = "off";
defparam \data_out~48 .lut_mask = 64'h2727272727272727;
defparam \data_out~48 .shared_arith = "off";

endmodule

module DDS_48_v1_asj_nco_mob_rw_1 (
	data_out_0,
	data_out_1,
	data_out_2,
	data_out_3,
	data_out_4,
	data_out_5,
	data_out_6,
	data_out_7,
	data_out_8,
	data_out_9,
	data_out_10,
	data_out_11,
	data_out_12,
	data_out_13,
	data_out_14,
	data_out_15,
	ram_block1a64,
	ram_block1a80,
	ram_block1a96,
	ram_block1a112,
	ram_block1a32,
	ram_block1a48,
	ram_block1a0,
	ram_block1a16,
	ram_block1a65,
	ram_block1a81,
	ram_block1a97,
	ram_block1a113,
	ram_block1a33,
	ram_block1a49,
	ram_block1a1,
	ram_block1a17,
	ram_block1a66,
	ram_block1a82,
	ram_block1a98,
	ram_block1a114,
	ram_block1a34,
	ram_block1a50,
	ram_block1a2,
	ram_block1a18,
	ram_block1a67,
	ram_block1a83,
	ram_block1a99,
	ram_block1a115,
	ram_block1a35,
	ram_block1a51,
	ram_block1a3,
	ram_block1a19,
	ram_block1a68,
	ram_block1a84,
	ram_block1a100,
	ram_block1a116,
	ram_block1a36,
	ram_block1a52,
	ram_block1a4,
	ram_block1a20,
	ram_block1a69,
	ram_block1a85,
	ram_block1a101,
	ram_block1a117,
	ram_block1a37,
	ram_block1a53,
	ram_block1a5,
	ram_block1a21,
	ram_block1a70,
	ram_block1a86,
	ram_block1a102,
	ram_block1a118,
	ram_block1a38,
	ram_block1a54,
	ram_block1a6,
	ram_block1a22,
	ram_block1a71,
	ram_block1a87,
	ram_block1a103,
	ram_block1a119,
	ram_block1a39,
	ram_block1a55,
	ram_block1a7,
	ram_block1a23,
	ram_block1a72,
	ram_block1a88,
	ram_block1a104,
	ram_block1a120,
	ram_block1a40,
	ram_block1a56,
	ram_block1a8,
	ram_block1a24,
	ram_block1a73,
	ram_block1a89,
	ram_block1a105,
	ram_block1a121,
	ram_block1a41,
	ram_block1a57,
	ram_block1a9,
	ram_block1a25,
	ram_block1a74,
	ram_block1a90,
	ram_block1a106,
	ram_block1a122,
	ram_block1a42,
	ram_block1a58,
	ram_block1a10,
	ram_block1a26,
	ram_block1a75,
	ram_block1a91,
	ram_block1a107,
	ram_block1a123,
	ram_block1a43,
	ram_block1a59,
	ram_block1a11,
	ram_block1a27,
	ram_block1a76,
	ram_block1a92,
	ram_block1a108,
	ram_block1a124,
	ram_block1a44,
	ram_block1a60,
	ram_block1a12,
	ram_block1a28,
	ram_block1a77,
	ram_block1a93,
	ram_block1a109,
	ram_block1a125,
	ram_block1a45,
	ram_block1a61,
	ram_block1a13,
	ram_block1a29,
	ram_block1a78,
	ram_block1a94,
	ram_block1a110,
	ram_block1a126,
	ram_block1a46,
	ram_block1a62,
	ram_block1a14,
	ram_block1a30,
	ram_block1a79,
	ram_block1a95,
	ram_block1a111,
	ram_block1a127,
	ram_block1a47,
	ram_block1a63,
	ram_block1a15,
	ram_block1a31,
	out_address_reg_a_2,
	out_address_reg_a_0,
	out_address_reg_a_1,
	data_out_121,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	data_out_0;
output 	data_out_1;
output 	data_out_2;
output 	data_out_3;
output 	data_out_4;
output 	data_out_5;
output 	data_out_6;
output 	data_out_7;
output 	data_out_8;
output 	data_out_9;
output 	data_out_10;
output 	data_out_11;
output 	data_out_12;
output 	data_out_13;
output 	data_out_14;
output 	data_out_15;
input 	ram_block1a64;
input 	ram_block1a80;
input 	ram_block1a96;
input 	ram_block1a112;
input 	ram_block1a32;
input 	ram_block1a48;
input 	ram_block1a0;
input 	ram_block1a16;
input 	ram_block1a65;
input 	ram_block1a81;
input 	ram_block1a97;
input 	ram_block1a113;
input 	ram_block1a33;
input 	ram_block1a49;
input 	ram_block1a1;
input 	ram_block1a17;
input 	ram_block1a66;
input 	ram_block1a82;
input 	ram_block1a98;
input 	ram_block1a114;
input 	ram_block1a34;
input 	ram_block1a50;
input 	ram_block1a2;
input 	ram_block1a18;
input 	ram_block1a67;
input 	ram_block1a83;
input 	ram_block1a99;
input 	ram_block1a115;
input 	ram_block1a35;
input 	ram_block1a51;
input 	ram_block1a3;
input 	ram_block1a19;
input 	ram_block1a68;
input 	ram_block1a84;
input 	ram_block1a100;
input 	ram_block1a116;
input 	ram_block1a36;
input 	ram_block1a52;
input 	ram_block1a4;
input 	ram_block1a20;
input 	ram_block1a69;
input 	ram_block1a85;
input 	ram_block1a101;
input 	ram_block1a117;
input 	ram_block1a37;
input 	ram_block1a53;
input 	ram_block1a5;
input 	ram_block1a21;
input 	ram_block1a70;
input 	ram_block1a86;
input 	ram_block1a102;
input 	ram_block1a118;
input 	ram_block1a38;
input 	ram_block1a54;
input 	ram_block1a6;
input 	ram_block1a22;
input 	ram_block1a71;
input 	ram_block1a87;
input 	ram_block1a103;
input 	ram_block1a119;
input 	ram_block1a39;
input 	ram_block1a55;
input 	ram_block1a7;
input 	ram_block1a23;
input 	ram_block1a72;
input 	ram_block1a88;
input 	ram_block1a104;
input 	ram_block1a120;
input 	ram_block1a40;
input 	ram_block1a56;
input 	ram_block1a8;
input 	ram_block1a24;
input 	ram_block1a73;
input 	ram_block1a89;
input 	ram_block1a105;
input 	ram_block1a121;
input 	ram_block1a41;
input 	ram_block1a57;
input 	ram_block1a9;
input 	ram_block1a25;
input 	ram_block1a74;
input 	ram_block1a90;
input 	ram_block1a106;
input 	ram_block1a122;
input 	ram_block1a42;
input 	ram_block1a58;
input 	ram_block1a10;
input 	ram_block1a26;
input 	ram_block1a75;
input 	ram_block1a91;
input 	ram_block1a107;
input 	ram_block1a123;
input 	ram_block1a43;
input 	ram_block1a59;
input 	ram_block1a11;
input 	ram_block1a27;
input 	ram_block1a76;
input 	ram_block1a92;
input 	ram_block1a108;
input 	ram_block1a124;
input 	ram_block1a44;
input 	ram_block1a60;
input 	ram_block1a12;
input 	ram_block1a28;
input 	ram_block1a77;
input 	ram_block1a93;
input 	ram_block1a109;
input 	ram_block1a125;
input 	ram_block1a45;
input 	ram_block1a61;
input 	ram_block1a13;
input 	ram_block1a29;
input 	ram_block1a78;
input 	ram_block1a94;
input 	ram_block1a110;
input 	ram_block1a126;
input 	ram_block1a46;
input 	ram_block1a62;
input 	ram_block1a14;
input 	ram_block1a30;
input 	ram_block1a79;
input 	ram_block1a95;
input 	ram_block1a111;
input 	ram_block1a127;
input 	ram_block1a47;
input 	ram_block1a63;
input 	ram_block1a15;
input 	ram_block1a31;
input 	out_address_reg_a_2;
input 	out_address_reg_a_0;
input 	out_address_reg_a_1;
input 	data_out_121;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \data_out~0_combout ;
wire \data_out~1_combout ;
wire \data_out~2_combout ;
wire \data_out~3_combout ;
wire \data_out~4_combout ;
wire \data_out~5_combout ;
wire \data_out~6_combout ;
wire \data_out~7_combout ;
wire \data_out~8_combout ;
wire \data_out~9_combout ;
wire \data_out~10_combout ;
wire \data_out~11_combout ;
wire \data_out~12_combout ;
wire \data_out~13_combout ;
wire \data_out~14_combout ;
wire \data_out~15_combout ;
wire \data_out~16_combout ;
wire \data_out~17_combout ;
wire \data_out~18_combout ;
wire \data_out~19_combout ;
wire \data_out~20_combout ;
wire \data_out~21_combout ;
wire \data_out~22_combout ;
wire \data_out~23_combout ;
wire \data_out~24_combout ;
wire \data_out~25_combout ;
wire \data_out~26_combout ;
wire \data_out~27_combout ;
wire \data_out~28_combout ;
wire \data_out~29_combout ;
wire \data_out~30_combout ;
wire \data_out~31_combout ;
wire \data_out~32_combout ;
wire \data_out~33_combout ;
wire \data_out~34_combout ;
wire \data_out~35_combout ;
wire \data_out~36_combout ;
wire \data_out~37_combout ;
wire \data_out~38_combout ;
wire \data_out~39_combout ;
wire \data_out~40_combout ;
wire \data_out~41_combout ;
wire \data_out~42_combout ;
wire \data_out~43_combout ;
wire \data_out~44_combout ;
wire \data_out~45_combout ;
wire \data_out~46_combout ;
wire \data_out~47_combout ;


dffeas \data_out[0] (
	.clk(clk),
	.d(\data_out~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_121),
	.q(data_out_0),
	.prn(vcc));
defparam \data_out[0] .is_wysiwyg = "true";
defparam \data_out[0] .power_up = "low";

dffeas \data_out[1] (
	.clk(clk),
	.d(\data_out~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_121),
	.q(data_out_1),
	.prn(vcc));
defparam \data_out[1] .is_wysiwyg = "true";
defparam \data_out[1] .power_up = "low";

dffeas \data_out[2] (
	.clk(clk),
	.d(\data_out~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_121),
	.q(data_out_2),
	.prn(vcc));
defparam \data_out[2] .is_wysiwyg = "true";
defparam \data_out[2] .power_up = "low";

dffeas \data_out[3] (
	.clk(clk),
	.d(\data_out~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_121),
	.q(data_out_3),
	.prn(vcc));
defparam \data_out[3] .is_wysiwyg = "true";
defparam \data_out[3] .power_up = "low";

dffeas \data_out[4] (
	.clk(clk),
	.d(\data_out~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_121),
	.q(data_out_4),
	.prn(vcc));
defparam \data_out[4] .is_wysiwyg = "true";
defparam \data_out[4] .power_up = "low";

dffeas \data_out[5] (
	.clk(clk),
	.d(\data_out~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_121),
	.q(data_out_5),
	.prn(vcc));
defparam \data_out[5] .is_wysiwyg = "true";
defparam \data_out[5] .power_up = "low";

dffeas \data_out[6] (
	.clk(clk),
	.d(\data_out~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_121),
	.q(data_out_6),
	.prn(vcc));
defparam \data_out[6] .is_wysiwyg = "true";
defparam \data_out[6] .power_up = "low";

dffeas \data_out[7] (
	.clk(clk),
	.d(\data_out~23_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_121),
	.q(data_out_7),
	.prn(vcc));
defparam \data_out[7] .is_wysiwyg = "true";
defparam \data_out[7] .power_up = "low";

dffeas \data_out[8] (
	.clk(clk),
	.d(\data_out~26_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_121),
	.q(data_out_8),
	.prn(vcc));
defparam \data_out[8] .is_wysiwyg = "true";
defparam \data_out[8] .power_up = "low";

dffeas \data_out[9] (
	.clk(clk),
	.d(\data_out~29_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_121),
	.q(data_out_9),
	.prn(vcc));
defparam \data_out[9] .is_wysiwyg = "true";
defparam \data_out[9] .power_up = "low";

dffeas \data_out[10] (
	.clk(clk),
	.d(\data_out~32_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_121),
	.q(data_out_10),
	.prn(vcc));
defparam \data_out[10] .is_wysiwyg = "true";
defparam \data_out[10] .power_up = "low";

dffeas \data_out[11] (
	.clk(clk),
	.d(\data_out~35_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_121),
	.q(data_out_11),
	.prn(vcc));
defparam \data_out[11] .is_wysiwyg = "true";
defparam \data_out[11] .power_up = "low";

dffeas \data_out[12] (
	.clk(clk),
	.d(\data_out~38_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_121),
	.q(data_out_12),
	.prn(vcc));
defparam \data_out[12] .is_wysiwyg = "true";
defparam \data_out[12] .power_up = "low";

dffeas \data_out[13] (
	.clk(clk),
	.d(\data_out~41_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_121),
	.q(data_out_13),
	.prn(vcc));
defparam \data_out[13] .is_wysiwyg = "true";
defparam \data_out[13] .power_up = "low";

dffeas \data_out[14] (
	.clk(clk),
	.d(\data_out~44_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_121),
	.q(data_out_14),
	.prn(vcc));
defparam \data_out[14] .is_wysiwyg = "true";
defparam \data_out[14] .power_up = "low";

dffeas \data_out[15] (
	.clk(clk),
	.d(\data_out~47_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_121),
	.q(data_out_15),
	.prn(vcc));
defparam \data_out[15] .is_wysiwyg = "true";
defparam \data_out[15] .power_up = "low";

arriav_lcell_comb \data_out~0 (
	.dataa(!ram_block1a64),
	.datab(!ram_block1a80),
	.datac(!ram_block1a96),
	.datad(!ram_block1a112),
	.datae(!out_address_reg_a_0),
	.dataf(!out_address_reg_a_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~0 .extended_lut = "off";
defparam \data_out~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \data_out~0 .shared_arith = "off";

arriav_lcell_comb \data_out~1 (
	.dataa(!out_address_reg_a_0),
	.datab(!out_address_reg_a_1),
	.datac(!ram_block1a32),
	.datad(!ram_block1a48),
	.datae(!ram_block1a0),
	.dataf(!ram_block1a16),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~1 .extended_lut = "off";
defparam \data_out~1 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \data_out~1 .shared_arith = "off";

arriav_lcell_comb \data_out~2 (
	.dataa(!out_address_reg_a_2),
	.datab(!\data_out~0_combout ),
	.datac(!\data_out~1_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~2 .extended_lut = "off";
defparam \data_out~2 .lut_mask = 64'h2727272727272727;
defparam \data_out~2 .shared_arith = "off";

arriav_lcell_comb \data_out~3 (
	.dataa(!ram_block1a65),
	.datab(!ram_block1a81),
	.datac(!ram_block1a97),
	.datad(!ram_block1a113),
	.datae(!out_address_reg_a_0),
	.dataf(!out_address_reg_a_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~3 .extended_lut = "off";
defparam \data_out~3 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \data_out~3 .shared_arith = "off";

arriav_lcell_comb \data_out~4 (
	.dataa(!out_address_reg_a_0),
	.datab(!out_address_reg_a_1),
	.datac(!ram_block1a33),
	.datad(!ram_block1a49),
	.datae(!ram_block1a1),
	.dataf(!ram_block1a17),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~4 .extended_lut = "off";
defparam \data_out~4 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \data_out~4 .shared_arith = "off";

arriav_lcell_comb \data_out~5 (
	.dataa(!out_address_reg_a_2),
	.datab(!\data_out~3_combout ),
	.datac(!\data_out~4_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~5 .extended_lut = "off";
defparam \data_out~5 .lut_mask = 64'h2727272727272727;
defparam \data_out~5 .shared_arith = "off";

arriav_lcell_comb \data_out~6 (
	.dataa(!ram_block1a66),
	.datab(!ram_block1a82),
	.datac(!ram_block1a98),
	.datad(!ram_block1a114),
	.datae(!out_address_reg_a_0),
	.dataf(!out_address_reg_a_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~6 .extended_lut = "off";
defparam \data_out~6 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \data_out~6 .shared_arith = "off";

arriav_lcell_comb \data_out~7 (
	.dataa(!out_address_reg_a_0),
	.datab(!out_address_reg_a_1),
	.datac(!ram_block1a34),
	.datad(!ram_block1a50),
	.datae(!ram_block1a2),
	.dataf(!ram_block1a18),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~7 .extended_lut = "off";
defparam \data_out~7 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \data_out~7 .shared_arith = "off";

arriav_lcell_comb \data_out~8 (
	.dataa(!out_address_reg_a_2),
	.datab(!\data_out~6_combout ),
	.datac(!\data_out~7_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~8 .extended_lut = "off";
defparam \data_out~8 .lut_mask = 64'h2727272727272727;
defparam \data_out~8 .shared_arith = "off";

arriav_lcell_comb \data_out~9 (
	.dataa(!ram_block1a67),
	.datab(!ram_block1a83),
	.datac(!ram_block1a99),
	.datad(!ram_block1a115),
	.datae(!out_address_reg_a_0),
	.dataf(!out_address_reg_a_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~9 .extended_lut = "off";
defparam \data_out~9 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \data_out~9 .shared_arith = "off";

arriav_lcell_comb \data_out~10 (
	.dataa(!out_address_reg_a_0),
	.datab(!out_address_reg_a_1),
	.datac(!ram_block1a35),
	.datad(!ram_block1a51),
	.datae(!ram_block1a3),
	.dataf(!ram_block1a19),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~10 .extended_lut = "off";
defparam \data_out~10 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \data_out~10 .shared_arith = "off";

arriav_lcell_comb \data_out~11 (
	.dataa(!out_address_reg_a_2),
	.datab(!\data_out~9_combout ),
	.datac(!\data_out~10_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~11 .extended_lut = "off";
defparam \data_out~11 .lut_mask = 64'h2727272727272727;
defparam \data_out~11 .shared_arith = "off";

arriav_lcell_comb \data_out~12 (
	.dataa(!ram_block1a68),
	.datab(!ram_block1a84),
	.datac(!ram_block1a100),
	.datad(!ram_block1a116),
	.datae(!out_address_reg_a_0),
	.dataf(!out_address_reg_a_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~12 .extended_lut = "off";
defparam \data_out~12 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \data_out~12 .shared_arith = "off";

arriav_lcell_comb \data_out~13 (
	.dataa(!out_address_reg_a_0),
	.datab(!out_address_reg_a_1),
	.datac(!ram_block1a36),
	.datad(!ram_block1a52),
	.datae(!ram_block1a4),
	.dataf(!ram_block1a20),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~13 .extended_lut = "off";
defparam \data_out~13 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \data_out~13 .shared_arith = "off";

arriav_lcell_comb \data_out~14 (
	.dataa(!out_address_reg_a_2),
	.datab(!\data_out~12_combout ),
	.datac(!\data_out~13_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~14 .extended_lut = "off";
defparam \data_out~14 .lut_mask = 64'h2727272727272727;
defparam \data_out~14 .shared_arith = "off";

arriav_lcell_comb \data_out~15 (
	.dataa(!ram_block1a69),
	.datab(!ram_block1a85),
	.datac(!ram_block1a101),
	.datad(!ram_block1a117),
	.datae(!out_address_reg_a_0),
	.dataf(!out_address_reg_a_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~15 .extended_lut = "off";
defparam \data_out~15 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \data_out~15 .shared_arith = "off";

arriav_lcell_comb \data_out~16 (
	.dataa(!out_address_reg_a_0),
	.datab(!out_address_reg_a_1),
	.datac(!ram_block1a37),
	.datad(!ram_block1a53),
	.datae(!ram_block1a5),
	.dataf(!ram_block1a21),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~16 .extended_lut = "off";
defparam \data_out~16 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \data_out~16 .shared_arith = "off";

arriav_lcell_comb \data_out~17 (
	.dataa(!out_address_reg_a_2),
	.datab(!\data_out~15_combout ),
	.datac(!\data_out~16_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~17 .extended_lut = "off";
defparam \data_out~17 .lut_mask = 64'h2727272727272727;
defparam \data_out~17 .shared_arith = "off";

arriav_lcell_comb \data_out~18 (
	.dataa(!ram_block1a70),
	.datab(!ram_block1a86),
	.datac(!ram_block1a102),
	.datad(!ram_block1a118),
	.datae(!out_address_reg_a_0),
	.dataf(!out_address_reg_a_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~18 .extended_lut = "off";
defparam \data_out~18 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \data_out~18 .shared_arith = "off";

arriav_lcell_comb \data_out~19 (
	.dataa(!out_address_reg_a_0),
	.datab(!out_address_reg_a_1),
	.datac(!ram_block1a38),
	.datad(!ram_block1a54),
	.datae(!ram_block1a6),
	.dataf(!ram_block1a22),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~19 .extended_lut = "off";
defparam \data_out~19 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \data_out~19 .shared_arith = "off";

arriav_lcell_comb \data_out~20 (
	.dataa(!out_address_reg_a_2),
	.datab(!\data_out~18_combout ),
	.datac(!\data_out~19_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~20 .extended_lut = "off";
defparam \data_out~20 .lut_mask = 64'h2727272727272727;
defparam \data_out~20 .shared_arith = "off";

arriav_lcell_comb \data_out~21 (
	.dataa(!ram_block1a71),
	.datab(!ram_block1a87),
	.datac(!ram_block1a103),
	.datad(!ram_block1a119),
	.datae(!out_address_reg_a_0),
	.dataf(!out_address_reg_a_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~21_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~21 .extended_lut = "off";
defparam \data_out~21 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \data_out~21 .shared_arith = "off";

arriav_lcell_comb \data_out~22 (
	.dataa(!out_address_reg_a_0),
	.datab(!out_address_reg_a_1),
	.datac(!ram_block1a39),
	.datad(!ram_block1a55),
	.datae(!ram_block1a7),
	.dataf(!ram_block1a23),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~22_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~22 .extended_lut = "off";
defparam \data_out~22 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \data_out~22 .shared_arith = "off";

arriav_lcell_comb \data_out~23 (
	.dataa(!out_address_reg_a_2),
	.datab(!\data_out~21_combout ),
	.datac(!\data_out~22_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~23_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~23 .extended_lut = "off";
defparam \data_out~23 .lut_mask = 64'h2727272727272727;
defparam \data_out~23 .shared_arith = "off";

arriav_lcell_comb \data_out~24 (
	.dataa(!ram_block1a72),
	.datab(!ram_block1a88),
	.datac(!ram_block1a104),
	.datad(!ram_block1a120),
	.datae(!out_address_reg_a_0),
	.dataf(!out_address_reg_a_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~24_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~24 .extended_lut = "off";
defparam \data_out~24 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \data_out~24 .shared_arith = "off";

arriav_lcell_comb \data_out~25 (
	.dataa(!out_address_reg_a_0),
	.datab(!out_address_reg_a_1),
	.datac(!ram_block1a40),
	.datad(!ram_block1a56),
	.datae(!ram_block1a8),
	.dataf(!ram_block1a24),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~25_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~25 .extended_lut = "off";
defparam \data_out~25 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \data_out~25 .shared_arith = "off";

arriav_lcell_comb \data_out~26 (
	.dataa(!out_address_reg_a_2),
	.datab(!\data_out~24_combout ),
	.datac(!\data_out~25_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~26_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~26 .extended_lut = "off";
defparam \data_out~26 .lut_mask = 64'h2727272727272727;
defparam \data_out~26 .shared_arith = "off";

arriav_lcell_comb \data_out~27 (
	.dataa(!ram_block1a73),
	.datab(!ram_block1a89),
	.datac(!ram_block1a105),
	.datad(!ram_block1a121),
	.datae(!out_address_reg_a_0),
	.dataf(!out_address_reg_a_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~27_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~27 .extended_lut = "off";
defparam \data_out~27 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \data_out~27 .shared_arith = "off";

arriav_lcell_comb \data_out~28 (
	.dataa(!out_address_reg_a_0),
	.datab(!out_address_reg_a_1),
	.datac(!ram_block1a41),
	.datad(!ram_block1a57),
	.datae(!ram_block1a9),
	.dataf(!ram_block1a25),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~28_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~28 .extended_lut = "off";
defparam \data_out~28 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \data_out~28 .shared_arith = "off";

arriav_lcell_comb \data_out~29 (
	.dataa(!out_address_reg_a_2),
	.datab(!\data_out~27_combout ),
	.datac(!\data_out~28_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~29_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~29 .extended_lut = "off";
defparam \data_out~29 .lut_mask = 64'h2727272727272727;
defparam \data_out~29 .shared_arith = "off";

arriav_lcell_comb \data_out~30 (
	.dataa(!ram_block1a74),
	.datab(!ram_block1a90),
	.datac(!ram_block1a106),
	.datad(!ram_block1a122),
	.datae(!out_address_reg_a_0),
	.dataf(!out_address_reg_a_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~30_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~30 .extended_lut = "off";
defparam \data_out~30 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \data_out~30 .shared_arith = "off";

arriav_lcell_comb \data_out~31 (
	.dataa(!out_address_reg_a_0),
	.datab(!out_address_reg_a_1),
	.datac(!ram_block1a42),
	.datad(!ram_block1a58),
	.datae(!ram_block1a10),
	.dataf(!ram_block1a26),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~31_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~31 .extended_lut = "off";
defparam \data_out~31 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \data_out~31 .shared_arith = "off";

arriav_lcell_comb \data_out~32 (
	.dataa(!out_address_reg_a_2),
	.datab(!\data_out~30_combout ),
	.datac(!\data_out~31_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~32_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~32 .extended_lut = "off";
defparam \data_out~32 .lut_mask = 64'h2727272727272727;
defparam \data_out~32 .shared_arith = "off";

arriav_lcell_comb \data_out~33 (
	.dataa(!ram_block1a75),
	.datab(!ram_block1a91),
	.datac(!ram_block1a107),
	.datad(!ram_block1a123),
	.datae(!out_address_reg_a_0),
	.dataf(!out_address_reg_a_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~33_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~33 .extended_lut = "off";
defparam \data_out~33 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \data_out~33 .shared_arith = "off";

arriav_lcell_comb \data_out~34 (
	.dataa(!out_address_reg_a_0),
	.datab(!out_address_reg_a_1),
	.datac(!ram_block1a43),
	.datad(!ram_block1a59),
	.datae(!ram_block1a11),
	.dataf(!ram_block1a27),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~34_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~34 .extended_lut = "off";
defparam \data_out~34 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \data_out~34 .shared_arith = "off";

arriav_lcell_comb \data_out~35 (
	.dataa(!out_address_reg_a_2),
	.datab(!\data_out~33_combout ),
	.datac(!\data_out~34_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~35_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~35 .extended_lut = "off";
defparam \data_out~35 .lut_mask = 64'h2727272727272727;
defparam \data_out~35 .shared_arith = "off";

arriav_lcell_comb \data_out~36 (
	.dataa(!ram_block1a76),
	.datab(!ram_block1a92),
	.datac(!ram_block1a108),
	.datad(!ram_block1a124),
	.datae(!out_address_reg_a_0),
	.dataf(!out_address_reg_a_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~36_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~36 .extended_lut = "off";
defparam \data_out~36 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \data_out~36 .shared_arith = "off";

arriav_lcell_comb \data_out~37 (
	.dataa(!out_address_reg_a_0),
	.datab(!out_address_reg_a_1),
	.datac(!ram_block1a44),
	.datad(!ram_block1a60),
	.datae(!ram_block1a12),
	.dataf(!ram_block1a28),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~37_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~37 .extended_lut = "off";
defparam \data_out~37 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \data_out~37 .shared_arith = "off";

arriav_lcell_comb \data_out~38 (
	.dataa(!out_address_reg_a_2),
	.datab(!\data_out~36_combout ),
	.datac(!\data_out~37_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~38_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~38 .extended_lut = "off";
defparam \data_out~38 .lut_mask = 64'h2727272727272727;
defparam \data_out~38 .shared_arith = "off";

arriav_lcell_comb \data_out~39 (
	.dataa(!ram_block1a77),
	.datab(!ram_block1a93),
	.datac(!ram_block1a109),
	.datad(!ram_block1a125),
	.datae(!out_address_reg_a_0),
	.dataf(!out_address_reg_a_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~39_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~39 .extended_lut = "off";
defparam \data_out~39 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \data_out~39 .shared_arith = "off";

arriav_lcell_comb \data_out~40 (
	.dataa(!out_address_reg_a_0),
	.datab(!out_address_reg_a_1),
	.datac(!ram_block1a45),
	.datad(!ram_block1a61),
	.datae(!ram_block1a13),
	.dataf(!ram_block1a29),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~40_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~40 .extended_lut = "off";
defparam \data_out~40 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \data_out~40 .shared_arith = "off";

arriav_lcell_comb \data_out~41 (
	.dataa(!out_address_reg_a_2),
	.datab(!\data_out~39_combout ),
	.datac(!\data_out~40_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~41_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~41 .extended_lut = "off";
defparam \data_out~41 .lut_mask = 64'h2727272727272727;
defparam \data_out~41 .shared_arith = "off";

arriav_lcell_comb \data_out~42 (
	.dataa(!ram_block1a78),
	.datab(!ram_block1a94),
	.datac(!ram_block1a110),
	.datad(!ram_block1a126),
	.datae(!out_address_reg_a_0),
	.dataf(!out_address_reg_a_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~42_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~42 .extended_lut = "off";
defparam \data_out~42 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \data_out~42 .shared_arith = "off";

arriav_lcell_comb \data_out~43 (
	.dataa(!out_address_reg_a_0),
	.datab(!out_address_reg_a_1),
	.datac(!ram_block1a46),
	.datad(!ram_block1a62),
	.datae(!ram_block1a14),
	.dataf(!ram_block1a30),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~43_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~43 .extended_lut = "off";
defparam \data_out~43 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \data_out~43 .shared_arith = "off";

arriav_lcell_comb \data_out~44 (
	.dataa(!out_address_reg_a_2),
	.datab(!\data_out~42_combout ),
	.datac(!\data_out~43_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~44_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~44 .extended_lut = "off";
defparam \data_out~44 .lut_mask = 64'h2727272727272727;
defparam \data_out~44 .shared_arith = "off";

arriav_lcell_comb \data_out~45 (
	.dataa(!ram_block1a79),
	.datab(!ram_block1a95),
	.datac(!ram_block1a111),
	.datad(!ram_block1a127),
	.datae(!out_address_reg_a_0),
	.dataf(!out_address_reg_a_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~45_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~45 .extended_lut = "off";
defparam \data_out~45 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \data_out~45 .shared_arith = "off";

arriav_lcell_comb \data_out~46 (
	.dataa(!out_address_reg_a_0),
	.datab(!out_address_reg_a_1),
	.datac(!ram_block1a47),
	.datad(!ram_block1a63),
	.datae(!ram_block1a15),
	.dataf(!ram_block1a31),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~46_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~46 .extended_lut = "off";
defparam \data_out~46 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \data_out~46 .shared_arith = "off";

arriav_lcell_comb \data_out~47 (
	.dataa(!out_address_reg_a_2),
	.datab(!\data_out~45_combout ),
	.datac(!\data_out~46_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~47_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~47 .extended_lut = "off";
defparam \data_out~47 .lut_mask = 64'h2727272727272727;
defparam \data_out~47 .shared_arith = "off";

endmodule

module DDS_48_v1_asj_nco_pxx (
	dxxpdo_5,
	dxxpdo_6,
	dxxpdo_7,
	dxxpdo_8,
	dxxpdo_9,
	dxxpdo_10,
	dxxpdo_11,
	dxxpdo_12,
	dxxpdo_13,
	dxxpdo_14,
	dxxpdo_15,
	dxxpdo_16,
	dxxpdo_17,
	dxxpdo_20,
	dxxpdo_18,
	dxxpdo_19,
	data_out_12,
	pipeline_dffe_0,
	pipeline_dffe_1,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	pipeline_dffe_10,
	pipeline_dffe_11,
	pipeline_dffe_12,
	pipeline_dffe_15,
	pipeline_dffe_13,
	pipeline_dffe_14,
	clk,
	reset_n,
	clken,
	phase_mod_i_0,
	phase_mod_i_1,
	phase_mod_i_2,
	phase_mod_i_3,
	phase_mod_i_4,
	phase_mod_i_5,
	phase_mod_i_6,
	phase_mod_i_7,
	phase_mod_i_8,
	phase_mod_i_9,
	phase_mod_i_10,
	phase_mod_i_11,
	phase_mod_i_12,
	phase_mod_i_15,
	phase_mod_i_13,
	phase_mod_i_14)/* synthesis synthesis_greybox=1 */;
input 	dxxpdo_5;
input 	dxxpdo_6;
input 	dxxpdo_7;
input 	dxxpdo_8;
input 	dxxpdo_9;
input 	dxxpdo_10;
input 	dxxpdo_11;
input 	dxxpdo_12;
input 	dxxpdo_13;
input 	dxxpdo_14;
input 	dxxpdo_15;
input 	dxxpdo_16;
input 	dxxpdo_17;
input 	dxxpdo_20;
input 	dxxpdo_18;
input 	dxxpdo_19;
input 	data_out_12;
output 	pipeline_dffe_0;
output 	pipeline_dffe_1;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
output 	pipeline_dffe_10;
output 	pipeline_dffe_11;
output 	pipeline_dffe_12;
output 	pipeline_dffe_15;
output 	pipeline_dffe_13;
output 	pipeline_dffe_14;
input 	clk;
input 	reset_n;
input 	clken;
input 	phase_mod_i_0;
input 	phase_mod_i_1;
input 	phase_mod_i_2;
input 	phase_mod_i_3;
input 	phase_mod_i_4;
input 	phase_mod_i_5;
input 	phase_mod_i_6;
input 	phase_mod_i_7;
input 	phase_mod_i_8;
input 	phase_mod_i_9;
input 	phase_mod_i_10;
input 	phase_mod_i_11;
input 	phase_mod_i_12;
input 	phase_mod_i_15;
input 	phase_mod_i_13;
input 	phase_mod_i_14;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \phi_mod_int_reg[3][0]~q ;
wire \phi_mod_int_reg[3][1]~q ;
wire \phi_mod_int_reg[3][2]~q ;
wire \phi_mod_int_reg[3][3]~q ;
wire \phi_mod_int_reg[3][4]~q ;
wire \phi_mod_int_reg[3][5]~q ;
wire \phi_mod_int_reg[3][6]~q ;
wire \phi_mod_int_reg[3][7]~q ;
wire \phi_mod_int_reg[3][8]~q ;
wire \phi_mod_int_reg[3][9]~q ;
wire \phi_mod_int_reg[3][10]~q ;
wire \phi_mod_int_reg[3][11]~q ;
wire \phi_mod_int_reg[3][12]~q ;
wire \phi_mod_int_reg[3][15]~q ;
wire \phi_mod_int_reg[2][0]~q ;
wire \phi_mod_int_reg[2][1]~q ;
wire \phi_mod_int_reg[2][2]~q ;
wire \phi_mod_int_reg[2][3]~q ;
wire \phi_mod_int_reg[2][4]~q ;
wire \phi_mod_int_reg[2][5]~q ;
wire \phi_mod_int_reg[2][6]~q ;
wire \phi_mod_int_reg[2][7]~q ;
wire \phi_mod_int_reg[2][8]~q ;
wire \phi_mod_int_reg[2][9]~q ;
wire \phi_mod_int_reg[2][10]~q ;
wire \phi_mod_int_reg[2][11]~q ;
wire \phi_mod_int_reg[2][12]~q ;
wire \phi_mod_int_reg[3][13]~q ;
wire \phi_mod_int_reg[3][14]~q ;
wire \phi_mod_int_reg[2][15]~q ;
wire \phi_mod_int_reg[1][0]~q ;
wire \phi_mod_int_reg[1][1]~q ;
wire \phi_mod_int_reg[1][2]~q ;
wire \phi_mod_int_reg[1][3]~q ;
wire \phi_mod_int_reg[1][4]~q ;
wire \phi_mod_int_reg[1][5]~q ;
wire \phi_mod_int_reg[1][6]~q ;
wire \phi_mod_int_reg[1][7]~q ;
wire \phi_mod_int_reg[1][8]~q ;
wire \phi_mod_int_reg[1][9]~q ;
wire \phi_mod_int_reg[1][10]~q ;
wire \phi_mod_int_reg[1][11]~q ;
wire \phi_mod_int_reg[1][12]~q ;
wire \phi_mod_int_reg[2][13]~q ;
wire \phi_mod_int_reg[2][14]~q ;
wire \phi_mod_int_reg[1][15]~q ;
wire \phi_mod_int_reg[0][0]~q ;
wire \phi_mod_int_reg[0][1]~q ;
wire \phi_mod_int_reg[0][2]~q ;
wire \phi_mod_int_reg[0][3]~q ;
wire \phi_mod_int_reg[0][4]~q ;
wire \phi_mod_int_reg[0][5]~q ;
wire \phi_mod_int_reg[0][6]~q ;
wire \phi_mod_int_reg[0][7]~q ;
wire \phi_mod_int_reg[0][8]~q ;
wire \phi_mod_int_reg[0][9]~q ;
wire \phi_mod_int_reg[0][10]~q ;
wire \phi_mod_int_reg[0][11]~q ;
wire \phi_mod_int_reg[0][12]~q ;
wire \phi_mod_int_reg[1][13]~q ;
wire \phi_mod_int_reg[1][14]~q ;
wire \phi_mod_int_reg[0][15]~q ;
wire \phi_mod_int_reg[0][13]~q ;
wire \phi_mod_int_reg[0][14]~q ;


DDS_48_v1_lpm_add_sub_3 acc(
	.dxxpdo_5(dxxpdo_5),
	.phi_mod_int_reg_0_3(\phi_mod_int_reg[3][0]~q ),
	.dxxpdo_6(dxxpdo_6),
	.phi_mod_int_reg_1_3(\phi_mod_int_reg[3][1]~q ),
	.dxxpdo_7(dxxpdo_7),
	.phi_mod_int_reg_2_3(\phi_mod_int_reg[3][2]~q ),
	.dxxpdo_8(dxxpdo_8),
	.phi_mod_int_reg_3_3(\phi_mod_int_reg[3][3]~q ),
	.dxxpdo_9(dxxpdo_9),
	.phi_mod_int_reg_4_3(\phi_mod_int_reg[3][4]~q ),
	.dxxpdo_10(dxxpdo_10),
	.phi_mod_int_reg_5_3(\phi_mod_int_reg[3][5]~q ),
	.dxxpdo_11(dxxpdo_11),
	.phi_mod_int_reg_6_3(\phi_mod_int_reg[3][6]~q ),
	.dxxpdo_12(dxxpdo_12),
	.phi_mod_int_reg_7_3(\phi_mod_int_reg[3][7]~q ),
	.dxxpdo_13(dxxpdo_13),
	.phi_mod_int_reg_8_3(\phi_mod_int_reg[3][8]~q ),
	.dxxpdo_14(dxxpdo_14),
	.phi_mod_int_reg_9_3(\phi_mod_int_reg[3][9]~q ),
	.dxxpdo_15(dxxpdo_15),
	.phi_mod_int_reg_10_3(\phi_mod_int_reg[3][10]~q ),
	.dxxpdo_16(dxxpdo_16),
	.phi_mod_int_reg_11_3(\phi_mod_int_reg[3][11]~q ),
	.dxxpdo_17(dxxpdo_17),
	.phi_mod_int_reg_12_3(\phi_mod_int_reg[3][12]~q ),
	.dxxpdo_20(dxxpdo_20),
	.phi_mod_int_reg_15_3(\phi_mod_int_reg[3][15]~q ),
	.phi_mod_int_reg_13_3(\phi_mod_int_reg[3][13]~q ),
	.dxxpdo_18(dxxpdo_18),
	.dxxpdo_19(dxxpdo_19),
	.phi_mod_int_reg_14_3(\phi_mod_int_reg[3][14]~q ),
	.pipeline_dffe_0(pipeline_dffe_0),
	.pipeline_dffe_1(pipeline_dffe_1),
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_9(pipeline_dffe_9),
	.pipeline_dffe_10(pipeline_dffe_10),
	.pipeline_dffe_11(pipeline_dffe_11),
	.pipeline_dffe_12(pipeline_dffe_12),
	.pipeline_dffe_15(pipeline_dffe_15),
	.pipeline_dffe_13(pipeline_dffe_13),
	.pipeline_dffe_14(pipeline_dffe_14),
	.clock(clk),
	.reset_n(reset_n),
	.clken(clken));

dffeas \phi_mod_int_reg[3][0] (
	.clk(clk),
	.d(\phi_mod_int_reg[2][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_mod_int_reg[3][0]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[3][0] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[3][0] .power_up = "low";

dffeas \phi_mod_int_reg[3][1] (
	.clk(clk),
	.d(\phi_mod_int_reg[2][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_mod_int_reg[3][1]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[3][1] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[3][1] .power_up = "low";

dffeas \phi_mod_int_reg[3][2] (
	.clk(clk),
	.d(\phi_mod_int_reg[2][2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_mod_int_reg[3][2]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[3][2] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[3][2] .power_up = "low";

dffeas \phi_mod_int_reg[3][3] (
	.clk(clk),
	.d(\phi_mod_int_reg[2][3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_mod_int_reg[3][3]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[3][3] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[3][3] .power_up = "low";

dffeas \phi_mod_int_reg[3][4] (
	.clk(clk),
	.d(\phi_mod_int_reg[2][4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_mod_int_reg[3][4]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[3][4] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[3][4] .power_up = "low";

dffeas \phi_mod_int_reg[3][5] (
	.clk(clk),
	.d(\phi_mod_int_reg[2][5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_mod_int_reg[3][5]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[3][5] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[3][5] .power_up = "low";

dffeas \phi_mod_int_reg[3][6] (
	.clk(clk),
	.d(\phi_mod_int_reg[2][6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_mod_int_reg[3][6]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[3][6] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[3][6] .power_up = "low";

dffeas \phi_mod_int_reg[3][7] (
	.clk(clk),
	.d(\phi_mod_int_reg[2][7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_mod_int_reg[3][7]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[3][7] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[3][7] .power_up = "low";

dffeas \phi_mod_int_reg[3][8] (
	.clk(clk),
	.d(\phi_mod_int_reg[2][8]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_mod_int_reg[3][8]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[3][8] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[3][8] .power_up = "low";

dffeas \phi_mod_int_reg[3][9] (
	.clk(clk),
	.d(\phi_mod_int_reg[2][9]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_mod_int_reg[3][9]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[3][9] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[3][9] .power_up = "low";

dffeas \phi_mod_int_reg[3][10] (
	.clk(clk),
	.d(\phi_mod_int_reg[2][10]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_mod_int_reg[3][10]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[3][10] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[3][10] .power_up = "low";

dffeas \phi_mod_int_reg[3][11] (
	.clk(clk),
	.d(\phi_mod_int_reg[2][11]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_mod_int_reg[3][11]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[3][11] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[3][11] .power_up = "low";

dffeas \phi_mod_int_reg[3][12] (
	.clk(clk),
	.d(\phi_mod_int_reg[2][12]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_mod_int_reg[3][12]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[3][12] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[3][12] .power_up = "low";

dffeas \phi_mod_int_reg[3][15] (
	.clk(clk),
	.d(\phi_mod_int_reg[2][15]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_mod_int_reg[3][15]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[3][15] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[3][15] .power_up = "low";

dffeas \phi_mod_int_reg[2][0] (
	.clk(clk),
	.d(\phi_mod_int_reg[1][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_mod_int_reg[2][0]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[2][0] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[2][0] .power_up = "low";

dffeas \phi_mod_int_reg[2][1] (
	.clk(clk),
	.d(\phi_mod_int_reg[1][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_mod_int_reg[2][1]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[2][1] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[2][1] .power_up = "low";

dffeas \phi_mod_int_reg[2][2] (
	.clk(clk),
	.d(\phi_mod_int_reg[1][2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_mod_int_reg[2][2]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[2][2] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[2][2] .power_up = "low";

dffeas \phi_mod_int_reg[2][3] (
	.clk(clk),
	.d(\phi_mod_int_reg[1][3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_mod_int_reg[2][3]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[2][3] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[2][3] .power_up = "low";

dffeas \phi_mod_int_reg[2][4] (
	.clk(clk),
	.d(\phi_mod_int_reg[1][4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_mod_int_reg[2][4]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[2][4] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[2][4] .power_up = "low";

dffeas \phi_mod_int_reg[2][5] (
	.clk(clk),
	.d(\phi_mod_int_reg[1][5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_mod_int_reg[2][5]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[2][5] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[2][5] .power_up = "low";

dffeas \phi_mod_int_reg[2][6] (
	.clk(clk),
	.d(\phi_mod_int_reg[1][6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_mod_int_reg[2][6]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[2][6] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[2][6] .power_up = "low";

dffeas \phi_mod_int_reg[2][7] (
	.clk(clk),
	.d(\phi_mod_int_reg[1][7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_mod_int_reg[2][7]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[2][7] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[2][7] .power_up = "low";

dffeas \phi_mod_int_reg[2][8] (
	.clk(clk),
	.d(\phi_mod_int_reg[1][8]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_mod_int_reg[2][8]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[2][8] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[2][8] .power_up = "low";

dffeas \phi_mod_int_reg[2][9] (
	.clk(clk),
	.d(\phi_mod_int_reg[1][9]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_mod_int_reg[2][9]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[2][9] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[2][9] .power_up = "low";

dffeas \phi_mod_int_reg[2][10] (
	.clk(clk),
	.d(\phi_mod_int_reg[1][10]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_mod_int_reg[2][10]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[2][10] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[2][10] .power_up = "low";

dffeas \phi_mod_int_reg[2][11] (
	.clk(clk),
	.d(\phi_mod_int_reg[1][11]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_mod_int_reg[2][11]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[2][11] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[2][11] .power_up = "low";

dffeas \phi_mod_int_reg[2][12] (
	.clk(clk),
	.d(\phi_mod_int_reg[1][12]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_mod_int_reg[2][12]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[2][12] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[2][12] .power_up = "low";

dffeas \phi_mod_int_reg[3][13] (
	.clk(clk),
	.d(\phi_mod_int_reg[2][13]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_mod_int_reg[3][13]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[3][13] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[3][13] .power_up = "low";

dffeas \phi_mod_int_reg[3][14] (
	.clk(clk),
	.d(\phi_mod_int_reg[2][14]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_mod_int_reg[3][14]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[3][14] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[3][14] .power_up = "low";

dffeas \phi_mod_int_reg[2][15] (
	.clk(clk),
	.d(\phi_mod_int_reg[1][15]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_mod_int_reg[2][15]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[2][15] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[2][15] .power_up = "low";

dffeas \phi_mod_int_reg[1][0] (
	.clk(clk),
	.d(\phi_mod_int_reg[0][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_mod_int_reg[1][0]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[1][0] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[1][0] .power_up = "low";

dffeas \phi_mod_int_reg[1][1] (
	.clk(clk),
	.d(\phi_mod_int_reg[0][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_mod_int_reg[1][1]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[1][1] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[1][1] .power_up = "low";

dffeas \phi_mod_int_reg[1][2] (
	.clk(clk),
	.d(\phi_mod_int_reg[0][2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_mod_int_reg[1][2]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[1][2] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[1][2] .power_up = "low";

dffeas \phi_mod_int_reg[1][3] (
	.clk(clk),
	.d(\phi_mod_int_reg[0][3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_mod_int_reg[1][3]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[1][3] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[1][3] .power_up = "low";

dffeas \phi_mod_int_reg[1][4] (
	.clk(clk),
	.d(\phi_mod_int_reg[0][4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_mod_int_reg[1][4]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[1][4] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[1][4] .power_up = "low";

dffeas \phi_mod_int_reg[1][5] (
	.clk(clk),
	.d(\phi_mod_int_reg[0][5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_mod_int_reg[1][5]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[1][5] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[1][5] .power_up = "low";

dffeas \phi_mod_int_reg[1][6] (
	.clk(clk),
	.d(\phi_mod_int_reg[0][6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_mod_int_reg[1][6]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[1][6] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[1][6] .power_up = "low";

dffeas \phi_mod_int_reg[1][7] (
	.clk(clk),
	.d(\phi_mod_int_reg[0][7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_mod_int_reg[1][7]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[1][7] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[1][7] .power_up = "low";

dffeas \phi_mod_int_reg[1][8] (
	.clk(clk),
	.d(\phi_mod_int_reg[0][8]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_mod_int_reg[1][8]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[1][8] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[1][8] .power_up = "low";

dffeas \phi_mod_int_reg[1][9] (
	.clk(clk),
	.d(\phi_mod_int_reg[0][9]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_mod_int_reg[1][9]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[1][9] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[1][9] .power_up = "low";

dffeas \phi_mod_int_reg[1][10] (
	.clk(clk),
	.d(\phi_mod_int_reg[0][10]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_mod_int_reg[1][10]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[1][10] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[1][10] .power_up = "low";

dffeas \phi_mod_int_reg[1][11] (
	.clk(clk),
	.d(\phi_mod_int_reg[0][11]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_mod_int_reg[1][11]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[1][11] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[1][11] .power_up = "low";

dffeas \phi_mod_int_reg[1][12] (
	.clk(clk),
	.d(\phi_mod_int_reg[0][12]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_mod_int_reg[1][12]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[1][12] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[1][12] .power_up = "low";

dffeas \phi_mod_int_reg[2][13] (
	.clk(clk),
	.d(\phi_mod_int_reg[1][13]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_mod_int_reg[2][13]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[2][13] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[2][13] .power_up = "low";

dffeas \phi_mod_int_reg[2][14] (
	.clk(clk),
	.d(\phi_mod_int_reg[1][14]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_mod_int_reg[2][14]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[2][14] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[2][14] .power_up = "low";

dffeas \phi_mod_int_reg[1][15] (
	.clk(clk),
	.d(\phi_mod_int_reg[0][15]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_mod_int_reg[1][15]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[1][15] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[1][15] .power_up = "low";

dffeas \phi_mod_int_reg[0][0] (
	.clk(clk),
	.d(phase_mod_i_0),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_mod_int_reg[0][0]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[0][0] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[0][0] .power_up = "low";

dffeas \phi_mod_int_reg[0][1] (
	.clk(clk),
	.d(phase_mod_i_1),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_mod_int_reg[0][1]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[0][1] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[0][1] .power_up = "low";

dffeas \phi_mod_int_reg[0][2] (
	.clk(clk),
	.d(phase_mod_i_2),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_mod_int_reg[0][2]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[0][2] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[0][2] .power_up = "low";

dffeas \phi_mod_int_reg[0][3] (
	.clk(clk),
	.d(phase_mod_i_3),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_mod_int_reg[0][3]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[0][3] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[0][3] .power_up = "low";

dffeas \phi_mod_int_reg[0][4] (
	.clk(clk),
	.d(phase_mod_i_4),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_mod_int_reg[0][4]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[0][4] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[0][4] .power_up = "low";

dffeas \phi_mod_int_reg[0][5] (
	.clk(clk),
	.d(phase_mod_i_5),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_mod_int_reg[0][5]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[0][5] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[0][5] .power_up = "low";

dffeas \phi_mod_int_reg[0][6] (
	.clk(clk),
	.d(phase_mod_i_6),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_mod_int_reg[0][6]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[0][6] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[0][6] .power_up = "low";

dffeas \phi_mod_int_reg[0][7] (
	.clk(clk),
	.d(phase_mod_i_7),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_mod_int_reg[0][7]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[0][7] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[0][7] .power_up = "low";

dffeas \phi_mod_int_reg[0][8] (
	.clk(clk),
	.d(phase_mod_i_8),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_mod_int_reg[0][8]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[0][8] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[0][8] .power_up = "low";

dffeas \phi_mod_int_reg[0][9] (
	.clk(clk),
	.d(phase_mod_i_9),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_mod_int_reg[0][9]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[0][9] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[0][9] .power_up = "low";

dffeas \phi_mod_int_reg[0][10] (
	.clk(clk),
	.d(phase_mod_i_10),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_mod_int_reg[0][10]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[0][10] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[0][10] .power_up = "low";

dffeas \phi_mod_int_reg[0][11] (
	.clk(clk),
	.d(phase_mod_i_11),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_mod_int_reg[0][11]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[0][11] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[0][11] .power_up = "low";

dffeas \phi_mod_int_reg[0][12] (
	.clk(clk),
	.d(phase_mod_i_12),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_mod_int_reg[0][12]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[0][12] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[0][12] .power_up = "low";

dffeas \phi_mod_int_reg[1][13] (
	.clk(clk),
	.d(\phi_mod_int_reg[0][13]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_mod_int_reg[1][13]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[1][13] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[1][13] .power_up = "low";

dffeas \phi_mod_int_reg[1][14] (
	.clk(clk),
	.d(\phi_mod_int_reg[0][14]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_mod_int_reg[1][14]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[1][14] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[1][14] .power_up = "low";

dffeas \phi_mod_int_reg[0][15] (
	.clk(clk),
	.d(phase_mod_i_15),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_mod_int_reg[0][15]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[0][15] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[0][15] .power_up = "low";

dffeas \phi_mod_int_reg[0][13] (
	.clk(clk),
	.d(phase_mod_i_13),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_mod_int_reg[0][13]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[0][13] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[0][13] .power_up = "low";

dffeas \phi_mod_int_reg[0][14] (
	.clk(clk),
	.d(phase_mod_i_14),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_mod_int_reg[0][14]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[0][14] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[0][14] .power_up = "low";

endmodule

module DDS_48_v1_lpm_add_sub_3 (
	dxxpdo_5,
	phi_mod_int_reg_0_3,
	dxxpdo_6,
	phi_mod_int_reg_1_3,
	dxxpdo_7,
	phi_mod_int_reg_2_3,
	dxxpdo_8,
	phi_mod_int_reg_3_3,
	dxxpdo_9,
	phi_mod_int_reg_4_3,
	dxxpdo_10,
	phi_mod_int_reg_5_3,
	dxxpdo_11,
	phi_mod_int_reg_6_3,
	dxxpdo_12,
	phi_mod_int_reg_7_3,
	dxxpdo_13,
	phi_mod_int_reg_8_3,
	dxxpdo_14,
	phi_mod_int_reg_9_3,
	dxxpdo_15,
	phi_mod_int_reg_10_3,
	dxxpdo_16,
	phi_mod_int_reg_11_3,
	dxxpdo_17,
	phi_mod_int_reg_12_3,
	dxxpdo_20,
	phi_mod_int_reg_15_3,
	phi_mod_int_reg_13_3,
	dxxpdo_18,
	dxxpdo_19,
	phi_mod_int_reg_14_3,
	pipeline_dffe_0,
	pipeline_dffe_1,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	pipeline_dffe_10,
	pipeline_dffe_11,
	pipeline_dffe_12,
	pipeline_dffe_15,
	pipeline_dffe_13,
	pipeline_dffe_14,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	dxxpdo_5;
input 	phi_mod_int_reg_0_3;
input 	dxxpdo_6;
input 	phi_mod_int_reg_1_3;
input 	dxxpdo_7;
input 	phi_mod_int_reg_2_3;
input 	dxxpdo_8;
input 	phi_mod_int_reg_3_3;
input 	dxxpdo_9;
input 	phi_mod_int_reg_4_3;
input 	dxxpdo_10;
input 	phi_mod_int_reg_5_3;
input 	dxxpdo_11;
input 	phi_mod_int_reg_6_3;
input 	dxxpdo_12;
input 	phi_mod_int_reg_7_3;
input 	dxxpdo_13;
input 	phi_mod_int_reg_8_3;
input 	dxxpdo_14;
input 	phi_mod_int_reg_9_3;
input 	dxxpdo_15;
input 	phi_mod_int_reg_10_3;
input 	dxxpdo_16;
input 	phi_mod_int_reg_11_3;
input 	dxxpdo_17;
input 	phi_mod_int_reg_12_3;
input 	dxxpdo_20;
input 	phi_mod_int_reg_15_3;
input 	phi_mod_int_reg_13_3;
input 	dxxpdo_18;
input 	dxxpdo_19;
input 	phi_mod_int_reg_14_3;
output 	pipeline_dffe_0;
output 	pipeline_dffe_1;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
output 	pipeline_dffe_10;
output 	pipeline_dffe_11;
output 	pipeline_dffe_12;
output 	pipeline_dffe_15;
output 	pipeline_dffe_13;
output 	pipeline_dffe_14;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



DDS_48_v1_add_sub_upg auto_generated(
	.dxxpdo_5(dxxpdo_5),
	.phi_mod_int_reg_0_3(phi_mod_int_reg_0_3),
	.dxxpdo_6(dxxpdo_6),
	.phi_mod_int_reg_1_3(phi_mod_int_reg_1_3),
	.dxxpdo_7(dxxpdo_7),
	.phi_mod_int_reg_2_3(phi_mod_int_reg_2_3),
	.dxxpdo_8(dxxpdo_8),
	.phi_mod_int_reg_3_3(phi_mod_int_reg_3_3),
	.dxxpdo_9(dxxpdo_9),
	.phi_mod_int_reg_4_3(phi_mod_int_reg_4_3),
	.dxxpdo_10(dxxpdo_10),
	.phi_mod_int_reg_5_3(phi_mod_int_reg_5_3),
	.dxxpdo_11(dxxpdo_11),
	.phi_mod_int_reg_6_3(phi_mod_int_reg_6_3),
	.dxxpdo_12(dxxpdo_12),
	.phi_mod_int_reg_7_3(phi_mod_int_reg_7_3),
	.dxxpdo_13(dxxpdo_13),
	.phi_mod_int_reg_8_3(phi_mod_int_reg_8_3),
	.dxxpdo_14(dxxpdo_14),
	.phi_mod_int_reg_9_3(phi_mod_int_reg_9_3),
	.dxxpdo_15(dxxpdo_15),
	.phi_mod_int_reg_10_3(phi_mod_int_reg_10_3),
	.dxxpdo_16(dxxpdo_16),
	.phi_mod_int_reg_11_3(phi_mod_int_reg_11_3),
	.dxxpdo_17(dxxpdo_17),
	.phi_mod_int_reg_12_3(phi_mod_int_reg_12_3),
	.dxxpdo_20(dxxpdo_20),
	.phi_mod_int_reg_15_3(phi_mod_int_reg_15_3),
	.phi_mod_int_reg_13_3(phi_mod_int_reg_13_3),
	.dxxpdo_18(dxxpdo_18),
	.dxxpdo_19(dxxpdo_19),
	.phi_mod_int_reg_14_3(phi_mod_int_reg_14_3),
	.pipeline_dffe_0(pipeline_dffe_0),
	.pipeline_dffe_1(pipeline_dffe_1),
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_9(pipeline_dffe_9),
	.pipeline_dffe_10(pipeline_dffe_10),
	.pipeline_dffe_11(pipeline_dffe_11),
	.pipeline_dffe_12(pipeline_dffe_12),
	.pipeline_dffe_15(pipeline_dffe_15),
	.pipeline_dffe_13(pipeline_dffe_13),
	.pipeline_dffe_14(pipeline_dffe_14),
	.clock(clock),
	.reset_n(reset_n),
	.clken(clken));

endmodule

module DDS_48_v1_add_sub_upg (
	dxxpdo_5,
	phi_mod_int_reg_0_3,
	dxxpdo_6,
	phi_mod_int_reg_1_3,
	dxxpdo_7,
	phi_mod_int_reg_2_3,
	dxxpdo_8,
	phi_mod_int_reg_3_3,
	dxxpdo_9,
	phi_mod_int_reg_4_3,
	dxxpdo_10,
	phi_mod_int_reg_5_3,
	dxxpdo_11,
	phi_mod_int_reg_6_3,
	dxxpdo_12,
	phi_mod_int_reg_7_3,
	dxxpdo_13,
	phi_mod_int_reg_8_3,
	dxxpdo_14,
	phi_mod_int_reg_9_3,
	dxxpdo_15,
	phi_mod_int_reg_10_3,
	dxxpdo_16,
	phi_mod_int_reg_11_3,
	dxxpdo_17,
	phi_mod_int_reg_12_3,
	dxxpdo_20,
	phi_mod_int_reg_15_3,
	phi_mod_int_reg_13_3,
	dxxpdo_18,
	dxxpdo_19,
	phi_mod_int_reg_14_3,
	pipeline_dffe_0,
	pipeline_dffe_1,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	pipeline_dffe_10,
	pipeline_dffe_11,
	pipeline_dffe_12,
	pipeline_dffe_15,
	pipeline_dffe_13,
	pipeline_dffe_14,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	dxxpdo_5;
input 	phi_mod_int_reg_0_3;
input 	dxxpdo_6;
input 	phi_mod_int_reg_1_3;
input 	dxxpdo_7;
input 	phi_mod_int_reg_2_3;
input 	dxxpdo_8;
input 	phi_mod_int_reg_3_3;
input 	dxxpdo_9;
input 	phi_mod_int_reg_4_3;
input 	dxxpdo_10;
input 	phi_mod_int_reg_5_3;
input 	dxxpdo_11;
input 	phi_mod_int_reg_6_3;
input 	dxxpdo_12;
input 	phi_mod_int_reg_7_3;
input 	dxxpdo_13;
input 	phi_mod_int_reg_8_3;
input 	dxxpdo_14;
input 	phi_mod_int_reg_9_3;
input 	dxxpdo_15;
input 	phi_mod_int_reg_10_3;
input 	dxxpdo_16;
input 	phi_mod_int_reg_11_3;
input 	dxxpdo_17;
input 	phi_mod_int_reg_12_3;
input 	dxxpdo_20;
input 	phi_mod_int_reg_15_3;
input 	phi_mod_int_reg_13_3;
input 	dxxpdo_18;
input 	dxxpdo_19;
input 	phi_mod_int_reg_14_3;
output 	pipeline_dffe_0;
output 	pipeline_dffe_1;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
output 	pipeline_dffe_10;
output 	pipeline_dffe_11;
output 	pipeline_dffe_12;
output 	pipeline_dffe_15;
output 	pipeline_dffe_13;
output 	pipeline_dffe_14;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \op_1~1_sumout ;
wire \op_1~2 ;
wire \op_1~5_sumout ;
wire \op_1~6 ;
wire \op_1~9_sumout ;
wire \op_1~10 ;
wire \op_1~13_sumout ;
wire \op_1~14 ;
wire \op_1~17_sumout ;
wire \op_1~18 ;
wire \op_1~21_sumout ;
wire \op_1~22 ;
wire \op_1~25_sumout ;
wire \op_1~26 ;
wire \op_1~29_sumout ;
wire \op_1~30 ;
wire \op_1~33_sumout ;
wire \op_1~34 ;
wire \op_1~37_sumout ;
wire \op_1~38 ;
wire \op_1~41_sumout ;
wire \op_1~42 ;
wire \op_1~45_sumout ;
wire \op_1~46 ;
wire \op_1~49_sumout ;
wire \op_1~50 ;
wire \op_1~58 ;
wire \op_1~62 ;
wire \op_1~53_sumout ;
wire \op_1~57_sumout ;
wire \op_1~61_sumout ;


dffeas \pipeline_dffe[0] (
	.clk(clock),
	.d(\op_1~1_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_0),
	.prn(vcc));
defparam \pipeline_dffe[0] .is_wysiwyg = "true";
defparam \pipeline_dffe[0] .power_up = "low";

dffeas \pipeline_dffe[1] (
	.clk(clock),
	.d(\op_1~5_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_1),
	.prn(vcc));
defparam \pipeline_dffe[1] .is_wysiwyg = "true";
defparam \pipeline_dffe[1] .power_up = "low";

dffeas \pipeline_dffe[2] (
	.clk(clock),
	.d(\op_1~9_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_2),
	.prn(vcc));
defparam \pipeline_dffe[2] .is_wysiwyg = "true";
defparam \pipeline_dffe[2] .power_up = "low";

dffeas \pipeline_dffe[3] (
	.clk(clock),
	.d(\op_1~13_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_3),
	.prn(vcc));
defparam \pipeline_dffe[3] .is_wysiwyg = "true";
defparam \pipeline_dffe[3] .power_up = "low";

dffeas \pipeline_dffe[4] (
	.clk(clock),
	.d(\op_1~17_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_4),
	.prn(vcc));
defparam \pipeline_dffe[4] .is_wysiwyg = "true";
defparam \pipeline_dffe[4] .power_up = "low";

dffeas \pipeline_dffe[5] (
	.clk(clock),
	.d(\op_1~21_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_5),
	.prn(vcc));
defparam \pipeline_dffe[5] .is_wysiwyg = "true";
defparam \pipeline_dffe[5] .power_up = "low";

dffeas \pipeline_dffe[6] (
	.clk(clock),
	.d(\op_1~25_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_6),
	.prn(vcc));
defparam \pipeline_dffe[6] .is_wysiwyg = "true";
defparam \pipeline_dffe[6] .power_up = "low";

dffeas \pipeline_dffe[7] (
	.clk(clock),
	.d(\op_1~29_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_7),
	.prn(vcc));
defparam \pipeline_dffe[7] .is_wysiwyg = "true";
defparam \pipeline_dffe[7] .power_up = "low";

dffeas \pipeline_dffe[8] (
	.clk(clock),
	.d(\op_1~33_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_8),
	.prn(vcc));
defparam \pipeline_dffe[8] .is_wysiwyg = "true";
defparam \pipeline_dffe[8] .power_up = "low";

dffeas \pipeline_dffe[9] (
	.clk(clock),
	.d(\op_1~37_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_9),
	.prn(vcc));
defparam \pipeline_dffe[9] .is_wysiwyg = "true";
defparam \pipeline_dffe[9] .power_up = "low";

dffeas \pipeline_dffe[10] (
	.clk(clock),
	.d(\op_1~41_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_10),
	.prn(vcc));
defparam \pipeline_dffe[10] .is_wysiwyg = "true";
defparam \pipeline_dffe[10] .power_up = "low";

dffeas \pipeline_dffe[11] (
	.clk(clock),
	.d(\op_1~45_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_11),
	.prn(vcc));
defparam \pipeline_dffe[11] .is_wysiwyg = "true";
defparam \pipeline_dffe[11] .power_up = "low";

dffeas \pipeline_dffe[12] (
	.clk(clock),
	.d(\op_1~49_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_12),
	.prn(vcc));
defparam \pipeline_dffe[12] .is_wysiwyg = "true";
defparam \pipeline_dffe[12] .power_up = "low";

dffeas \pipeline_dffe[15] (
	.clk(clock),
	.d(\op_1~53_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_15),
	.prn(vcc));
defparam \pipeline_dffe[15] .is_wysiwyg = "true";
defparam \pipeline_dffe[15] .power_up = "low";

dffeas \pipeline_dffe[13] (
	.clk(clock),
	.d(\op_1~57_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_13),
	.prn(vcc));
defparam \pipeline_dffe[13] .is_wysiwyg = "true";
defparam \pipeline_dffe[13] .power_up = "low";

dffeas \pipeline_dffe[14] (
	.clk(clock),
	.d(\op_1~61_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_14),
	.prn(vcc));
defparam \pipeline_dffe[14] .is_wysiwyg = "true";
defparam \pipeline_dffe[14] .power_up = "low";

arriav_lcell_comb \op_1~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxpdo_5),
	.datae(gnd),
	.dataf(!phi_mod_int_reg_0_3),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~1_sumout ),
	.cout(\op_1~2 ),
	.shareout());
defparam \op_1~1 .extended_lut = "off";
defparam \op_1~1 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~1 .shared_arith = "off";

arriav_lcell_comb \op_1~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxpdo_6),
	.datae(gnd),
	.dataf(!phi_mod_int_reg_1_3),
	.datag(gnd),
	.cin(\op_1~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~5_sumout ),
	.cout(\op_1~6 ),
	.shareout());
defparam \op_1~5 .extended_lut = "off";
defparam \op_1~5 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~5 .shared_arith = "off";

arriav_lcell_comb \op_1~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxpdo_7),
	.datae(gnd),
	.dataf(!phi_mod_int_reg_2_3),
	.datag(gnd),
	.cin(\op_1~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~9_sumout ),
	.cout(\op_1~10 ),
	.shareout());
defparam \op_1~9 .extended_lut = "off";
defparam \op_1~9 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~9 .shared_arith = "off";

arriav_lcell_comb \op_1~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxpdo_8),
	.datae(gnd),
	.dataf(!phi_mod_int_reg_3_3),
	.datag(gnd),
	.cin(\op_1~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~13_sumout ),
	.cout(\op_1~14 ),
	.shareout());
defparam \op_1~13 .extended_lut = "off";
defparam \op_1~13 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~13 .shared_arith = "off";

arriav_lcell_comb \op_1~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxpdo_9),
	.datae(gnd),
	.dataf(!phi_mod_int_reg_4_3),
	.datag(gnd),
	.cin(\op_1~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~17_sumout ),
	.cout(\op_1~18 ),
	.shareout());
defparam \op_1~17 .extended_lut = "off";
defparam \op_1~17 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~17 .shared_arith = "off";

arriav_lcell_comb \op_1~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxpdo_10),
	.datae(gnd),
	.dataf(!phi_mod_int_reg_5_3),
	.datag(gnd),
	.cin(\op_1~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~21_sumout ),
	.cout(\op_1~22 ),
	.shareout());
defparam \op_1~21 .extended_lut = "off";
defparam \op_1~21 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~21 .shared_arith = "off";

arriav_lcell_comb \op_1~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxpdo_11),
	.datae(gnd),
	.dataf(!phi_mod_int_reg_6_3),
	.datag(gnd),
	.cin(\op_1~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~25_sumout ),
	.cout(\op_1~26 ),
	.shareout());
defparam \op_1~25 .extended_lut = "off";
defparam \op_1~25 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~25 .shared_arith = "off";

arriav_lcell_comb \op_1~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxpdo_12),
	.datae(gnd),
	.dataf(!phi_mod_int_reg_7_3),
	.datag(gnd),
	.cin(\op_1~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~29_sumout ),
	.cout(\op_1~30 ),
	.shareout());
defparam \op_1~29 .extended_lut = "off";
defparam \op_1~29 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~29 .shared_arith = "off";

arriav_lcell_comb \op_1~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxpdo_13),
	.datae(gnd),
	.dataf(!phi_mod_int_reg_8_3),
	.datag(gnd),
	.cin(\op_1~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~33_sumout ),
	.cout(\op_1~34 ),
	.shareout());
defparam \op_1~33 .extended_lut = "off";
defparam \op_1~33 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~33 .shared_arith = "off";

arriav_lcell_comb \op_1~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxpdo_14),
	.datae(gnd),
	.dataf(!phi_mod_int_reg_9_3),
	.datag(gnd),
	.cin(\op_1~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~37_sumout ),
	.cout(\op_1~38 ),
	.shareout());
defparam \op_1~37 .extended_lut = "off";
defparam \op_1~37 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~37 .shared_arith = "off";

arriav_lcell_comb \op_1~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxpdo_15),
	.datae(gnd),
	.dataf(!phi_mod_int_reg_10_3),
	.datag(gnd),
	.cin(\op_1~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~41_sumout ),
	.cout(\op_1~42 ),
	.shareout());
defparam \op_1~41 .extended_lut = "off";
defparam \op_1~41 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~41 .shared_arith = "off";

arriav_lcell_comb \op_1~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxpdo_16),
	.datae(gnd),
	.dataf(!phi_mod_int_reg_11_3),
	.datag(gnd),
	.cin(\op_1~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~45_sumout ),
	.cout(\op_1~46 ),
	.shareout());
defparam \op_1~45 .extended_lut = "off";
defparam \op_1~45 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~45 .shared_arith = "off";

arriav_lcell_comb \op_1~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxpdo_17),
	.datae(gnd),
	.dataf(!phi_mod_int_reg_12_3),
	.datag(gnd),
	.cin(\op_1~46 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~49_sumout ),
	.cout(\op_1~50 ),
	.shareout());
defparam \op_1~49 .extended_lut = "off";
defparam \op_1~49 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~49 .shared_arith = "off";

arriav_lcell_comb \op_1~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_mod_int_reg_13_3),
	.datae(gnd),
	.dataf(!dxxpdo_18),
	.datag(gnd),
	.cin(\op_1~50 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~57_sumout ),
	.cout(\op_1~58 ),
	.shareout());
defparam \op_1~57 .extended_lut = "off";
defparam \op_1~57 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~57 .shared_arith = "off";

arriav_lcell_comb \op_1~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxpdo_19),
	.datae(gnd),
	.dataf(!phi_mod_int_reg_14_3),
	.datag(gnd),
	.cin(\op_1~58 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~61_sumout ),
	.cout(\op_1~62 ),
	.shareout());
defparam \op_1~61 .extended_lut = "off";
defparam \op_1~61 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~61 .shared_arith = "off";

arriav_lcell_comb \op_1~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxpdo_20),
	.datae(gnd),
	.dataf(!phi_mod_int_reg_15_3),
	.datag(gnd),
	.cin(\op_1~62 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~53_sumout ),
	.cout(),
	.shareout());
defparam \op_1~53 .extended_lut = "off";
defparam \op_1~53 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~53 .shared_arith = "off";

endmodule
