-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
0ul6qmyd2aACXyxLiZySlhDZBZKBXycWBTLiwA0o/m28yORvIpNSqH0m8QnG4h5pLhOiqEPtQYXu
zOCRnUADq3JwDwfIDieOOmFiXfM08KlbWK3Lkd4X3MwDXwjVMr4Z1ntglvTSKqxxze7DQwOBxzPK
okYtZMeYvRHl2TAF4XQnPRWspaYCF8WtR1vMH2VJkCjfB/zKE/TI3qQMMrmYRyB6HNgIGRWM/BYA
oZ8B9o51gXzU9Kf5xgHUz/rDwa/eF8ooE128e8sRmLCGx0DBZwrGGvIHIyxP4Zz54QV6iJ55k9Bu
fyO3cfi1cbuqc4wdOPDL0w6pCPg5+w67crMYPg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 7296)
`protect data_block
977XMAwHoeZqmnyIfP/1LXq1OxUiBkeMRMfUmCW88NtUXhgTvfdBgNGOECQgkdKVXF8wPCdRGa7P
hIsmoWSWhJUDGqyNHUtebIq0k+48ZY12HgIDJ/v95Zocypv5aFvo6VG9yF9TQQeH7h4zkURXcigm
asegb1dPx33ArpS6ufOKmBlMoYBwg/XrEwKK4AmQ+MzuuMour/T6U061WmbxUNb2C8ewXJEcmBH1
yLzkrwbMkXGXyYPKluB88Jrbvt8jrZtnCXiRK4WNCSFeVe0DoKBLiRp3sBmaa+xKveemWCRUTx4L
erH/RvCANS6CN5BBUcTugIU6ltPzOmxg/FqD/Qb5ELFNesyDR7uaQyfVISZtfBXVOrRdWRV7t6ug
nrMUvorBTTqnC9a+A72JU9Tasq75rT58rGA0Ytrtt6nH/bSRJPLZPTR/11oRgsDDdmqZx+hTrmRC
roz5nuS077sGnq55bZRtWE9UCKVvDpoHmPYIk917C1+gSMAAY/yrzb3kXFUd+eTBFr20ptgVmpBo
fKYsK8B0TPZX8Kpm5J2SmBVZbu3LqBiceDlkr3F1RbaVim08sxTYTJzLUG8Iqv4PaeKD/uHlRAU5
U8RZil/dj095W3DKXNyXToP/eSfh2l1SbWANsa6HYBxC4yXslANoyma3m3FS65SD0eNXBwnUOmBc
85Fb36q2UzGKc8z46f6H2BANavDGcPSfGSuvTRREEAxCFBz9OYfeo8q6wt3DeYBHTeZCqsomezlC
6c0yDRN+ONwY8KznrJDJHWMS4Fnh4eafUwxsxfaUyYzq3waR3jSivS/WcoyX4j20lr+U0op6Znm6
rBldjBYc6ROgYTI46+1epT9HasKQSCRv5Y5SBl7PFMDmlQf+0dCuX+Qgnm4Kcxjeea5D2iys1xwO
oN9DOu6eHcohlUQenRMPm4+54U0Vs6qlVX0avzUP2nFkgky3TM2+RJywsWZUs3jU/DuA6P37ptS3
auMkkIlxl8Xbs67xd3OotFOTYDNlRKXqdPIvnj8O3dUzL63jmhuZHCtoAZMwpHP+9GqjfFlsqdhn
216RwQpM3f2UpFXZWGrj52byAaE5kPSs1dwGRobkXCA0+KZHcslrr9wRRlITVe24R0VmCxGpcwe6
IftXwjTqCIb/eQwWa1iRMIW5hHH8PPpP3buMLppFjTcXpct2m0qVo0pt2AJ/jvGSKFeXogtN0ljb
tsftMTMWW55jn6/h1kSfnLPXBPHmgOvENJ7pvXgj4P4mlW/ofEpua3KonwfIWoX/L/1AFGEV1a/f
+FawioRb1fvI4Ov8qM1t598W1J2u6pv8Wu+X5jWjRXqvRihdLAoLb3vFQhqpvYWY6BSgFvKUi9q7
ECFfJpz3MWpcwr4w7EygDn2ZLSrtH1ezR6i7nBuYBkK8HHKmt49DEWvWXUxtyYil6LZ0zk4dTnNH
mls8GmjRl8aml4VkRi9XaPpOgT7L09bQJ3dBRmAhqGTO7Y0MMJKQL+ZU0eqxvAb6kIv517x93Pgs
e920Cx4H1vFmkVoE/geit0ucQw8sdp9L8ODYcCT3+8xF1LcsqY46YTBgjX1gToURB4mUHB9qF8e9
FlaSuUCmMo7hATOMFBlsM7eXJX6dRk8YE3YZStg8fIMEn7FqA7sdAk+zbW0uP+BrC9K/oddMZGbF
1t77Rfsb955inW5n68quuXcz+rSkwWR/aRHFeidIxRb+tKnqyIubJZWxwX/W8w36NjBslLKdvova
SUAEB7pMkVklTJYEIkxoNKfdQ4lbRKo3QZktrak3SZiM/WGoIQd0JGDq3ccycftSP6DNMWer6z7e
7zjUJ1kqalWpeT0a7TjZcR1CjIpRHn6GSIYdbcBYVMd+eKGJOvsZsLWjw8njlKepNZsIbdbxAvsa
3b8+8Q4cDILAUQWJxrmIJ1h++DUVyFX6Ti8SBkt2hxQKPUWIBR0yBlxmnvTo3ICsDYT6/Tt/X1Uy
+7xzlyyHw+qtbglYMdoaUWwJ1mJaII9488JTO4ggs89gANy/dsIrieqmZEfMfi5Rl63TUYvvQHIR
NuxzhXOOCtNZBUomEGkFrCxIopclcqjOTUA3sDeylQPvVlPOAxCT0uM4R6osM59x0QbxRQ/k88Cg
TgBtGTCiNJyGyoDeISj+GMZar3Vziay6Fz8qYdVO4Zoq2Pu2HQIs8atdD5rwJdH0iUg5TSZav51g
WFihtsNHxT9wMrFOIjAlGCbgEdYbpw4TVMzR8IipF4vHkDHkwSXe2UIq52KD2ZpxkEEeyY4kSL1F
HJ01NQZlt/ZGWv1HH4oUTjCAArezShF3avK+1LDK++qlV1BMgFGsskhRrmURRY9bxGR6Dit6tvdv
WgcpSDMiTpcmx7vw1ZU0plvx15j/tiQlrKavjkBK8hdtYCSOjE+InSut2E3XbfgXcFeWy66cGgHK
ZxRsy1CwPNDvcHQGww2serVYaOOgIMftigEQwh4VlwDe7k98gM/DpY/MezLK8F0pGaT1DiErEYrv
TLx50vNf6HIKxeQSMAr/957gs15E/QACEydDOE4RziVDjlB0yrCFksiyyHAOM1jYnNjDoS5It4Bs
XJ+Bc0EmR8njhUUZDULbHKin/pLX+N+lYasRQ8SKJOjR4eRg1dk2PJUvH4JE3sdRT4OtxXspH44j
87VWGArc7SeYrdcV/kUn6kZicJlbHhlRetoQdwWVyyFC3GQr/N2xXt1x9Gbfa2b+8bCyH3IomDlN
/IGowhitICZrB3MuvrpVsgKxYBPUhJPlWg5J5YntRyObcPzsWPsyLk+H1noOIsMpPjNO9SCsXJgu
OpVoeV6lgx/Y0rBe0vRViQxDc1WTauK2p6wRR+ZLXaVFTRn+/nCVUTHBi9RFeUEFLISI1C1qo3pD
vL7/5iwxmXaG+ggineWgvafPEVlq/dqcM400zaD5EDjru6K7BQklnXZHIgfRA+F8ZxcDxO4fE7aO
0puk7KXSOlInOu7BoDvYVfQusoe1vnAKDA65pRfJPr3Q+qqxI76DhsAUptkBO2e0R4KYm9Pt21iP
4G+9+kOgimKkLjF5kT1p8r/uHlJiVK0byVqgbySzJ/dl1U6AOmQ2OWryoVpfoxZBJpVyNJA/X+fN
Ru9ASFQakgazXxm/hF82yB2UyjkXln/DhquAB3js3gP+IsbRlvxKI5vwY3aK3x/KzrZ/MtdxnEvE
EzRf6q9WYJPtAFus3z0BcshkQNeZR92dzHZajuFRkEuFFONlVJo2Tr7bKtUPaEnH0xuItzpNEqw5
IphLztqPFxw+Q3kG5y14bmDAA/q/yjRJqTvi/4T7ofqgtuVYVGXVwRbIGGSr8udSR1+P/qx2ZYh3
OlVpZHHGckidQsZijgvMzRwT4657+hvXoE4Mj8mwNsm+Xq7WwLPPfDpyf6KP1t5u7JS4JyusOywB
6juoyc0sRD/2P0qm8PLTbOwUkES4TmmLWYk8nhXDGkL8nThuVV1iG+KSkss42FuSzgrtuxDMHweP
O9CsciGwdgf5JpUznF2eP4QmRwSHLr+JEFv570/O5Gvu3rjewVU40vY1Vd97PDTZiCauBrAnR98H
KgpJ2tyjXWVv4qCj4R+5LXtLC2kxRykqP3cGz7B/V+nHjLNhMycuXM2E9Y+WXiH7XMjIwY0AB23G
ljl3qmmdQInIj3LKsAY7gWOivwJN30T8GQf9S1Gcvv/VOxtBIKPWnOYLDJI2AmYzEVvXkitbnko0
EpzVSXZSeU+yFrAu8DK0wXwSERUuti1fz3eWb1o0VdwDPomjsOQW9U9pdqqA/jLVb32Gwo+AFntd
i8UDsuCIrUTabHIY/Y2VJ3e/7xpBeOvU5vNZQW+hLRi6AnnlV7wTX7iMRUSDNeoIsXhGSmrTMAxm
wTDq8IfNtUHemSsYpXYwSpxw+CgrsYFknJKFt0gJZ32gASC+Kn2Kj2FvtQ4/79hxwI1lJ2GFgYpJ
bioc0L5wK6hActPk7bkq8HwUj9w67M83qSt5XUnnec3sQ6HydFkUapNxmSl7AHXi4VzbqTAq8Mqu
Zz7F4N4q93Gom5T6kiJTvjJg63BS13iIAfQjQD+rH55XCCJ9cZMMDLp2vQ9cKjsWFqpDwzD941Rt
qvtA+WGmDs4pOA1C9Wy66dZSlB5PJsRCx07hwGhXO41UBEBtTA39u4MvM+qQYNzwj1cIUZPpNJlo
cSVOuAi5pkRy9Zhp5b+u7hjkTSoTryBlNiEZoJUhqPmJzrrsWJyUDwBCLjrCbl8qXAQmyBbAptsY
PxQr2urdwWcsAmHo3XXnuFdl1B8gwCr5CSHa8zJkGbwwaXKtywR3VCklc/KjgnKbDF1ZTJH5Fc3P
t0fBbME4iCH20Web2SHzPUYN57nx+Sg8ts1n8RoqqUvVpC8UVbmsTVB363mYx0WlcqJrcULNP0td
zAgt8sYyXTykX1NwhEtenlEmI3M9/8m7q80gFWdBf1BMcyVaIOtq/mC1CJqlPhH9+Xwm67z07VPg
hWbrWkfG9tLXQtKmjliKUACeEONefrWKcyDlDvndgnbofejdEsSkOP2MEwabdVL5n4yYCi3Mf2vd
UpwIsnidqFxVeYp0PLObMsIZUB5u8sllKAz31Dp9p7iu/gv7NG76WwfdGDbI22WI7VUSJY/jwh3n
0bbZ19WUfRnGiQcYDBuhTXIsP7ZDZ76WRYvsN3hSkzkQch4fQcBzuJmrRbqc05PZ7F9A8B4pZ4tA
Iho8IG+6CLpv4pSrckY+gw7vdHSlwwVl0HN4R6zNTp+XxdH1ZoSEMp3nZBoksry18qqJJ54ylf/d
2lkGnmpgxU1daJkwdp95KkH1a/GPveNpy7LQNS8k/1RJPfPmffusVvA0EdQewNiO1Sr8gLinllD2
1rbVyCHoGJw/si7pXGdj05iPE2U21pnVj9biRzrHQBus4r4aSJWdTda/FUwlxbpenzxprTT3Ryzk
oxNARMBkQ4xBiDddNmmoMiJG6x/63CIeFbLUjwB/OfKN4NNV0xvVCPzfOJ+rkC7KSPksrWUugmuR
BK7X99Kw9z8xLbWUNx6sHQEJGISgluH4RMsG+jnkvlQx6Y46nrFgIpsuOB6Q4np5ygH+1CDEDBF/
jPY5rPwRbtGpKZkEHI2jEx85IQfqfv1FlVO64IgB4drL00jKdbbbAfjaeCLjCy7ReV8Mu4UWwkwH
G2z1zUf48ziQqE/QFlLvLh9Jym5KIkC2J9o0ba1sJvm/oN+HctqC+YAhlALrxwCrLcWDyKhT+nLW
6Vq2lU3Km820ckrOI63VrL4IhTyRkjdFHhkMS19O7JbbfcjMKDo8BrMbxy2Uc+anqJi9uBM9Kdec
IP7nK9w/56ghNWyVhv3vAih7+AhcDn0ospzmBSVKuNuhnCJncP3HQaZgbPGO2icZtWlMZ0YwhOqb
rCF5IOQSdyBM8OeZR18iipwuiWuVrMapCK78g6NC5XrICmDovgac0sR+E2gIDeszFcqMK4OrKzQn
1n2KpaQ0nFscpYd/99gTMkJgv83uhSkVEOBtZ0q77akpZ/5//hChn+HRRsvcMAUaEngzD7fPrvUE
7qpxj2LUtjKbJUKfrjcQgQoNhXP/MlT0yhFdkbruFyd78agYV2NI/mFx9lBCxoLrWUmtbEmPTESq
15DrARrweXd2zuXgPTonlhCEvhp3JXvhsIzeBLJ9eMeuqtpduDBUjTQyfpDwkaLI5YESUmNheTsh
ChTg4YEvxVG+h2Yt1WXVOQmHduMoFZhfpRJmWW0usuZe/h/mutPIoTcK6MwdFPM1QqUOT46IZKTl
amqxiX7aHwwoSfqzTzZRtasCQwnTPq5A3HnG1t/aPQND2tJeSMA83bw9Dzz4Jty6bx5H6SQGxoYI
ASX3YUf4qa42Zt/wTUQSShqbkimazkJciMaWTrGln0x8fzA0CvuL5g/6BC01Z04z4a0nU1RLUA4n
CtpbuCwwQ3oOHxrcAw45HXmB2aLfydLlh0IKnKDfXx0mt1DrbWAMmhcOzrjyqu4+FnUprA0+GvwF
U/M4V+9E9c8YMMjn8b30ulkMsrC6hT6XZ0oDO0nv5XzGwoyK3aq33OCh081/M9pxZRSdRexaRrs4
8IeloVkxo2xbDbWnJvmFDZyNTtjvZ/e1Lr1u8X+XNkDzlbm75NBP8JoT5jC6CKLXq67Mt9xCbjqj
z9d5Lk84D/40OXi9Dd6tGJmfQ8a6AM9vZYOul6aNMsfO1YLe2XDT9e16IS7CQavk84pGMcpUuQ/I
5wFwE/Mrl42vcZjfDV5c1vlb3DxunnL1tkgdrvTP192zU4Z0IH7SOws8GlWr4dYvIpuidIqABEXB
oPfoIGNye0H13+0Y5wySRR3A0CMdUy11oZFMrCWtwpUyjRYoqO4dyAB8yqsmbrPM4M01caifN9EO
R1phrQF2qG+lKlfdonWiQBaPo7BlWXdW8/LsikLb301Atxy8fF+LmFrzaJGBKxQKR7bEXuLV8n/G
bigRWkifRYMXKJ/tX01tPvEpNYPUdR2/J3F9MhyTSxLBQ4TZK22DkrT8SCJJncOWvPgv5elXxEru
bO0gB0Y5OsJ0NM+6eEO7E9muZvrHG62U6EJAlzhJQ8pGs+jXsbGKILuL1lC4gXclMR0apqU5mJXQ
hPvLmSc97DTYugyumNGpLGep7bvu5jUwIskIUBdsClfISBpWY9iEUUHad3cCH9f8nWmYJRCDOQj8
nd9xZDWsCmUCqAkQc+nMLj1jsV/lAzW+d55Lhn4DcuyKVoIdMvg0wh3SrwAkhS0IYNNHqAjlDc7n
HAReldGS3aVXLql77sBHzHZsTKA1fMz3SMZNbdlHRtpSIoAouh0B3pRh8zMN+zhRJoO7b1l4UwJT
+GIAjdd7cDE8bQl7K7ipGVpUtKA52BeqUKEJbCpZSjfvtrt14hmkB9e2uy7n3ynt0C/34z4aSV5w
KljT0d/4jy9Xf4Zk+TC5DHsZGKgMQNaXqtljthrpn7Us6pzXO5Uqc0Bq0o+nmXMOBDUQwSwQ1uhl
+ZiRmGIjD1YSjF8j3Pt1bEBPoUCTl0yYEj3q3BS6khLI6kjPkJM6q43GFOgMobLkEwAVtkKvjvRH
G3YQJ2KHxb+NP70WVFq52v44fZPWDFz5xgCl4iUGO36VshzMRmtonPzqtihe7LcVRIjUTUkGFX10
+orFsoSbusKbhOv7eRDwI0NxcWYpoKBQhXM2XTbNk2Ge+Kr+ipQpZg9hSKDuOkJFjrzAX8tde+OQ
bBQ2V6NZYt8znUgZ2Bj2PLtSUUW+7OKOpU2dRyOmce2AP5MsKOyQ+Q//e8qQj/ooiYBecGxWGcr7
RzTO/Ug71qFo1UjBa/g5r8heVUkFQqHzwxsR3GQx9dsKc7ihMnla4EiQ7bq8WUgaqQpyRLv6x7mS
K4tCtAhNELlW9yrZYiiIIVek3G2SN5gWZXNff+JvyhKn90yRviCZpoliaDbiKlYknVJJu/QWWsIO
Mzww921EfT9U/3LHuUKzt7EqlJcrchbKnVg5nikDCs9uFksKuJqi9/6KEbwCvZtvk3+hEuDjqQEp
1GsnDyq6/KI9Lar2MSRod4e3QJaPq+iRgOD7PKQZ6qL7QHxPms4LExHR1Iq5b/5ymy82TdTkQZa9
qGo2tKMGJiLyGN94/LVOWj5TxPszxD6yyiNQz6VeAIMxexieLt8/zfNz/smF+mMmDu/VeG+sOXJT
8vlA8hZhGw9ngTuPqXd9E+MJ2l17muFTuiQJ+IC0RgKNOdo1BZmhi/7/PPKGH1giJIWEgeya6IoT
KjBR6D7n9H8AYWOFyShA+W8YHmq2RLmjl0oo/nrcM9wYk83WieKaUCWbOJo2sPeBeWts2gWjman3
PL2UFW+O4lMsLSYyKc5hQR5KG/GSnC/7vOZpetPHLw9cTTXTMNTMzUP2euq33wXsI3rfWDFlWGct
lloLGheYaZyBpaZUI+I3w7qpNzH8+cTvYpwlV33auQch8LC2NEkLgK6j7dS/tf9/T36cka+WlHi4
QycnN81A2oIRyrrQyzRW6SRgYTsLVOi2lZ3AHg/FaQU7rmz3ePMYVbS7TT3zhv5JnqL2ruWWPJSJ
UO/0NpQxmUQpMztV3TpfioDqCnDd65QYRxKutdjkDH9DxeaC14lNHkthrmj+7tinE1GztUIFUvUZ
WeshAkcyMtLMzgjsC7RcD45pVbZ/rx/+n9Hc20ebm3x/UvhJKyxv+9ISWJnE4rmjdyPKjYSK0BcF
9w+1JC3Xlqqe1KqlZAsL4pXPtoENpRodvyrOzBnq6RSGyvI7E+O3ASM3oJEoqaolm+I2sm7K8Glq
FIgJ5VCwhVxiYHtnBd9/i021lGbgHFC5lIJxfB33J06PY2y+STeYswiDB8ztg5YN5+Cab018u+2p
geLTjN+a8X/kWR7lm3I2Pfi0Une2eHehkFqXQwgT0peIX+2vn5BFMMi95I/YZg0EN+4phnZa3ACU
cb4T3nfWvPiHV5eZOtPE72Bq0LZZjp/HvhjwvzOFnjGy0tGbNbn5mIfSOu85V7YvHOX42Jy5Ir5v
WvQu+DjwPrEPgJa0loMGM+LdgkQWyRXD0Us6mPC2Pqy68onDf1sX6YWEwTHRU1qyUhZJ3DvCWlcj
IQyJWzz8MjTBeKSyLaouSnEbbjEquphlJUsUBa+AGM20QYka0dk3NVFj9a9UqbFSKNTPrZR7kOEb
EWhJufGiIXhgsNAifCHXKq+gqc+qgHgvbmmoQZe4eq5J/s0cmRuM6QolOJNRPHgSNbZBfL0Dsp62
yA3xKPX63VD9uLqIU+39Lau4QTRySQ+eL/kh8+ckGJudDfjGDgRm727/aoEIPTw79FWZWrZSEQ64
p99GIhq/lpFrWXxaw658FmdGT8DQYQaOqr1x7fUggcLB8buYI7pQHTtAGN+FTT+RVDR4h21RqE49
EvSHWDzwj22zwHbcKHZwncVmKdSS2AFOZcHpRjim3UIFfL9+iG+flAp4aPvkKrX1B6aQs4TqPfzX
jSlbsyzZ6V9Kj9T3Gv1Kyu8mYJR39dobxVGnMFMnQMMVVTwuaVVWH8gygdUR3waTVZSfD5e6mvEu
hWZ6XjjBCyKB3/wCQJ8lTHl0Yy5nq10dsUCGBPX0Cj6drmHR/LskEl27OR+YtVdH3/O97CxJAuPs
pE/b47cOnGVol3BnIcsir6ltd4nVLjLNwiL1SgEeRQg1x6cpMDYiEcQeAutWP1wvLedn8Sz/idiR
UPxQnv0sSd6YSBDrArUg1YgPjHovJ58bJQM+ygLrQifCWLYMYbfoE/ziyiovxg+BSC8rHtAYd4O6
p6AHBTAW4aEhcksj1EQtv8rVHrge+2l7SEKQg4PYsMsG0a3RPuOf6xOmKezN0a4+DO9XgLl3Lh9w
18o0LdKlgh5ggxPW0MyjJsdX/pDYvlt/X34hBkzEVw0nSL+0p8jrUk+OxYKr+Seyp7W9DC4Dt5Yh
Q9VenZTpdYVXkmRCRQm6KWWYdUIoNjGrHeAyLcwCy+OQ13phLTduoo+j63402g+2H3gDaCDG3e5T
nsOdYnR0b3RDQRT+aZtYjQUh/qAXeLCtgrYcw5dk4/+6CHuf0n0uGT5jt+AOyYRmS3FV9ysMu07P
XUVcS2cozUzluZz8t/nv/V6433haPFC6BSutcnZsOiD37utCVSiD/0QrXGw3pLokoU4NRVsTyyEi
ayKDXjkCq5b/k9FNIfQ/CIa/7eT4DYzyyWeff5PBbdSN1Q4dwcM93oNSXny8pxkt9zKKSx1msvsg
`protect end_protected
