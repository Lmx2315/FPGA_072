// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:37:06 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
G/hlyswqpUjsQ3gy6Xm5eD9B82c8+RCY++hFMksAag/c9t66PUVCrIk/8GBZA2QX
oSgwHpoYITf79lfspbT4mm0wDgU+toEBBT6PwwlsgBa/Z5Q661tPMWbN46J39T1C
gcT87GCE1MP8M5hazeXCRZaRZEnh5txvv9/vemjTQdw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 14080)
llmPIePGd3Qo99DiEPdbmm+F5BlEjbCtOgJhtJNzgHzbwct9pmvCB8G8dyF8pawx
Dfaf8jIFeI4/2p7XNnnopi07xZ5yrJudwQA7suojJGA99inbYtldmvITAArFFf4W
jmCCt2DIrgaoj6XOcKjQJwuaTDbZ9fyUehUxvosbe6T3PT/tOKP9tHS5HD4nVYwh
MTwyWSi9yG1yvtQEYmNn62BIYbhwZxTGUMollMHlHKkEnJO3vvB3hH6xvL7e69iG
DN4Wjnojh1B6c8TCiqp9LZ8BndAdmy9/woR2EE28hhT2tOvqMCwmQp40cjmDGP8r
/H0tRP5DtSnuP9xXTW2na1TJg0wB1C4oc57i2lQ20wkjtoCxwje7MNhK5kHZ0kjZ
StnZlt60Fr7WeUKpgVyaYvvYZYpZgn8xypHsYY7HX8DCBxZTJqZ6gQMApysRrHM0
mCp0VM9QAnJbGRR/b/JB5kKnjdSKEpSJkKZyY0mYhoTxnPrXRll0o/rtyn3zFumT
sZQlQ3fkKRsmHiCq0D4a9QXNscIYlLEJmBP0ugRlLFNZWACMpRXFn6UAYuab1nL1
X0Bh/TiMsJTFcjle9ePfH5GrY0K8XJLr/hZq2AIlwO8qVvTo/bujwC61JXzdyInf
6i4Bf0THPutf9Bl0/8UKJDfi9M2lDqiIqR5OWB6V7+QJEALl7o5KlQKkzOM6839z
cDfEx9JQBME7qBimN1u72RnJWKvx1w3M+sZubwvlhpsOksmuTL8djosa3KkE4quA
fe6w6G/iwsfNPjNNBQmvQ5sxOphNBVvuSGUheFIjo4Q+GI8kuS8KB/bL6KNkqJ1O
ohenSiT/bOyoOhphFmgNQRCBBekle/C1H2CU4rOIIm76mqIrUvQIx0TVIvwQkERT
B52QAeHUcu/Rcc0QwbNr0VxzQo/e2i6BUGpPtTzbFivQ9uYu0Q7lWCe50eBQcUZR
O33evVDL393F8H/jeie0Iqa4tYNICtcHCRJ4elzrm1fYHASA3Jyvc7a/go4SQAhB
e7mIG2ztbA6ZOOCg2YL0LqeogjY3hM+DQYwJIwJha//slTrs35u73OieWvpnlXIl
MIlHmUUB7QmrcE9vsswPyVEZzP+PbnHytlTFIqARKC4B9vpEZZgn73/IK2yjBjHH
v5WoOrnOAKcKDse0Yb826PqiDpMrGA8bE904O5yvPzbRCoEPwFsp+4CiH/XGOSjX
f4MGUgeNqguEppx+YDFu21fBa1akynE9nIhLnCKlOgNkR3JrwruSWe+za+PIpDxg
L2ZSWod1Fu67nKi5+PcwD4ePTqHTRMyObGOT1IC/GSFBuYquNAtqGsdUyree8cTO
hb5YpkYhcc8W0BTv7MORCYIJs6NSuauEJmu5bzu43UOL1wHScWzhiU75vmkRv6Db
LYkYY8q5XP6mVAURgGGSSuDjBzzOfzWUXybNlbe/3MDr5qGAmK6G3+CMjyAjmOqk
Q3TJyVL+yY0omsv7XA4eZI6KvqG9odnghFCtaU//1XqwGuIdefAz9pM1WXcMB5A4
B5kaRX9lH2XtS6nmyUvoK4C+TMx0Lxu0AVEpHh8C/zlEeaZKWnxhspLXnj7mhnqz
gICC2TQ+9PkmXCEzg957LDHEcCdte3fuvAVxju+orrb8Iaek28jdUMk+Gash6xNj
bczs/IZK5OCag+xrQPYljMOgQbQUlwlJlaQAcg6ccSZSbRNWTY+9Bv/95WnnsfXS
LgkpRTyQE3WJFTz2Z5vUdK7dn2kzdoWSY4c/0Jgv9gK4gxsGDHXwQl4s/QUOePJP
XElFtFP04j210Ng6jM2DPTck7w6NBp5f5VBzNxAMuJVU1qCOub8fA2L0TFvbtvM3
cKYA6QpS1fdSskfzHeaIpiVm+sDh8gAHxkffL0GkYqQhgHU6IztEtjZZLpzetmMm
AtjsqHxNiPURsBtQ1n4Xtro7+ANspUk0RlaLuOByWYUB4Tzogew4icadXQhR0k8H
W1oJo9hsEkfo2vSZGRy+GqSnZNQYl5+98/FgEkZtLlPWUTbMWiW3MwzBsn9rJWOp
XklAw+b036zJIcwJ/CQLK9LzsDXYS+lLygKP9+lG3WPj8d0kS2IQ1Dj+PoYxE+42
a8ccSDfbTPy+2PQHgByZ1icaDycD0r1T/dBUzJxvWbWAiVgqZp3vNJG/wuFjmqtj
xbSUa/B+WvkXFvzaQa6+RPK5ulskVU2uBEzPdQElpRtm673O8JdG1iXTITZ/+L/o
GJQonBaV3ZPbgtxGJgyyRpNvUfYRkVbKFBfi596U3MDYKwLVWGZOmLOJqM5Y8+NX
lTQb+pryY2vrN5n0xGfm71a+dBogS9wO2eoMBj/1+mtMgrnZ8KuspNTVuOh+ZeBf
d6BNFpV/9Uo61OIHYIBA1EEu5AT1aS2aH+/ZOkIXH8jRBQMKf27S17hj6/nA1CSx
gQp3JgMeMXHKG2bKUZwg4EAuI8PD+sLCpd6LKRvdqpsX/aW2Nxwwo90wbkrEdHND
A9qE5xegpgn7epR7Z1cGtCMQg+r+USqQ2zGZNmc2NwDYNuWy032h51h0l1f6v/93
tYZ6ipvXsc38bqo3KlCKWsEDORaWTqw9sRQrT4hcvnVvEo0W7p65HhiP+TABmBo5
ST6Fnkm7AOMXOu5ijdXswQwoaiFyLU46qcWBhXY6y81QavsIz9HF6vdKkNDDaDOj
dxAsPPXbKvMVHYXrpwT0Po4eDGj7d4vCIP1d3Mawi+mP9F2smOm1LavVgEMisRvR
G4jfm3jWWTKijuYhC3B8Dk8xWnjeZvMnkHpsvOPvt6iqy4qkiSxfcfM4Qp3+eAM3
NpBviiSUxdFLLR7UIz63Jc3Reg09zhUmnmom/1o4WYdHm1KyMJCZu7J9kMXL0b+6
ylp3I2mUdMbBKuZ02fK9YBRcOAzSiu1AWGDVCtGKlEm1cZYx3orz+TkNjYDsus3W
Ths+XWjW1h8TeUpmYLzh8iwXa4gdBRX5Fq60g7RgJFFD0LEYekMgDWP7JRbsfACl
i2PDiQ7EDDeaVNM9FMAEA0UDs5fHPxyj/AjpSiz6OgHd5xp5UFyTRF3iP2JFYD/5
TUwxrATMT1gpwOJE0SJsOBOefNnK65RHIeQaon0i1sS5PI2GCN9vAQZ8YBplqWZr
nFG/uKCMF2U73lwOh1afGgpthxbSV1uxgCNqeSoy/rvWjYGzI+fLseT1x6XJ0a/n
NXouvYf/h+Do4Z4UYXWB7X/3arxumKIHV5zxupHNk1rxNNdnK3I+7NRfMgazsLEZ
U8zs5S59eUx572iBNaR+6l/9/CrczNNUHA32RZozfy495qLBeJX0qh/UxeXFLPIv
GNfkyK3oScnL7FrOvpY1vYPMwyQn3g5W9z3BuRwCJCZtTJJXrVUWjHlsV6exX65B
u799lceQm7Vz41fSJE7FlMRRbFZsttyGCVe1GXzZHgxaMGCWoFRJRevz56dUCxTR
IWaCyCIKXsE4OvIVpJYl6K7fu0WvXyooffqole1JjoGoLEv8B14n59v87KFNMQ+i
qGOFhFS7R4dxdH221Cd18jsGW2dCRGAOG4k1r4wvPjTecplWGEOEwgAhCXCbDYxE
4qY8ZiQd3/PCul911FjIZsEfeRsT23No/IdUb3VOMIPOUiHHtqOBMOnMYCuIcF8O
XV3pdvVSQDASlsVlY39ljpiqTi5HIUvrUUGru5zyKmkQu1JIn7pD55K6gu5uY+/t
NIVsl8ywubrCmg51mvMTpMdeYI0+6oJx66MqQfmSheSTXdl1ews9CSWGZr2l1aIK
L6k6XGmkslcbwJDgcNu+23F9sBBx72Kj8f2XRp+A+bIPa6JjUt3TVO3emiNwh4O+
yK0he80iuuMOJ6V76Ta+kEOnDc1Ic96XtUEk+e4kNlVxnuEds1CanpgN7RNpn+tc
FSg84w03jD5bM/hmXDuSatMs6kM2eYy2xkuNiSqfeaccklgV4eb5Syq8iKmX/VhK
FchY+IUL+fXHCKFv2RPCXPsh7OS0DAgCQWoHqJEv2lDu4P0xjeeipKolwCxWPehU
V8I7rSOS05y+ZXUWBlc0tKKO5U2nAGCC3feF4DQ2bl8tidVCcyxM0Hp6XtHHuG2k
dcdX3ViJurSZXbb2DlOZwf4Th6Jtploo7ZpiRPI80Ecn5MEQcrSnXhF8yxJ/jj8k
ZHH8Md0Skonk9YhsXN1oX//neQPu6qDaA3XY3whF3U5t+96O+oplTtNXfKjGxmiV
doq4zepFkVsfctUyYJMVhVK7POfqSTok3pLHu9Et27EFeunFawsVB+aXQVhUf+BH
Q5ny+5dLGGIDT7516a4gMVJJEEgRs+TyD9gJod3o2cso/Ago6M/1IVz7G3dw/YD9
9S5cyLgk1mUmsOYMSZif2dHYsscLrduBPbGutH1PHlOmb5V/BFEMuwl5mrzEBQ6P
+/JbnUFp7IPiuwbkwaZpqR9VXMlgd9P3Xc938emCSkYR7wiNFEhGFOd7LptGsfF7
a8ap+gKr3jpWFQrp0bWKTxuMwuSroTPfMCkJ6mzXcADVypRldND3rZgO1tdJoTP3
2tBwkDdyFnN7kDcNkbumAb19jmKKRyTa3K44K690GncFFFZW/HomaIjJaS0TgSt0
l0CT+Hb+Gbv9tfYAXMAT/95pfdlspajHicI2ApCXpZwjV7WBNxDUXLCeCdWqExut
qUsh8800n/AMTdjlCwinwLa/TT9p6BuHgv4M+RzlF9YGWpvGNYX3iSjjrzNInz+H
sS6UnC4H4uC9ho8BDKdCFPx2gyexNXbL+vThAU8uGHrZkWN69vUR1JnFF8dZjo0s
J3B+6uH5GfeFa0nbhvpkMUsEF2TueGgSFntWe6hKkd2mC/nFYvvnOm7wV/Tho5TN
9AfMiKWZCzXocr375D5ewuJa7H7W0GbxlFkaxDTzoWYEsDfiOQVnt651QV++XARq
jEL+ZuhUqkLbqkfxHpGQyAmJRcvuesHs4tJ9oWmcfj3QBeyG1ZLP8LNyGcYJnDYD
GsCtfExaNuIGGwus/8woInwPo4fNFGGfGr9+I01TCwNUeAvHkuXw8rYZ8s3Z6KXc
kAgQ4h7IPzcxao5kJwEcRvXMvoscoK2t0jgBMm+6FKSUCoG3QzUQ6w3XA+OytMZi
bvIW86R2OlmrwfOH0r/KUPiYIbAtWwNrZOO8PMO5+h4tZKm6eE7hIAXpNAZw4+9l
CbZyw8P/u/pVgOFJQME1OsICk2vvBN2XkhHIITCGuBy1MK3yOaOaegTXEw6wuljb
xH5ZWuHX8nYBNHehSyPT39ek6cNv4eop+Gmn1UY5xjvuhtKhhOuBM7D3U/i4G6Wp
fPcagHSkYdH+HL+sCo34ecKYWwvagPc0qfgahmb0QOfxgoHhxZmv+7Tgta848pSe
Z9+6uDDBvCQ9wpU5BDEuKG7+sNmqJUiZTAeFYGXrVcQGChKaFzz5vZXvGV4k9AOo
1t4BYFr7YDR836n0pMQCW8kpHGm9MKT4vJLE1r0pzYtQsZaswCzcOCh8PsRhx41v
K9xvQH8ZBneerfnNnN/OxqIExV1NZgf0h0Ns7R9Q41bOqgbaUyAFSlxvaAtk5Dxc
y2yQLMDT1lBX5XAhcpoAXoRJJSnjbT9CIehBP7ETeckZKRBd9YRex/jIIgGYKiKn
Liy2dU58fYoK1QYh1BuXs3llpXgUb+5lXItHlcZohG1WF/IWt50EEOr0CwHm7x5S
lSxGlfOtIgeXjGREPHFNNa5art+CLq67UtO7daw06m6iqWhI1JFNd0GyyzSySjKH
rQtYVn16yEeiaJbm+clEDulqlikTvlDHq7kYvx2b9M7gmMNIciPgtBOTGjnZtQe0
0QCud6ptqxlbMzAQkvqrYzb0T57j9TzvLIt/+stjOdp/+v6Ws39cVO+864svMEx8
MqyD5q6bnRmd/jlacevErdj4q2ORNlHSlXsQ8D5UDcCMmPkiLwmgqVTmuv+wmHi0
wmmfoKntuf54HQFjIfCa6x8/4wE0UYl3AI96e2pRUpUtAzgKfWECqffbEDYfna2W
/YwaP0Jll+DuNro+KS77aWi3iqlpXq4tGh79/rNrlPRS/aDYOoKP9B7UxIUB+y1G
6v3e3ccbq9Nr74F6NtMyvK14Mv2wS2gX52UXaFvQcINv6TtRea3Mqjoh+UQZaRhZ
E2FWazRS0Y6R8b057YjTJS/6WpqM6WEAqIuj7TK/n4wJx9FzmRGuJJ6q/lpuTtMe
9JDJEfCocjXiKrsQqtM0oC0SQGjjoUruYd3wsHW2ivVKR/VC3NxUwXnw37sOSPbu
jyBhSKktuSs998zoC4gEG/nEqjn7dzIGz0mgm1kAB1BPx4r7faeRwDXAGoRbe3ht
rRAuI1PO0d1VYNLFC+1U60ncpDO0D0RaBMCsBrBXrQx368TiwiXdhKVlb84ZpZrN
HzZWzOA++R8yd2KVfcfaBnkIH9vJfp9qMh4I9Uia1ahIFuC/A7ZmlePQgYYKIt2U
i4GVevx13vnbQVFVFm5kE8OPO1+iHsIwAWzOmCkk6+yTqu0bBZR5DOJ7fPGuVk2e
YjQ5zfKEWs6tkWbC6hjTo7ECmMmnALRyvRlt6X5ZtfDUAbvRSVFNXgHoK7hyggWC
nqc111+h2pvcxW7b3Yilr1RX4yxbLISqR3IKBwxPRm5G8417oMOIR0MHb3v0BivL
YXvY4ef2CoufvQ5d0hGsXshC/s4nOxJWtnq+PQ9yPLOr70MAWaZab33MJ/CmO/v+
Pr9s14wLAsSSwCRTtWSld3LoQHlPvDfsYNhFShD0GN9a2Vz33Kjl58eQAreRwnMk
gtHjaeDlKrxvoAEHkGjkMCOdhO+jQatQUGgbMKNSzxRNQ44rFcbLD19LFHRC5tVu
SPAD/61k3KMVYXTp0jarfoDaQ8QegmZpTD+Vm2gis48kzFFFyUHHt9DFvWn+yQHq
n5R73s+13s5WFjmF9NIL+OWKIyKhlYli5u7+2l6RMtd9YDpjczOH2IGZVWH4vC96
a78tb4e2NqXDyXmjady+Bp+nuHMrlI6c8FEOQ1XcFFU/ZpmsAo3lzqGvIgCRAB1P
dFAlsb16qjYsw3ovlQr9sjcOeHwzNU0943ZFXArzXv6eumBpj58aVi0fcqBcZIEj
hHSPagDjAa9sxAQM/RTyW1ncBfD/c2cgd+0MgOieAKr+fAqKx0KaemRhSZhloblR
tOAmAthwUEPRnnLutE6gmmADL1T0aY8pAKd01qk6D/diGUEo53KBxr4PmuchrY7v
sdG7+mTZr2nQM5NoC28T7d0s2aIAeFcDandGIK8v1iiivXSbpRYOkx6JKVqbCJxu
z3ohU119baFdMexrUz/CcEpns8bk11XKp01T0GHuNHUJ7RxEKLEsfLTGVFEBoKUP
EPuTU5kiq5pBPrCr5s8zWZXJKXpKnR9HyvHKj8LTC3W2v9T9M1FeyovyAvUTx6l+
+TdoQ1uuZHPUhRf3WeaRj2s4vj6s5Sdas4P/q++r/T9QHMKwf9gl9ka3vimORsUR
T5KlwQmHvaXfLviWRyWlogvYpq/K6gEko5JtqWevGkzJqzdM9ISMCTs5JuaaCrje
mRlWhBNQSHbDxoIo4VCg2Hc701lDzsPSLVIijME4hJs0Hx9bHhy31h6qJZ9SQ2Sz
TVoSA0Rt6V6kudLkoBgpPg4RTpWKOkMKPbbNUOouDBr+ELobV9Mzj5w0K+PTDs/7
3Qd9s5vpU2AQzBPrqyxqmipU4WPp1jNXvUN7C5582xp+8jjVcGWguSdyK2xF1qAv
wZBc7K23KBH9RlUGmuTvUWkUkHKXK4To5FPy3rmRDy3caoRYgNe56LVUlj1OueeD
F3zQTNWdP0UjsYp0QuiKDPje3i+rssULh2kb7Y/ztO02bpb3eq+pFgv2g9V2qrmV
62icxkioVqrDt5Qu8VK9j7NNwkcb3D+gr6K30Onv4ygqzedar1Y2+5u95dDgVqB9
3A1RkQJnA034y18tb/IAGW0JB0lCfVXcbn1awhUoqaEE90W36VjCbVzhP9KmSWJg
HYsD+Qf0ggVWS1ftf9wN71+c6spsmtJHvvxMJXkyJuwX7NPRUQ/V9rki3z3aOB/O
/n+8zifixEvN/rxOQvaXqBuF/hjaxLLBi34k2ooFb4kjbBQuRxCQ09XfwW8vws7A
WAAe24vD+SsNNVATwDGs26afeJWxzZcE1ED8jh5hBBatUbbxrzLXOB9ggj+/gafl
H0bwv6+J+oJpzMLVn913E0oTP0a3SpcBH+QjtD3DYutph/mGr9diptNVkH8Y6Ttu
UvsGWe3RalZmpgqy3yEIAShA4Dym9xKAPRsVROQrEiTIf41YsRufZ1pNbDXxgsEg
SyGD4sy464kF5pufdxF3oaoqKneFnBmY8ZYU51WJZulzVeqrcWt+i2ZTLUjndlnO
Lm3ajH0Z1XofcKnDZFQCeE2SMRHfy6ldnr1ZYgKKtow9fY+OJdYUfaAG0wLbXolR
F8DHpjB/uiQOdUXW7OyvkvCgaN+KXTz2fGrDwLBxg0tAi97MkIKxJPWPnIOzQNRP
t+f1km7Q+DUQiOcapn9rAhAxmfMau01wXQBi5nhRQqGb7EKBK2PFKNkfVjgiV3R9
cUEbV5EpeFHUiFa8K+aBrg+Eef4rjaVnDRKZRMPEG4QrTi4kmKnvb/nHD+VqpANz
LFYmbsKxwsJB9bXxQ7EGl1I/OGSx3uNicmrVXkVZiYBI/i/BFaO6WUBi1jQSVclm
ZnGbOgBEpP4LaM5AOIBiHfCcFdO5yMyWrca0tgNCt6n3O0iDruaBOM7mhJR7Cloi
bToicg8DPsnB4RL4p7IN92D3KnXli4liVup+HdTdjfFWv3W5s6MFWKS8RYyFTs4n
+gwgbTx/3AAqeXob677Rq3Q+mr+rKU1MaO9lcrkpXKWQMc4TYoRgTRZLSaOrVmyn
U78ssFZYVod+ffHTW5dJJevhHKYrSZP350kmyeT4BDhCcwmevK7//Z0rhfYfpRN3
XgdvfiQJFsmtGZMDy/9YO9aLaAvFLoXnVpYK93h3LjLOLVy+Se4gWuebbGMz/vi9
29elSfcRu1eOZK0N7LyKlXf5W1bSpw2SZmixeVcu3YO4M7W18nwfUokUJ3B1qGP8
exuZIBeUy9YZTuY/FnxSbL8BWSu5AYmfWRaATJZShYKMuIibfGtT/+SLlYwoKcGd
HXK/CJDdODk6awMH9KfF5sjeeqfyCR1r5FPMX+ZNM24UfpiTAXTI6M6y7ZuA/v8d
PPjeEegxQDTeaJ5Dy182sLauDJVLFM1BvJN9B5heymmPHlIwqlw83GQd43U43uGr
clq6b9O0bnwH4u+/2Cwnog+ld1yItu0BmoH6HoG7l7nsuQxvx1bjqBPi9TuyXudR
58b2FdMr1u9VkrO+Nyi8/uhhyV6+rVHlwgn5z8jylQ8wOqZQq3Lc09foqQcTMFra
H366mmVy4O2PAkCb9SpomZ5OqRUwJRRwHzDz3etP74sMEWofioYC4EBgF3UBUD0x
AZhnigZeTTV5YtXMeltZIANTG36nrQAT4kV9AIOz0IeNyJP4Mc/KEjenkL9M4d5v
3f19BsTAc4bl7vIqd5CcGWCBwVgNABxJOam2gNBRCNmQjxmOtwvXROLhMWPTn62n
m60gXWJGXJugVZED3ptI/UwlbVS5HHpGDWPXLNv2P9daOChcbEoi6Botk4hItO7H
VeX5DwtIfTJNCJoJaET/YGugO0OgRDh04jvXPI9RJIEiMKDwaYhrVl9ezseROTmo
EhWmBKiXrYkyn/pMom7QxNuCd4Xk926hA2jno3cfd4RAhegAhnPNtvOcpXXQ6DVr
BWIb8OBsYueiIAarXSmqKedQqIxNowzKAu3r/8WCWofQtRRrUXbHFJjmoj0Rx3qE
LT304F7ZLiIO3OcmEcbFj+IJpDnYrj7EF4Iv8tlUpofmxeV9so3/fkgShN8olpO5
yQDRhk/otoYZuoe68bWZl27ZSlDZ6MBICcxAkFcaPKB4MzzjdeHBbosDOJ4IXjZP
7DHF2yalmvINE3P3ApWNYPPXtA9Q0a7SZUvu1MKePAYrvnYtXpnIbK1iDczReXRA
lFlnJgVb1a0rQ+EAG7SVPERZ+vfVZUlXOMBL/UFPgzAR0ff1pQO2PxhGdN0Xfpl6
QRygnQLNFxxaqm+U9nzLrH/OBiOTeVuSrEkLW49OHc2bcDFYBHk7eP4VE+Lz3wR1
Edf1o3xibx7meVZbg9t4axQA6f7gPOzaqw4aFb2LAvNIN5vfMZ5xiWkgoEcJj8vT
Lsa6wSWk4q3RpBTWuyJFavHfWrZAklwciuTIFNx7HGXq8ot/Sd5fTdBJXRnCz2Oz
Rn3vy+wJmD+Ashbbi1zYglNpL7axKITRatLSgn9DqKYG8HERcWhhbvcesSmnUtX+
PkT8Y2BkgvzP9Vdmg9dpEx1GOoW8nKpvGQbX67xgR2J6618puX+13KMmJiYG2QsH
Fq/ISJlltQyjr0KAq+anLj4eQklRoH6qUcNHrwsQwk6DiE/Q9o99EFtV4JDwWiLT
bZtwUuFjMtFFkBm4DVPhOy/hPORUZAeiyIWXwNaOZivpEZYuLKJ9q8G7SSkkDaU4
N++PNuLCRJnRfHSjE3TTOtfkQ+zuZRYlV8P9QXRnLxDXmYoCswqnsiu2utfzaR6q
Ltn/R/3MbAlN35dvrXwcyAWTfxJ9C/gaQ1fZOEpFlaM+aSyxGQnBzemprekAz5A8
w7bt9+QtjvsymxfkRCOH5ExORmk14WqWtyJHWtlLeUnQjLv3JNwZIWXFHzB45EAz
6tgKnaR5P9TLzqD9Uqx87lA05x8w3igshxiZHIwmMawo8HeLacFja6xLWEAU2JRj
TkPdA9RjywZ2GSfBOsvX2AkySyHpKRhRHKQxg7HnLlv3zucbGWhpqH7gyehDzEgx
D9XagoIA9FXm9p48eaXT+qh1cAmlHNNs9TwKPdCrF7zDORNvEr1FBBXlzWjipI8c
Wij5uzX+S+hH8B2O2fCfckdthafhA83cxU8H8hZcW91V60FISIBbE1bIjevG0w2J
zrUQN0dRMirfhdjP6ClbBc5igkXTQZao0WuL+uT8gcACPeCj19M36ZS1fu8X9DJD
yC43nM7yMQqQ/LyEpTB1+b9z6m2ETm/NRlpYYc5K1q0a15yfx3AZIPod406pp2pt
7EY0OE/vyt1ZF3U+SQOmZrrpdVgf9b+0nJfFQDhZJem6uCJPNqiaCT/Yoc5f9nLN
D9cVIEG38m1+oqKrNvzjpdWyGcq59kZtVJ+6zMOvvOLAtm6yO+pCX7epWptKHtV4
itcTGRpy2fkTK/t8Z01aidfPWPy830G8V2onnyYsIx4FnYQFXw/016VnwYOdkFgN
gFP7yJ7erCLqh0lGMO9cCaWtTS80pEK/lPqcwTc9xxzLQIFtkmBH1lXZmZXX79Hc
rNNJSCZosfj/GavGV0h+HEdeOxMzNO0QlZZUse8j2q+pgD3FfZs7aNyu2Yao5V3D
cu7+TuT4SJ35CGbpifblkfPKPqrZTSNWlF23Ww4ZH5aMt6EPGrM6PCWSGMyrnahP
LCUkk1nbYhi7COcKqQqUtvrrW09NcgF0z6Qbk2tK8rVApZJ+pQQUKiTSD1Tkjss2
C6xzOA0e5AuF+6jyWHo9yBCHGdTxOueGpPbBJJ/6l1CY5/Gmet9r8irOUjmyYnY1
QSTsafo32pSL/vVLIqzH+y18GAhwUFXJ+SLfo2LAu7HY3vzwinXS1+XYGuKKzKND
0vE44TznzBvmVYpscdNeQmasdvx3jlcJlL0QJFbyjMubmVGkKTFdC4+FgMt38/SF
KP5iN0P336JHGHJ6TxRYq3LknqaIed+7ctkMAWQJoIDagvjwrf55wUmMN7y8ZWDn
0bmA+WxJfWACMY1oxeeKJcSCmup6jGoHIL851K8VltmvtdBB0LzVXjZYsmsmzxyp
cUyMwCpskGsUodOIfPl8iXRK0FTPWu8dGi/vMZXB1i34JhXQHmWBcwfr+Now8oyA
akASI+F3L96nCFIMjvLu79awReNabqZ8F2z3P029SAc7qPO5zNywhQmpQseKWj/K
TqjKbePqDmLTqjgqlgyHu4MaRKL+gvUmxHK0DhE0AVrqyB8RRiBnpMIuXQhQO/l8
VB6ZywpeFYSOX4w1zIdJAeEIe4nKL9jeSSlejl8h+IckGLnRnYNkYlBvom8gDQG3
SXA9jCCSmEE4B/9DtVdlL8nATriAaUcOPNo4KXQ0d47DsJO1WXVGkWqOzasZ/+qd
Ko9fVkJ9CXsI+eZs3MqQqcirvCb1XGO/Uuu6nyLbvbfcSjSI8XVeQBPXUw/Orw6x
K/MCvjYKpQ4FlMjhZwzQMJ8FHrLQthwnlYU9nOONSyJQlyeodFxjEkdD+vmqgp+E
KJJl9wBS7ZSAc5Sk30CIqlVX1kX077CfxktmYOn8aKLRcK8LEUKuFjxJe4n4TtLf
vBSZDYHOktp9BPo6nxvNrJ6yY6Kz2IkDLbAnnnrZBj7S3A5s2RJJdbHc1CWqyqyp
vd2aD58SijoaeJ/82YFJEEa5bQJypL2L3BjHO8E9UJJJ6HZNdlCEe3OBIgD1QI+y
mMM3JKbv8yVczQXtKFICu9opwPd23LmN8Z/h4PaH5lpuUVUMJNN/iFs9OdFBJHAe
F7PM7eDRwrCxsZF3eChqUuxqdOTFqg73rahIhBkacd1t7DnKfPsnU7G2WU0M8Ft9
zL+woGTVpGRg3hfLus/wPuEmKqNyuvEJbJZscHB1BgyDt3vfP2/bE6Ug5efhtygU
8g8LOyr62JynnNIhaQoFrHrJ5V5k6GNB5lbpAlRhVZqEcR9ZUHMy08ROuRu5m+0a
7Nj/cTZ2Nh7PQyhAVAg5oyX5yRUcY8vLgT6Gqm4A0Fhn9FSB3enmUfeu3JATvs57
RB8+5uDztqjMXVaUC64r8sun/OnPPayq9wq1ky8v6Ev1awV3IiKUGMyAp/ybow3d
KPyFfOBYCVmuZ/5v0obbrSY/eOY4+ShZXcc3AYw0V1CHFqN74uEokrHtfZQjA2Da
U5fpek3nyI+qHgPPnvAbOWjkUzPBLK+sX+/4HuQLaUncqUKGJ04iSvY5Q++gbILk
CZAZYrrERdx6I/LdgRq3AG81uMThyuOKY5jp6SIu382BT/Ro+H047EJ462IM470D
Ru03qWYBiowwq//nqvcfwzO1uolIQD3N1Qpk+CAREbpdms9A9VtEBHMe1GL0FErj
uXxPzZQBZxpYGWaD7wc5/YD3PB0LPwm+oo91DXbdrjOUBRdOYyYymzXA28J5Txbe
CKEf6x+PBM8y8OjwwqgTtjRY5afRaD4iNzADHRwi6bMUYYNR25LXpm2wAmxG224b
wldeZHu7FFIpPba2ir+9GzJu+yYysxd7AVUlKPMa/8/0ooLJrSVftsGiBKl4r7SL
Q8Pu8YPCGBcrTUYNL4F13L4k34BLJpgkTa6959oM5nwuqPfelQJcr4UY9ZTHFE7s
L4ja8tQj2Bsy26g/c4wiU0llqrb5r0iQQbN4b0fGqCwfXcZ3FlMsq0kyFhwLhdY7
wuMqyQqQvX5t2J9LEGmdLlEhyuK+U8Ptu+bGCJCrzRe8IcfEOueKpQ7fkA7qEI5s
iMnT08vyD/5cQ0StVR2jj7mT6mo5Z+DPx1+Bee5MHNnER3dDST0qRVvJknc4FcCp
v4jV0bjfecMBNGO3FyXH+WGMx5S3XuJD4nDsoSkiN5dXVJ4BjZThIyWmU0o8UmEV
8HXvirj9sBJtgp3h3EIB7kFvRWggySOapUvNqd6KmuDk/sDcY83fBhlby9Ynn0im
hAdPkbQ6VCnxjbUS5hd6ZJ9R+xvCBhLWmRA7jLqRJdmALsFE2mX4XbRCkpeAkt5w
BNdeqwr7a51/YUuiYZOkLhNXJEcj0STW/abcEtQ6a0JUz1WcatVJeU5emx5owy6Z
xadCey2pYAzQ9KcGgY3i50zepDm9X2YutlW/p6tekKrtd4PoaxAC/2Hrnusd7CQK
f43Ha/hxee17vo0sA98h9XB4W0gNSatEJgdB8dtsDOO0hQ2qWvgQaFdm3F/0I8sY
yt41+L5vou6ULW0o/MxE1XORfLggoCv+F9LIMkrnfg2ELtYbbTlPJi4QXzxq+S0f
hXJPlkgK+AcQ/GQ5XxOr05vkHTBq0sdUA6cmmGrnIrXcUMOFNv0w4g/42YBX7NN3
gO1iX/5gfGySbxBgE6wHQWp16xm9iFVDaP+aLO6X3Mx7ELSl/ltNUDC7D6uqb7+K
0++PuFEiI/enhN22LrVjxkAeeyOPQeX1rX/MEaYVRT/wozmHY42p3cMH39TcX8PW
HwM2qDqMfGFKriOJazmJACFJ1T51F5N1IhY3f1EYx15aQ1Pd2gy96pKpyQifKOJj
djqCcsTGbi4iVPmsIAx91GXQZWUKW1ksnPKyisLFIapwFW1NMmC7Z81tecyEmZ+Y
fbUdw4SbKISdW7BLt/8Aeuy5DlJFOQ86+rsFyChgmWMGlbE/8rCfDOYAY9VE/bex
KnV94sGFgaVgcmUxlDC2bVqGLn/QudeVrZHqo4oKHVVD5Adllq3jWnnFHvHbfkN9
gm2i7yT2hHCezpd6bkVuP2H0zBRWMQG8doYuhZaYYMD64vD+IVgJhyD4L8SJa0Zf
+AAYhOz3izN7+bbVi/spYMC7d+BHitWJtXRSggc3YYkm24Z/025fUU3Vwj26Ou/1
FEvDm1tNsViLTTMyQSwL/rJyDB5DE5yikj3vRtPWNtOR2vMIUBsqcm75UKJyjd9D
2zakZlcKSwF0MkFtYI9dSrs0moi9w/QT6aYBGRn/w5yMlZk4+9DqlUqrNugsac/i
D9H/XdVXN0JWj4SbqYsDKcXeu8JZnBBRRd9CjuHVKUzr+PJogDH/N+Q1Rjm0qkvk
lamtinUO+cuFbJwDVP9IZj1q3dTmna3YVROwFT9OxNt6eAOsrN+YqWKMfkqgBt+J
FspRy+3jI6I+IubkPXfK+aU3IBzNE/lNXngJBBW/V3K8Via02PwtW19vUdaSowdI
nBLRz5V3z6xNFOZSJaF0kBgarLTTbHZH2DI2AHKBJQn5keDD5JHZRGEOO7Nju+9i
E33Pl3/+eaG3Oqk0Cb6umJK+CQ4NtBuJyNnVi2JOCScyLOvcFsLZC/wBm3QEodDt
GB9jKEtlLBNqKpbXQqE1cJWbsWFgnkZc1lPSCsnX6YyCs5VK1Ul29vD8Hrir68VJ
1owJrunWVYIuEfrq5/3Pjjq/QK5R+QitTZbDAStfXjW+RVqm+lyp0pZNKFNR5FUK
ORKgosJB02vL4m2v7tRFUffFw+fIHk4g/08zr44mA0zrcKMntxpnc0KbqOJjCoWE
aKC+RCPgThM9lko6u72UvaURhES48UZLOQiszrAMY/zjqCGriItZKd/3Cqce008y
xDpNcR50rdbRmh/OHpx8q0fSRE1QgQtjO8W73atLPs7yQ2RCXXE2OvHm7V1kCRGx
qjIBW8TFBqrfQdnGuQuyq63M/ecmhTJiUdAsj9TWmj3Y8NPB4NYHaQ9cf4E1YsTP
rLHbJsddsDXmkAIlfV7BNPpK0n3a3AAmm/loZHk0vf3IFQ6UnCEV57YrIbgNTVq7
vZxgTgEdCloRrrJHgG8B5PeuBxg3QqPcYJSb4WqtwOCdflTRi+NBXA30F9rt5927
O+09Z2N0X2zVBXrLpXV+anH2aBFdXh7iEov+12XTx5qWvlyVXuNN4US84I9jkrts
H+vXwYAb34a0sVKkOYud804P2Eu+PMdQ3Bvr4kugZvutm25+a3ZxnGX94pZRf2L5
kHFtByziLiEi2SUmRk6EwNqrHJAiqBpGX5JGP8VzDdzwvlhniqfZLt35rOsiZXGe
pwfyBKraRK9h8o43YHTSI8MjvMfYPOyy6nEr/VzXOhs5OxjWGHSGyG5jGVMqw8Ju
mJp/qCGhWmH/SNrz/2KqQFJOH6XF0n67MkYe9YGxKAFyQ8Ai0I6ad5iYmskLkq6i
PDixmtro1GVDpkxAm6C2l5uyNnWNo3AaTIe0MzxgXQ2oQDvHxoguKMn1BUgkP2Yj
QdcUhATDM3/l0U/EKP+In9irOT+4AEQp/m1QMJd8fpqXrpc9MJ3xHYb9ZXZMM4T5
Z+gDCusmFtbp1ON48fRmXkvyduVVVGJFtWyiLMKv2qLlMTBKbyfv4uvGH8ElJ6g0
tvM5xsduEc3Jz9imAQmychI+jaUDKmB1qdv7oyAUdSBwok71UaDnnPDOZjN3EqYg
SXydwB+UIx+ESCEUSMHuP2mToKYQuBFAbbhXqjbItRCJHd5oY0pLO0N97StQpSWx
FtL0z0kXctEYfHxQ4X96uD2hDqiqANb3PveomwFRFeuZa3gbTUUxo4QnYC74+wiX
CFMzRELrZpMcFAKQYONRn46nuEcgvkDSylSlxhR4Eb0ZolyfWkMQoNCaWQoG3x0q
kLjpCkp5Y4ht0XvifJH/rSQre0g1FFZX4yoL7a0HLmVM20m1f5FumAgEzdyvhPAP
G1wVRIp/Gt/jPXqkdVPFjg7ELmr3HcMqQBz1XuLLkEmmo/+GNe0H/8vejrukDzuQ
S8JEIP14rIOfbsgGwS+t+6MCB4DhqGABHtgKj2y/cW0OiZ0WrsTkDZEhOkMOLR1c
1ai0ixjALn3CI0zA465+x2gGWaMsC6r1A2WIhJYyrYDs+Mv7vTkgi0ERxs0OQAGK
pfiGtwQFk2IBnXg4k0TeFqxcaIXkWKhnmcLBFetQIXXyj/gBOQZWxN84p/0MW9Lr
0Oz6ierNHSYZYYpz++4+IKpmoL9m70jwNfUrGY1uJRAKJRUCftE9WM/NdA/YsRtw
AU0tkMFTRW/PmSldgUNQU+7/0S0vEwOPxUJuN23GM2LetIKysEyt7gsMGHAi3KJR
NtditQaY9UtWVoj+BVkfrBaY6zcIxrxJ8QYP567ZrAfrg+EbniHEPByuECSd8NIC
AHxa1ns52vY79+a1jN6HylHQGhUN4V534XfaoC2ssJfKk22XN0trZ9hIvuzyZh7L
Nq83bMDJUJTHAY8iDJavXJTIhG7Xx5WjfRYFit4ECwDI+0Wx5sos8RusOUDHSTBV
pih1sKBXkxezrcLqedXX6Nzf1/JQWQ5JJRIRwpNQ38A0eNeJIE1ttRQpYoVcyKlH
dei/kPwaxr5ZJOwHhIjJMMML1z8z255BCpllKbJ70Q3ZggGU93NZXQO90zoVwGqj
g6MD4mzeqx+o5LcPvDqwI24vwxwLUvoUw8cAllWKEveD3I6PeMU6Q7ik3+lZI99U
cXuL/VSY9hq2lctqSWg90ZNW9XPoeZCuqiYnp0fzpqXgpYAhKz+OmBKAL17kB4Qf
WKQY93zEq2xcvkVI09n9RucUgUhGMhj2I/5lTDsD6jvpvYUGI/d15XTUQo6H0TGB
5kPZNI37j1ZebRRxjZNqzNfoMJHX+QENHriVlFZe0WZTz42p16AiCE8s/kmJrXw5
31A6NjfouDnyi62bPNWmvCyA1BItuSIwBZU57bLzLj3ayfaA3ClzyK1H8CcvDX8d
2qv0A35u8xXGekiAzaEELzTR1NQB1lIqJ2yL9wIFOkJgPUhfxraNs54gajfdiB1Y
wj4fuHOPaGEMLD6Ad1QUFF9WH9sZ8Nx6YKOMRNd7bPuIb9OyJMipPQDB2kzjD4+M
IJaN71imS7onN6ryP1tm1fMpLwCDQ4JJeFoPiI6Cb/5afEr5yhJ5CvMSXznHzjKW
Eux146qr5Qrv+SYl7nd33WSymxyPNIht1F0iAK2UuUpp5Jtwv6widPEyZqzZhrQZ
cp4y9rfMCsDkJcjhCAsPUSIK0ofC6UaP++UNLsdVwY8t/E65AKsSoq9mm3OCj+wR
19uHPZwrtRh/38ti760HS5t9yTp6OrTRTcdpK1Y6mQhDr2XeHQG4wAQw4qdQJS2k
29QFOJt2M80B6LqQH9zAUXJnFKf0llqu0EGgXthTMenjilZLIWbdCqlPwNsmIV4d
9fC/nVOEIlzoEFF7S9zRo2D3wbHCoBGyj4uineqUkljcEWbscZq8VawX4gvsMwFA
l9YYPhTssnGilpQXLRLRqg3TFhUbJJyTZDUCDl1bIPOHbyrFSstYrwfWzUch8yIy
a/y9hGes5wbuAEbTdyTfJAy7EqN6cfexdn7m1Hc+ogJ+QgN+GmjqjPPed8IEkKAI
1YCjBCd0f84hJWWigki0d5dwz4K6kPNE12Kk8Glm6QyD8/6J8Qzrl0dMt/+ASIdj
LASIsZ9rL5pO4Ml9FjK1deRq49mLtOSl/otSUeecT9DT5K7NWM5Z1W/henZnCnzN
weVoCHHSzERT3KofX+ebEhqKsNqn3Vmmp0trp1pioYwXddIDk590XiVx+vodFr0h
qt07qVFd/EFUgbQCaqjUN2+15QemWQvqvf0dZlRai4ybf6koTcbZv1cbgZZWyF29
PyD6H4mmU1agTFP/PUPIuK06mMyTLZpkku1ia6BCmpkumQqQGphBpj+/SosZYFIR
YNjOgBbUVTV6v7k5VdVM5ie7WE1D615wldHwSADOVOpqpq2WGrDGmJShWaq3NoHh
0CUR4KO81qQNR6ucElCjPETuPihgMvtPzTzWniMy7lxfSS+KwWnAUsVvCNbCzxEI
SRxanhcM3C66El7Q2snEHMTDxyOEh5PDGlVjjEXDQpccNeSvMVe0IweTzQt0x+UY
KJ8wpc6Nx3LN67U62G/PmyvFKEqUNv8/wTxz79KyX5fFuWgt3NwtjQUsiMH1YucK
om03Zwp8vXKOFvRGgfuD+MsbmZs4Lde3HkZIHBaW9j2iRgYRrR4MjggC5s9gYP4v
Tj4LASL4xErUvPT4moIXzg==
`pragma protect end_protected
