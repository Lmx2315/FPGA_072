// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.0std
// ALTERA_TIMESTAMP:Wed Apr 26 13:36:54 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
mq4AO4yoI+nH7+ub3jicraeLRlp1VkWhsI7uxLLYMZPbcMiwHnSYhHNI1BvfoVcM
CPYC42Vb2cVrk2L3EwvKUTeGM4xDAT/4ftP1zvtFB0Mz0Y0LDwV19VsY/sLmFJ/W
nd/D1vEXfeDJ50PZN5RW4ngsAAu3B1q7gB3TXgJrV1E=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 21920)
3DUBhtYek2YtFQvQdJCWjyum2CBuSx2n8bgUmohrhsmY61uBwJpJl+wHI5ydrkZP
rfXQERCnkz6yaxZuuwQJwerfyH9t4VETj/vktVQ9yHpjN29hJLo2vY1+MbXBx5KF
g5ORTJOPPsHoCkpMFs1IFuzRXjb+E/wAR71HOJNep2IE7HO2bGVjD5gkIMf4miky
yEaPdcpuZzdxYMyyKDOPXlsddyyAnalNx2BNsvhvUApkbyqKqZoR+A0k06ZKPYod
afknrXnlCYiqUtZtXo2ArqJFbTVRhIyvZWQ1kjkJ7jDU89xZa51cIfHEFFfVbQiu
mh99wKCMHqVVd01jItN6oli1UvxQ5ocee1XqS+dJKn8bnN0Av3HPkolO9V8aQzha
17/Go9kbDsET3VfDXaxt5uwoV932RAy9AQOkvoQZULAkNsLzKYYN4adXjQegF57d
Uk9in17rjFI7HDI8fiAqKt+fAlApvMbp2/7rB0TSZ1OQUXWv5RMgNBXPZL0QxjtC
yE//Ub0ANtOXxsK/qO9vRAzmasi78FW+7ddW713X5zA6m+H+dW3jbPY3WSaGeJRk
3obeaJGwwKjI7CiwGUzeyW1K11CJe0JQtl0sLkzROLnD6NFY3aq/aOfcRfYKdM+6
jxFDwAvXqKiPHy8hNpvGL3VuwKMICKjgNxOqywRMxcMWrxslhX04TI3Lubt56jn5
dW0E3jHaOdIxAvWmw6WUN4/vZEBnV1Wckha3/JXDFg5ZKcQKMg0+C/F7ug1JmFHj
0ctFcbtGfu1h55AT/5Bv5/Ja+x21UytNyg1g6VGXEgxrhkFKOlOlUvxVjgqEj6Jv
ENdRQTz8HlKHOY+p94MuUMkKz+iklTtaTp3dFhmt+SDUm8oLCgXfjNDI2ZIHO6vy
ClMG/Ognr8ZW+1tYBhWf3AsOT1J3aE2t5W1icixlTLBa+k+kucoX/qsnDjiYOqyG
BnjFxWceYEDzdM0fKy/Dfp2ZsUxj5vCyWsD9Qiz+FCuOS8P+wnXPRGMKLpl8A8Jd
AVs5hOWmuh0WtYFhgcosyIH3/BRYrXVEOph5CwhuE63lHNDD305qn2ry27vgIsv0
CutKEH7CBxiBJnP5rJgWM3matXSwETlnqGgMIOcVvQ/bktRqbboX3GZE0sV6jmzJ
TZf+/i4FGOaDux19MGOYx3ry8GEm5lzoCVRpAmIhEV11SEUha8jtxP91ckoAvSCq
6YDEO5QLAYgSezCe02t3eLVs+2iCo0GQi4xU7hS8XsVa+TR+4/pgkgt2J9Pqp6Yf
7jTrZ0q7v/2RmdE6xjXitclbpJ9+9VSvb1givfsmDU8OrRybL0R/tCFz3aojTCLu
5hTlXuBAdxlT5F6F1g4PI2WMnjkDon6zA3mzEPOz+IntyDvstkHxNJqlnoaWqoyJ
+cdfT+hbwBinH6RyH7JRLB9vBFnICqZJerQq4T9L+MY4y7XVyjVyBhROnTEiZ5/L
1GHGXMumYLYxpwz49yv7quKqjtuVHfJ54QHP01rzBEzpg1bzbgH57hgJyYMsy6Os
2DuMkpFSNcog4s81GS4SXbk4nqfcsCMbylM8UDcGkhU0krYAsh1F747yWw+aDamV
ncqkICMbsd1buDY7xANGZvRwfc7snuvhaQ/peuEyXFoFPdzSV4NqrdpseaBLJrU3
Bi7f7W5XJ9m0WdGVPuZi5ET1a1aCXLJMuptkH1dMgtXExJgQMaD0/8Rbfrwq0Agv
V52GnP3J+lyiIN0YLb2nFLghXlIAiZSyxAbOWBNuG+hR9rPrVlolFus38lTaSl25
MXLBU00ae3IZOHbjx2PrEuHDI7guszKbUJGF5GOL83HDX+Fmkd0FqpR4n/Y4d7mI
HaweIKH4mZkLyMSWB0rtmTGR3BapYjh/EF00uf/fm/uBQ3BdjNCX2IxmbTFQestv
46kVyIROGSCVcCrXJAFfjaPr5F6ugm/AnRn0iNQS7CyvMu7UShOGkFlbAZ7OSU7+
8gnEwJ+jKH4iTUsw3sn1U83r4bc5rGprSp0jTd1b3YcVv1QM+43EARx5W7XchvUn
Z/1OreYOws9TpjtLY3uggQUze8oLUuI4bbyqpvxk9K+tjABx4vJICOERt4s07pEQ
I7ymi+/8PTr7/vGpT04O7HyT+3SFHGZSQRk4aZ2skcP/DlMmYJ7gOHUMzLK5OHVV
gJZseFFQGnhw+JI4C1BBRzX1Y5I5a+y5eKTsSfiYPDkPBaHR+27lnGTcJO/1Z7Wz
ziUaNCs8x/HeMg9fbMBnp7CbR2IcAVFMyy7TjcNPd5V6rod45XQhIeC6WW7Tv1dL
wVZVs05a3ZHEI3xXQPwlJ9DBFREMdXBUFOcp7ez0m78Nn/r4xu+I8q/D09myjfW0
PZ18JKNIMs4eejQyEahMsvR2Kvr1x+E/4vCGVAvQinLCXX0IdtQ+M82qxQoj3BsI
7PX8HIt/u6iJIVxubib+l51/qosrpfOxIrzBdVkubb5jOXfECZdGW4HktDuo6xz1
sg8ktIs9nf/p8dqzfBJQWbxhSq6Kk/XBRloAAs82i2qULIyfGlqyUohK9NXa/nfu
qZgMRGFbYQQVfurWCaw2PVQVEDYOjJJ30/SSl9Z6AIGr8L1blGAcQqt8/7HNlfS/
5puvcOFwBiUSkh+8VJyUWxDObRh3f5h6IN+mF+GwbUJemGTamQyCS1UqK69994DS
I4X3Xrt6WaWfeZMB5m98SRCJL7gOlwvbvX3IgYZGnZ19lAZEpbRaFwsFpHidOdR9
dtjUZ7eyvM32Xua5Yw8kZkVRnjLRgO1BphpjPzqD7WzbrwwZwD9RRm0jcD3EX1vp
oD8y4d7sXthlVENLyUl8mCNoksjmXumzHKfvfBPtCHXM05o2q3Z9jADBlum6ui0J
SCZ+Gi8xS8KfuCgpweTmwjoqQ9UP+sqISi0aB6o0iv3xGMLXlz357oA808MRT72v
pKocRwMYBSpwVz8KnAusLOMeJSi3XCg+/c1S6/dnb8JAz3inRE53xVs8U8vna34p
n78+cHq+LRcDcAg05gthOOBPW3f9Rw62pxqpeSgICQKgGu1m1R5WPnu3wvuRySZF
MmD8bLnBMgcQM0rVxA9wDmdye5tC9q8Cn53bZ399hiAHhhcrBbDs/Xo+4tR55tFS
FoePHMsxslwXo/RY7v9RJy90bfWtfrC91QJ29kT45+qcuCejgbLnUgQbrZWB6OAA
1j/D8rJpqorTFoNRUxh/SRJRHnoBTEahuYO82RUr62antACWtEuRLJPU3J7qEs0U
jovPCZubBUWk5GpTnw3SV2PrNDoXbmIxNcu0yWGNydLphVw//PtGX4PPCjzVsJaE
/KtuQe8VrgrHZBWYTwkJbrx/XxDZQnqqmlwjN2V/2SnQPyNg3DFBJQsKSPenaagm
1XstHdWGYKOL5BE28p8a3rkn4XsgkFY54SJXBlwQEOuzVuVh6WATW7QCWv6QSIK1
KurMEQwCG8l4nQoTmAAd/b2x3YNKnN3v4F+IL8ZrlAXhIR1Ou6b2GgQ4eDfOvnUT
IPY8KXOMn9CDetDVHOTt59dZrF0/QJVtUAFHWlgdQUJeJtKz8q0qqxJtEnLFqFH9
Cafz9Dc4J7MvvmUN5JEUk68HP6oFjcQvvFUU9qIZLdij6E0SxdPkUvNenUvt4VnP
LIMPKkQ9+OWo6mR4nvfhz7BSfoHD7iPFNIC4b9x9gKRUZ/WfgoBntb/knMR1smic
zIKttNWgIUOO9wUxvIJwjjFTGqnvIpBiXEd8mRSxCRgzGbBviBMMRGRuGO6YCce0
8UgYV2AP61bgoSTRqGQsZKJeN8BPznHPPnX8UV82tHAAOvzzbGKmYt1/ggZ39YUK
xj6wBKUoNzNsVxx6he8mT74GZFT4758wqkJ3WBZRIZuShzT4AKCAkez1ts4GrjPs
4vBGWWczpkLfYMmLtio8ArG2BInYnSSI35wk4pgU6YPieNKkgE8iStjxWhvRaoLJ
ElQMIZROmPUN1RQFWKe+ZawC4QlNH1VRLW0D0H3PKFyj3jTvOoPdveXtSXZZpPOZ
tBkq6eScSAg8L82g0Z//yIwb7+Melbn7ccG+ZY3cngukimoJtHoOcJyGe5H3VmWX
N0nEzKxB89hXSQ3W3p9+jpYaRgisaqNZHzdTQJg/u8fZAsxFrRkEyZG429EMs6vS
r0H1Jzi68whVOVqJ9Jry2UdwY03IO+hBPtAk7FlSk2jiu9ouR8adbtX4foEMfDNB
fWQxlHIL1YW88hjL1KrxFHH866hFgCy7PWXw94oDSGXY2LCB+EziGsudZKxCu74J
3y2mqmGlPGk0FmJLOAta0MjBEi7AIS9Tv2aIDwnpQRSC+WGXcUlqD+hfL0X9jyR2
2pbkGP2JIPhKh7mMZeAggnmmpUDBTglPPb9zPIOx6xCljp3MYIyAipX7Nzmea6mV
nBOAPesWFiQUuwHEv+SyauCkRKmWgRJu86YLGyUBPAw44KU4NRDgsIZGw16WSfZv
huYS+QXk8UZlMrIk9ezeovYR0QTAl4xrygU/EvcnFOCP49pYsm49oGKmjfRNIxHf
tLtlMOIW39Pnnwza9av6eKTCrl3g1EoqY0OKumnadGkwL12HQDi8PZuz95VWaMO8
Jj0CJ67bAUsPCxd1JhGj/uPqee4renxJnikjX/VSRYSByO8tnrGxf2iZ/+9ZJfAT
vD1zY/uIW5cz0zb3rg6Prg0XndC5TUPC6AFJ4YI7xg1X/DieWEgRvhFiAt3flcXs
CT2HBvOdBid2QmMGCoNn/N4SPmteRGEGaPzzu4TLCoNlUVzsnwgnaTD1R8cUlsut
7ZpWTzGuuOcI6KsWv3PtiUMQprRPzTdGZJhWhLcfMjSorDKSavFN+O++dpv53iIr
SLDXbpfubF09nEbmiYcTW4UCF0eWPLXcRBinG5NyQszeajlBhyHFalG7aKTrITuF
6APIsGVHiOnfFv+Am7V0kmjJB6iThMgkNJUfBnsljo2dtkv7945EZZjoFm12GSBa
cjAGmWidcHNdZU5DDiU1t4290HZs78o6+j45/YPpD2PYISoz5RzZ9zOIx3yITID6
7yAnLVN0Zu7lbXfRuyYzTMqWZPzxrSb9Dhnsgy4qJOJapWsDlqabrzRmMsZdH5Ek
iYZQVt23VOdphx/Q7UV08HYkj+sVbOeST4Z2JvaChcTPOOv/aIB78LpBrO8aK4kH
lvwO1O1GW1xMo+1j6DY4rW5U14u+kwjbZTBK8f/x0Rzx1W6nYPOJFd1B+wwIRoWt
GeaxjU8Iy3F40BGw3C3MpCIKGecC5wAHWD7uEnJx6vq2KHFgdKWk+HGXD8IjAy9E
SRIv9sMRxEFFYLyOYS2VeELfjRbxcjWyNqLlyL5EAeN3Iao3ZgxT1swzvd/3DTIo
v9NQ+AcrM93tTDIgCO3HFhsnSxa7oupp78Ic2EtlO5FtKgZVEe0hPYNgCb/9XkYB
5VgTv/R1GZjusg/4rgCU1v8TKztgnxQYJPe3u9Pj6oBh5PWueMlhsHLFgl1IORcw
XYhu31XMvapzTOrIurFreiT3Bf/SZUjJw0pGaawMfDXItpnRbmhAAkveHwEBggNC
AtXQ634BZDjY6UvwS3nDEc9N16BU7McWKEmp6HczstWCd6kd0mFP3lwNN4jhB6jG
kGPqDFpPDkzAgMSvcmTeySksOJ4o6HZjSrQquuoI+yEeozA7v5u2h/sgYfhU7RoT
tsftoylVVAA7fhSht514VDYH1pfjiHlSRgTNSonUbyEDeqipGuF988QQopC5YLtC
DTS14xbd6dPcBfm1Ozgofj7OoHukZ9DTpuCIfAoymY7BalP67kGgbVtxB5BTl7rs
zRsgFcb5AGew7VczLyB9daeyCnSOnvc1rRoH1UVjhrdmg767HFxCZOrkCpR1IDV6
GqP7Eb285DncRNWEMbw/rYG4p7EhQHdyB4SxKB6xcB0+d5FdmyR42Uy+3MLDWaAP
emY/ByOD9Fq1Do5WV3td5dNRZMMzxuMBlgQLHN4ZVeycBAX1BLEqxzo83ijyrnEZ
igCVxgEiDDCT3M+jLK8Ol+yC4aVDieo5YJWNCOH/104k/NCBYYP+nSi5S4jxJdzD
q6FGo6p/4sePXTD/XTcskGPfJQUIMMN2cj128JSWWAnAfQqu9DgXCZsd2BitqXQd
nuiUcyXZu5afZbA50iwHUZ5ST9Qatnv9B5jQX6i7W+t7X84FujyX47iANKF23NJc
T5S4++VqAV7hdGXsJPZjVY0tQP9ulBjApL8O/pyWwuSaEQkREbs7MNAiraYpbadQ
o+9MQBWACtibiB5QArIXTQQph8OzpShmPnzJP8Apn7PipiDo9vEmWxMvExfQNT3b
6drfWcDyVTY1fQ44YBRsdj2HQT5KYK5pWiaq3lMTommoy/32hKKP9Nu7kVM1/yTO
PDScNcWKProfTPbhTJ3sgJYsDidzz8pEk47Yd0b4pSPLzYDWHorG3fwBV4wwC4PM
nMT0K8YFBmmbGdUY006j0yKfpWN3OkmNtp+sI4xdvQc3iYvqABMjE+sQ2GDuOj6C
aoJmObPlgKh5WhF3M67p8/PEl97RwUlI+DD4DT8urHJk716OqQN5WHHD8W9p49gk
WrM91A7iolqd0v2vGIH8//2oZ2mfvj4rltGusqsGZKzZFobIjWqlIy+jXl0t59Eu
SLGICfgJFJBELU4ygbU/9m85Xha6aPTA4iK9EN/o1DtY384VQsvS/5EAgs9uP4gj
wlLc4qGc9CHwTTX3ZYMeVJaKVVNTgSRGXW+qadgEN3tRbUZTcPDXWOur1hbnwzxB
UwIYDWe7CDbhP6Zo2Ew4eruhjIHYKrDUJ8fIdNTXLe+5mxNr7lrUS1voLxpVjjoF
KN2ZQqdgPEVMsDb0Ybz5dr2MK0y5MQYTI4zu87ctvAXfOFJNclrEYH5yeD04UXG/
vfE6zaE5GYs+LxfHLqBtrAKebUBJ5QBbZ2iU1xWPGyLeaQiF7+q+O8FMdnA+WvGC
5o/5oDuqJU7jQgaeIVWtjXRuOQCBq1a/Qr/Hocu7tvHGuwG7UQZijOzITamdZXG8
bpYpFkQYr0C1a3NtfnZIDCO8sO62LW0zSA5Ly/Z9PnW+H6SIKY3QRoDX/fR4zSOz
QWZKtrL0AFbDHL4RjKynI7cKXxdzHSsqbwN/Epe4SVcKx8dY8hFzmnW95HqsrJAb
NjPTOrvkicryZ5V/5NDFCcJaGWn/6euR6F7S+X6FBprBavB43YzfBMRb6eJr4BZq
XP8fRq8TZT1ehvXyT8EOwfGJ1s8i0WqkJjybeh7RpEjlXKjrMA2ARUn67j/I8uY5
+PUIkBzHjLzW0McX2IeGAwfgCbFran4fdHE0IGIvIVnCXDIn2lzdtlAJZE4PCSIO
jkN+iR5aLIzwB1bJvuysAlXTQXMzwB2A0YoNc0j+bACPpJjYVAFnG3FLFp+H6xev
6mz8/XzDNp+GUXQmA6Bda0/mlBOmet0rpHU3xsdo45B9+qj9BhsxivS8649RpW0t
FMvodqKmDRBreAKwWd54mjT3BAIKSg3XCrxVsbX/HvAFR/r6pWU8x6MZFkPHBRyS
hGh3iKQr1HxA4s8wIhg2yFKtNsFA0AwwqXRVCbGvQ3/poqHwz+j67jr8h5U8LwfU
GIJp0tXwyC+webSG3S+6CWUZHfhE45vFwk1MK8GH4dCxrLaiYgmrE2t7e70pliva
DZBjBXU8aa9rG2KMiPjoQotK5GEXfRWp2zY8PzYjLdx+2amGIpOs7O95j+TSCxK2
teFU9YVMgwIIdlQ2/dvsBXhLr54oXXwmc1hZ4EW7dlf8m5pvYyuAANyiwuT0X/Cl
NLBaEJ61ryiRccMPWZ/8KS/hz+NwddqOWXU0xojvqTvwRHZxzVH5epcGQMOMv34v
OPBKh55HrrhIkHwO2dauNHGY64X6ZM4wSgmBxpI5M6Oww6Ept10ULPRueccGb78Z
RXqd9H9m1rz8QvSFTCZ2n9HDdHI2kLchESXtPgnDOU6VhVh/sjXbtkxRSniBWL0A
EGsjc7H1xgqHkLMNDy7g9bjI77C7GjdvFnM5qUvAgfONZY0RbzOOpicIG0iRsA40
URyxj7906+g+AWzjeF4HYQg3rrIojXL690pF4aGDoETPxVnl4DyeYhau7kItVjWI
9AA5G1/n4pXjw4DnFTaCeoi/uUvwP0q/Oy8CZmKUAgLgqVTXwnavGvi+gx8NwKtF
b9B747Q/7A9XPDrXg9TITY2mB3zgx3xS8u+yfh4zIr8U9swldrkPfNdhXJtm+B1Q
PcmqxMdNpqOqeIM1ONMq+bhx2F4q4GmbcASaVH1fsDbYnnNxe2cgYVJIiFY0FIH7
TtK5Kfr7LuPo4XYNDtg6AC8EMCMF97ApTHus9+1SdJxeAM7KAAeg+swKbJmFoCsl
8lTIUn2dZ1RZrRsg2SZTepZnAgVc5NUVJlxSpzW7D6JU5QYIOikdqiPheTvVOzvX
15SQl//BZFb5/a3FPc3WPMJuDt+PVKYMRRXziUUl3wvEpBZ5Mez9eQ/EinanJUAS
jVBm5YMZvGXxabMyZvqUKf5e2cwTkctgAKAKexXYm+Vvb2Ighjjt7F30xlqj/GyT
N5UvjO9lU7PX44flEeTtgr6Tns+nld4k9gUPnMtL9jT3NkH1x7O/6s17Hejli3od
B5GecORoo5sn+wcbdRzmNjE2DHMQx5P1MozfqxcrUOqrZT5OGAqcGBzYSzSyIi87
cUDCwSaUSAz66X+xo5b7Yo9oYNdS46jesRELG7aw0q0m/PuuVTSuyU/EbENau9ew
KHwjKdc9pcBw6BVFFo/1XCRtvLGn6DR2LQWxZeA8WlwfoHDM/hDNlwRAA77WIuwT
XZ0lffQlaVHL72tPooj6aWX9IC6Z89kdc9vVxOtFvqIyrDl4CSjM3AerKsv7w1FM
+0cPM1z56FdRLmYySnQP4ZkOuv1RK44t49tniWfM1IYVGpbRh/x/x9QoHtrrWg62
FN2cHYKINwoEDmU/c4i6MuneVqfuD2Sntz8IXmB4/uBFPM+X5CVwQfggmuBKZAdB
T/tqL7In5rnDi0+EPhux6S0sGcTxmbLrrxOLf5ddAeMshT+IDR3YloGKRM2awMLy
BAVI4HqLv7FZhU4XZQBiy3892LPVpmKfXHZDDYpgARQqD8JceE1Thgd3/Lt1c050
Zn3nZGr31+bgzXpaHASUAC+6RsEi9Fz6HOKBq8cVGc/aOMiAP7yxtjfGRIC7CRpe
KJ9J0IoFGHONikzyHWAhA+7nhvWYwGF4VzRYPqx+yr6ZxavknXN7hSbQc9DWYaHD
JL5az2hL8oTBihQ53Ee76FEStpdsT+xPzhZrJa0rd0/r4ClqKP4y3ZjJexPISypQ
fWNinSV67eEUUoAIIOOX7RhIU9lWZ6tal3sCz6uxUob+1ONLJO+kNcHAtWH1RhUw
jba2ocFIsseY0y6c6Yi6qcKx80diPf72yGvvXr8iUX2gX06w5aC4XZbui2HT9Dwb
GyjyqYDqXHtB4PwkyVMJLcdtl786HqJ9kXpKrdEArjR/WD85egnK9t+qtoYp05B+
8dHs38p0Y3jDc1ohDwjotzS24VhSQM1heCn+J9KDI8+Gj7xTmHXXa1g1tJKfEM5n
ojCM5IMO02Rn2RrheNfFUgCTueV7ssepIdo+40YFXlipkxneSq5afx6U2CY5mnJK
uyM2TYKnYxys84VynSJweBz4ylYAQkuX7mCJCxNsTl3aDknSZRHEdy53AWyb9kPO
06qCMubE0hig5gYaqCXZXVQiBUW3CrSupLFcAczCFjIKR3Edr8L6HXxGyBpd2rH3
ggAz0IsdA+HLKF1nbenXevwHUCa1J4nC4b6no3QDnb2oKtWrfwVvjvnXgyIuXTlq
cDEBKigBpZ9A5VE2HgIVfyUjKBrruB/pwIAEIpfb5+iz0W1aHZJK1H/Y2xhrv0Yw
N7lojZsI5/OQlAdMRqmNZ5fP09r2B31/vIF1p2zqjPtlSjvRS8H3DkglBm8MPzt1
oeVpnDK0YGplNhmonGEHcmuX5FIhaE68QTKTXs4Cx1Waj6b2HGsr/Wk5ymc7FzyT
fDupBvhLbuBscjepF7VLSDkCdkDgzL5DNYXSry2nxifVKdCY6w1y3u4aKyBu3jBz
exD74inAzXh7EybFfLqhPLmq6bhpUMXjU7SbO5MaDf3ucVnDmJLzCWlVS32WxaHM
/0mguoRGiqY3LM26AL0M5iiuW3e4g9TBAIqZME6sofV7yQK5XkUldEBZdWyXenX0
gxLlShqSkqe8EhUsV/WoTfajXHQ8rwG0ShrRYEDAITgbn/ZUw4NIlRIAzNrMAxl7
1B0h4dWuFwcO0I6dSvVBadR6pUBg4GGdlpO6EDkZ1m5dGhytekTG3XtyhhYruuOC
x1GYdpP2LzrPVuB8YU+yC7m11xqRdkWJNj9m29XmdInRKFa0YdzjAYMXiATehAiZ
HlptHV8DHHfwB9ZoVI9QIrV9SBhZz+ilOHlsM6yp0UK7iosmjKNkYjrlxpG3VEDq
9EM6vcciDcMp5YXdqkgsDV4ply29mlKwJcwLmFs270NoptbkgRzHuC7/HBn07ICV
SMLBlBsdURhMUoPnJYCr94Qp3bs6Ba0lcWnQmCNtwsVjj+XYTYroedCsbZRHvdjt
aGrM8nte2whU1vSQa6QB9gltNLPJFdSJP27uqVaGOosm8RyPYwdTQHb/m2i01nPB
AfYu0iLHVCIizjMZLa9ga7Drz8mQCzqm7jLbpGJQ3YzD0x5xx/ofoa7V/nkfS6lg
yBsF+gQ+/VzL8NGWXAY0LWDdTMjnhr8h/7JPEHbLKWZFvONmDsQAEe3qi1z/zAj0
LxxMW17p6TeyR5iReJgW5b6yyU45dnC/FctiR9m8lV5OFCJsMcuKK4aAeNVlE8S5
v7/zVojwygknRmOkbqoWiogy0TuvpEvINNuQFUt161dAuTUj3e+SjXIm2djCQlJC
eTVvt2CsnWShDWCo6u8uV9tB9HDVi7qQgYo6UXQYA6yRfPIKBs9jY63NH+2TA/9h
FQg2EkFzkkP74maxWL0HktOjZyNnBQVYykdX7d1j43GTt2OCUIGd2QgnDzaiCcUj
lpRqieYZDZZAhP4NU9gXtlu5cyrKacneiaCm4nJpoeOcfZqyVClKTOjvGPCjlwbm
MB1GcKBf920CHf0PVD6NjT3ULNVRdhH9M7oSE0vrzEjM0lZw3RMVW6uqiUGpVx/u
T7Ciqvqub+HWyX5eq1vpgOamiIlTxMDypC8OXcDC2L6uhIK/tGCyaPVckdrT7/ha
atTFu7lytFclt0kmYz/L3GSxol1RaQTBa+0vs5VQQasf5nsIQhKYMC9M9VlJ0i6o
iRwYGPCo/a353h/kb8banSFpDTfVN6rtI7A6oFUik2KyFceNEWE3QAs3ciufcp+T
CdRwFbNv7Gpq8uP3Icpi0be9plXc1y/3s1iNKnlw1EeuqXh7L4suamoFG/pQCrjU
TjeAazPxGEz5/t0WRzihyPKZkwIsfGR3r/IHPXIG2g/NWrsaXYWfQT6+hccq7S6y
ej3g4qLSeDdWqu4oMVBWXuC0D7OcDGL2q3xI/6CQ8O2Ut+j1Tr/jne6Mhg9kMnY/
i/YPLM7UhgeHExm3B7hwrkxwIv/1HhHArKGwI/hBYFEPqu8vHjZrHV8T399RiC06
5ZjXWIisOtnxB7CRxtrbpKQ2P/RIvoCozHZZ3shrdBlj26pGAWREVBOHycR95lP4
rdI+3M56tJnJcQudLyi8/ubCTDPDiC3SO/26+6d9SyWjc/LM0iOKdTx3oGhsIVdO
nfGtW5jPn712pKIpbrN3HXaABeo5G+4G4GTwtNYLyJgecnuPgoTJ4KBakUS1BN9b
8AqfYv0uzrZYLB5P1JpEDbfKNfEmzJIL/Clv/X/Re4CoLgcYLIMX6a3FmRfCEpIn
HjA5uAPp2dt+eHp2q/fuZbtA5qtO0w4TaI5aVWNzSlg3X+u2AfmEaO6IMe8xM1eT
37dF6wA7wKy+wJxwAYclJuRNFTbAIgg6eF4niH58FZGv022rrRrpxXWSObt0TixF
bx/hTvkyj/AtQemGwS1pFpzaiO8/xT5kgNGVjyxW3i/98o0Gi52C8PMCOqHAjFwE
QjZFRwVTpspZT7aveRbMbOr0eDHs+uXlJDseri8WL6C/lUieAV6v4AHsLj0TDihC
wa1HzwaL8Tj5LxFzXSEihzYYgRR3nDI3be5AyLv3pIadR9a7RWojmnwsaKGzxKqi
9mwPtWOQWQ1kcDYV3KoJ7X88JM81S7xdxvmXZE5oWf2uRRodz0v54FxjXdos37S9
KB5K33nSKkjV7pDtADH9V+cu1YAKy6AFWL2wpYRo9t8r+00hEzIx7swBQea70EGZ
DSYKxhB4ppPPVnHFeI0ZSegLvzt9Cx304fGZ+opAE2z7hmjgBQ6WaqpLSc6EA4tG
wj3ukCms0eM+OWb3uEwMdfPKBBZ0zqJMZwPcwCUWPbFrHZcQvuwOPZ6k0immf1r4
YIoCanK+z54s35r7M1bhusuyQKMVGceX/+SBHirF13Cn3v1lOK0mrgxJMOBtMbsr
Fmxhs8j32+24a8+GxKkj8sbzG5EHzBrg4KpcdvxDcp2qeKEKYfYH5aw06Np2QW8l
oPd9s3g4izkWGaCCwKzjfsDpaw7rcAGxYMBIbc0kWbnBipLCpd1YCO7OTKqTrV2B
uwU7CSHYFltKaBGIKPAnw8AMLT/j9T8QNzevfqbVgw7+2Wt5Q7u33eSf4e7wo9G2
iPLQpN1g9JqUZc//TCy74NNmu/uTGZCT2iQNUNOzRecFghYEWNm81ST1ke1Pm9m3
SSR+apiHLvU5xZ+eUfEWJOuTMKPRc5K85XfA+uS7JLA8gNVBCpXnjd5zooIxMd9J
6UBQxTzQCIGEmW4bmbb74J38XTllG0JI049GnAkbk6ZkPr2Duj3gkDkHpDcV4zrE
Jk99iqbekQ4tOVWrA56TDnkS/NxOXVz5iayH8WGJ7yUUOXAeukAT9gnvXYvqhkPf
0vGfl1VzGmBsQ6HgRBC+3SiuZjjO7Z3tX2LxjMt0z4DffkzBgy2KGpLNlJiF5D9j
oKroK3+2W1aoC5vgEqezeRmjHq/4YoPZW3jnew466nOttNc1SnOEBszrVKhWXwBW
6NkUSQtBcNrO5cnEpKKZQZnj4z+RX0ieiT+1fxCmXS/9UrHAcj8Hyg4kDRYKBBxH
qmyi79TksxO03zjd9GKnzNz5x0UJ+6xSIp2+N0DmUhPvZDuau+av0dOx7HvuDyob
nS+U4nyy1eqmiFFf1GizNaQ5eN9rbzIsxllhFMVSZ7sVYEFmtXvDVl+vqOuIqUZD
VfLHpSMMQ/NI3nrRWqpcE2VQTP48IZcVtsGxbub93tTaPtCffysRPGCCGLwsJltz
aYclaJYd2ZYpLd1TGyb8Q0Fa5Y8ql9qQM4O9/E0TaaD0G9b7xu9Zb73krghL9J9C
vCDPWrncDjvDkGpyyqpiAgTf5FGqwWw4InYgEixWx3zVvYv3WDlGVaaGh4gqD1Oz
pOXy58X6UXwO2SLgrEWPw9IRqdD7jtnFnykJ9zJywsUr8mOm3vE/0PhfiZYSwAju
H4rHZwTgE0IIOoX40ROcmoeLhtbwrYXkAJTrwJw0w67VgP8JszfTujkabVSpE2qX
/Q1D2kKXDR2D1rRuhxaZ3FOfiND2VmEyyEd4pWZ+pyR7Cyt1ZStEmHzYDoUaVVPV
608JPsNSXrh/yDCeXsFR1sh6tGXY9bjeoltY6yNy1ivtREHGMMMdWUaFVJNPYB6K
0KKZsOjvx8Y34DpEasWjazarw7JoiRI/nWxTdFtgZKnybwqy752W/52yXuJqnIZK
E7RIEK7VIJd/kqsu0HX1I9/+oInKICRrMizQQCRt6PcfNKxypgNOn5KWv/dRwrl1
VpUK9trUeToWOgYXrWP8Wce7UcnjzucZ9I8XjY/H3UMl/virAkW2SoW3t77UUO9i
3zk28hFrMk2Dau3GNPnfcatybkVBQ0gF76qavybptVtGXBRCO/m4dvz565dsledr
U+uSRwOe7qK8fG7s9aKoEw9HS4H1nbGusuI5aZBwN1iZfZ1xIxBO6uoZTrDBCbx+
dkb9jm7fYFP0IQKH3yKeL1/oQndlxBqd2ZA2y6E9BOQBPcPPbDixjHzsd3KSiyWg
WFnk60MHg174kbr+BX587XV2xEyDWCEICnrtZiM4JbWJxmeUYV45hgQmni7GgLud
eg1qdVxLP2iZsaq8DJnTeowcs2o35NRhw/2WNIha6xAMr29qWVY5mlubg9X5173X
BXNVbvEgYskP3zUJSZwqbXj2TLF9MqeQhZsLZCnO19josFQyxOMguouTZnss2/qr
spmD6S9S1O1YeIiHnSLehZHioRGDk5188xjeKKHPmcYqGutHiRhG5sAU7SlGfpLy
ygIeTBR+SisfhVAjECti0a0lZQ6SBZrplMonRUHhF7tUE63gCH2mv4rSfMPTqD6H
NxfwiJ9O4l4Kh4bFgVloSYqciUGd5znTKYeBcjt89zDRR/2Dln9x3VcOlNi1VLJ8
jhHfs3ukzjNAJb32lqgYU5W8n7iMDZY4a/UMecq2dhBGsVp6yr1IOo/u5uWKvUiV
dmveRb/LSI4AW/4gkZHcjkD/bOobxaNQ3vHYvpYuQdiUmH4l22tz6icjK+wyiCcx
Ap7d6TFWOvB7dlzeAG8EkUFlBU2vdzUu1pfWEZnMpSZhBPLXO+XFIFaq6dTsR+Ba
mj56csy5K45Duj+4JBogjHWfvM9BCS6O5DrAsx3ZjmDzsUVla+gg53ju9VVi23Qa
z98XJ5679wWXTECg0fTpz0ZGi7uMHuswBH8qn1Yos/jIB2bAXoX6iTc6MQ+kRqQA
gROUizR4+qSFvKoek/3UCq4Rv4CKUarMYkWQPAd0CTbYqVQ8N6NUjhpExAiATwTu
9ENLN4LojpKYwTO+5ZzqdpRak6wyJC/2t0S2Lg4BMnzEK36Mi/j2qFmuzZH+JZtf
30Op2hjE3sfRlztwsNVimfGaHI7Z1UQmxo7YarkY+hr1OaQyWqqCeibqXbcfl9Y3
2rvxX9gzsNzlGkRrqIt/xs44X55OF/h8jAxJF+DkkSdepQrNBOkAywBMAR/ynOaF
RpGNzRZKw//H6yKiTaAIwHAA1ezj1SCmlVdJ6UBXbJC2WhlK1J0oZKSMdckKGnaT
iehiwYSRWIaPvhGkdWUk5eiot02SXUDEYaE0CaHbTziEbDhLAmBeaML0p2EdwJsA
iiY7ND7H53sQRgxCjpTepMSV6/SgNgGYZjQOxp3Iy5MzEPxz/LHcEupYKXAjE5Tv
IbL/dDeAPyoqJ9eLLVqOw+lOK0wi/sSRvCiCAKO3Sf0K5mZs5dlaQJQF5rvAh7RX
DsbzxQqrULeWZXree++BmvKBPOX+XzOO4ZCTI68yLUqfhkeKQbtvrDZXh2gq0nJv
xUy/uFRRlbirBLWNjvsAK3nlvsXpZ00CUiXiSW19Aeo8Ek6Rs2s68IPLM12o0qPA
Nx7f2ZTnJMtLzPwRb29N10tnh4bTLXVa5zAC6K9dyuBclhlHp0lL85J7YMVN75Z4
sZ0Q5D6AptpnlYGdR43tdeE2Pec77EsFWkm3aAAIE/t1tPuAY5uYOrK5VLea1axP
Me8yuAGycbxNZBHss4PosijTBD053GiVAHIG3ZQvgXP/K4fL8NbuFmMCkCnU3hNz
b8cAfQBYOkXzO2cVZ79I1/ARMuQty19L0RxbOgnikr/5ca0RTXhatYNWq7qn7fCs
JqGLtq6/wq0s0BJnFTXBYa6CER4QtSVrLINoctqlea4CXm4wMuM+ie7H3K+I2NUN
tYXwf8APtCPDXLQbXAUcnBH968VhWcghCVF+FG7/zaibyMqlDuGN/TcXHDsnU417
U6YqXmwmAyheIN6Z+Pa6be4Xy7jpx1R4xnDHeKHlfTh8NDuoK9sgnD+upFNz//z/
ffvrn+SrikkJe9G/QQHjDH744OxEIHtPDtvCLlmLaVKxHqsXZKb4QZFFKpz+06SE
2d0MpHIfBcJcT0Mey8e+YL+pFyAH8rdH1/SSakiHnSDSzL5yWN4HAabZ6ieVnXFs
IZiyV3l3v7d6scpgC/xja1xF+ewtEbNuP+7ufcM95Gizzs+QJsT8STgMyV30BUEu
MZraxGfEDK8p9R5iWSodbbRef8/PVHZQwV4CNrfwZ5CBoVhcl1hsnf83c969sdHK
xl5h0jcl4zd0/Uz9V5hyJWnAgTT7C6flOSF5R0WI9kQBoWy07KKvxJPsKP3r89Tt
X6Vwzlo4iQ2Zcp/mBDRG4dH7oZ1Vr2vRJ9gUDb2L65qt+is3DLNR8h0vTcR0DFLJ
H1l/XmC7+1C8z7QdiZxOojh3f35vSVl1Lb210leR3U91Wgt3Rri3WISua4QxwIsk
HpeSGazaklUahNl7hbf1KDLrx86n9SgIOcyGhnXKIk+KmuCx8UoESE31Avz6UlB2
tN+0xmA8ufsUmxAO7Q5lvZ3QeM19Bz9O+Ah+7sVN5Dba/c9kcoS0cqce8X+8nCh1
Dy4vnoyzUz2GQi4Wzf/NJegzFSAvs270nUEBR2/gZy6NYNfsd1U/1EpJxSBsbagx
EVQsQfR01BArmk6oOPpTaAyetBT7uyH1k5HiD3AF+qNb73+FOG3f9T5T1VtPJ1Bd
Yx5WidiHv6C54pIIusnyksns0bQ84VqcQf5tL2gk9AV01KZjYAssbLx5K1Ngye2O
yAO1eZFRBUIpHwD3NLUMo5i86EL0s35g0lTf+5XCWAMqFCyiO51RJ73EKG7z9Z8w
Jmo86EP6oJtNKTRWxtVBNnbH/uZZ9lL53JFctL/n5+hFcrNRz+Br2k7JVV239aEZ
Btvr7EBIAZieks4jl851kYvl2Tt4jRKcraym9smyhmUV75YdH7RBJTPog/vZU42t
u6hRj5kQ8ZTA9xjREm9BINoySggaIh2Z8N2qS9Ylfi3gjzdVyAPB7nlp59TuW6dI
Ef+9cbvas+bVzJb2z4RBqNQRoy7bucYbXNQKyGF0pF294dkb+qSG5gbl9Us7Myqn
WOjoHVqN5n61e2r1Q1dMpv9flX5psBAYMM2Y+P0FPAydP+ZoXJQXpg/LLQCKg5gy
zqe2nWF9vHWF3iiX8XoNvVeZjB4T4IbRkJs6hd1q3rKPF2tBIlX3nikkRie+zNfa
d43+zxEd34uBXa57mU2/LQ37BKdFB6kEaRpx5x25yNklkSjqxCQwqi4vHg9SE/4g
aFyxd0x1zHKgcum8cONcDeOezU1sPIhmqAUcUjP1Bhy2M71ywm1kad5jRNiWFSkU
6lY0HiXW66Zx3mAFe2xOpCFmjOIuDP2t2BCEaKQGgceKBjuzeCgLpTpU7ia5WptW
aNlkbmAGKeZM2Z/U+Q5h6huoXGwnUtVvFh6+G5P64rbY+5iGc1IJ8x5iu5946gvP
MieD1vmvIAO+rfgSPLpJxg+oOxNks6e/e7OYeOev4JkJTMuP1jPJgHl/8AQ3vkYd
Lt9g/nPviTHtV/hMJd8NRFZ010O2qdKCWAFxNjQCFEkIpBynFHKGPIkRWJ0gegVK
uNkWdsRqCfvqtwLgq/3PE7AjBjXmBTra9GeYGpWQS6dZ5eFq1L4frvodpNwPs2wM
rWTqfAcDR7AhcKbqrv+yUZGs9/rc5gzwxUgg7LXbxcB/NxuYkOincpH9zNlr8D4W
UKMWE8DY2UNh5hITd2VFyBocc+3W/3/TNlSjja1jPCMXXzL9PZQbK6rcMdvonl5I
Dc3aAMlAP9sHK1Ijk2WeqKUSIntHSWwlImKdAYhYDTbXRs/JRIzeO/deNIIjew0M
OLCkhH/1LHguP3EFPXj0ZKEpR8MVNuOC1CtHFwOpcr81IzRY+ZWwV406BeYhclat
XUm99TLa2s1j+XiHiiWW71auGl1OsgfRBSyB7N6+ARd78ivkRextJh4w3tHmGreF
8ypvEy+itbTvievtLVTmYZ/6Wq0pkY+iL40HC9/bBnU9XORgLN5efqO5L04WGBxm
WsDS9b3019pYJO9KSMzyJfV4wQdFOJzrIFgI09SmH2UwjJ5wRqkqbCwsqxfCSEIm
onp6+Lkxrljbv1AelteO+ZAddnU7mfgpzSgjYMEE4e/sHeVoCRpBojJyXzIvoRK5
EJcL9fiR1/mCn9BPeYCMw0olQl6lwFksUHl7vk1M1qvxHSeZBwAQNaDeXnCdr7W5
1RfZCnQ1B03lvvtPGmDZs04HNP9x6/5FOM/0rU5n4nUpCSb6bxQbk/3WUyIpNrUs
E9L+3OZmxUl69LrLQN8BcpFb+tgWOvVSkjdiHqmau1xUh4OVsb6BFkldAh8hdeHh
/Gs+E60Uw8mmHZSf2c68JOjbYQN2O/8Ov69tmDkgX7aZ8uI43dzDfBlDg/RtcQGl
fTPk1RL/RfIkLg0hJlSECgnPYhCWJaf9ku8IvdCDgTRqo61mG0+NPTGGvqSPOwzb
MSXj60e68ydKKBF720RhHhZvvNulo1TuJmJYGhGaidT+koGxXq31Qg7Ra2XQx752
Gx+PqZ3OKyO4BKVsnO+V2Ki9HYrut+7Af/GbXkhb/rIFX9YDD7tjZ8TfKGP796L6
M2bsiAfRK7v8gCHxxCwbTgcn4lFNQ5I48VYaqjd8/a/n6I/pAx7hKvSEw7k0t+rb
yMs9Roq11PKTVlTNLoxuh61zyyLovwluH07x+3t0eZNlVYNvCycYyC4iPR/TKthn
8kUNECqfTqSIQP6tdrO/o4a8nlyaS9Zs6qe2AYc78E9bnPqs7EVkJ8Dr3X+foHoN
BtrGgMHAUxBw4KqsOKC7Tjt6cNOQSczs4/Wasa5OklYDD7bxK1Pmd4t4J7Upp6iC
jtV2Y5EkXrnORZNg++tw94jLfnfr/f4umFfSYFxp8FgbbBRq7al+G+NMB6XlakMT
3c5q/7mpjo9w+Hmu9fR+g9srGS4j+ly7eiGUvAV3trJg8wXJJET/CyVtQM7upql1
RGNjngFq1A1cGAKMx8Vlw/gCzSkCSzw6+KXq3yzHgECgAm0vUmoHDee7TbwV6v5Y
j88M9h3Hh2Dc0+VoCaNKjZnJlkeeL17iglOBN+1/pSB0IkIYaSYFZYGCYaFhug9w
xDkz9RiSbG/AqYm2nou8UIenFAM57TztTKe1C9Afz6U8AtKULRdjSlHaYhUdDvg+
3zkY0/JCMcECj73UHyPGtAojkBcpbfSev9LcPieEmIPAZfAYLLXvAXZ/ZfssAc3d
rep1WhkXa7tOHp8U4SlYlyvQB6VcOJykQ0POwkHxSL7FfwSdt2p0Dcq/JvMYecSx
NpKgSTPT5MGJvgR+dehqT+Vj1lrGyME35UABW90stkK+qvbvWEO8/anObty2M4z7
wRlugwUdr+PT8vyZRGsSgPaaJB3/60qme+kWbcAJzFopKZoTwFwdIWzED31SM/N9
RA9fGdPEvTkVWPyd+Am7oGNoC6O+q2p66HKOc8VPdLRwn2zpGi7Jf5UaV9hiBi5w
DB/s2zuvJI8s6sGnVag+BTwX7uEsU5vdOjtNsEfQSPJ+K8OtOulIj8Cr+NLNRSR6
HSilMtwY4HSTu2ndrAMJHMSH1ulUU0OMeKcQRg+iJj/QXtIvcQ07k7t3ySYQe/lB
O0flUGemCFcIZeyYAmaG5ceHJg0SpW+gIewky66JzcXUUHxz6wetpfzO5biz+Ewv
+tOD3htPND1Dd1JQz6BOZCroH92l+uOHZX5pZMT57JWieMaz3vgD/C8sBgR/Tz5I
9ocnUxp5o3KYXdC5D8ukKuMUmlywjnMhwSgvVZcbQ8ozBMBypdpZkjJB7X7GJ6XB
y02IeyK48av5ul7mCd9whDZ0FLiC8FmybrEKioKcI1cr5rfrRL3AOdtPc7lgCGg7
o3qqdRuZLUrqyx07tD0AfqDJ4GNexDPTNq/nv6uLvjABt9iv56G48IiORQImnrGb
cHHXyk2TDXXsjMy6C/+L5RBX3lpA5A3XehzKZsxIo3Hh2FGz0JTRrTAFSaIWi+O/
hEYm/6M2yijanIhrJ3kmDc2OwMusNL7AUp8kpBStOe61AkDKqSdXvEVEKv8WYQp9
GuVFByGJZqsRkIKpTBpPsces/0l+9lu+fRmCSg7QjqWI6XE9cr4te6JGfQ5Tlum4
Om6QHdB64OekQOVuAHW/EI1oZ6xQwVWf/IX35L2Sfe952rpQkHwEJDeyd48kArx7
MKriNul0nVj+ao6uc1p+cda2e1qPe6YvU9AiVlwrbEcjkYtUviW5hMDzqz4oUHS9
lLRJUsXRyTTCMuBnrQjEAFH7RjztsB8Z8az+hQdLvKVQxZz4w79IGH1P8JUOkXQE
RAZXgz8CI0J7tIigjoHxNRCduEjvCnKEBzUHJU7PjjX1NK87l3es/p7NlBBh0dVj
JZa8m63XpAv8U3NwLKUIJDJsOnKHC5ObAvJ6HLgot4joMmhbemNeWpfl6e/1zM3c
QeEPs7U4AQ5YTR9rBZ/45ELD2gpGBvlA4MCHWN0xzne5aBoysj6OB+w/yaAQ3iJw
AV0OYM9t799gaDSTgTDDUq4v6sC3AYmP244eGK4oD5oYBAKNuTeVxz0GUQ4lKA1c
DKk4BqxXKZcPLUTLA5g59Xvzs8nqEjdufj+U8lWMbCcHyEuQW5zkaNatnfKmk+pu
yEPRt7FO8cpR47eWGo5SP4z8cI2EyRZUEKHs4qeW3PZ1YjB1WzlEI8k+2zbvjm9i
EiVNVhSfUX5gToPsEttcxyFlA0mzp5i11hcoKxUrrx/RzedsUzN/fukydpp43kef
kXM3lXnvKOo2HqURMWdtRqATGfk85xf29WU2pRvIcojPHqax5P5vqX10KT558GOn
1jogp43ukgSRvC4wZImfK26XmG/x4A+ncJb3B0gTwMAWiaxMw4/Og7Har1PE7TO8
iK3CEtTTwKUf6f7LCX84zTFFoeaCSuouMikRYwSfhwBSJkBsFyGX8x6VDwAcIAN8
0pwW1tMu/BzsYdegoIxyYWiJGeWMNamawf81s1Q7pUw3LxFPQCw+r9SWmoMxQO6c
YWAABCNDQjUfUW+MatubkhFqzzuuRiIhmdLvZnx6FDTP1vTaQiu6rusyJdbqE7Ue
snLDH3aE1Ojq95lhRRhkSro3Cyy6tuwDeQya5HQV0EltBaUY4EH+c0RAAyvgEsNV
xMbl5A4vVGd8AoQV0XyhswfrkFsQDeXV3jP4Wt1zU8y3ezVKyyrOENgu4eSrYrsr
9W7Z6a+n7P37gq7bY6v/3GoywduYJLRH+rFdeyQuMhaqidYDHQRT1BE/VkhXL2fj
TpcFejDefBJchjRweVDyyaO4QX1D7nGsehN0uS6s04s7fv+xgoayDwIH7ZlsEmQu
CICRMYBhdRTNBlb2epeUKxIIpBvPLtip1tDD/zcCQy7LQIhio+uBPcgBLfDHdzkl
or/dW90wREb4egdli194MRLl0G6VjXIExRsgTqm8QnUdihwV3MA0ws4uegRkHbcH
ZrqIRFOFHlhJENE5r5FotsR3E8Q8J/AUZXo3prel2zYeSPlUstkO0s/o4Y5kWeiI
EpNSUdJ9pNEmf/CbZow9JDDQpkIuJrkZ7qNfNVUc+tYk2tmDlQknkvNZLaxRZ92G
4qoa4h2yX8YQGqlSlLKJQhbD6U2G/RCv+n4D1HgpVtZRHAiVUF2MQEwZ9RvYaces
+/IRuicfzBWXhYALDvoFSqELu/EHhUEVBxLRASGmN89cloqbHd2/iohxwzBwfo+Q
EEXcu8JF1XPPumUso2yu2ci2LlHzN3eeLOPAWXi1vLFNOiftS9ebGi0oLVv47Gef
hDja25YBiFXmIHZ0Opg5SaaKZOS4F3liovzhZvXGDW12ywMKvkTVYy6scjvgk5SU
g2S++GMJTFX+PyF2x4MmCLzHo42diPi2gI0FJaBpP129/rf1zwuXnrmgqVECFuKw
ZS2woms5x+IYW0QVVvyHLzXaf04z3tR4LstTBdcMWFbKTj7/g1YGoEzBXlP6gcbt
ExlnN2voyxp/1HEs9zrpTllys/Rg5A04cRqmWOSeD0u3DqcuP1X0qoQSMZfDje1E
5NcEsOU9vP7EO1Qk7T5nkXm5dGdGUT70qEf3FQWD2Cik087KVoH0lNpwptI8cQZ1
fTKGyihn0nOJJPoeyo8pv/hzwKDkesVH62sAgGrGAVgxSmMY4VQtCJuc54ERyAWu
XCCquDUK2Q4mTTkUxGkQyW/++4Ox0aNp3tZGC8GgJ16h/X57kHwVmvMJunUtfbvd
1a7Nuf/DRP3scSR/JNRdV2Ep2sw8t3JRC8Vm9nKSTZWzqt9cKevfr1aE9nFaV3yW
eQFcRHo2yhAXvR5x2WgAEh1y+qZV3x55rNIebyOuIcVN23k0jb6otJhImRpZfb7D
LS6/RkRzfaoYIYjQUvhpxVGMuKb+XQUgWlpfL0vPmc0U/scM7ZwMqHVmcqwznKGp
ox/lv0GKKd2ky8hDnSo+mFQyX0d3UXK4AQtVA4RV20/7YpEiYOfbRv5d/MzNM2+h
UaJ82vdCzexjiYCeKRqYiUT/A5OyVFOyJVty6EhWw3QulXk6zUznUQh/gPFVhFSr
O5F/PGUI+8hADtcZ3PZpkwDWyrH2B0z2+ODyLiQf2GQ59I1nDUfi6UhoITmgDX0j
qe3fmdqYlJJu4m1o+clvbjcVR7Wc45mXlcYKDdj30fPRh+8KJN89kiCa6yP1eQtZ
F8vhD6oPb3Z5lI1OwOC3mWx46zFKu54q72kOpL4K2gnIjYPWg8U/NKhlbRs4GVGH
4OCVD50wCLVNYGiL/HtIclETSJb2vPkgdEF4Wsp0F+p6bBLZkUQMHDC0w+BZiypR
wyGnuptGMhsZ2EW3mVsI1SK2Fiwnzex2834tpT6LvLbxPzJaURZtoawpQfnyUlEj
4MIsnpPkG1ef2qLzJLREF6uO7cxzwiaWL377zjpODWUbcXoejGepmoal9CrOdYsB
xzdXXbqr+/n3eeVAz8SzVNn8+XFZX7AbWJax+g127/rJl6QsbRPtT4H86EqISYpg
cSGRH3pfx/2VwNueJ5jNZBYIzVNjRuF72t/ZZjS+e99mMV2j8qWue1q9VYKQgqGM
JICE+sqHiE2q9/1vqXhRbAfykp4EAx63/fk+h9lg4b933vyIJU6ncZB8YIldChzK
jfiYyg6OUMBr55gEv2fePa2IXA9Pbk/TnWvKRGEoBVRIUwZwoJdfWSzDX8Nr9VX4
tNnDI5UMBtzvqi7ZdDfAMq+17lwho8qpC5Ud+pEgflFnk8KwSHrtWJPEpjIjSPYT
0GY8rGujblagA3G7+7RtsWpluckizrGhR6G9Ig5sus5M6USheB3nGcwxXltPtkBc
cSUNBn//Nzwdm16yVrSjY4hX5IqhQDvii1LJIVhusf63cAj9wWE7O6YgsnbbsyqY
pm+4a1UMTKvCxuhUm0QwqVZvAAloNy15o8oYm9H2BtrHEtajJPl7aii9NyBDS3KO
kSzaNyPmmcSDe/t8L0FSugW2OJI1lhIzd12uvlxAounnOtS9PH5iEEg93Jn+JqnI
Wd2keppZTXCBNyS3CeE8ZSMd/JBFseRASDg4LukqVrheBnImAYE9Hxngissb20xJ
1KH8i3vpWLlIvo23HasFeqHl878mo3Fa9ChX9LXbgpKNCv/+Lx9a5Ekd+Xa35twY
PfFSQMY49mrj6pKxZVfVdFS5PyuxFyT0EO4pjO77vLyw68OLrCHzU72OSjeCUFas
h6sShu91kVloFULu6q7r4tq+YW8yqBtgdCfllN1jYwEjZbJXwOkE7O8XO2UuLXeY
9ZcAHgjJlYV3hn+t1/yJ1hCg8FfGRME80x78WNOisIAUzimmV0NzZ0brP94UVX0T
K6S6dbmiGNMa9b4hFyGJrz6an55fN9GNFO968fKxeuHYL3QAp70e1CgIB9BfDfuY
Ck64N6TIfk4KS1bL+2J4jVo0ryfo9JvApUOpwCImji5+qBYOfCjDlynHNfN713c+
9KNBcmn9NEXg515xLmm4/yMAeq1xkqrXgPfxSQGGR+Ob6xH42yZqaRShoJZeo1S2
JojqGYdauw6yo276M1m7N5twJ0f+/iyUzlZVR2ssMRfohES9QzZBYgy11RVKq39D
izCxwwG/X2KpyvfIDbaFr8wQgTo2jn4YScV0LtdFaPYklM/XOTYzJ++HJDRsJUWf
GUk7ruLkbdkL6MKAoPX+6VsPzeboCiY8V79QFarSrn7qwqoDhdXVQ4560p1g61j4
qY0shp30ydX/AceO3jZW+pB1BO5QjDbJKy8d7+GTRhV6X1+W4nFY0QGdTVq66srn
9dPy3ptx/SzzrtzyvZ2fWAlC2duMfOH0jYSJJ9RvUJywZVKF+pXhpBBZ7Lu6xWPd
1A9MMw3jweA9CUd5ffQuyrQM4KNB6zv50fZaIufmaGFgh/m6yYdy5VFA0eRGFNXW
f0mtA4GTWczAVxUW6Sxk2bRG+6G65cZKdqy0JVr8aeYtHUJWswKOxJB6OrrGkDBi
MHHLUHUz/PWrl1IVd4ZcBmRZR2/HvQbTA+QBodslv3BcHPZUFuhtvx9sXHC10Ejf
kaHqgfLUc2DeFDDxn+37M8Id/RdlC2f+mhthfTovEPPa6QadW/s7yywZuEbvSHln
XG1VBhGxHyFrpc/Bqy0tgfu50ogsFgyyefpOemaQs8c9AioknOT+NCxIClmsarlD
49kv67rcsE+rwLCsGZWQtLbkr5TWKhH3mlf+/K3SLEC0BNXFqfDIz96k/R5VeBGA
gJXts+SxZC5E3z1n1x1ChUHJqsaYiQboGK9D2HWV+/IsK2fmaJjL0oX8g4jcC9F0
ISXy6Mfo5F8A9NDmYh6mH2eTkOdmNyi1AcrbxYsW02qXmUQAZ25WdS8ehD2w/knA
RGKZaws5blvutPHcCPlKQVNK2QlgaZT9Q9AnKNDY7NVdnE4RNQc5KK3iPLxH08Xo
GL0YGm34kJbP9pe2wNuWA3hJeLspro+IW6R+eVBP97RdYZmvdx6BJrIlS+j2tiHb
D7lRzEHifmpRSgFyzyMyjtvNyIw3JVj6MExxN4h9dv770kM9vO8ApN7XZoRPgHxD
iqgzvFesu/twAIFfPZyk4nguwmh1NKz882Opbna/r947T55f1ZhAXDBpwHSgf20K
fwa2/Tc1gD3p62Mmw5Q0gJxbu5C561DEueiLaOjXZeJQB2htzg/Ksl84Qo0PeS9z
cA9Dobrjw1m8DM6viCCtoMasZGzvp/nWacXNQnWAjsNdmWznKcNpBBwOB+tfA4sS
nOkkriQSp2K0H5KSxiOkbGSLYmUFvAsJZubVexRQJg9/yOFNXpmRZM7meba3CxqU
DBZqJ9KXg2d9HrJcSVVf3fc4/Ai877IE057bZ/Hr+IJChbj6e79tjf/v1iv2VZIc
jCx9i0XdxAxOJDqSxFRZ0lrymh34/aEJ/+K/7ShzcMz8tSu7rJRze3StnhSQmJ96
NQlCCko03V2RGhGnRmBzdFssRRL7GStgD9BwmD3AO47JnONIq2p+p/tTH+VLaygZ
mquicEbpDzgKPNBWn084R42GG7cn+A+4Sc4Voc5nh7rH6xotBr2eURF2cKRB92f4
8rYSzw6cm+FbtkY9e1qu0xWe5Ig0nXuPWnBZqe4iHAF1eT9Fr3R78z44NGKMsQ/4
pVCtyjstyNTSlYfL76dj5z0EqpJ0Uk/uf1HPuxa151lBCmCRS5XrdZinYceicrBq
HPKztj9+V1t+XtD/Fh+/ufQujw2HXZ9+lj6T4n9xUT8pDatGgPe4KIYZgB00datW
UHLbT+7lDW1DElk4TH+2KxKNln2r9K+1Gg2+6jiolPWGlMc7v5LKfWR4tbcdCJGV
ToWWOebXMC0BHRynAtNhPqsHeYdJS140sXNiSXqsmyVUPOXeb0jfodlOT+zsdn+l
usdOdH3XQLT/bhdc5fw690Cc/mGjpS56DokxA13FCcD5VOp9Yc6ZeDehloluFpIP
Ow8EL8yMnNYvsz6iXhPCl8Z/luBX2wkC5a3Q82LakEIW9jIenqb43aDwP0RPzKwi
fIofPo6E/NxlvmeawGmfiBFTuWaYGW1pJ+dZtYZz0pTot+7JnoJ2obKsLYxprzzF
Ls7VaRF5b/GNRm092NVeignlwgjsWEAc0jJpCD/xcvZa1+Ol/5D+5e30CNcAq6Tw
J3c+Hw1wCoc/I2hP+1gXKPLbTNiDdbudCv2rAccW0X6JvTN6G8lUBBIxpGoG5KbG
qRHPaZixJG5mSQYAGMQVCQQuY7+XFzki8+l6Occ0V9wNzrUcw8Rk83r8nEmpCAla
ZQDNrOaQoe439VPwws1ryBwSzGHsXuCsT4gvY356OAqjQt8YLj1B/zjaZYKEMeMx
oXJnkpDIoXP3Uoa0z2H6GY/2hmL3J0fOAHoZufF0KJm/KFaiCECJqNigUb8Xaq3l
0PRc+dLztK9K7zdML8UpMXtpCJy915MNp9dQqXTJ2vhGc4xHwl2eyRcmRD/Eqsn2
b3ESNALcZPpeoVAHe/dcH11nuKHXcc6jS/YQR1zIW2fIOqzD3qtDfn2M7x2vOYF5
oIoOL+QQC1ClTSuTHJir9l3Tmntiiw0cthAvDV/YS0cmZQGbn7loxxwft3IRyYk8
YDyfVKOhyw+Wc57q5nT8Fnzp5u1gTQnDUcFcBQzK10aGRYlOjS6tcdJFBIWcnXtE
Fu58Iuz4aObU+4mCWh3SDdNsHogGza98cEDUYCy5hkkEJ5crgBrSUSj175Dbxy4X
RvBuEx9twtJYqdCjsK5QJUMINpH7BdUY/NbgYCw6SDPs2CT8QydzOF2deLT2lTDH
yvI0rdLOMIswaDKBPYxM0VmJouvi+zggZY/uLyjr/k+wHNdvPwbfH5AcyUkjaWW+
7m/ZFKT9O9E0ITRTR+8Iq4l2f64Gx1EP1IPajBMExr3csGOr/tyZVogqboesvi85
cXloV4mSFfqiK4if2jCqY1EZwUtdK+CGtheUVcZeiGxaUlpKbCOnjkcSGNNEZIWh
VhAqcBSCUDRLqtO8jtb2X0Q5zWSSEfq+RST9n4lBx603REG9czvqZj0hOKZj1mYG
c5t2RoL58eBxpJD70bYelAs2vqRRtyOEZkcRMvX3L0qP9E956jD6zC6OtcPb2FzB
f6jgwnRttXSj9+iiKwV3EdOvA2idy5a0LLc9NmUiTTQ/I1xMhLIR9FCZHdDydc1o
TWVrDTUxvglZfv/HAztrFIauPIYJ8NPwn19Db4B36w1cy6k6MGPViJ5e7gTD466m
5wtNZs9YpJ8lOdKWSpLl7Wd/YWHJ1R0eo38Hk9Pa7RfErngbZJRSdVgipkO7eorc
kuannRx4lAIN5mxkVp4E7Euki0sKTuh7QTodzskwpF9lR+kUGNCs0dHuHS6/mPPr
YuTEGwvIvfOgIuoxpZf4WxMiaa2oJnawP361JmAghzTBRKPrk2g+BqGs3N81C78A
e+Hk4jRtM0sRT/l6V17zotO48gE7ur2K7Cz+ZwpcedI90JO6UTR7KlH2T1xJaK7s
RHYerN/kP8L1+PmH6TYGk78hTf8tU9+Z5EGMXAk98ZRHA6dBTGOBkDJUSSx8bZwh
d/OXANTEYCB+WKhB/pfpl4GM1J3iUOhdzv7nPcaPborinRidUZqTM2C+lRJozqds
mD7BHmY1igPyJsR4k7JIIHKwy+nLatvQi3lCDGpy2zaFtWPn4y9koqs1Yw85K06v
/IbksDqGRvZIaw+svIDAPPKOFCduB8XyW1v5qcDqCxZUe0xO1+prqTBHTt2hDPeK
7zT3yX+oXaoY0kiFV40LqUW3MJG1dJqCC1KyW3qZDVLAv1aSvK/Y5LWZe3dREPQh
27Y7Tes2HJbUZCjAip0zeikXhLq9GvENu7YPat4pixE4yW8C+Cm5h9otr3ovQwpu
CUcZz2zE0vzn1eUB5Mdgw46zVMyCkWo2+QxG/xcL8GUwKSuY9etCKU3FkydPqk7r
qKnLoN80ihE6Kor6BIX/hlGjt8kwr0Kq235UVYvGsj8pKmbi9/WokPHWlQHgg6+V
ih/XKheIh08YxwevFO+fvdxLm+3ykzJiFIu+eVmOZlOyh6lJjuo0r4oGr5QmwOMi
4tDFPJ90NyNIcEREWmQG2PBdS3WkP/nPRIxqfPyX2dtDF7xAug25Y1CvNS+FG4DI
BU8YBO+bVQ6yj10XX7P+qEjl90hWbOLBRzoIeoonpu0UaMJ23G/3n3Yb8Ta90Oi5
6sZV/5o0F5wS14sODGyvV/UUsIZ6xNJtxAULQI8GGUi6n3egZYYQVOVSSzYPQZW5
hDo6GiF1a9CpGm0jlQTxEXsrFm4i2ykt7SYXGCjrklnoDTtQ2vDXDyUov+o1RpsM
VAS+Gbpj40QY9SfYaz7+IIMsiEe0qSGr/KoqmS+kbO72Nz8IHcCcckGbSYhK7xxE
xWwLvdZOtYNHqXHA1SV5QU/9f/tGiDx3QDkHJH6+/DBOCYGCAv1GC7fuTlVy4qfo
7PdahrxFvNEhJuaq4JXdLIWG4F7KqvwO07vrWAe9Zd2f4QWDbSJjBqS0AT+K26aL
RAjVGCnCyNA0vlf6RjELyPMDzDVdqbb1K0/9gvFX8Gje7Vs24MLueP3NwhuEnzMO
8wRenVr4hrxgj4VJ/SF94w+iEbfBbF2wWJO9Ivk9nLDhZRk6Wl0DwgJ3AaZp5Tv6
s6HVEQVJrx3h1HH//6oFUGfwpQtlwzsRDXbVtrroxWFq+wgHhFl/LqtmRQfk/ufr
4NlqIfQa2rS+ztrC6Q+/ncjV6XMdE6jwtO3V9SuNjKHsBrK3vyBRe/yavfaU1au3
+6ozgtmq/PsFXbbyyKVDnavbpIr4L8bhge3q61rIvfITl0xzw/eGepgErFgveieu
Du1RruuWk4IHvmTPkCgmqkTTud/QYMwVL1Y0UHOm8sNAHYoWIeK22k/GZLdhSQkP
55/Z+uP/ZIvCrKcjqvXVO0Qt6Zk9LwsKbX8W9ibItI4OXKUuloDaTn8FaqawOMPs
6C2wedkMqxTqQFL/FxhTXfOuuoL+tcmWG73TAXtFobBiF42bQRi5BqI+sdszfWPT
i5UO4q56WBuc8Idm33/RHklVJ8llxRG6B8wwfdtICtHq5Ll7Mlac5OSszn22K+GE
DJor17wM7U1zlp2v0OoIC2lI9wBt/xAQ+hbGDUWOLW/YQZkkKHFsGkOD1KmmUNmC
As0VyEOjaKyNsOXYqTDJSR6hSGqTAYScyLK1h30pArwqTV2lPizYUf+nVExUX7+2
bxhTGvgSD0o5hubXCn6yKWWMmL7b4tHF9g7Z4huC6Sg=
`pragma protect end_protected
