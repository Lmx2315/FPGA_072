// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:32:44 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
qqVO3IotGmJZlZ5WlyjYGvHtb2y3oB+luJ7e1h8hx3V5e3TJDN9qUXU/0VIVJHD7
eG3e0ktuYfJuJgzV0Hc3EkT2KT1Z0OOV9uNuHHXu4G6FscKn09SbUZUCWX23BRPF
nmG0g+ULVuXZb8TQmhSkM1iJB1JjcBxkz9gfvpCWazg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3040)
IL8AxHGmI0rUGFqQIPfPt9mpl9hU7jvD+cbKJpUY74JrRnJWnnLh6evqKgmW8bOM
1no4NKQtHIRCBEj+jP9/1tiHruUefpa3rLk7FJWOBpwJjHaWh3btRJ591tMlWsGR
zsIP8OiQZ8v7nllXC8Zu0QpR/SCz2rEs0ImGpXswgIO9RdtS04FUPlJEU7yf2plq
+efB+xAUTBH39DNdO17tLaf6ep03OkgsK8blg0Y2TEK1u98ujiB+INqdR2naJYNi
KC0pxeP3xZ1revqpqHhhO/8j6kKTebLMHVqU2W60knqr8AvBgf83YsBFVAzNUApN
ahS7DXe9DOE3CFCg0IIsHRZ1xZhh43JzRame0jykttZ3fhejrjQN1WPqwfwO58yJ
T3HxoPQyESpozatC07S47Fp3uv1emth+rGdSyDwtdfPuZFsJycp5G0dywGSde79/
lGyjIwd6GPeaS/vUzmzrGtdTY7Swf4SEureOal4S0UKAsEVJfRPo1HgUfALK6uUb
OLMwTIfGZ00k44Kf+01hrSMuTm7Sbm89LzHnyLPYle6CdE8mujkEhNO07z3dPGAK
eq5Vx0+FVt3PeOn+n+eDcql32eQLAa6YitCZr6ggh4CQFZ2BltvBHEpqx7P4VaQX
nKGIVceqm5+sKcFaVEId25weYYwE2aZkP/a+oIzISkAyiw2KyR35QRblTc7wh7GA
CWIh6gJQE9fD5MNZwgrNuSbJG2hptettdKKYtdeZfo244Ne77Iyfgat+R4d0EcP+
EQiR2UqgdbSFcRd+LemVcQdYqNmzj2LPgijsBpLTqK18j23JAhlr0bYv0D9N8zvT
DJKJO09lZAmfGhsEDL/SE5rVxeKium46CROYasApc8iVUjdJBqllSBoS/QOEfeUY
wQS6mEc/JwjIMwoCBRwy9KjOqbUwApFGHQlAeR0eWy3A1tCjOSv8uESPvEsEvr//
Z5Kj3xZ9ZirZSNphCu8/r83rlnjK7QRmVhU/4auxA7eDdrphUECR7dNpOUHjkbg/
2IEtEOWMxh6T3+nLGGkFW2NH+SFVlA/y4Aiyi3/sx3ravzFFdPw0dydTsznH5eFB
llrQ206WOBL1WfQLL6F1fsJ+Qa0aHYfKXMfkv6SEFfNDFMDaftNRBDqH0cuTPsx2
buyeLbeEc1GiUlOQdl1j1LWfmhqenxha3DVmpYyK9u/XBulYVhxSq3ooH81pXLI5
QxZIxkCIAan8DsbrUiTfdWxOB4GCdjctbAqgp5z/bWNV40N3hAN9P4TNxn/2ula7
3UR3KHpT5Yyn0fkAXxUxae1JyRcHEmTuW4tWlBTEUOz17zziVxRFGYKIGzINpoyO
UV/rgl8nRaw5z0Fgw3Iqgo+KM2/O1/HuLotF7U5SyRwflYmnVssj7dWep4hzqOUB
+FIb3N7P03vFzv7VnnQdK11yEGCsbgghkgrao0TBTRi0s51WSAn/lyA4Y0LuTtUa
9/qAooZIqc9BNNDUzE5be+xe4ULJJCcuGYtuRVbcBak4qh26+SaowUKYaqnJgDJw
v1srRcxnMidlkbr00kpT8YX3aSy3xhtQRdOGdjDUeNM7HrkRXT4edFiTR3lPidnG
3aUXY3UPXr3e84Q8uzPenFNFBqYIz+d11BpMVHKMNEiB1qPsOuOyCZt2h3+wl2ii
Fh88cVLBfZ7Iz1StMadqD2yJ7uf1fgXbgQTKZ9ynlDWa9QB9OBlskFdQDSG96meK
5CzvMjAfebiCVyMQq3nISrykVikF0C9sTw04YSFiwZW4tGEwglou7or79nHQ8jNW
URpJsoQir4bKwNJNKv/EOVyJsUJmkQQBwUM4sRfp2nxpmJsSZn/sftU0cBfauwMq
Rz6Nvij1u+Vx8tDgZFUD5q7oxpPqR/oUJMwODSZTr/i3yllMEv6zLdLaULV8YFdK
1JDVN6G05Y9hXSU/9W8cCSfQBORLGw4EG5RWm4cyoMs7F0QR+uSkuXzGDvP4NflO
x+US14QkiWOirqzLZ2AS602JV7HlNZ1LHjDlUyevaZRs9hOtskpwNEQERi9scG5R
PU8dyeyFRfSYsZBQR5U1oWELLm9LaGRc+vS10Y/SnEuiazs6VVm4u7NuuemwTbhD
ix7D1zSWyuiMs1YivCV9VC2aNwM8JVfFsb6wBgXUv3CMi0/i2sPFWdiXKZJ7wWcG
Jgfls9kY6fnSXJVSz94uqoFYvYGnmsEdEJfQO0mT9HvZOxMV36BcxvVstz1soqS8
MH2fcImei9XdIWgLN7tPLPveAc329yoa4LmeIyacY+xcqepsfuwVw9N9I/uQtG/T
5WaM9RgOyWFrVVQiLJCqM4wavZjGUUexx3HxKJMYRS8Zl1GqmkZQe/gsae/vUV5O
XZm52CQ2EJ1zg4N2dFPG+qd10lV82/OolX1ZXtPYqOJ2aOeZJKPZWp56LZFYwnzD
jJg72I10VyvMzmzBPBH65qJtynTNzH+uTZJw6miMx63mo2kG+rCh1RNCQRvVD+7v
3We7GiGskHapTGCN8fyi+bO9Jf9bcX/fAtpVIjfqDHanVtrRVN9HHsC5z1SJd7uY
PiqtPFQNQaS3goMFCmtX4s/kwrPtVRCPgcMya5cuyVRGwLDcy/P/w6+SmDpZSaVX
eghT+f7vJWjDr90or+7jy6i+saRfCSaW9uBaQyN2lncdam25uIkYfN2YQBsUhKyP
Nd8ThzsF8OBff5oAAU6h8xkSwApMZsqvlZiX+v8exv6Ma9Ohj65s1eePgxBhMc6i
R2W5U5sQbweogOLSbG+trwn/ACy9OGcgPtFXSYL5Onac6GCdQoMGI7eT64FlfKb/
jHzXxKRXrfpfkI5e0gqOagZ1vTxcydHal/7aAMJIAbwk9R5Bm9wkWllbdryBNP+W
w4yN+u4iKVBycdzHfqlgdoGByr9bOJQ5vYUKzjTxBTxcScCRg5MDkCQ9bydK+QGo
D/w2wgKbxEYACon2XzZX0VXGq0nuJMtiyADYpqnq+KU7LGoImI6WUo7ZIje8d1bT
3hgzHRq0DtNqluyPuRpMZnZPH+r+vA1OLymT4m59yMQ8+J+w3BgOJWH3B+MgUbV/
4A7jBueesfciBoamkSJN0FvjRl/7U/dqCJcQeNdohxJosWMOW2hBWSl4MxQgGAvQ
xFL1Ccr99DwXpU+P10Cv0GNk95+Erf93SXvQQTAqb4iqJUr4uGtkr07jBBNdvHgp
eEOOVwKVZfjoBnvBBkja+avTydnCu34+rTcyd/xzF8d0Fm9c/oVx1X3+T/b+J+tq
tx4mnJhZsm/sT5uZND1sAg+O8g63ZtDGrIUXJTENB6liJZk+gI3lAdV0FXgWOOeG
nbtq3i2zDiRfgNVbMlpsRMe7rjWfgHrtGTj/EkS5byDXi04b/WOFfsQa8ic6zW73
6OfKDjqf0aYJqMLglSaVDenijCOZ2kYNQjPoDJ1zV/ZtNwm8Rjuzh6GLgTG2emkJ
AAEMXk5Im0VwZIMS0RR3fed8a+j4MIoo4HLGH7AWBKOdNYND6LCd02GCrHE1EZWw
rMIPmBcD0THBo/MdY83jPkt8NXKD9WgnkMSMWVVPdbaO/PkGa2IOvq3cAFfDd6xP
+U/wrr9aSkldBMRX8xkBuFAoP8huTb2rn1wJYcX0N1LlZ+T03l6c/7TJTzT5Vfym
Bb/aq2jC9KMQMmed8eOC5keUi0HUEkBi6f70vAecc28PAi34thhBRmI2pIO5x3ug
gFycPY298lsf6a4L50xN0UMxcKiQG/0Iyn7+w2PXf8UM3bgr9h19op7Iibzhe7By
sJ3cLwOdJYJMd1nrnYD5veD9yIWEne6RijyFO/4Q6xkClKdPAbU0Pmn3P2AbH6sw
25jMLIvUrfrIhTPUvxyFb5RbAK5F+Z04hEl5j9RxAqFSoEWr7W59B+xfFoHqL0ta
Q+DkaF1Une2rPi/F+KdLfkpkk1Qn88IV8rtQY6/FwYQi3EwawEBPM9RQmQ2L1PXD
2Qkb5jDKYqSNnriRmfqm3VUlsju9O8vB415hM5AFX0uoQhxglF0KYWRtDHDWJUim
gHc9j/W3I5cy2h72hRSoIA==
`pragma protect end_protected
