// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:32:41 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
XBusMZa5DXzfnxvJQCdg3HEXByQCly6HBQo417WVXuChxOhjmTM5dW4Ph8HoZdmk
JtuiDDuL5lZYpeUgpUSG1Im1+SlO2jJHhJYMnlkYLHvGnkblE4dDtV2NPi2neUML
oYpaFZ6uI9s405YuBzaRWBfQgjdM9OKuSIHfHsRprcA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3280)
cHesCXq6dn9FHPyDmnTj4iDmLBHXJeyHGPM+SiMDcaDCevhy7s2ZP0R9p1p9hl1X
nZJZoTH8v71dgBn0nztN4MVzdJc6RKbqrEYskqsenp1tc828WDejIlSRMh60XHKG
9EmTERg8D+BTVAEdKbGSYjkLBsZbJxl7ZLX8owZQR8dCQmuYYlUrL9v1nCcNnMnl
lZ7emX+5ljd7xR0eJQfb33mlhqPzQZxI/8RZVXwxA4U5Jy9pxiaVBNLlRpALnKj2
8el5F4ehBF3i+GmsdXBRKlxVEtgFcAaRzC4bMllnpFoQOg4N88cZmVscmYxRUDHQ
BKJXLW3Wd0nOtrvw1Wu7duCl7P9LDkIScUhBXBCbcMYAW7C6u/aHNwYoaJlHfzsD
lqAAdxknOx1caaj6b/+15DFAeW1Rr2Sxy5B/T5sPRqNg7RVo6yhSxnjkmGFVRdA/
N4HYjZZd+q7YJhirooYtidjqR0JTD6A9ddP4IpY3n5yceOIkeUFLiGVnS/T5fDtn
tk3AiyT6tWlM2nhQMurDSaKvIjhNqQgmzugrYk+o/f3TeyaNT9gdM+2SU8wxhrp8
zd9JFz6vEM4hUAH4DgnIuTLMoT+OCvyQnDWsMLBBzbjchFgt9TSKJCmO5FHh488y
DxKFeH/+ouCjaRL9npdA4a6Wg6oNliOKh4woTo9Am8H1BxkRBrdaZ84NvqLIbYC/
NJS/nWze8i9eV7y7HHxKWha4FqR3P/qhWPwkLOoCxvcfSSpYRI75i1lRBqyaVFW2
VSIqQsEuj74BQSKBelUiZvqD5CeAjcxtW1FUEN3jzkktEc16XMa/AftnGX7j2ArW
ZrH89o8CqSDkOZ0wtwrhSVtVDtRaGqYDa5TBY6XLyN03FrsyAXHafefOF57QyV5r
ZZsfKfPZQfr+t7+JEe6zkGab7e+rYyOKHpowjazOMnzIXT+IXl1T8ieqYVjqLqv5
DA5LSPIoK9MNPEK7fuuoNlkL7vwpo2SOqQnTyg+0SocP26heiVXMg7aLsOUIsoND
wLItLsDxi7Y5IzdyGOtnhxzBMAezHZfZ8a/76kITwgp0RGf2lk0DaJNO9QNZ3bMt
6wop8VvyJLqj2vRF8UtIzA4qlK+raPqpXC4tEGPLd1IuKi2rMslN/ykxapwLD/Iy
IdAkmOBbHyxE5+ub+TsuD0+wkrG4Up7iWraxax/OC/RHa6V7wARmsinW1rLdUQix
Aw/RYsbQ1SUwbQcAxHK1zs9UZPB0GJAZ/69zI/8iILXdWSlI+OGF8wLzdtPdo0kd
230N/3x2jHwsSnrSwNfpVpQElXUqXT6g+5jMTQo/z7Rg43AdpdlYe2tdiSqXEbZ2
gXRNPfvQE3rB0JqfEjk9tfCOLu96tDhOUCl0t5UT/0afFgzTialGbTXGCwZpX5Gs
KBg8Zguf957lBcWzzHM0RnRT2x0lLJldSX/ANPveWkeDHcNvJuNJfEtR872rUTOD
t8McDkrlnZ6T2CpGUgPlMg3h72M5aUWED+3G1YSyv0ZfFSgABm7CAoSP4q0RP9oY
HDGhSf0fuldDCI3ekC+AHd613PTZRFLUrvpvDJ0ACr9S1KPFs88Muqd5oWKtkJns
osZgGGqpbjNbPS3mXi43HnpZ+mKRprAOvyK848FucBmDzgo3cJFrE//nSCzaWpxQ
J0HduO0S0zlmnwECcM7aLl5rK+coYOlt7fI8Ywf0LPpiwfI2GFWbmwQRdvX20LKT
4S9IYNgmigPLgUKxdiMyZVa72qRKE4qRsDtRf9JT/07DWbVAF62H/AakMyI7n7zZ
8zHYOndv6CJ4jix/zjxWSgqIARIiCUeWTnVHNAcoPORvTSeRxh15MqtELGB0A8xA
VAwD3C2mpxk9GQXQkZfzc6QZLs58QoL/bJe+ouODioj/Fj5kQcCZe/Tie54yL/Wr
9utQNw16ADVPH5LXxER+996QGk5ydIMgysXPAOdVXwzWsYLdM3tyFgKSzxbIrhdu
STPSdCBEJXIesAAPFP690mMe9hJc5Ibl5LueKlGeeUhaQbsglEz+PXJOCZQh/rUp
W+IT0I7y7uSVn3vv4Dpduq/2EY+T1pmHHPihlAtxdlDyaRmmDIvo1AOkIcyUBm7t
4yfLR0yRr6UWH75dlgfQa1bsCxmNSCujqu4PN98659whNDE928st61HVTaTUnr2j
su+7NebbdEzPVZF+gEJqmt+p4PErYByVjsclm+kcSoGnZc10AqLHnvbzh0ewYDaJ
tYdAIsxJmSaIRm/4PRbyyhkE43iaeGr2+dBgLEhctno05Q2m/aBiauBFXA7XeRdC
utGmoOe2IS1QWnK8Y8XiQavQwoU4wtFZZHpr9QR57crHuPaUpuY1YEbDlCPLo7/i
7qS6iZrVdXH3FfU6rVnMBgtJ9wOOeF5Vpjxv6ebeFt3Ts8cm41wgf/S1TqO/4wbI
kHEl2HIjrtfQ7ljNxrWKfFdWXFTikyhyrAwPuKTdokJzhaiUO2wZ85O0BMyGjCON
/CimIaN4SoI+6rQf4Tn5Ht3hxGskGZ4V/avZ6TRTXoQEgWKorZx8h5BPlD6Y7/77
0ZxSVuQ/kCnkA/+rgwbrKg2CC5iYPU6Ej0fD9Z6cZM/kAId0rTp4ruJcHY5jC1+w
OY0UqVuHpk4nyKL1JTOUHJHfraAXCqbOdceuPs3DmH4Ux6lr54PK8JuCCsrCRyub
2D+nGfoNjJBU1sSTBrlgGXnFjZYRNlepC/ZqP1KwZH/wT1SLoKTvVz5TnM3Aucn5
9Z64YGMA+LbgxbduVeqxcXyStOOVdLAVG0+oaumpmg4t5hnFMmNd9IhMnxX5pJVp
uoGxGeBFmf85DX9qOFnpoKnt/YpPRypYXUf464zj++Gq0x+ItkXIP6sjs2/+KjqS
DLSfaHZ/pIwc6kv5Sutb8poVElmhiATraYgQc1o8VDwxyokuuPywPK3ol4B86KPX
BMEEDdlzAgnQJFzYTlHI+DmbP7Y8znbJf2i9d1kZe8L26qA5UQj6YYq//yZNbf0H
e7bsZkbpR38k7/yN9pviPRYW5VqF50E9zSoH/WJWZOOlsOxX8k0CA7s/sRxIzhu2
yvGifjlAB4lNo3MvLGYuM3WfJUHAZW9eVMZ42wS0ASxJSsImgIQFxX+D1uhxqu/M
mQTMol25USHAYc8E5QP5FMZ1K3AMtYmtosgly1VepVl/utxfvGal/rN6Or0UfY/2
NC68d0ugWLYzPQDOb8/snTaGrK0NzPpq5f6Ua4gmTT0fKDQMlz4z0z/8/I/9gOPk
/ImyNQEXOEnYzA2kJ9AVOtpXwo3CLH9cbeAbgIxNUHmenzjG9U+9rtyZO4A8yj/c
+8eaPa8XXx2SjyeNFwTiV5kRmEmNzccm+jxn1SwkaFXCkO4k7H/7y2rKDAhCs8aD
6NvdFIw7LDdRj0eax2Au5xnM8pFLbX6S0HIm8vW3nmX9GjfBqKOovBwhqgnKeCnR
Bmyct3iAsD5ZbGaO9nRsvbimvjC9GrIYv5FbE422ShIuSZSN2Wv/oFb8gyMecBzX
4p2DP8Sdg0rw7A454zaiiitq4iTC0C72D16yUj8sYyjBDwQp4zrxPnLuBPFgbrA/
+bMfJR7Zzya348wdACBW/FsGaCXBs2rOcIFUEAncXibrmzIzh8hO6b4Ae5aXu5p7
jsM6ItH+cIZDRfKmUJWJDX2KrkCay+ntmqTgiAEqhwwAuW/Y1tqWwbq6fhVx0hXy
uYqA+w15rK019LPZVqD4pZAJBCVNjATLobOh3IbEeVJ9MCYvAaoQPiUqm4Ts+d7F
wQGo5ofpy10Vk6xq9yAy/rNDgm8etq/TZiJOR+J2oGWNmA2nlHkeGZeiNua0ePiM
d2ogIMAxI5lqcwN0x+4OtaIk2Uz4rH4nAGE0yvKqXgTj5I7NPSqVWdu3Zjw5N4sI
ZjAGFGA2pzK5UsHu2qGg5kU8UENwzs89bGnhHfP9JiTEUUahHahDUHQkz76oDpVV
V5z5MFMa+dDwRDTvGhoOiSn4D0gNc/KWB7vJsNEX2QxtQFXRstuTxGw7VEpGwPZH
5Mo6Hbe3UmEiY+UO4MtprrS+/8eXisDuOKaLfdCcW3vHgEnrJC3Gzs13jyngbina
cp/OxQWKqk/DDHwFmkNOmjtNsMCZb5y6+cD3Z6RXIPOCOE+0liy/usARyE2kql2w
URC3Rfbz1nVe5LLtZsWjthBMpZI3RJ8GK7Tal42y+9bsvc4f2Ge5yEeD6bpV8bmH
p/NyU3i88bZdCl5DLcTn8VrpL9NLPOGeTl9QcubcHD0bgbr34HcQw9SFDCvFCijH
7hqUh9beBWHeAPStXnYxnxY6Q2kFaSMRtvHiBS4eY1dDHTtxcEMesCzX4ZRrnCZO
Jfjynbje0CHTDcbyTuWImw==
`pragma protect end_protected
