// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:38:10 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ASYN5TTjEuai/1RkZ/akmRQvLbQg6j2ZdRAGApJhbIcHcTxyi+5N3/grlYXpA9ga
RM+eNzpvbyT9HOU8MZ2rdDnErRDN7Fzh1R5iujhaqN9hdTbxCMgUwPmGXhSCCrNy
W2WfzMN0/K2PgMsXtzsZkLDimqzEtTh93EO9k3/yhIc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9536)
UaasDGL4YaK7XQq/ppBPlvMDA2WeSN+H6Yk81u3LhX/2DzJx8M8Wwa94mO/JEKO3
YJN2T/GHnlKS74ufi7Kf35rOO58rZBbgz/wlMN0L/sHmpaKuHSkDcFJaZUkaTHrB
Kpr5LaI6g/Rev1AZKTyK5AJJXm7zR/X2NQ6HdqJNfrlwUjuWCwkZRbRYQgwutALs
eWvLl0ww5JPx3ql0XBGoF6xcVZB2huZ/eh9DMeFBEn90RcIF7abiNgjJqrlPdFjw
5pu2ykqdTe8QYBaNwQLn7tqCytVsnHJ59/Dw8kAO03TUvQ5fclYY7WDaZlJeAMZQ
Y/0G1EbRe7sNXwKGBtmRGhz9GDO+v7SIY4FG6O4Q1uJlszTZ7139yFh1cOKnQaR/
XeDDS+NNfoJG+Y3a4TWtVpxiyQckjtcd15yxLaST3inRrlnNzyuoZ4qNHOZO26un
81uHxirTYQQz6QmKKyYK9nSfQ2Ry+E1Oywp+ipAGSn69julOAcgbdnJBIwcrr2qw
5yByAFul1Jw0+d7oz/vtKqi6RmQ0WeBe9lQHmc+/KgJs0NWi7auGL/ePbeUVnrFm
jtkNwRa0yUjW1cMVp+RvDAA2+vqu3QU2X8gPwsWwSX3aK/ooAMrkYYYDGManJCg0
1+Xq2OP8+O5NioxV+8/zt2tJFf9aLQbExS6QLDA8c/2/STOk8cHDuthAHpPPCupD
71vqNAjB8XdTet5BvT19ZFOsUuUwP1m/lUza53q6VoevplWX67CAyDO+WmlFvAzo
KkYRwxAL0dKG8EShVBalTpE7yBfWmTq1kAXyWkzC+YlciAegK7fS21hK7GnoHGs6
Aue1dtH8W0zOUwzWrsgTMtaCISugyLIpJFhWXOsSISe1EIIZoUhYWR/V7WWHf0p2
rfzBTisSdUmID8GoD3HjLNLDswJMA52L0ZNrqMJzSi/OLariAIPn6Lw6OB/RYmCt
UwbUJGGOfRWs+kBm6IUPLSka1n0EujmuR+ppp+XFW5WQayDV1T0Ge7oLpQAenDfN
tLeun27/YxjwsdfGlEN5adQ4Ur7CKFVcVYAQnlSsNyR3X/b7IMM+FTn66QSK0uKr
b5mCaLb+q79oikejHpWmXEUgxZX3aNoHHYSeeU16N6OHAFFdyCBbA/8VjXEN7Gwy
12VNCRPWMWiYPhvyauytj0pnQwaz1oeqnc5ZyypJIa3tVX7KzXQ0X/+TLxrPcYBp
9Z69XQy1wQlwmFwfNpQvWSrzzZiIvgXNDIFiekUPHBLXnVMubh4Tt65yzGSmOEcy
0uLzmoupqXZ0HlGnL/mT/ODFJldFI3K+kQJxxOyubYxdxVIk5AbzHexZ5MLHdcbF
g0B8jaEPyiBCE4BrJHM2K7RsTHtSEhrQsj9oxCvo15GiaoHOxsAWFIV1zvN5Sfb/
+FSQzW9bQ6ysyFodP/2I36ZvubU7G2OmLsPBHng6nOJpsPgqIbkcnHr2O+l3yRAk
0+t8C0Fk5HcnbQcE4qsfpSwSUvswqh06qdDy+ONpVpwdm+jVjcB2klpLGkWWxstb
tAFh0dr1922188BJnLrAJy6Nobnh4n61Wo+EGVCV/Dfd76t1XzVDo+M2jVCnXRfn
3IAEh547JSBc/MMvQ620abED0reF3Qdcp2roiHuwfl+G3ynsMVeWfCN9OGcys0RA
6ZmO/ACET6+QqvPXtP7uhYGIMOMXpJlqhgY4rak+zkdfNxJpDmYKHPLaljRrH/t9
KqaSeH/YJnirPuiPZDj2Jo+4cv+RHajn4zcSkQra+URrg3dibz4L3aUi7WJr7VpB
qmyGJ21G1oTbgCTHV6iA5nXW0QNQcd7UCpmrCpPvxQcn4r0SzCRJzQYMoKHrIjd3
Vr43ZgW6iKIza/6FQXnmNtCzmf98b5Udm9di0ezr5f2Qn11n6eTWgliqbYuFI6lN
qTKBybcJAapx0Acf07J+5cYArQGChWMfQD6R5MOnPO1d44ZgddmIeLeiNXzOuFn6
hy+JvJDtC4bp/60Eco8iKoFKMF64a8xrLlnqsOrPehjA9P1j5Xxm77pz0xG7MO0O
isfbLn92GKZDYEUQSGsEAQH7QW/jiBTxdPK1L+50Jtplf+3siddegqGFvzuuxrFO
xugFwrEMt5IMEBBrF5wsPU6LToKFao64iA8/7G/lG9LFx2WZaFRXwPWWJHzgc9HK
V7TrhvF7tX7sRTYOf98T89Dcx1lhnhfWnzJES8ng+0d00s1xMfs90zAzQB/mg3gF
SBh6/RG/AOTGnF8o8w+GjoGPzlrVWhYLICsTDnHNqh22Uo1kKjVuUi3GFAkwbPpH
oqGYY8GlEygFyLihMWtXECvrz3b5bAgfPMmlsmbJnPCa+oJQMS5uBnOWmkp6DDsB
LLa+JEamokAZFbzqF5+Fn78d+t0n6MvVEDrmXDzf51CAfHx+X7fw/H8SE0+6RZ1t
2t6ciBbJDJ837Hdndg6D4WgaQfdbHzD2k14qdd4cZOsJlYPsOC/jOWZk/1NKpVPQ
ra5y8Kn8E/rt2rDxwA51D5CuUDB63CHtkgUJcNoeJUa7zInP4VQzttT1iuXJTNnr
YEXPnlVAYCOGoRIjNxv7nne7+wZffA8Ltz/BGvENKVaFsnZb4YnhcHxccPvmQg6P
znOpcJZJ82cdBiuKg6PDBB7k+dqS47PWO2Hy8Coyit1nrPWEH4k3ep9cmIgtPNlk
QgU5S5DdMw8pZhvi6CDjVDgN7F0R0863+7ZLuav0kfmPw7c6nnNtk+CfxREtaxaw
RtlsmWfySN8e3J3TYN6HjxumfODJgRth/ziwr1kbEyaV8vreTsJ06HdwsHBQWs77
5yCt+qxGqpEIJNJhaaSxoazJkoWBrjSBlhUTVGkjuyl6RPSWojuCSRGaayqNWmiI
CUAH6QmEXQWqwKSIfbCBrBIQCgeO0HyIem8fdFXE6o/T7xlFVfFheyylbPrWV/zc
njg8hn2OCkicesoyHxhFVSBA2MNEHHZu5LQTEI77CQFe1KtKiH+X+nez2RI7s+Df
k2P3I4o/k8hrxRggQChefRaKmn97OUmIJmwdCdYjA2CvptGDdF4sU673LJE9UFgh
leagvbsdwG2n+i5Dx8PkrmNFP8bK0R5CP4FFNDLbT4we+2OWqCVXYDZzweKeh6H2
BG0kDH+QGVFQRyAOJ7xZu89eo2YRuxuSKL01c+00HYFm2tFE6Lfu+JqIANFD0zuD
SBrDDTqK0ANq5bKLnz7Mrz6yqNtppM6CykX3WqtIA5YwHjrkZ8j8zR+4zMvwVR/Y
60VSJKgJc+T4O2TzYcW1oY3gcmEsD77TGnh0bNZIrhXgllIpbSISSPZCkbpfQQNK
jwd8mnKqNwEu3Y1v/PNYv0rxfi9mqYiKEnkVSKcE6BbK2hCF73SjenJp3YgRW+7B
FpGEwCGn+ZdCCEmCgTv8XjnlfMIYm8lLG47AZ7lkP+5MLI1JVmS94E6sPCN9qgj5
yBBXQFCn65aR43lOlNQQFEQJPKpVtMLT2e7DG2V1vmbAblUswuP+WqaspzqcQMpu
+EcaR/1AKQWQmiOKTNKrTFxHZJIHAYQU5rEkxf2PrVAWoz0Ji/gslpFUsx4dof1H
QCunhwhSxeMjtJLEGPnha4NssAFKTKVey6YHPzx+WsIBQqFlAsQ8qPqfX9ubh4rR
LeyA8py/YqDqRbmButQuaCzTTQS7AQgzuKZ8qdb72uBVmZrgeCkcZFM4yLYwPfHL
pmBK8+8JOkWrbVXrqhRLODWEo1MIQ08tqEzxk8ZALtr00y8Y++QR4lHYsVALMB9+
eJ46QxLDNHuEbUXkHiMUoPD2DHXDsmCBYN1lAJjeROMLRyWJU0M7il7OAEALmJTK
G26yLaukJR0bw6Jujg0xsjLo36B0bmdXDsuS5qakd27chS1omORx+ZKKPzNWmTb1
/2nfFfkFQJbeRy2HGAGBX68h9JDHdF2/pM0iKitPPsigMoL9D5oZUQtx7uTY4M1u
N+MWMksrdguzwWWJxiqlyqOON+xi7ZulBiMj2C6TrwQMRhS/smAAGWHhSyrsCFdj
JQYX39iyMIKY9tFH79irmlPaSSU+ccnFdVLScVJxg9++pKYIELmzRQUpFy4qlCtU
6/JfRWwsgTgdHpjos9GQUzEm5kNmxwh2yPFiexRSdcfm8UqEvlSXnDC0WI6YHxOQ
gWSaKlDFhzhb/z0OxjqDdBZJCteLv8B94XRhHFrQVad2Y9XDkzAN0dwqIqDycOvB
EA2MGgKuG50nAweM9Fo+Lp24uGzmcfxrUL/k+0grrYlsu3MEIbjcPjDkRIEtcJfc
h4fZkd8TVBfFl55asiuSd1jvzyELa1Hl4D9Z0glj6adZN5PEPQ9y4ih9YQTzQS02
2XnZDBK0WmR/tczOXHaMpA6giT4RzFNhWuxkH1D9unYAvkBOAJxVyXiXVXtabc62
WVaoJKXBblaZWpU/eYgk9z6jpZRTUFXPpRuwFJG0YGRui91V/3mwBD2qYvvBXEcZ
pkNIrwADyvZJTWEFgJ80Tcsu6twFD0qJboq0WjjhSDOpK6JqEq6TPR5Ed95yKWpn
Bn4uuV39XmIn7wVP+hym2sM4AJWazYK9du12k4bJ8/7apq9w0rMohdx2trgI+jDH
mXeRSqlOVI5LxB/4T2f9EuH7I5J5mnJpVRu1LGWnKGY3F9sqSkBHNGk1hQTpQbyC
8y568Mb/41M/OjO10Nfv4Lrv6PI4HEzsDMRpDpQZx/54CCjP3kiPIxKP764zYRg0
RrYvUzD7tADRTPnONtJ9Wg3qdFiDcZGEAftHUhzm4SpbmhTPvAkE8878dVqtPqGh
ETmsJg4QPPwv7ctUzFc2LaOregATUkyUyuNCQt82z0WQVjjBGg6zXyzezAzMwehe
bKdiHQGsskrBTQaVRHWsaOyuwbUcgKPf8iy/anjx0ZK//3O6FcJTtpZI1RyOFEHF
5emKdaXdV3MXofQ/fbnPZLV0awiN1pzcQcp32R8G6OlRWBzDytd1iSc/WL1/c82l
vO8X3QHtn0esAvXnvUtLT8IeovS/E6fgh/49upK/hhRhorqZFsrh4DnXveTP2RUa
5LdYtKZyjlYP/FTBQxBfzPUYKHzbwO+9jnEOtx+u2q+PS2MgjVnPqAoCgb3ik2BJ
KR3UWgoKHMMtU1XuzEGTePJ50LQMusl7l+gp9rF3uHP7n5AI8O8hTBRPKyt4pzHn
djJWAZNJpEpd+OghgaVVtyMaUABsougz4pruNdOyCN3hIBlfHh0ovIQwTcEgO7UH
CimIZ+vaoTChWdZ/gltBYjV0mPgmmQNokgK5i95fQ/73UHq+RZVevMSSndziqiRx
4c1em4vKG/++gagky4qrA90zKYaHS7EC0HSNdSAnRptB/25dMgvKvx8zRtTeCN1M
HPDFO/CdFkpOV/4law0DvTWXaOEF8dmEBF4v68oLn/HNFQrm1HWuxWpCxB7KXP/+
T74YUlpdGBo7k06zyRHy96OlLpuVuKHduUgROYuki9nEf4WteyQIHb5Q1aan2V51
rJwbD0IjIDrstkcRN3s0sRqYr8A0C1gETmLzjgXLeUuG4rC7lbmx3MnhQgYH+s8o
0ZLyVkvDeRV/9nFq57OgbMpZHiACE9P6S3ixteQRxNOQQev+4J5XD8CAFxRBYl4K
loxRnH80P3XyqkXakoNYu35rrPTpzOfdLjLkNC6tm3vgMCcJo24BO2HnvVoUvxW1
iRjvLB5o0mXGLbMBqYyMsyDiX3Zufy/e7jzKjcfUoPG1o8mIVbl+mAYxGQqOQ7WK
ADxEP4sCoPizF/q2yVW/wOQ5aZ7P5gLd/QmJ158wrfTSokJ/upAd5y/DmBNuC/4f
JhfoieHDbeH2GGaZa8Z+WohZDMcj3uOex6j+TlzleK1TNWnnTcZ36995NxDu3ypl
IKBl7cAjpAB0UU5EYOc4sfJUEn0CGyhraNAiKl1Thiw4nKlvbun/GfhVRg6Vji6r
7t0jLCg4DIj07FFfhXQCC66xwM/LG6+bWHyNUH197Wq3xWGqqRC+24Bfv6QAeLL5
ZRCv8fvGpiRoS02+7+KAgFnHsTXoq0J4pkwo7JNEAWYJjUR0WMOPrd/4LTr4j14z
QJy4ixjMSyGDB6uUeHZBlpVlMK5vVHX1gq/BcGXSdRyYOVkfKwOvvT6Mp9wWWFpz
8KRXbmgCgn+VrbA86emv3IIi/iWywZWvl8+u8wJBcYxoaOcLuPxgB3S7OKUamCBs
oAjJTnw2mhuaEbvv9UvFME9EF7A8R4X+4aKY5jUGOCa+MZ+KLKJ0zwCHhVDke+32
XwBgjOAuIi8XlaY+RxHSPDnRzgjhEruAkzVcCZMSedfa9wgLntz8xN68ZBWPE641
7DoVDoDmfSjcwbN5uCOyl8dfDfI06lxZe68meNii3mMXvjfylAWMSBAmUbNNbDo/
hFLT+M/nvrBSyw8gPZCyyGvS/N287P67J+vUOHNXuB9JcC6hleIPiQvpOpKxWNqz
/nFQ6kjedcu1nbBLJqVz1+h3y11Q+zYQKVmRinf53SniMVsDjqTv/mXnscmzxF15
2yytqS4NvZNXiBIVx8Ly9kO4Fsl3RU6JmPRTdw6fah2KhcBZ4gHBVz5zGjl9Gh22
evTsajXMvQnTb5EetFFyrGX1Mg6q6+Dl/7YL2b41BoOczePcuIfIEBGcP7uEnP9h
auMe2NKfsEkogiG/9r38A7gX8r6PAGyrCw+Odv60pPZjj83vI4ILOhbPLxgMyuv5
Ez6RQxA1swA+G3z9bO3A4MDV6xWACAtDGugXWYMENw3zoWtBNx006zzg+rhFGynb
LrlFyS+Ny5m76lZ7FxBY2yvh0FvUJ5inrGwcUEJZPq39uYz5ddzCFTmVx7HP/e2v
Chz+9fblmp7/4ubhYnK8RAlkv9w+ThEtSeKpLWZhbdKMCeSCpMSiSjRYvD6oPdrZ
MN9izGB9X2o3uBQZZeSWuzUxConKt5kfXUAXBG/z4YsifGQKApfNCq+aBzkcR7at
2a7W+3yHMnZOBdQuNPIOp2S9JKJ03YE2/mV1JA+cGSonzKw/MgVvSxkcjNAn/crl
If9som8uj9xfO0n5CBrc4L6U61ecUJNVYlrRjwCC1rjZxab80x/y3i8mKt8Ryqxq
h3SkvvKc1nAD/GyOwWjdL06QPLOEzjTTETRY5FZzOG3DPVvyVZb50liQ8mSWY89B
sK80LWD3N1ktZf3zJgxndnVHZBlmF6+cAKcnrTnpYawTnw6hW+GiInQJqrpV2+Ip
156LBUTbM427gozryzUMV2DqFYa911+Dk+ZUAH9FmNMQGANzRBHWrIj5vSuZznRo
fQW5xh3JRFjbfASyrGmBJZjpRgSHoE3tpqVCMjbDJMYBt6yHGXfjoWQ8BnlA4i69
05slKXzw7jCoVaiERUfOHwGBxsUEa8TWo0scVYLGw7bcbJKPpPnSb1pAEzeQvAwc
R3EzToXBxJNKtLpFLTJOkQ40t/IaSVwGsch+lIDxk7TWdTmUyiSA/pYkUaPDdmaB
kgh4vC9LgKgx5riVp0KaLBDq3voaPhY3eMRX020L3AHokcU5enLbcrgSCsP8GTZm
InfInUfcivUALnYXhu6eiJUHXYxpd/fO548OQ5AHN5vOpZTsVS1UivZ3fRujaPRa
jx0rmSCqmoKpuv7BjRqKv965BJGHwGK+SQuXYYGUZYkVxURCqGY8RhzDgxHwz6+B
5Cd96tpO9qbprg7CxsYXeJFxzykFav7/m3YXONRMx+/lO6z8u5+Mjo/wrK2AvkES
JgkJgtsNZaY++ufrjCrkyUTjOJ7FwitdGD2Y6N/p+35ShJnVUcMIXfKOglTThE6X
NZgcK4TZ0JMob3ON2+pVrqA91zgoZF16pl37WuH4/6hhJw7FMLMrAGln7iupNRjt
nQxr6IbOoB7CIio7f428M4OA8t7Ax5rxk7htQWGfGb+eqymnGqBVKqzUXXN1mozg
cDI/qjP6KeZa+oOMDQney2DczVU4FJDIKrOgESYFxmBOuR7Da6KwXMjVkdquvkUM
hLbsTe+2yfAwpmS6u0D1MDi3lt73CfBNzf42o4i/K2wBddbgxUF0lDQwwxRilfyS
NMiQJvrXOeIosj9vhk02LTDEFXyrG7hkXS2FAZJrGa6IlrWFI9/H1ZLqHTDsNVQk
Gebm9JUOWl+JmxjSrD31zzcyorGSncmfNOKKbDPTNgdhsjorzlNvXjZWAWjpvY/S
/uP4ofTeECKzBZAqpasGRW15mLx1Da50WUgMQy3tU8VB9EevbDn4yD3rQKWjMROp
oOhh7k5NxcDzF9iHa8Im7pIMWBF27mnrBJzx3kEmaDcn0Y9eSTzUvyyjiP8VUHEm
9tGF7mImuwfn8ePinumOrTuL346gw2euFpoOXsZsfe0fEcTHQupIttKlaMlIAkoX
2MmoqW091VS7sSU3uiK+cwL5piC3VTNaUYM/D3/P6o6m1cpwpswMkG1APUxF7ytM
wW0hQ5TMx6m3+I/uP5xFr0AQCvyWm76fBgPHKJtI81x344S1Nc+jrH3aNUoJ2FLm
fXhF4eWk1PwyXe7VUowAGqfj+Ml3IxalfcayHU+FdCN6kVS+3bFs06nTEVLURXcm
8gslFDkdHSC7uXg2JJldimqvqkAmpGZuhYCYIKAoTuY+7JWl02FvsP7/UQkWviVY
sX13fn50RUSE5us5V+d1OLRo0UIGt/iQZzC71oQkGUZgyoQbhAO1epWAtpMgg4dC
gmf8hxjmSiqDpsgLDm4cUbwzn2yIHIigS+yO7E26Umx1p51vo10JjHvSjfMss8Af
Bn7Fan/P9q54hc8SOHcPMd8I6PgLqI2xNK8DdmqqYGecWB0z2Ovynla4eksPxpfB
teC1i1QqjdrITi/332r+yCaRkhJtFyInOUYU6JIZ3XWjflctxvR1rqNHJOA3EN8F
4i7Rmt7lDRN9HZQYN3+xpPNJEKkoPMFoaSzfpRMo0RLYMKFsYIv/Po+zPrgnnHqD
zf5HH9xogTlxDJ3QKCfEqHuqHMVqLmOmh6idHAaqRfhaIcH28H94zj7I0VpdvfaC
nY5NGN7r+zQw/wKklc5eVPvi0bKHYZMXUzL8MhpJYXGr3e3cd9yVFqLdDDi+cUpO
dOpDGSlccM2x4ZuY50cJs6jGP71Kq62V0gjGHZvDJ6CKpwntXITTZu0kPFxKAA97
r0YWNIwvzPXA84VN1c2hVRaTlHyv6VHEE4v0LyaCODOy/1Sjc3k+xbqfGJUNCSFz
tH1RyUJyNyvIl5Xmll5u1oG/kccWpXqzhuUFPXMoBRl/HOwulalD4zFeX8c2sxqa
GhiTbU54H1ruHMGjw/rAN+STLj0K7gkoSVUoEqFwDTo5SvcJvicGDzVFJsMqltZB
zj8peGcCfQ5EGXm8FL0j3ub1pH7ftE4+HAMj+7bLZgIiuz444cjMHiaf0PApgmBd
dbGNqaBNmcdrbedCreFGEw4c+Sqb8uHwSJATITFq9IOGRwWEtj6LhWtMjRRm2lTA
Bn/ziGP/gWwFJvuUL1EpxEYDLgwWcsq4S4bVdjm3Zg22RayB6tSy+CWC9LFcJ9/X
mI4MPYiu0DsF7HKTUiwXb2N77XIHyuvsQPV48NQcOTST1p2989AKEz2f6aatXOVJ
5oSVjSLCvejcSLX8zHOnw+it92IPMn3awOgesDRyC5mKLKkIx0JkEXQnd8zudxxV
tiuBjUiFWfv2zQnHEL6NzarGOUGSVcvU5o2JX1VcpEvgEvEryplJEkjEtZAo0uLb
WJqgAL/kiE5oLYWT0+T8BUlEetJ65cwu2FiScqgdcFp9rHUUmBWTK22dO3YLDDeY
5+RUGrZwCz9Ovt1r/QdIbgGAqSCwgEO3vj0korZnAHgKww3HDZ2M4hRDc8yNjiOa
scSlen3wff63rfMMX6rWqnSEJ6k0LyOXylg80estc8ZNHQuAcFHAlH+x7IIpJf1P
0Dhvzfi9HCsTtjHgQldUVp0vMfU0A3xtZOpOrtx8Bvy8me3jXAvjPR8IXpkHwLH3
KK9SkAQxZbanetuZFUgKsb1+7Inw1dBfNfWwN+PJVo/hLuYM3Eo7yHkHGvK9aWII
iwwOUyovE9rMiap0MIRD22y0V3ma2mj/BEFWLaZStFmgEt4vLTVpFq2/itIquFK6
kgrUNgOGuq3an+0W5ZFC9L4OzOkTCGBE3BKNvnrEwM6Ya9e1wWPDUc0s2FllpCEY
kqkiu6E37aI6snlfYdWSdUALz+7V+BYYk9xwtA7m+Ew7sWu2fhloCyu2eZgsgMp9
WgU8Smb0t8jvsNsdZDBqySdGSKH/LHxUvHkdL7R5KAr84pQL4HG0xWy5e5RfDqmg
xfjEXHZ2hJGCK9Ku4rXHDX8ycC72aK+ichrAEFPS5qmDD7vXE6OursNZoJL+EgbS
csYIMwA3wbQrefRpOC7yzm9FEdBv3wOBsZGcTc0rqwW5enw6fAvxWmzUjyMyUgLb
LjSbeauAZghQfBDPQ2VXFGdxl0usXYZvqTfK2zC7YQm+fDzRl/MFuVinO7cD2U4Q
Qr89FgN0JlUBoyFOfPbsrHa5l3JRrBQthesR5f1hf0qcDWG61/mxeCx2GxKfpVxY
3iBlJ3UnV+RtrNPFojG2TwNjhfuKwUY/Dk4sWRFt036+nXdlWUYarvblQG9wpEZb
UTsLROuQoyp6a9mk4gfDXT/TRZ8Da7rmpHTdJ9+xL74qgya6a3lfHOWS6fWYWVs3
HGayvM6wgehpZaig9cffq1YcdblWTcikUH8J5x5P9L/44L3HEJF4NCjNy02J/9Pu
h6/w3b/bBiYfb3/WQTO5TY0BkDMzeR1Ga3ekzLrfLpJR54UgChasso/cOtK8DTD6
0WNkPzQIaZBtvucG5aBDhX3S2HCKvF+9de6zJ2F/JrM+8jHYS/UcSgo+BIWLQfu+
8ldyqzUroqttnC/rs+2Yp5KWqQV6bLbS9+QNADeaZrf+SQHvB/2RXXSXgqPqdmM4
hjuOBQZtLIHJ9sW3q/fDh584cQMHMwiTTMmFdEvak0+ksuLi3a5sY0UTqsvM4lV9
YuJigSXTB94Qj59VFkbssag35TRQGoWCYYiSY0ef9Apj/jEBF/fpB+QdNAa9cAlL
fUgjgu4hOa+xvyurlIS+jmKQB3SFtLsLekD8FEkaANnedsHXhhcxO4DkfATUrj5M
3+LxjCo07n6bMi12XuFFM9W7TX1H+TBMKn0Lq05vWX+vBoXdgDjCBLbci8To46JT
PJNn2UZaNnuaZDop4RCBdUKGXo7RZao9uEI6qGt+cy6M2kKKyvAXn61PfHo6PxLJ
Zpnk+eJEVfQFOfXytKO2SNYnKQU6E+ZN7UAFYYlykMtPldSq8MtA+6bP9ylk+k/O
TT7IT0Ahyyz0KV0BCXOAvl51MgGFbMc5vhOkOfkgy+UqYkAsBBvOnLR/rbgCjpXX
KUU1fMwVDVMA1U2BTaT5LrXxR23kUEJjz8fw+TNt+5cHE3NrLlmQU44LRCNZKq4R
v0coS7nAwt6uSXbWer/LBFHGPRNN5kOfyJO9WmpDcIURzl4hucjtggSSueRopmNl
I0WJUJWkxcDvCUbReBkTPsh+ZtwDiLjQ8EMULhYPB00VyfJgxlxpANCVvtlTIEZH
rh9Tmf9oBVW4lrIiOgoumYVCxnmQoYiyOH49UDsZSre4epDKSw/mSVyHw/Xn59Di
/3A2kBPHq/jYdYwehyDpAb/+Nf5YyhJ0oIwCwaNs81L6OqfYaAB1wwWsW2scne3R
lrVfD8mLK4MJ1eZoCPSrUzHSn6jNiDegVbIkvMzFxWZqlvMjBpgKeho16h29lgin
QUMCyAj8RMAx4QyrLfPwO5rDBA6nEWyuxPoZXC5nk95iXnh6u/fzf2W1XDLqHNYH
RqanFTfaJfO+QEwSASOVyJ/g3Kz+/wd842NybDE5BNQaGbEhXeapscIDHQddUXPY
7j0FY2crltM/TcaEQXu2sMuWtcjVEZBUk1tsYKY3tSrM3KSSIGBLryKWmxJQdQ1F
j1VIqzHc24sz9q1byiiqyvtwGhwV8uigEDDxfWbIRtA7oYzR2fLvyQ2nIBExP1KD
6iCTepBQ93Yg6K1JN2nL2a35Rw8qvo1yKYaY3tsHHo3GIsBkNrImRcmGC/faO4a1
bEjJCSKoSX6SBh8Mk1z1A2huTiolSBNGQkJQsz0Tr60wpjdqMuF8F0SMp2WY4ldD
YI8xpO/E6tJEDSuWWekVuZW3cRjAZLVCoyfAidL44KXPrTxUfTtMMtbNQdzHiOLV
i6r6lchE/m0d9aoggtNsjHwJDoCPDKefhSRnXLZxPeS0WRJrLltllnnhtY+BlcuK
9NSgRIXJ3mb4c58H6TO+VSfB3yXlyXs3QTy4MPTMkL13L1BU4yzGyIwFI2aH9/Lg
noKP0rGTu98Wmy0DcvCJZBbJvLxJvXhvyMGsBezqvuMjyvpnKuKZy6tXCh/jx2wV
SzOD07/bLahZ92UJ5bPNeipqV7890hQ3Vu5JCc19d3VWaVUBx8Y3Ssn7uiTnxhq2
slMryeSwJA3dIH9v/iW6aTqt0J+0XcEYOCJT/C5LYcHU/eFYIhMnyM9gD5v02ZL7
mz/tVL5yOWnEGkWEqL22BGh0/cpvEDvyOWFp+ZQzBErzRj8yip7RpnnWs1xChTFE
/rZYDR7r3UfeHDIaQ7HsERmqZq9e1uxtDt/YvCUSjq6umnp8DtYq3lyrUuhT1YWf
Qo2WHSYLC8/IxrNhyZuphNfvmNfGkGGlcosOJ440Eyk=
`pragma protect end_protected
