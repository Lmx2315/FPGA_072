// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.0std
// ALTERA_TIMESTAMP:Wed Apr 26 13:33:40 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Qg7OyoBOsfdOivXIdWI8JAccMzOLRNtCcVIzasrgENSkojO2ZmvEYAoSJv/6pt3g
T8FFzW5nocE9HeVaS9SG2FdW+JhOu9NAfc+jSkE9IHAIKAZ0PflGvUqRZMgHu3od
29GalnvmETps7WSbpaTDVY24KFX4jnhVl0MVhnZq7KU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 18352)
j3rGjFDrTjJoVtxIKzKqWNVOkjDwK+XgxfuFrqKRSEjCia2LDcTQ6nlyfX/MPyze
XusdwyCAQBYi0yTqW1YF0zLj5cwnitCsh1Rex2voonHTvfZquWcXLqnoXZriAP2+
ivkRvf6LwFR2nmBx3fzy4W2jo/Rn/AcPE5Y8jtModarNrZuxiMF36IlX/LdIDQEn
9F3+lcdD3gx8rPMv1LFv+QML7xFgEEVyBGqEiy61Vztw/Cuw2g99U0glj3QqYCZF
HBBpEOHBONtB7jI9WaA6qeOYp2I5XrHbfhIQM+ntPauuED09vBTv9dPjqSo56cwJ
HzruZuW1j3+m5DStxbvplRRXhz7kJk3Y/HhBjecgTzKFCOvqbyMJNUyOWEdHtEi2
DtHQlpGyARmuRG3L448mRtu9sFGMG6mEFa5SIdh6A53x6qKvWHAUpXAMwTU8sCU0
6qnMXgFr2s8F2NzCxhpcHty6ZqoecQYcg/Z8EsAtKMYhiLq+JiTGxs8WYkZgmN2s
l9atzd46asYmoYJ791q5n6Nb808MF17FVXHUjfe/XhjylggOkwJbmVNYPEY8vKjq
vQk6N3ag6PzMMjR4O1Es+iZiniTM+tYdGQ2lrUBbT4gmwdRswVEMBlQQ/zlGKli9
syhr1KTfG1cHG5uo10TlivRh2rZOuuTqfrbPfqLSZZPDAdhkFfdN3gP/ywxQo5qR
4AIZrX6scmYs1PspgM5QMeroNx5EHBo5qxDwcaSn7RVN8iCAJHiRMKmeNT6FCZ5m
UkHasnHkQ3kRDW7SoTJmOVX92Aj/U5HSd4yvOPg/wd63qL9LVQrCJ6SVBP0EB/fJ
5ORAK+c9FlvXhhDhaZwpyDX9jLC18BWDc7f/ZQ8cNMp9hCJwKyPUK3F8Bu4uvsaW
wr2rt97jRP1iMHCStewoqsYvu3opYErKU3WxurpFbDZ4F2IEkUxLYTJ6spbNHQw/
QcLi/nPJo7Jv5yggVeZBQwHYMJjOms8X0dERSRykM6YN4qkjuJcBhNkSI7vstJmG
IYW0XZMTTDjHjGTgeDudbsipfvFuAdwP6E4voCfNJcSNIOiEmBCnTC7sCWBlfKnf
LHQXOJt8QwKDbtcB3XZAwm4ek8m+cwvI0CYUlGuyOmshtgjgJhaA6miiZ96Da1x8
3WF7Z/r8GE4QEvdW01982qOSPQbp5zRsSz2dDfiWDdLbaGIjRAaLYxT/thpcDvVp
3O4Q4mpWxy8GTIpPHqQeZsdaLBG1kiuOXymcBSXdTEc5h12XMN1aQkkf1Y0dSUl/
xirJM1J82ft2uZ8XgWnNQmUkZnWjH7NwUn4fSOpAJjBaRcPDifQoy3RGRDmVTTMW
JEDH3Ufe8qeqkPc60b+L+eTfnF8Li0E8Ht09Szpyhofd2eHgd9wpQM4/6+ywwBjw
NAPxq/IqeTO0vAokzYfARRX/7yRuOrvR4TKmzQ6Lk8nFzlF3U/TIpV76AwrI9+Je
1zN7rRRUXsg6BVxJeLxtPrYHm8SS9aoSQnmDeLOpPbHmMvOnDBczyVAgwlxUxVb2
yHz0mLlXRR8rb3AXpVZ+h3bjBeUSLA43Q8W4PebuwWrSk6YrIxi6h5grNHmNOLqT
irzCNtafWPXx6xqCabFZYyc56TjF34FETYHl0mh1lbHXiZZ1wGhXTpNocB5DKkaa
A8LLJB1ALNkhevvMnkmKAvL6t3dwTMlvKDEI/tMbQBwjMa9Nvu7SzFd+EFrVSN85
avzhtgRaDREuDJDM1pBofVFX6wm3xnNUXrLdH5uoQXv0M8RTymCKwBdpduaj0Bw2
cig6E6OWc75nhzdY8vbHqLj/aOUTDjfZI84BX8PMbiZQ1eV/4ECeCMqCqksu8W9t
B74bR1T429Py9NRPummBbRg7W2gvd7EaMIfY5da9FtzHwiW6GadkM5d6B0v++fKW
ZzcYC0zpDelI8hTvjQWisu6BCLq3jfhTeHtO3v59YrFklns/0+V9rHmWRf19Gykh
BtDlK6t4bP9NV8kwljyVB/iKVFUZRM+7wowB/nPn/pCsx2X+eeVHQrYotKgoeL3m
siYrW8dfE8hoJx5SrEFpprbu698CK+KZDC+YIBY2V+2VjnqdTTu7ouguLhQJS/Bo
1+8mEpgUX2j+gJN97oYt4NZDLh0HnzLqF0BG3+MsAeOhGtFPqOta2H0SCQMl0Bvv
fpPCxGgmwAfg9fYj/UE4i5Xo1uWelSGNBi1muqwmwkpJqiftihLO9Xupn0yrOWUN
jOz/W6L5oPGepnst7v20XCXcFmX7OM1F2Ui4XwCX7VVqby1BUr9I6SklVnqbCaF0
tln251ZRutMjnFDd//2F69sFkgIoWZCDruXzuRpFRveRzOhH9SyIfs4RxD1/QRFF
reMZx9pVIYYPCFgMc/pRgQxUVZX7JCoL2ttMnqnaNzi/S5lRE9+zmgDyT2aRZTmi
TKnZ9VYmXdBd5afiFSTylHqvwN0+wPajnkQQmcEB2bKhNSQPJzy53izo9MJmpPkR
NmzgnV33Ztb/HDtInEKW+cuJz1369Tu/BSvMJa53ywuH/mJ5rgcYgy92/wYzPjZA
QF09Yt4Eq4m8QPnhw+quwMVESOvTK7zWKKqQ47zqpMLNNEF2dy3OzClZI+FYYKj5
J2CBfWOz4sKpaTkC9bxCFGLAxtxCmGY/f3H0VZT/DPDWLQyeNZlknzfPcKSjftHl
cUWQg4DR5UhVTX1SNSfAaJbI7oODGem374OI7XeKStSWgS1aJoqlNAceU2AdH6qz
4C6OkWckVIlEfLR/hMy0eJA+EQwMqWNwAVh0Wqe2DFWfoNFKI2bXFvu7+1UrMlE5
L1jqRaO6q6JJAT4+44H9VYKiZKBcd3xW0QF7PV0/xIJ66kVvsqPFXAStN9gDrFnY
SF5NqvEHcYMpotHZ/wqOFXwUdntpOuiXwY49s678ITv88nT3sN5FUUYutMsWgOAS
BYOPOkqLvHfFy62we+M+t1X81ExC6jNF5c2V629CusrHQxP3c4v0++ZAPjEKRrRx
ZgLA4wq9asOCCM9DrKEXdtZF6GfF3UvyGPC7zBUKTlJyoCzrCmvHEAb6NcgdMlKV
Onvas3v613N63/APhWCZgbxcVGdl2AEAcdYoxGgGRohnd6+Fkafmooe2m7peicei
wKwaFt1nRH06xfHX4/HsURK6YhrZJBF5YnO46C4HhKWZSDOOSHFh1snOWkjvJdxG
0BXdfE0DGZYaBiRwepof4BVkoK8iqhRmefNa8hPAswWrDc3pIgPQGyOHA4uDD3Fd
2yxSlrndtM8LNPk/mqIxPPvH7jSem+yASKCrvPzLkSybphH89h1y8ASy5Ntfz65/
eeDb0xZoBt0/tFgDNKlxJkyVTv7u9fjsyQYPAdhwOkgiSdabwQIPZdAvHjOa1iX0
u/Lknj7HX3SiIvB2ujEU9Dhj38zKdu+ZJphYfUGU06S5XQc022WCZS2OeNY13Fa4
OV2zD5MR6ByFs2TXj7xmlmmWNIV58eGinftvcSFRt6qLTQOl8uCs9hohMvUMWCws
CVHYul5fOM3OhHxR5QrTOpLOqWeuVTr7zs9P/NI0HkrSorcrqAEt4HvF2G3C2gE3
wEagb72vc0vrZ86suoQBUeIlOwGq4gZeKxqvxG9OHgHxjFuUwPOH0htt1tfQzbe5
D3lCoA0Bu35Um52CNMHso4qQQpwSB/uGrcJIHdq+Qp6lSb9TsgYzT6DKlS/nTVRX
7VILVUbE04cjpQ+/AycB2I8SlrVY2OIk48Tcq96EJB5UDeH6WIm2AdNOAt+2KatS
AsZ5TUxYlyJ0OU6yNjPJKFLXtMTFH4v+EEBHt62VIC9D7WE4IHniQqSgzr586JWt
TpB5twjei2PAtzPCsuL8vGVjWnt7c2unUgVHip5rrzjACYOIbD3G0UyC12ryNi+u
ZcXxNyLRdbiEqqfnINbGzTYm9LbOADej1VqHf2UTOtfr1Q6/cJX4Y/PGn2WUJMX5
6FKrpcnnJi5ithSAEN5cXQmpMvrRhnARx2uUjA1xK/stkB+TYZjbsqOeDlmo/J2j
HFPctzpd3lXxjCXbXloY805qXT5sCQ5rKV4Ig6+swix28/MVQJDQoQT5WsdkieMl
h4J8f42WUDV7fsrPHLoruvdyBNVuiwAr4fAg5JQX4Aea6oMrtoYm1jddr08ru5Kj
jhuKdFCsoAAIN8jm3hBdChUoprU0DB49U2DgCcgc6P4Qv4XUg+Em9ixCQvtcb2fv
SI9d7+5T201vb2kQ7na6JhiBrPiQ8UQhYOpOxaaLXAnZmbvO1tczHBscnDLzykjO
HI4CJM/XeraFuEG2Of177gi2EF8iHm9fJ42wriHfZhgexCxNYNqPd1lncRCIhf39
J1333HEhLMSRS08rx6svEN9OWNeE7jVqxTmtuZoOXCEoFp65MCsbGrxskUEHoGr7
nYfLXMkeofpdnvX71+IOzOJHOGaNQnFLLCo0h9msoTkOPzwGHshPyxzPU1x/SBbQ
1BvP1Hh0LBPxLeJjqNiAWF2w1A0Ke+atjVf+asGERcumMbQxMq+FO5VNU9TYsivS
UpMy/eU704b6E8zbQl/yB4ztm7ta4Lx3j2+ZEEplwhqQINYuoSJc3sZIkU1KxTOW
vKoqZNtVv/odmGDLjG3teoRnvg4K7+LuK7QCoHz4A6dK7pJnFJK+ZsekFCeRRkxo
a7fK3nflVsROcJYhwRanm4m7zd44dbsfN+8mBgMcuEvOIek5MjmvOGcIXOatoSh1
TXvAWzWd5dkMpg70ohxi3yTcr/p0oLHm5wtVL9SvSZ6tYWZfkiVnT2kmGBxnO8Ot
thwtJI67QMQAlOrjKcV4/xZ0NRAa0F5zKqzXftmKVfYqFmz8IAmxVP17jH9by9K9
pioF8I2cvGUBxImkFIXp61G3op1J/eoNqLWsNDAlOZjgaHa8T3x8QFqf4gCkkK/f
C378cIeO8rOsxo/ZUhT1bLAwY5uBFKvHfuhKpDmDnSKcTWZulKRLcmIUsa+dVBAy
2Nmqayl28Sk/JeJrZU7Bcc/sAhOFU5MbBJFSRSTXihGUTn5tLUA4bmJRhptHp9ph
0mRAQuybGP6a9cYOP4vUZiHZEHmpreFcJt7Bp/q+YoeNDsxkDcvWurArTo930JM5
hCt+c23Nl1MgMq/L2iG2bmoss/MXHyJMOOElEg8dToIrytQtq8iE7pod39j37MiO
ib4rYRBVCuNZOLeXBieaLGT9cH5lkfksMW+aRv8/5PnEYSuhFpcWU0yH2zlg1WvY
sV2J0qbJ+iREDi+l0M11503Wf6P0qz7S8uhQFPleW03ObC0BRYcii2XX5WgzOTib
+xn90G6ACC1Shpp4/xWfcONQRnc0Z9uVUgjsIZGT+apqXMzxbdxDnACVZD14c9js
ZTYjfGLto+8PDN/cYLPDATBFhSDZc4bRjHoalJIRQswWwGGE0mDWjNg8hF5/MLB/
E62pjkbWDUOVj4kkbXGggBpfKJDUJ6nR6VQXfmFg0KIOqPavhcUZFaCUFk+WV98W
KDzGdcomrV35X9dMjliMewrM6Iq1zUfpRkqCE1qdODkQ0BrDoVLdb51dBjHnIm8B
za1aunL4PesG1s9uSZkXQL16re/ZwpolYHPWd3GR9KYFRMg9Y90otK+/QM3cmsMC
lMr82VN0TbnyFdk/qNnDIrGof7sfFtjYXcGXzlrLoHRMIIYLbZ6Ttwp/Fjp8LFMf
/oFMh786Bl3xTQSyT5j0VRyswwAMQ5jhtuLLj3rHozDklbqldOe6A1YtNdBjsoAs
rdcaZ51x0zLqPg4Yb7FwdnRGmzRbivzfFYXtqAm9/+EEi+imu7QtL7JyQbRVO/G5
J1mjr/j+63Buxo0gwDEQI07n+HioXrWh4nlHZbD2zBn6/Gp18kONQWjHcJd+Qn8P
7bgOC40r1ODpNjTa9uOVqx7jpGwR4vdHJdH6VMQnmktf2G8KYF8gCc/3qQDaHJNe
HW9owjWCGo9b2yc+sxGgVQRHk9Gc48Z8cIgZjegrEchlET2Be2teUPLg4TPSB0cU
Zq7e1RjkxL4cw9ttPXvcV9BjnBmk8EShASVWlE5LMGLctWe4S6UT0imr3dKlaVrg
7AvYpnp70UqSD6fwF2Lmxr34z6tKyDAM4/8H+sgIIMWmEr/wJTbIKbKxG1/10BA0
uLDBuR9iAy7Oeti9UC4xXwiD2SlSm0+XFTIzZ7JZz9c9rnY/QwnxFzLlVoItoe1P
506B+8AOlS/nmplL+oo3pcFLg4N79Si6fhABu7Ehc2qVFZ2xGIZuSo08Tv3UqoyZ
nhREY4gB7lHHnstmWOPQNn3DADDFAADv83tmHu3OqZjnPtcb5bHK5XpgqtpN75MU
k0DdaOvMJEu2ggwchiUy1+jnK8E8YLWFVjjx1cO0a+SFsyFVIJ+mpy6qoaciHRyw
puAdF8nKxpcUIBGnFUhep7iCpAUdHpjf2YieVklMYJ3ku5/jus6lwbSsZZstNweQ
BkDslqOvwgyY/pDq7OVyXaI5a/UpGKqINJvPcwUvRrOrYIMBLPIQIPq59ca4dUv7
/6W0b1gc9RniFw4ZabZzlrT/4WkJvAejG+ns62PuAgdYq9A3SoD0ayHRZghkTNL9
Xf9gdZjbqMedhw1eayatOh3OeluxFiofvJ3vom+TJ32AtHNVBelvrRyHk6BkVaqq
NwYKWD19qbFPVznM1hkz71pJ6FKpyIPMte/AkcPuCF+/kj2VJL4ck3whToAT4G5V
3EYJmLbSd0xa+0R5/xNT8yWvr9Fv9yWF6ki2BSm5WV2cXlukn3vXK1OIEokNlhSv
WSdFqYM3hGpmw+JEsVVxRtg437x+hJ8z6Q2J9b1N6vm+XQwXwE9CetqoII7+6h6X
8ixZaEIPjx/kw8KvDR0n81UoVuwB75ItHgpDgIQU+/jpW0bdMD5EjIEA46klF02u
xKoB0ZML+CRFJ5zFiUXI4FryVQlusoU9OT4YLC8Ng3a4Jk90SMR4/nf1bofSLTBI
XXWKiy0VNastAIr4PFB937OF/EeGsf7kjFk0n4PCfG56rfmkRmHMi2U3sBc+mBWc
THd6eCbGl0Wfxv2ENJDRpjWxzr0v+n7h3CWnRBgNQazonP+Gta3E5ftK99qHtGWd
DVxcSILnpbpUjpSzQvR8MhVNw9V3TwFRv/5CpA/EbCP9ungmPwWsVwkHG86LKiBD
cEOIkK/q/E3ANH4iXqfDJNQx3egFOwciaoigN3LNHkwYwojWFvtb6ppb1AEqVYkj
mPOoV6tdlQKA/Xjw1GIBjNAfoVy0wISHg+3xrdU+lIc0nsDDZjtsXCj4GHNYryoj
Z61Av6DxtQVUVoy2Cg/2TeT/+KgE9yOptvZo0xTlrnmPmixFwuMLxekBiijGYocE
+oT96nvj1iBsw8PhUpyspBtaoLlaLl8TFDupBSrH4Dg3R8hp/OhP5N/EGea4B/La
dOGA5+JLNQX8QIQvdIL6n/RqYT0GCXbYBNcK21clvZu7uVnY9LFojspToYiVMohH
Vq3aJAM4V8jN5TGO1W+tqSvKKJibRFViJr9gFKZ0SNwAt1xAkRqxUkJ0y1zAMUuC
tkqs3nisazZfSR05FKfpXeSY9sqy+1ZjTrX9GnxYFxNlOK0kfICkiItub9ZB1t8N
KwEc/MATElXvLHNiqMQMUoDeBbRmgpmm52mn6WR6DnkW+/PYhkI2r2BDRSZ9Sct3
FsMYYZcLZj0rs2k5PzIxmlIdE1IuJkcu3RbPtTvx+mwFw8Xjv2UBFCqY2q9hdniI
XjRZcMwrzp9Xbb4rJuO7Sw5mL7zVHI+hshecXb91zAUZC47/k9KcsV2Zsv0xs14q
BDm6gvzpk5lpdbZ+Lws+zn9u49NHv8/MFxSDEzh+dhmTGbr1As0SgF7aiR/Aankr
gtUEOxM6JvBEUdeGGhU1LnCv+Wi/J18iPrAkc9r0l6/8YMWGvjIM17S+bs1hRmk1
jWxTPW/qBTUS6GM+bMgMq1iew0SQ9BBf8Qqx616UgFlNaF3vg0+FoeNM695271/3
aCndtakkvf+00Wtug3EY/WpnuGx0l9ApXNpJMTfxhE+DeNKgHNsi6tfZVu8QogMn
ROp0aet5pPA7QdS4gOGB3pVkhmDERE3lt2b/2q9e7OPktMcyf3cWvgTb/6gASaZ0
XSoP0hBDuR5q/vl0+BCwnK7eLgLqaMfrbkachE7r5+ww0e8ssriH8FS9dDYf794f
5S8Klrqzb5kcs9DMB5Tjk9Oj0zwEb4Uf8KKMCN5c8lYDoJTVodYdsVhUC8WDb869
CfvfAgjERNCI35gALbGnFkZon7p7dOu/ecLA98UwhKcFvD/hlKpmuxgveKWSp99N
rJvg/o8Be2Si2wIRLD9iFiVtSAXYFRRFCUD95ubWUEuZOywg9L390d7DQum0ag35
oOFEu3GZ/ZLqgl5WutWX/q2y9AatL2o09s6+lsBmZ53tDnPz8eVTI2sQxZc+iJWq
cRLQ/9bUbqJHVGRpUwhrivS3XftVh4BZobkUq1xNx0o94Axo4n6FSOaW3IX5WUtV
A+63sHgI3Y3Vtg1UaJ+QoOEOUpSKioaoiNU29ctcpo4Ma13wn9EWWno9DOYuNq21
abj0QAcZ9LAUKiAAodvDUW+qu9HQz2A7A7qJKkWGug0/S3DfMf3gbKllPqmEOAeH
hoyqyu1EbG2YKr0kL8rLyElrnNXnjSopbi/bJtjQ4x0tCBObSWfcJCSp/xlpMXDy
Kk2xezKyHSpTxA695YGRgyQ8EkOHwiiJmmB+Kwcp3nQHdTyzNR+tXc9gf+4p/vue
H0Yguq3cASP0UvD1F1ha62tPKX+Mkk32l9qLpqXEYqQzprtpFL2okXz/o9mv7MrR
dxSm9TRzs1MrX7Zq+dCldiF2XUgA/UZejFAbEW7h0RwF7h5VsKKcOgxzHAT/v+sP
6n1nslEDH89RVZZp2YdGwHTmP65BbUJkFyCwmGPrX5rZWHPwM6jbEjI2SN7nm/0u
DfGbAA1eCQcAJDmPit7gwvInKOlY/oedWsUzijMjyXqRFqxzojZUuW1+hYzAVRdx
cABDyIH9lYOsEpq+PLx7HEV1i3QcSFdkRh84Ba21PAo7h/zCJHzjcVEEEBlhxKQv
T3kyiUGD1xqeabkZiT6Bm4SBowNv3g8juvCttLk0vV3+RkJuie96ToWXqIyDArJJ
k1V2D9zA0/fXtj4wCGSWkdsiB4u8zuV5oEJcXL+gAg9QyecH1Zo+G9m4bxg9/t/U
qs5B4zp4AbSjjDLdz4+ibnUZ3nMZxPoapmrmZumO6nuh4jkbbDDzOj1OixeV5FD0
SQp8pR/hxtLaOzYkpURp7Y4/2QRIb3pcs0AiEmLV2tyhLWbNfj6cHRVaOfJP1Lcn
IrKjgKk4KMGLrzmHxzf9zw6DoOR/jpXCgsZs1gTGttJnnn/B6XhmIUdPWEyq2N8u
943pXpzeY/eukH2lpTvNPVK5rHePHD0FM4E81aAfUfeEMoteQl0gMum+rvKeFX1l
gG6S44V/tYXfQVmCubWBEcwjzZV/IvIo9+HueFhwLzVjIbY61lOvYc8aLPwIdKDa
SiwHtkilfNWwjNkWZSaqfBbrb/v4AQaesNNlKwkSSQp75NqadqORWCEXjh2jpRHo
yP8Bzk7heZ9P3m+9Z7WuN09PbusAdioWYXrt9B58gkDA+SMPR0drikQ2sw4dYNzJ
aMeLiRuoIeqVTdl53RH/K3hOIUsydH8J0Lsg4jZ1t0SddyW25WOqGONzlojfOpwI
oi5i6TIDLEVtNLz4heLK+zFVXeUJbSp/6aBo8qKg+stDo8pAUDP5Pjcvv/bzAJay
s4VFHPqWG2/r9isOc66O40nLlEbrPEAxb5/NWzattZsOVkkdcifwz+tT8FE6mYrI
p8tJzDC1Yh+cvgEYmBsNr/nXyN4UpBfCcIxcps8t5yMHELe613JzEz+1n9T2u1+t
5+jb0J2AxBmydAafjd1F0zuzFUT6Ey4RKHHoYAdOOU6leB1CVjktlPFPIQkpG8Sp
pYl507BnSluzg5yLuEZ8xkg8u5JZmy2pQ8J7N6S2SOPypmKHmT0c1UyP/I1HJ4j6
rTOuZnr65JOqYeuccwgKwsDPbhxvs4A78Q1SbqPK10lJyUTBG3hC4OxHlciXtT36
Kq7x7pnoamuOfqALIRamqXdp5pv06ZwBjJbRpwA3vTWAwftvRpfxUhX1RMgic+uf
JTOjzS8zwAfV0XY1/IopdUXD848vZVTFN8p39myXUamdhF7Gdv4r2Gnxrkh7aLUL
qUZygvJmvXOvitlfFIey8FqgJEySjowcQIoUlgB0DYTjEfJWWynxiHcrIUrFULV7
9tDuSeh/eqwGMuoK4dcOcrWSW0oJU1vjvoZ4oSl6dtCDqIgweReOlMj27ZBx9TTL
Wyl7ibUCLQm+8dbmZzYnyg05HV6x52qC6u1sG08X7NDxiSkUOx8u6WUWjJ4LXmG4
bdxIwdJsZ2PFLqmIFb6Tk+aCZcFWc1ZaPLZz766mrTnS8O4dPTYia6ijQTdYAPLl
qCTygBLLAHEXKko37q60fmfR7WrIl5fXuKKZUAZ8cJ5GINwm/Z+vsFsd4GyJyT2n
1J8f0TxI8Rj/klXAr+NXQJa/xmJ8FmZo4mr5PJy9u+7emaRCkik58WtIlSMEbzoc
+5RyvBCt7HcfjLkU/YeD51JzXhEyszWmaa/vHYeUcR7Q/9fXO00MBwbw2UZG7IBq
zgqjHX9tEehKJBqDZf2swV+EhzG2HKmNexmp0dQAwrR0wmwRfRvUKOeEke2/60+w
fKXbFUAipMvyxp+3Xyl0cnQpBk3sn/Qf7qnvCoaz8BhfcAzHbtU2NR7gniaT5Z5S
7ODiFAR+KafLD4S3dsoTgg4NcUkhq3q26nDCTnp8VZUxFA7dwL0IM7IdA06+2wed
Ulgiu6D8OYOh0oZ6f5KZCyTX1hXu0HeloQQcgc8iQ3yWojh11pX+yBreTfkV8m7Y
2cdiqI1TuBZ+1yyPMQnWu2uGCX79Uqp5OeGMjRMhoUxK9RBcW712HpJuEBI0/SaS
bPhu21Zz/dWabQfl1HgdA5Cv5Pgz7RMzaEc0GKwvxI7GdANbOS9xXI9z3nb2d8MY
UsOFn1io65VJhGaAc9LRszXU5tPo0AtTWQab/sAi0ETPO1CN/E5/DghuU+9YYdcq
fd+Nfvo3xtrTaIOxDF/YiQYM74PTc2BJp1LQ7++v5s086HDwsXyNbJ3gEJSbyI9F
cSVAgb+OC3G2arZoS5X+aqENebAs8iPNGeshpQ5JCrpruHIcL4Ghwj4nPGuJtGIE
CR5odiZ8mt2Yc2z6v2nu8380JCCHoVyCeARhJHgMBl5M91exWaK98wMXEz8+wfM5
UCjpPgUkIGJ8yc0vzHlB1pUDK2K+7hoTjEjSlKvbfKBequpi9YQNMIzUNYKuMJ9m
NvJNKQ7XiuQ8eYM62PeJoFYLT4P8x/syoFN/tnzBePm9ylLQda+xfhem1yH3Hzrf
sgwbQdSy5Llp+0KlQC+rmj2nAkW3gUjf7HZnHsw7S7OcFGvfHU4BdTi1+mi7g5H2
MqScPaYo2h96puKSWyQGHtqXOaR4991hdloVviQth5Ahuv59+9ECHFOi6afyICHo
0bvRbV/go63DrldivS6YTWVkfcZby2zmI3b6xO181mpVyuJJF+o5YiRtMBZoE7Ah
sTZvqqkWUlTqj/1MG1jpxhl1oMmLrVQIX63I9RffW/2h+qAHHKj4wBdqmlvT0/AU
neav5VAaHB5JVMrP2JrueF0Pzacr+9Gf9z0yxnYKvGrOjStZvT7JRQ7+Uze9fjYC
enqtsZ3HgmfA3Gv09eyxwQStVpMKCkaoZjw+pnreN9KOWdV0rq9ZMk/YFGQAfF7n
A52tjDQrUSOjJqe7kdvZHpS2YRhCDWyhj7aewXMjXJq5XVznRdfFwIdJW5SycGnQ
EIhIdZintNN/NOhD3RJkN0ocP97epaSs6iad9UpvEG1isG6ViL9Y8MnOAdjtyX7K
JjtodDp3lbKxrqCKjn4R0fZCbcUACj/aqr1WVo/Q4UgCNUxGZMQXH4jkDJ2l2XCN
sScSGPjd9QRCxXeCllOmK2MjZ737bAvl6umx+E6rQk0riZ5P4WvfFZBJt9RaQLh9
gpCq5+/hV7znE8EfCj0Uqv28OgdNs0RgFaMM4eIIvJa8Vf3FUTZkNmiPK3CN7dRB
KXCQYOfvlNjNA9XF8b90dMuAjaUuYfNiIHoOGnUTy0FJwdkTRpWoMs/T8uDhavzs
Tdz/Rq8dYKG48wrm5yDMlDbYWMJ+HB8TsQZSBpUbdZX9p5AkGpAY1AuVA8+Uo+VC
7DL3lQ//Owx0zhKpDURTFlsR272/mbRoHIRlcT5skybK7cG5jYDaqpZed7M/MeXa
cz+iKuWX7AFaZppyFOBbqe6MM3561x1Xi61MCq0fu9DY+h0/JYDQjDUzQZQa49Ru
vqCCFJ2j7S3B0oqtHi/3Fc1A0horYVfH+3Q0ad4LboVjN+IQSWoa/J4NRc7auOI5
rdqZTAhWBz2JbyWZsvj2EcwtZuN8glaYPte+8B/xECbOdgyQ3sVwIkuT94exvXK4
a8kKFaB4H5/FArKeLyD3j9njaghXELag5wdrjUk6ELWkbohn4UUvjsenzeWR3eqw
4WsH8kzNaJfodvaAStH1rvVhDHmLAj1UPZuFgfCBnpyHqf8eM6mtreb7eZewLhuO
nENDuVfyzXJv26/Xjf14EwxPgPrbCT2KOBhHtnhNMY1ggvdQaFUiQJxg11mDk6AG
QgyCecBpbGaxk+Nrj3135VWz0CrlRbjSN5vPGdTq0LaCQOkoYI+xIJMhwLiWwkp3
ih0nF4P9NWteqwztBLdrbm9rrIdvGjGxes/WnQkfs+13gV8kQN3tkReZZvwGxtxx
h5xNUsM/FiU0JGqMWM3Ai1qwfPSwRiePYcdwtotwLN5uNCuj25MyDrDs31PaPGxS
7sRsEObV7qyT4t4//fd4CTWBeM5jBsIIt3YnOFe+Dtx9ycwQhNsYvybe1BJasOvy
/3Lp3H7WPNvuGijg1wOd1WXcokZ+Y8KEBoL7QDDTlDIHm4tGxSmvJB3f41oeUgJ5
AAxGJzu4h5CiS2HpF0OHGVJvEvcYjH5PeXRfANTnmErvPh2/ya4fo8BsBbPmXQG3
QNLDqq1Y9XbwlkDnuKYp3YjAQw/g2lfuTjVJVmo74SQMPIX3aG75popYJDP3Sc6R
3oTJxGTJ5u0suX4xp/lN5QbboCH2l3EafKmzMbuxOy3mu5xSvzCzDJ14PA91lNk2
v31OtYqMWOnSiWE/0P/s3OzbJVIdI+g2kUJQKwyv75xhJreRjbgTUpP0nRmu7XGe
EbLxw98+SJDvogx0fz55BRnLiOBofxVXtcz1ZVTQUCQMs8/ODBcedTRnfBOEBLTY
kyzbZSimhCbjJ9P8xFDUG+XFbuPlj8p5JdAu6/hFTAFAjRt1iJ6fzPUtR5cRcr8X
T3hv+FEn5XDAo6MiYvO9Ukh7JWo3De5fP19zn409snkoPDeXsRlO+RMaZEWr9TXl
HLUZBwjrvkVQ7WkR8vqiM8C1l3OgWdPSsn+zNpCRuxX4VEbJlr2qVMSFpkFRUUkW
O/QrSVAXxDecx9kmG//eTAd6+U5VXWXCosEg6YYjkoT+YVNCAw0K+b+F8IS1F2jr
BCBu9rhxXcWp5FUZZ2F0x4sUZdK7oc79vV/BAD+rE1IB/sDJnd91r/s7UfrDDPhS
vP2t7gRPGNeWNMTWkrhigRHBz2+Osvl9rBSDsM2ulfoCj6Qm7rXJHsB8DQboSTc1
piExGTk10i8Hh5P1zsQbHlhk1vTdIVfdjmSGxeTzk+KQNCHUTGJQlsCGAsAZt9wV
B8p99pxp7MB7QyrnJKqFXCnMt6V3IRHzQ3Shco1XoAH2oNy6GgvO+TRJ+TWhJbXp
qhlCBtvmFvqRBDhqOuEtT5JFPq36xqs39muSU5klNaux53RecnncQ870SdJxpRSA
3h54EVuZa5NoXqH8h9jnetAhvQZZL5RCbicki6yeWH3zGsYONPvundQdSbJz1kES
9+Qo8JmXEMMAYN1cU+QbO0Hudf6xppBGs8W3hyTBh7utdRRRT4yRLuoQFgse4F6d
VB2LFvVaCxqXqbgDgZRTOEBUd+h5m87SZrtL/j7ykd+RV45vF1PEOEUlnTepoiNq
4Im+A91jZxK63QWPmspSrj4sFDodJc9Ogm9FAx/34Uf8hGoMrTaWZJT3wAZqZF00
Q5OOsvfslGMEssUQ6KNYfSMHm0IIxmm3P95f1IviCU61eLhgfOr+/7ulu1aY15jD
lDhV6Q0YR5ygSO4PzqGiVtGZr8PNThmYODnjSqW/Bqgxj2DFSEHKaJVnVXL3Qzs4
713NKl/61e0YdXVNip5YgfYfdWVDprKwKES05BEpL7nRMQJdphZ3vZbv93cs7fMR
fwsRsbCHI6U/1RTKWeWbAoui7rbaXn+JUuxAkgLUAFRiIK0SI10gmEuJYaVi6+sv
v5g9NoByP8jvY9v/8JkjZaxyr8sQkveyytQFrL68JH9GB2PolSbXA/2nFidwuk/j
QMn6vOX85N8D8o7bjQTGLCCDPfDR1kg103fU1sfGu45R+Rec6kO1S/PCcInTtrfN
+zLUSCLVbxAN/UUf7Mz17tGWb2oSY6Y6Bh/TZSHU9buRUabwjf/T6TmFkvL0z++u
Bw0X/IgM7ddVprLb/D80VCX8KrOmtvwwg1jNJ4xPXlcevywnkjasEHUQubx1pBT2
JuMxBDgzerX7mutbNisqmboChrBZ15gI0414vK++i91Q2Zik3vO1N0PydaSuxGPa
wKDw2rEQorlzNvktI3FjhuuL/ur/McGnRKtPLlbxo69mi2kJvN6W8VDJq2wUAljN
9LG2B/iPXGZbWTjqLb4tmhBaJMwhvIRSfF/nMI+Ps9sPnQ1sudNs+Kt59dSvOMwh
wGuPDID7NdUU03gk8so19AqQHrpgglVud09t9wAI5cTtB2wzfdERNGMaQrulL/OM
VXr6BwNAN02DmEJoGgwG85MwOIfHByuMQ/oEpyTeWLK+pdZYjnJuS0TN2bzREDu9
0y7rsyQ9Z5pGqM5VO/TaPiLTnR5HRHAzDRmdHDsZp3STbG8L1HxOMivtMznyqSbW
Xu0DTF+Nz1kTRXAkLt6i9ZwQa4gLEidADCxOT5d/njfpZ4ilVyWv7MHd1KqVRQI+
0ci0On7z8ib/bliyCZn+CMkKe6yjyShdhr2hksbxtO/FLHL2+s23i1hiFYm/47iG
gAU7bQSisz3Y0Inh6SjsXUAl0CWBWaP5utgYsQ6JWXXC3GpSC4xn91zh73qoB+jV
Ec17/cCxdC0ByZdKVhuF6/1nNDLyiNMv8HUY/lFDsedMfgSEKZygyMPLS1qN8vZC
rOsub6/UXsawUIjI+hXy6z/tTD3gGvQAj408oh1th2Ki8myJ5WSWdlJ0suNmIdxM
UeJRnhS4vY0EQ7DDN2YDZUf/iFhbAOy8NH3R5k4RJJk6WOurxwYtitXP9wIYH8wz
N+JXrsxI8P3jEi3cmr+7rPHwt+DSEtAx2tNjT/7+AE8T0+Bd2UNaxG90uy5pTv2z
9rwOunwrCYzB1JU1PtbAg+7dNsybQOw1Oj6lupS7wr6hKF+74hsq9E1CLby3a8BG
z5HiHjts8W/U03KBbI51YmfCJUG95q/+46yPlKEbgIgfpLgsSJi/tAm7S8TxXeil
1eyaFvOSW4U7AjpwckmrFR5BGzmefT/oQIpcO1HslxZsqiqV68WdKOosuUuObVOy
Hw82Rg9l1PxgiMFLwTM7oH0wnnqQxKnPflU2ewGJgb1sBbkdPIBSnHKz9AnPdGC5
dUyfRMZoTMPffT7khVpTwIChLBv22MuMNpv25e14fjiyzey8sDr3b7p2bph/CJd2
pxj5BqFLxz+WJ7w5dYB1etWCGsY5pPV6lNeYD6L4IR/9RMI+1jFyidFXCH/Jq8If
ao0PDOmXwHLFZVSk4iBrwvWSzPwrY1JaUtm3ogll1r9xsliLRx9IdXo4MIkMnmq4
UcCQTOR1IWxz9LffINyFpHPaYLO4JbU7T9jqgr5bwGQswK62VYD5NNmvdaBI+fhL
c+ixq0vTGpDx9iEyEPkOFGzLfAwKoXdEqemf24PID7MfxYKZg8sK2RMIyrWuXMjA
Zz0BgmBzN3sNSBOx58Hjt1Ok+J6gDmwWelLbzy+6aXD5qhMd2T+hTaOyRvL7jKh2
PB5ZFlyLj8+sJG0zMn/RsBsJ0RUWD0Qsqa/EvbhjGjZOXnNiSIkwy1CaArfgJVlo
Bc/VPyXwaQtOmPGDPv6+KXn2GGQaoEla0FMufs0JJSYGjd2my3Rcz3npsA6qsv4k
EYGvH9GyCHEQUJaRfSFm9Vdd1KrW7hFlfrOTjZ1f9b3RTd9JfLyiOqZDZK3KYuXS
u1zE9yJsCkyK1memFxhbEfy9qmx91wNNzjVy0AlXoLAzdvcI674vh+wq6QO3qzgk
PRtE1zwD7gpMO6ngfvRVVgCsFkaApFnfYsgSYOhFuI+qjL2BAFc4lnjJ/3MsrM+N
z8iEZAtJ2p+fNRs4+XUyvz8UkeNj6R6+YRTUOlmt3Ppen2MVSflG3TWcck1RNvmu
d1vGmm999HKJ5bTQbCPx7MlG2/DtXFi5JoQe1NXdgypRG8T9lQcViWIgYiwacGko
tulFX5SJSLBSmz2l2WrtVdLm7BabtbLSFIsBmTABB3XWiAgs3wKAA+v+LwygIztK
wMXCJdEfMJbH2KpyHSzjvT2PUfBnNeSKMqNnLn0GOgYKbawP5P8MmliA7m/49GH+
/XbTxmFxg4N9cNzcJR+t51nFb/BhQ7kIRdb/qQg384kups9Dehgw3mcNGJEOXneE
BkrdIICKFY+2dAYqIYJcrLXEXFiPUgZoyR7m/d8f/HmF83IpPO8Y0+8GTEDqVgAH
5KXIe7JTRHaesTz8C0DVkKsyPqrATh8s4ZSLqhF8VzJjFDxvu0OMPikCqIcQgNw6
XX5zf481B4UdmOKNunKff+MFiUYyRhECn3Lxpru8cul3LPq1n5UGrqkZb5D387hn
rAateVCiZDyKID7VoXkrGJnZQNA1k2RTNc9s7CnL+LkaXKVptLQlfZ9Q9VkHePm1
bG+G3qkRnj4WyfBidduJmAROBsODgzqrUwmhOEqyQ4gFn34Apz/riuNjOVlvL5Hc
l8lkmdC+LUdWuwO+EULxRjzqRUozBXrzq4FtEtlTNbSnLBbl+j6+17qIEzNmjJRY
YwRHyWCeBIFyd+E+u0E3WssQAKRz7c2aHVuNK2ZH1WRCbHZC5kNB1Ia8v80Xgn9R
riNZujz8LPSsczad3RMVxEIIodNtHlVoMqwBqm9TMHWzaqACgjCe2TyxSUL45PZJ
Dv+dFfB7R4ap8X6wr/CSE2lsJnqbvS5mSZI23Zkpt6UjTjbsfQ7ACH+K7omE44FD
CH6Dr10T9NxmwkTqPK15As5p+wfV7R9RgnfknpqRZ87T5X5BIeCgqcp46BpsUCeM
9mYN0wWT4JAquN3i0hpNfYDRqBG1KHrrZWB2f59yNiBgQYcRQqEKqwOx6vf4W68T
JiYP9PD8lTHhs5GN0jdlaNYA94EWsdjmYwlne6JRLMBQ9NxCzIbP0EcCqYARJgKx
W01v09hIJaVhHnqDuV1AUPYEIXydClD4hwOX8o7S1FZxTALBXqy/av+PiNh1sDFD
Q5gh6XTjjKoK3GZuhtC258W2LYNhyU4NcgFn6KeMStgVc2aXN1r2Xj8HozQ/c9oC
lyqsjr5YxsB9K/PFeMLX66I5xYWY85KyNuW4369sO2qdFmiMEusjv+jTXmHtBqES
NNPH+fsZLyG1gI5C7yD2IaWNu4TVhFWkRcvceKCNkPYnfI9LaoookBjR7LwcwQYp
hnRHweRc+R8Ut/sPBwasN49d5iuA+Fskya9H8liKkCDl8jNOGOlNVd+mDuj6d3X6
dDMzRTqfcqFxQegQRi7gAWsavkE5rACXttPyLIbWFBDcL2JVGfyH/A1MIJ8Wlpo8
KTnknWoFAShD4eG9t/85jtLEKqJ/G8fpXTdwDEN1z7jgSWe+kaEDzeJJ08FbF2Dq
dyztIOsgARO7kbC7v8h8GQL3YR6/2DIRFDLz4kGmhD2/qTJIfJY/rcuKrp7AENoW
J2q13nhUM8VavjW23nSjfe5XNLQf4NK1UPSut1oYm0zT6VMLnr/WaLTbAoTZzf1L
vGEzeDOjQaPfwpLTGPWQeTfauyso0UMt99kwN97vij4KUAis15gV2kALt1FPCKjy
pMEdRqDtL+XAONLJqcjziAK2Dy7ovo10eHF6+LKvvgEjwCEfv6SCkL4ha63s7XRW
tNLy4CP5uVeM5Ayx6+fUvIZMQPc0SI085jmfkOYxONbk1t6MOz8QPT5U1EV3FDUX
Hil2/WXqaelDRwmeN/K5ac/XOPc9LuPO1EZEShFa1+zqcR2DHHv9lZONP/PD+piv
ztcpB9HU3QKlnj54aLUycEJgp7YwiHGOhC1ma33DTAo70KYzX1F0e0sBrcYorsaN
ieTFATlWd4VIaSx2O7ylgcYI2Ho5GnQkvPsPPfZBuNCLamJwcDiNV7pK13VklDwI
n5eFwggqnr5mTroC2ecY8M9OLWpE1u9EMoe3i2T3ZuI+e30Q5MCNBW86bY5iNwn3
fs+43sK5EF93zqOTFrJCh8dG3MURTE/0bY0kFRQScqkjictoTrupZwQ0CAFKB2pn
ATIYrLb1kwSNVDsI9TOM1t55B5QJb+B/VqAfloRCL7WumV9J/pY/Rg9jsKyFzq2l
javGjyV2VsFFNdPeBZfzgk2vppHzHbQ/O9vmGCf3EDm5lq1WMrN7e7Yy74qLvA2D
dOdt+Zb3Ij7LpJz09xTKOT2cJsvaUxTf4EEyNQNkk9A9gD5gUihRfq+UuwQcj3I9
L5N4bp0vxvmwYizZO7nGlg7sWOGx19m25vmbi1133XszBUDdkJ6C8K24TjbHA5Xw
2bwzRqipitsgsY/26KlwXMv103AHMJbEVi/YsY7/MkQjZDZCCRzgK8h+wmmH74vg
lz8i8b5PCLsrTGsfAMoZ1HzaWG21MNNSc98Sz/cUi88haIY02303p0GCQIBogy4i
vOPjoz0soR6hSjI/wNE0+BFFpvx51uhAqsk2MA4z6iBws2ruU+kNiofiZxBWoukJ
iCxOxPR8dREJjr6UxhY90SnwrnCrcw4VbeGjCsrkTzx5FLwbgJ+d/QQiuWMMh93r
PdQpg/Kr5Px7jSjaIz3c+UQLVvcGb4L17XOfRuAPfksje35MpsCkh7x7Q6aopdCJ
2FbYpwWX66bGgzUDN2InTQXWdrCQ4pf++Q2cDeMPMYife64bC0sKVYQAj8CdXu45
jBiAPfMNiMBhLwYYwus53EvMqm9CDwMScYsJcv1Q1PAJGWDL+9vONlM84eRurGZp
NvKZdktUNXg8HBCbuMgXjU3xHWZcvqBKaABRilPeGwOmI01T1cWrYmKqMtMgJh89
z4P0GaxizxOZMBY6sYq98AH/Y/YRDMX/SyCR6+X+H2DqJqoLXkMREYqgtCOjGDqG
pMLns+oDPunqOjlfCQMojwUY+eZxk4HK8TFit5JA83NF+MtrF5BUMQrHBjcF1LCJ
97QveY7IMsux8JWF19ZB48PpDF/py9piPbrbfJl4I5UtSTZaYjmDl0HOBjtg/LLN
49BBxp3CNZAxLgtd8BLN90BITTZLabdVrBaoRnvWNDBK6tiBg3KggAT5P/gL9kRe
MfI9Pt+XZgs1Zkmv8bh8gq70ncfBx+7nOcFuK5TMqUYdDV9si+N2qoM8uEWgMl+Q
XhxzEdY8q5P3kPCpv7sS0/0RyZYwz7agTTL0nDWNYtKbdRp8nf3m5GY6MrhQu0uc
Jp3SWPZBpaFbBmxUcAK8gulUujoZMW1FEqel9gIF48TRePf4gJ5Axhe0g+skrtnv
rEbl/UN02rdcxOj63ymeMotvQiY5DMRvXqrOcuewH+3j6Yj6KNBWURmFXkbeObpp
LJAvsihDuhQBHcLwuFp2CjCI5hTQ+m4xNiqN0ZYCs7HKVzQXCq7SqiqkXG4Z+x+k
OuxAFxfgbih5endP1RFVGdywM6x12Df7mPtgBVHch12HB4BfaxESFVH7GUeuvT8w
y/A/GJ8ceWps+rX9iWEL3zig2uu2hlU5wdsu38SXvwCD9uI8cjxlVuqFwgVIF23Z
aAe7yOZQPs4MTVAJuAgobqurN7h6SkiN+aTzc6ZZNpAT8jyG+3fl+h8LWXFCOlcO
te57HgxkduVD0iuYlTWQwljVj6DgaEiBPIu72InuZfCL/lUhCNNO+GtWAXx5nrh2
p0Eo1ekLbYJcfKryR/U5xYh16c53D7Fu1a2/WMPMRVaqQn7PwX6sDuZdPdJemZDb
zKL8NRDcDosBEVL4gaYu+kRJQ+YY004lxBQfJtPzOmb76RZLmA3Vfj3Qugm7VSg5
13cWDZKlCWo5ud7DYIaIaZH0uvmSx/Gibaq6J7tG2UJhv2+dx4pEnB+o+/UVsIpE
248dzpCc0nrO7m85WfENNf0XoGIdbI6mttja8Y9Sb8vhvxmNaFM+oAGdOniR+PqH
m366kfizd7qZZ0mtVYw8sxq2Pk5zihPAuCQ/xO3FycJxtjDG+Ik2SUO/iAA04CwF
6CaLoQ85JOUcz9lJwI50EG6lM9uw1ZoNMLLDuxBQwS3gebneQddSgwJjYL1B0l8r
1heLawBz1KJ+AKVZ8cFc00JAh0vVg9J2gqIe314fH/CASByvw3Wzw2ae6py57yjb
YMJi7PgdJeQRm8MCR1EyCmYO6ZZmaNT3mW0cZeEvbxKS4wT7/z9Mk7Q/paw4bAYG
ymuhkuHvwRlNTeV6yEOIhjylm3fPi5tKsMHWYH1137R7R624WxJ6LfC+pGlWl8zl
xIEiTkvABSsh6ERAHKTb3Y8G8lv2kFqkXuVkf1NPyFqQEQMajW97h1db5vGQRFaM
3WoVJnNm2y0B3LqRHJqIrr7DE9k/0rt6+M9I2SkTyzyeVIh0lEqOb+8+BSaXnxo4
g3fEKUc3gbetKrBLdmXFyyAciToTjPdrGSM2lkWsxPyqxlYhZ/uvhdeXln8JcrBG
AmV4Jw5J49EaaDz8e2OuhddBQlVsylMNkbmL6J1KiMT4C74aLAQRh8ZORyCTi61n
hhvFyrCYf2k7iF42ipzJC7klH9G5aiKl2hySIfv+lk9eTScl+D0+nRLQVwyTj06u
KD5iNq+IQUBeNUaaOjCsXhf6PTmO35aETdqNoKbQvUYJUcWLulhFHsUGZuaiXUyv
M/HGXJIId2hkgBl3zsI5NrmkUwfjH0v2khKfcByfgyMb1nVCdF3OqBnmywiZB6uR
qI9tS72eCKcF21Zyl5xBCAftpQOANyTXjz+iakL3mgjpyaIa2kQ2e4rQdDKGy3j0
cJnJeDQATb6mEvR0f4w5dycIF2hzfjzyQty6yXRM9jIbrqdTbaFheVEJGmzXm2uS
hvXXJPC3goSDfv6ceZaBNhctExDbflj9iOp/P9UT+tKQnCZCf039UZ1OIMOd2bNz
3nxvk15Fnfm1XpiqRGfnwa1g8XK3dqD4XICiuDXg4bBakgZIQ+PbnblLk1HaFvdD
EGidp3hgGFfzhoLmDEkzvroupJNKTodzLDVzKp4GZbYfmFKBbqtLrEr4dJuzNMAw
R4/RCv8Td/Y7DPPyOjiFQxfkBmVUdOu8IYsPEU4Qxhd9Vnf/4g76oc7AwLAWEopy
bCt0fortBS7fRQ2ZZb7XSHMH/pTk1sUiXLO3KEC52H0cudzeGqubOB88+SS+/v8D
/P+jwhgL5qHreQkr9Dh9PNgWY2Pkq2ON7vBJjxdS3RDv+4kHmPlpxDvx/moDu1AL
1iY2xwnTzNaUpcROQRHJbn4iinFzcQyt5A8gD6gW0fK0AmjLDx9zrDiJndEr3QRd
SnpJi+w/x9BWYY6fPyLqVkdikTHhVUTzY5HyCPr2EdZIVgzdrjOu+W/4Qcz9ttdy
F4qxh0n7vb0KvET3u1c4+NUzif2RILFloVryNtcUrf+EkuV92bYr6nhAtkH3rYIo
RLWmjOoH4cJ1CoGh6qilO99n+oxtNnwOo46svNOF/6HFmESaYh1ZeQ/1NeeUgxc2
yZ1eL9TkpLOGl/ep/dO28qPq63edZtBIu7e4Y/Q1r0Mb+ARHf9zTRdA3osnnVwB/
Dj3YPnDcCExoIBCgqOwtDPPy/WDD7CaKXrcV+KWOpP0bH738mT4fF3LISzCnw7Ds
9o2M7TVe87UhXKasiVGnj/k04na8rfksoi57qMWw/rcdjM2nOavlQqucgT0wueTK
EVBGik6P8FF+A5Qgt2U2tMyh8ZoYBgWwyY9v8Xse/Ma3+txCQO2lE4l5XAjfgIBc
UWegJ094jT9qqZ/qfBFepyt4aOhJr68cirUvNhURpFAkSYK8d2x7WF3OEB/JXkoR
fRIZIZM5NVlLHTTg/BVHqaNJpjRT92uEWwlge99b1PFWsI0BAwlR5bvRjHMt8RC5
2zImkrDzKUQ+wOHpjIvkVf1PPc7N50tGcXXfmkUY5yUTiGjS/7tHT+p648+uz203
Wv2rmCdc/BKF2U44ygt+6UYBKeBJt52Eb0Sc1EnSVoaJ1IoxmZbXZUBGU8HeVw2U
alKdmtkteNvs+KoMTvnRVwUgxFy85YZaxPsavz+j08iXG29iV+sn7U6YHCJy44VA
AnMOerIUZX8m8dqULiFxAFsUgICL9TkiaOfGjynLHapaGZFiCWVnRXejIEdsYJQv
LCDEV4EZmI4eMXxoH/pqgUxfZ3sXR3Lsc7LyuxS3ugP5F1DwHqwZW1HwvsvghhGg
FTpfZ7xlulK9uORNlNmeCff4TYLKHZZGzNSKzF/7AcRsqCYbaLy5hFlib0fKDSqf
ceX0oeQc1WQb1XHiGAgWB3kc0uenYV7J+a4P8vtrNt4AzWt/Qtdu5qT9h9yVKlHr
xauD94mzWVDvgOxAmI6OHabCSYeFKdRU2LgdjTFzzP2hHgwEcIG5k9VnlQaBbOEY
KQgviBn4aztRFAIPS5hyTOLxhhaIw5X5R3TsE8MLSt1JaIG8ut5AEQ+kM7qe6T4J
rw5uBQ/aDw/+lRag9Tok8tzJy2yADTc+Ae3zzaN670Ypdn1leWAf9uTKVKdiySOJ
TH8KRK3GtNm4hT+vKoAXiCviBzgv3qBhTgYWl3Us4a5zwqRCwEVy/o6RYcBX3V72
I3FxYj5d9cKE6/yzIeH4EuXTlV+Mn7mpzGVHMsoroNaT6J6M4pQz0QgfoY15uwtv
3n5awxwTiucF8ICnl4LqjvNGobuhiNhIXCJWzDsrupdJdJLgIy4sC3TpjCDNAy0e
iWtXVTqbaoA4fvhut1HWyvgYblouDKl6Y/2W0vwjWfZkiyivSNG2/u7Rq4LOMRV/
3w6boQAPHP7r/yuOPDqm/SSmbxZIEioTj1M9cv/T38pTAc0sBTrWDuKX0zwTRSku
fVs9Xq75fKQFVu3X/xlPLMnBMRShvk0UxB6zvaCpNinfFBW3IHmNextZ9Far89y0
A2JMGQvZ+b30Fy7nIveOQWBE5J81b/SOC5W9YJk0PmyDzu88E1g3CJVcWILEKZ08
g8WXqddwcW7HWkM5fvT4hXd9G9lcuZb3OPwUAZauQNoMMk0OwLk9EyeNz9+mK764
qErlUOJMbPZWr+oAeElsiYnhV5b965Qgna99T0EvKVQqAXvKPEVUs+kv86lhnEn7
CP1sZVtgpuwPq1aajF0ZoiIK4Gd2ZfBaBkSP/l7z2FPIaoYTB4bTHUPFAFkRLHs3
pZ52BEU6RDOFhgt/tzbttjmToycbfX/t/9DVUrmTAD1W+oNnyykedRQ5aTUFkYzs
kDIpXEcg41P0+wh41QHyPepZH31fCG4W8/p7kKHOz3P2+VWPfs65zt9HITsoQbbP
jlIsHpivbZNpVbO4Kvw6BktgzOCDy+81J8rPAWdthR4hED0Yhl8JNGD3JJ6oWbih
XbtmMsIvbEuw2xUKfMIiKFSrMmdPXKcrqzbTe2ZzwjHc60Vx5b0uVJbjMhsY/GXx
d1pA7ZyUfMk9uCizt0WIc4Ncf6N7X5UhdVUphFIsujd2fVTm0fERU9akeKR8u3IE
TEvWzWaX3fDQBzQ/Yp1q1g9eYk9TaHZ1x6TRknF9FBfVDFgWz5401vy32jSGu37p
MCbPbyA4U3hKL3Px46e60QpLjRFFmGz4nPiiMvjWgbZm3SEv1IjJOMC/OR070evb
4JIf0lvVl4jtkCA3agIYag0UHsoviu+GfcmrGhVn1AXj83P+DIdKTY5Dcz7qKtBN
NRxiR+7EhGP72NGp/tozZyXfXjBjIClzMKtjhcO977533kOXPcc7VKtnmpSoRsmh
rlHTQ06hmjy9Qvg7Y3kLCrYHWKlPtmiRx2rAkDQCWSjWyirm5L93she4ALWg9Xfx
h7+fblA4YVUd/dXRWD7Q8wUSwesSWG15bBUZXfcWme5ZfoYEVDct4qp+34PVn30+
cQVe5EcrYcz9/zwerWPT9A==
`pragma protect end_protected
