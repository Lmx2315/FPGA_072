// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:36:48 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Jv0VL7sRG7pD+suJa/Toj/ocXNCOHeFAndxiilDUCwMGcPr90GqD4I99Pi4TyHsj
/LLGdpnyvx8w918itpb5/YUybH1M2aLHTM1pfSnJXu/ud8L8ayePiprSlR+qkvBn
Wr0nNqDxnnTyvcM+PmSSiRLxDpcfO+94l8g/FLepzoY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8144)
P4z8aEc3UP0xr9NHkUZvKzLGHf49JM1L/3JM4gIuC3YCTf8mDA6DBQoXEmD0cKCo
9sltNQn7JOlXlcFbxOM8q1M79bMYUjsswMKVyWKemqEdpjvwQTMlZUI1qhQqomqI
vo2YxT9FCfbisjpxKKIDWB5ublT5fEMx+If0gl7s3CknfklIafcviUcv/EqAxw8v
WxWzSB/GqoPJIfR4mICWnEz4nTd509wj5gmLqaFWeLgmta59BG7/Nl4MzlRQxDG/
k51WE4ZyCc93hTUTfgW9m6SZS8uYcAkWhmfNkbi5Cpba3H/CDB5Tq+ObCx7hlC8n
I1zehUiWA+u8gAcMm0QCWIujRJbaCS73Aqho+Tj4DnJ4uXV/bGSv5JIMAFNLhC2q
wnhGqBWAneCef4tyj4w501Cw1wEejyrluyAvS6VmId6wb9IOWOYEV7UuUrbJIcGM
TthFq33y/G4op0ERu4OPmGPHXQSgInWOkjdZokDyoKGcJI9oP0nt2I8zH+yorvVd
k8t4O1byMJtD/1cdBurhiQSRXuq6tJb8bxFjDFMGFvV6cgX5ywvuSRrQE4Fgi4OZ
937m4hftGYEHRQ+Lnth5kCFiBiYFoI9llDbDbvvgthhOKCWTiclOX1U6uUuSevCw
jgVOVbjRUvMadkg0uxNGefR4k6WaB/X3kiF5szBB20zYLpyRS6v8yT4RIg39AReE
NFOJOlxIli/uCuNuiblHoC+ctpXYAab1c91SqTXFqNNKILls5HAiF4uRwnBsSh/R
ULIv5G3swJ7AqKCTXwIrAwjjcLAW8RV+/yhxD63CIcztOF2M0NTf9QROsaoddQuO
RVhakmj3huN9xf5V4vfSEyyLdnfQGBXo9sWq6CksvJ1oeAlL7cD9Vg2V0gCzFhRy
oNVJHjzX4IJLXXBZEF7fugZE3ujJ0BcRkCgbbwrF0SdutccfQzCu4Dw2ZEL4Hh7I
1K4F3ACWWUsfkDuxEinZqQrW6jNsS7QzjFzImYsTK7aeb3K0veCTWPUuDFzXHPM2
KC/D3Nrtgx1Tfz9pWHHo9/Zff/Q7/sgpYasS+0vHZ7QBuqCIxKxhksyMlfexkcQC
lgZ5iAMM7FZh13tzSWsZznoPT57qIbGdmk+KZ/u8G1SUN1PbjBDvbmgXHAplhZYZ
eFFPe30fnyZnxxuC2dhvu9z5ounhoH2xkEPDYQ9ukxCrL+PXjXwLoKYRKNJPMPiV
+vUxQ3pBZdCvvNONDR7RNlekgEtmf23nLip7QM+lK1mEFKcapkpauJGdBp7/IVKB
7e+aRv3gopN8LOx3VoGplssZnUGOpT4XiCBnM/FcP3aJSHCRrL8zgJtfKjA3QIXr
biKStfElIx5gr9bND5SK2FISnqmCntz4NWWnUtvjihBCn+K6TxfSE+okxojGQo/D
RJHETKb/QpLEXUn+gUHldPHQSRulO3PnnOSLA8+y1QlTGpmOE1nFo+Z5qmE6Us3T
DM+9Z+7U3uWqaZ3gcgPhqDGEQotjoACH/HKhdoLqWq65BJtYiQhATiEtfzXFJG92
OLN7qUYpIjyhacc2eaC2dasdFLWMM4yaJgO6A9StNlbuxJL7mEwhM94OeN/4eTRz
ovMG3Ff60tW4IC6IoHQkwu+3S3taEpBOHiWL49of9pg7X3eMtcbzhrkGF5PPVSt8
7yOPTnVOwtfAkNbR14aguc7Q451g2pd0SKwKwQ6tmLDkLHzMWcoaMKO5cecSULJL
+s3kh90bfRRL+AtSJIoZzdLjUrDwo0lrflUzssaBqwqSvqYKTeQpf2+4vxwGolHJ
eyXyO0BBAgW8VIi4vwqATl4BEBOixFPW+OI0a8UxgJYaXOT+TSK4+tYfpqSXv8Y9
62+bgQyqTTW5d4n/3oWOTusK5rm9oqty5Yrs8/0iVH0Y8JsW6MWj+QTM1++6v+Az
XfU2tcqVjmL5vb19kXpmVkKjswyPtqLmrpFXdBWk+8uJarZ2m/ppLVsuiDyDiBZe
15XbWXXyw7qzrWiNckchLMQ8VZVT4Gjxco2Ab08++sLRb1QSsqNlJQnEe3bqdOsH
U9PXfH5NEeDAtws4Evw5XuXcoQ7WL/xDfvBBXcDAVBAMVwUMQnCh3U/vihdnTsES
mU++WjROhbg0Gon1v280wE3MdEqj88CtMmly/JhREAtXN5/hlK9TeXPIhymjxtKz
zvtjojWXYLznJdcDDLZ0mn5ZVo94A7WgtCIBmDzPyyi5nkGf3LOHtKkrXEhVIWZ8
he5fxTnYXD+WWiGQ0/YMu1WO/0aLThdUsY1xtnrNCn4iz9pM2acBSMqzNXPuYR5+
/SdKA7BwwEYiZyXVL3rcjMkmsM550kl0Cg6hwb8jUg0MuWOfiYwWUaZwi2o3GG3M
NwYcogYBqamW7Ag2YZDULygmwY/6YlWqeKO9gBmfWqxpmEJbDwABKdT+LvHtI2Wh
+0jaoQmzsfFPFQaWKpo/CaNLH8QDZZ3c2/CbxyJu0v7QruLyEN6W5x4ekK+ifjdR
/jgioy/RElofCgihVkDAexqqL1TZUnJdhsRxVuDNyOIgvqAztEWTVJAex4Z2LjKX
NvO4cfG3x8hxAkGpeMDuW8xzkk9dNpnE54ttUN3YJOBSfNF/UiOWcMfow5oClQfl
72J1fcOoKGuLYhKOFpq2F0hsov2qfPVyLlf/NzN4MJdcSeV/jJT3ijz02ET8zfGk
uO2WmXpZUjqscAFqypM1oxk3jZVG45oU5byr07MmPgQGW5jMqvHQcwdyLhV3PXd0
gv8Uff6n9uf6zaH0r1Kuzuw0g0Pn/cN0LBUBt3sUCtndDFBwG4Vk6MFbTvUT3KRT
Us+oUpA0/EBAIorK99siiAEEM/RcIz7YHOlWvZgWSBxKPN8mYePyS9OhXckM43+2
aG9zA0bEg9/M/K2yANKs8DLilJ9PsJ1LucIIxtj+0YXabi1aGNMzMcLNucakGaDM
lGpgfymx7SJMUZmg6gA9B3gm/CnqcWKxPsdpd6GdFUzJ0pSs+PmOt84CYwzquROY
CSI3fIRb479wbauQClaR9R06jCu18jrpbb+oH6LWCO/NxEjcHulmLaLep+Vx9FnI
f51QHOwT898I5NnOLVBeG9UBBe/EyjguFO7t4aDowE9wI0f8tkV6I3KNoaH3AplN
FWI0DkAUpHlFTqS/XW87Tm02objLud5a0QSD4zzqGi2AGBvNNuIpigRTtvfn5VKX
51RKoV17BNRUb7htMgzQJUYXwEUyj/OGXwwNdCNxY1b0mg09D7h4CZf31/Ra2XYd
TJa3R1OjR+cHIQYMnapfzpPnqogAdV2Gg4qO0I0WNt/+iziwYN8+V+7+NgpiLe2e
HEufXc3c6bAy7XFa/mMbkIwElbQ9G4dDxSEHyYE4Jfv1ZOIQicipgWX7Yxd68+eO
pXt81OgGS2ijsR2dH66/tgrI19hMBZrcYKbTJfUX/O3dYcTvkZNEovoqFzzX2Tci
Hh/Xv8xjWRbQakjNsbBGuZB/Rp7SEqFnka3zE8lji3hClZ+JixBRbNNMtIFI9k4m
BJ2TZUxR4CCBp70KG1BzNBq0sMB9meyO68N/U9OBcD+uNg1HxSp6GucFuC5JBza5
FoPP+S50LjiP0/MBHDJnl6bttj9WsT69oNCAifUMRB2Spq0D9GvY+frV3b4K5lS7
khtPkPF+eoRRy7jBGRN2gzmHewry1frla41jaFmyplyyFVpmOumb4J0Ig8vkD0QR
ualp7ieBBt2ITXaX8el51i57+SRub2zqV2sB16SEOL+I4i/PX/taWWi8X9of2F/l
DMRr9/D4EXSoEaxIWEKjdqFoWZP0xNi0sfpjfRZZ83+5mTLZOmmpU2M4EEkfsm8f
1zXz1o5UkyRXuhHnx6v3U9h26fcJ3I1wo1R0iYEFbJfQoHYq1kKdDCAB9D+nohIF
H396E2MMrjC34poCDPYRC7W75YCCRVD9D9cPSotUSOYavC7hxDvJ0T7h7I0luoD3
k/8mQfxUQfk3ggnqE/YKSkp45I9hKWE1s4v/SNp1j8UXFz8r/if08vDLZDj90GfX
6FKCTA5iAD7/DKY9Qtxcah56ngglUVIqIEHFphlikKw3XJtQ8rF6530hGdsjAV3Z
3GlXHtMUfH7M1PQob5zojqNfy0609/M7lyJw2WDZrsDvhZbD49EhvnVTjl5woFu5
iayFW8SgEa+tq/A6J6vuVwhZhOT3zL0rspxpfN6CfaN1acDCAuCSziIfvAYelDat
bvnhyMsRXEqcc6uAulOVYnfr/46t1/bMzyY3yy6h8aw4ckFJdio7BNeu+pEDr75P
SXoHCl23H5HdVXvnfKdFy1sa1I4VbIFIX5hNqP58Yd5JWvtCxb//dBR8DA8aqS6W
haf+YOTxbsrm4UirryHIxJNPRmn+Pz6UA4tBwaywKpKDu7eL+HPLaqJTDuPc7KSL
3Eo/EuUVVFTf8Cs+XbZjWJOyvhYsQZ5Y86ZEj5qQ8NoDXKl2/tFxns9LPHkWqFBZ
5+zo6i6pAxXLdASNzxHNyS5+sOCrJ11H/S5y0SMzTfJYjSHua6wcYcnBSKNIW5kj
HNx0pRj9FD0+b7Gb2kTcppPjGx4kTsh8nyv/OXg+aeaaYzBICSC0To9M9QhvxpgK
g6PMS6ser4fGE6eMh7zWWPKA+sHTG5NdhZJFDhWzCSqz2TgI7bkl3iF2CA6mgQVH
yfxRmRQejdkNsBzIeLVznqzqsbokSEsqtvfFUrOvZSetzrpyr565fkrVe1fgaQeu
r919D/lscZWLpGoO+znlvPIz+Wr8Nnz8Xozmu3368BqOmTDIdlwqMJUw5n5eu5qh
0LvSXHnK5MR0dyUT9z5MqAmjysMCiYL+cFzlxzHSvfkAbwoxb4KkM/wKhPEA3OHl
wzQU3tz61btwXnfJ5iT5/BvRqVSgZX2pe1HjwM8LaArB+csKe9y4WjPYiW7FyTUW
V4xYC/Fkm5VnqQRSN1MlQu8hwubvWhE0Ipeh/sX5zQMg0dy2RxSmzM1yq8xPKZM5
OWw3b8pqar28p/UtU7PL1JWcfnNOyTkoVl+dj3u2qU8LfcKQtrPr4ECLvseb454G
LpnacoVaaH6kDJLLLW6UZksJHbAcKWXr4omUU7LAFpcWRZ7Rz5WuvnAzVni2T5zO
7vE3ifFc7RGZC4Pt69YRaUZ+XLXLe/SgqnWv7ckIoMQBguenMTF6rvwon8e3bk/p
1fraDN74f7cdpvTbT1js1HWCy1tn8kb+uSIpUvVV5+cZ1YJj9F77+22Tt8EIoTNT
9Lq/drWfgSs+nH3ppmee1QlcotI6sGzNWxE0rAVJkKTXiokjo1ao550Jhmxi7ouB
1TP1upNoq31+I2aB/zrVljWrJNmG1IFYp9XOBWJSs3Vn7l6I39q14ymj/uX6ynq4
IOP+YCEKL8ZWXeOjzQx0iRiJGucFMWPCx4NOvtcWu28JMWvn/i5njo9wUrjoQ0xR
+QDVCcwOTQ3wh3KdzvSCs6osuV5dH1tgurlg++muAHjfIbaa5VUx56mraEpNcflE
3R7it3rCW+S3P4OuAQ0IQjXry7mUQlmzUaANBrEnq7ltelYq4xBEZDaw/JsuCBPX
b7EJJLkqH5I0WiqkWqMvuDZzixlKwHhJyXvK6nJaBbb9GdSs7Yaxf7QoTyqGQWdC
uekZ6bLnn/om+4MYuWR0HoydXKe8Vm9IeqI1NK/nlF3V1zyZ7IpheW7JVtIW3/Un
/C/t+QmU/rgmsBH2oakOzivOi3t7mfyIrnP6kxyf0jmS7k6xCMX+EZSoA9xNgoZl
+dO55xVrC7LWnq5n0hqmo8OXXv1XRW6DTshYPg8/AFtktJ22Zj6RrkKSzyNZoD3A
2d50tNU3CY8HK0i8K6rneA3N9hYaTnH4ukaBWtepwXnn1LA3PJF95BmlMmMJ7D8o
0UmNlfv1KOkhUEhk0qzCayMmlTD0fBADyepP3TOcLX3f8bTtsOhpefncLV5zBktQ
mPR41ttYhD/UA2DDe731xgMeZLah6gY2sYUxj7NPx6RKhpGsOP3GkRS5I4DcR6Vf
OC618zNrcrIDQYQhXC0Q51eS2LKvp7F3or3quJhGUqVFA+Nhpbd56WBiieU8Uo1I
wWhVcRMhDukrpO5GwhUk1Zg5HGiJzdsPfXhL/jcSgDFi9I1s2uWhpRp8oAra4T58
TYQkpRCVral5EL47NOv4J8yJa5JQOEkFwB+LKUvnyI4hwkbIztwL8e+lR1+eLIhH
YLc6ks5krg88sP8FA04T8EJF6VLgqlSwJ5KHK6rcCTvXkL70h2TWKV69rLEREaBL
WyOBllTx7IMdooCPUtGTGDxd5qkTjJ+GJO58R8dAWXHxm5Tl6iy4PneA7HDoWBnM
Ft5yjQTTW9sfevDjkau1LbIkUetyhAkao2nWoPEdXPnbYukng3LFf9og9Dhorfha
3MyvuEK87p0xWRY9fOFarZWr+E2hBt5++orY19XOj1m6goE5FeDRNlCx6kSsDtLT
stjKKKh5aahSoXIR745nVI3WHNdRO218fNbLXkqXBaKijOtYM3TCqlipB2v2tXr3
tG5DVykIT0YoqpSgO2Zjn6EX/Jejw2qUo2VpM4M65iRZEm31Zq0XV3kygKVm3qn2
zOeqsaCb/vXHeIDsplMzGqF1LDJWz3PjfaV83GpnhbJDE8Fk2syDxo8BtGAlnvzl
Ewa79UZv/h+iDZ8peP2UWsqpQiYbd+/zBw7FNZnE9UBKkS13Yv5mX5YUjQAwbjNT
WuvkWjR/FSWkPignQBxqWAc/ugFk8l7TvEDrI24HAVgJC5d9xf9TcnIE4kDp/yz4
AKH6E4u2bWOofm2aAm9crix9WnCHA3NY1QIvwzCveuIzpBDFz3j4WVFs3zqtG/Zt
Np1BH4x316PmEgizDJeWH51J26v3hmff/QELs1faAJmXG64Z8pFxkncrJUV7yWBQ
JtLp8GaENLcOYrDE6MOYlt664CsADp7bArNNL89nRfy5vnu/ABMFoQ1SQf5dI3I1
6A6mStcqC5IS/CaPgrOe9rLg546NukGowCaKd8mTgVN7XgLmIKBDgfNjSuwnUZ8W
nQIwjSxugpFsTMUtG/uHJ6JUr47z5V/LECpNoBzI5Kg//NsAeZaYbcYDFn5UT2pN
q018rIWV4252BX5XOw+fwwVE1iacF0yHBz8/rDO0NUxMscVF0nuNHrVJSuaEvC8B
psly+9YUXSxfAwFrskiixU2VPAGH6Yr12wvteLx6DzwzazK9EVsKTdmlGHg/jhaO
CvWQ0GzXxHpORX4KTkdLCaG+2iCStDlnpTfqYQ3ukFn1bC061hvzrwuJvX4mLzRa
Hz4/Jda1vFIHoYj8YJyPsLcYEzRJApAw/LLDNYZjIr8+/zV0OlZrHlyPoF/khVSS
Q4xE7ewoEbvJGQjBb6buIuI+bRPvq7SujtmLne9Uv9wWIVfiP4Hk0H8ijuiQDgsm
dXAdKvTAg3WJ/BVlC6VWyAMdh75BtqXjdR/qj+fDkmbgKB+1lh8uJaW36MOVSpAR
5RamwO1NSLWPLhygzMtIfTqyO3BVbAkY1p9A9hesrUBHuTiz0/Z19AzTdCAmqC7K
9OY1tLp7qmJp64/QIYMtBsLgRCOj/DF+7Ap+Ti5Mqdp8MkbaJDQo/NEtCI0hgo/q
HyqsLObSIDTJe/xcnwLNNt3BF2MbKgFDJfSCBliHT7iTqkOyg+5XQRHFMGJ/Hcy7
eBPkv4Di1bV+I7el7Ce+vLIYsCSE7WdFKojiwsDbd+H3ubtaO2u70yRu1xaz1VNW
fZcWCp0jj8nqVRn/T1tkARBVJbylWpF21Zrzzo3xcLUQEg2/D4h5mEJmbbt66VaB
Xbi85gaYfs59FCGNsoceskJ2MaZY5tKmPt4aJMOLBEo7V5qzWE4rJ/JsqB3hrdPJ
nrjvrXvthd9hf4/BwQ1Dt+smgxX7VakUyzTyPvQWZFhdGCogXztO5wNYc2KG7uXr
jbZtmulCWaoOo+xnkdM+iZcH6SmV6O53OnkF0zuIoB0yJ61ke1G0qnvQCVd0tOvk
b2WgApjkiIk/W+wIlNkJRZrrBZ13r2zw7nSl8px0a7rqSdQrHyl3fPDGDGz+icBI
VQKXHIhBjPtXdQXblRbqBa66BqjrAmaI2U0EmBIvz3pp6bdSXrk+f4MMC8w/81Ib
44Px+R/ckwzVrIOw8o8QeZWdZJbRAzHvtQybMgAEfNdFf3nQY1YR3ZNBEO3w3nvK
8yLGqmJPy9xRUoMuznQK1gTx/ISZxzUzCPXd314kvosGyYg9GxdoNr1rVz1SoSJm
qkFcqIyvQqSc4eOLQccGOMNW71eng0FRoE25RntdcJbC7RfvQNoh/+p0bEVcqibU
pV6bSIyTwrhbG+UQSFpBuj4i21VhhKSdB66fYPYiZheBJEBASRV8QZiHC30iA9go
XcXMWvxlxZPHH0l6FdxVum8Rfv0LnAJ66ykoaPVY5gWnvqxqu0KZ2sr11PbPJnM5
gYWtGhYNNgdXZQof7hb1Qf6+yG2y+a9jUlHFNdwsJNg7Ik55mBVw0A5FnkqiJF7R
+blT7d5BrUf79xMPI7wHeMQ3fhHjS02FQnZz3nEoWJUTrbuqjw2uWBaufbA+n6TN
yL3pM5qJqNorvfEhcLZA0ZY0dB8xRLkwx3IUcbEgZoj3wnexCF6F77BgWVZqp83h
sNJNJei4IIl6oiuEtYRIAr8ntnbQqlMtGyYLHipg3Z0U61D2OdqVhXBNO9yQ1S6a
c2Tb7gGv+prnJ3ZyNd0h6JPhWUHVqSvC+Mq3kQcXmxCzKUYZSUm0sW9gMpjZO8pS
mhKPIxd/DcajsXrPsDYnphEW5Mf6dmYbvlavuWGBXMgUAVPsrw/+dI+1vojsVqtz
vCI0ARqHJOpoXJr1CSG1R2S2ez31Ll0rdrIEjy3UEABREF8zP/3W50vGS1GLOItB
YDXBqYUTGrk5uq6kwXxZ41izna5m0wAWG5wa+dkCm2UQRIBgnczNYYQK0IKYs1/U
PbQI+0+F7k1DNvWeWAKRACdhqrQ/C88fNmH7pz8sK8sLrA6mUNaX7RJ/HjfGR+X1
BU55tbpVIpwSIJYdBbH64vjkrzbGNecvLajL9QgY02Zc4QWrtnbT8XL9Nh3/KQF0
1ngBwpvJnMbCFYh/DzqIImLxJhGJ9+GWsNIJg2/aUSOU8/CehJPY84XnraP1aRQS
RTiWuKnDILU4chhXPh+78IX7H2JIGdnVZgRQtquYdbV4j/VgBjvrTimuHobrPZOv
fWnfHZeSjVsxSpHsosyTLH015arx+4PGT4vjCTmFepIu7wcUkHcYszj9HrBPWyJ8
NfPkN/jVm4mCTLPGmWdbWJVEBnwT1+ymVjQ8ezUShMt0l3psprWyR1laLU7FwRDw
AjGMKPXHtqTUcPKD97b37RyLXiInBmCAPlX+H0nOU+mVRI+AFL3QtmJ1lhMadiw5
Agp+A7ocTcokYdrYK1607LJvRudCMWbuzQPA2ZZjDO3pY24807PD8Y2Ss/Pycnm2
u8fbV+VDuqAjQeVKdtoU1YDoCRZGRwy6n8yhMOK3h84X7F9LbBDt650W7mmXQhTR
mtwnK31ce4x6uNGhNnzUh2K1nzTXoRf3RRpLKrXC9Y2Y4R+2ZmCI+5d4LzCBELW/
170FtbdnKfqNEgI/UwyvNNZ7Kasw4U1JmZ9BBZmDfuDfsaUh3X+PRDYhhKO1Fvj0
F7E0+IlFh1eOjrpzzzst1+WcQ4LxS9PnEoCm9nqMEXkCVyKoSGnUi4itE8/xgLAo
UiMFvxISGRJ719cfCPxsMaRPri/Z/P0fU8Pl6EorRSNjkC4ZyHvldAxnTod0xReM
+ym/QS0KSVjAWA8MG5BwD79ceAwW8cNxu8mKWxYx4P80hutSJOLuz6s2uoYFx3rg
IErQQbtIs5fEieJvumv3ni/nY71Q+sB0ft2b/UEehVJ7Sz8pd/Cdu+xtewQ/lbr9
o6fZf6VCbnTlZstgKAY3osiPFFsAtHB1zE1LFUydgvf6c8tp2QvV1rdN/8HHScid
1dDeM3a/VXUZXxsRep/zZ5xcPdbRNvX6c/tHoM3027W/wxIt0psb5+6IMsV3+K7K
MgoA2kfQuJqq9Iw6RoO+M7szezoG31SFYfhr98NCo1BGfpN99x2SHUhNiHOJRfNP
Aiu9TymY5PqvzBcG6/3lcEmKl80fp1+poVDFKgcMC3vAt2iJJRvko/jx0ytfKDcY
We18YrMovl33cWN9x4kwiXTL9koPKuwMrdFn4ZRtBKy8EOy3hFWLCf12cZ+9lCjv
jaBGV1KD1Iigno9FLRd2RmpHUgcuAV4lvtp7HuCWcStznit89B6nNluscc/7owwI
/dqFNZhL/6GJuUjMYEdkwD2Ll3wuE4XatbldsMYDJGKdJB+i7ZiQqjds1bsyzOa7
FitYqblHM7gZkbselfcOdH242H/9jpGre6N/0waQoznt+eOiRl+z1+84OEX0mTjx
b0zls+2cHc6v0TZyUFmR6qZe9dFzDvvrsOTijtqTWzp6qJE+we/jZAK9ZLf0WpEw
Rja1ym8NQKYV1ao0YnF1msf2T0fySnJiXRH6urawY5BFihJr0cG3amLsOD5QMJRk
rlbEVY8VtIrTUqZPaWMTrhU9kl29nsiaxy7s8V7EisTv5b2//Vz4dn1gkoM3M/PO
BvM6ABTEvsnCgwi96UKKYB+Il3iemzb2aLGQLHGxDdk6OFn4wZz+ikNUisPOuggt
8uTOeBnwH9FRGgBQXwRyWcstg0z7ZTu+IzHyopTW4gnD6uxAHgQQ16pOBKH5csCS
2xPJtd9k7E76HfRKxFQMFnHtF0zULFfTy3zmhXjZXmx7vUUJwTWXcxUwC9WK2sSP
7Anl5Uf/eFoWJaY3ozrOIsJS3Gx6cS/LMBzWARfMZ8M=
`pragma protect end_protected
