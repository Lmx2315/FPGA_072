-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
MQ8hv3XIc+Ywu9RSL9Bj6qNhVpw+WIKlZn/r1jsVe2P9b8L/EGvz/Ehf6rZiOgCFuWXDAiqYjOlU
4MNlvy0Jad5HjOytZsRe0lw2DqXj+ygTLU4eH8kh11LrrHaMQEEJ0B83Qik058Y4S3dKZL5ArSSw
tabn/oQSayuTfPs/xHYb/NkrEB+BWF2w0qYIUZGwwl0BmY196/mOwx77gTOeKkkAvSIeYGns8Y6c
9dMLF9F1ZzZAxCw83VpM86kDIKzAe2W0pyk1A9uYmT7qg6q3IaL7kvqi2n2p5gYE8dGO7nafgThq
t7FY1jQ7JxBS5ff6AS59neYBwp7ugylznMrpqw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 6672)
`protect data_block
4F5V5ExA3e67i3BBpY9kN+XlGqDIpZzPenkXmdazQ7/CGVadLog7Of4aXofbGwbNjctAz8aqf4We
PyuuVgdcvL/0B9czp1XMBQ72CY8JVBgVEP95pElN1f+MZYPBeGzR/nByjH9vFoXzETYWdDjCoejC
4CckqQjZvf4/oj9zh0vHRQ3zWfW2ZiMssiYGWXXLivV1UTZfGxeewdlLuxG55x1HJzNUyNbPRMMU
Nvj+JkAJ4iVk11LqkTqkc/0Ep7vZ1Oaa/wnBhU3fcburOIbFyksh7qBEdXm9wtuy1PUfoFWY2b7o
pGN2ArhQa5RAJMkNxfZEE+hvNq/jAjLuaJqoTXR/Yx6+yMoofiQ3nrGjEBl5XPrCJ5pi0x0aGwwh
3XS5JPdLpqXB9QMyM+mDmMrWxVMVVr2JauNd5fOkRAsUoA/Ddc+WjWzvsl499K1aBCbHJsxQctwG
mPcFLlskHdeSdIhwYmcm86i4ECHyXJZqzRnheBIsPDF4bZERH7wFDxo8pb6MQINvprLQgjH3t1Vf
04D4LJVczS0m2cQCJztYFisiEkcauCPMPQFwEQxmLOuseU1cKNVnxwzciMJyrgFaPfCnmwOY0JZO
7vEBo5xCkkSTD3LARMQ23UnLrv4bAtFz2eA0R7iZSDFFt61qbR83zUC3YH1OQzHBOYvo7rOOvgPW
FjLZsHFmXA86DqLmaVos3PsZrPXJrbYjyqw5wJnE9EGodo2tNxQQ18bAqKyGPxt0WSSF3KqTEpMO
h+ab7ySazL3xQJM7UWOdcLpRld73S0hozcDzvFOz+adR4+OxSHPtriUW4nhbbpK3olJ9VhLTD8Gz
QEEC4/U2tMMHRQ3tKqRTINkf7xaag61H8z5Tlxw3Q1XPL6yrzojJjNyagGbyxk3OpVAl1cP6HiVq
++cdqESSiE+nNU118r1XU6GHRmkpLesAEqVAP7Ewu5oCB8DHju3zxeWKFJmKMsevXh1/KDXTs/77
J6mQiupfCMIfUHSVf/1604U0pHYYi/zFf5ygLTA62MtTK4Z6RHoUe3GNrDAajpp07R6uYxUiFmhl
zaYPGvieEf7d8GLAhrzq/dbj8ImB3P3u11wrDE2rEshkClb7v3udYt9DoFVP+D7byY6J0Y6ICqv4
fUiNWBjGQrUioXDTrJ2Ew0tY+uzit/dlfxXGcwNUMVhxn6JAqXq7VJW/tulRF2DeIF4jdBcDtxVC
nf2aGI01ehFP/tOr+USkNyXOvH9e6+QetDHOiTuFD++6ADNSbGmttd2O6nlU6RCHxE4azG32Lgin
RYgApWOVrmbNWD+jDlEyAeGLfBH+zy5G224SFWsEYot7HuVSwEFMZcU/7QDe7UYTiSagnvDCcOJx
M3HH7bZrqGbe3RfJxRAwrwomI7FplQRdQ6q8sQalaTCguKuG0o9nbfFxk59UvhazAvHy05otoEoD
9L34lc9eoTuFO4+p5dTec5f1+hvH/QU4S8XURiV2YwWAN5UYogbI67YyWidweLUYxf27vwoSAdfh
R57doRxLDf+Qfguvr5fJgk3WAQ+yMdkMrsrliqvxuZYp1MAp74nTPymWozIIB03ZK0hbEIw+MC0i
8uro+gvUg9verGeLTikRjGwsdJbQBvyT3kV59mXWjhzKyDOi3mx3oVb0OMolYcKWQaKI/RJ/H/ij
1FDGS2hkxmdm4dMEJeIClMuUcyylxaf9RBJkxXB9Q5cVlJcqdLrvkdiiYNWjPg+D+27nw4nnnvqk
1buInwEiH20NFPqdidPIIr8cNi1lUExTV83oqqzYhEXE+vR0Futn+z28hulfRIOcxqIheCh0jTpm
DGJiWXRstW/uGyZYewkO1DIGwXsp9qkvfUeOjCgm1NX5Oi8w7S34kNDvkKo4JEDjjBD9Bjg50goS
0HpSxLxfk3Q0i6bynKLt2dDM5QhboKxmNUThfPS6dQ3yed2ihEHcBVKPd4DZz0qIjNehPPg3bqyB
uy/2qFIr+0cWEPHMK+OTxrlV4yT3p6zUPjB2icMsbmAn0Is+namE5zSMU6eufWGbWZaiG4QUejN9
AdudT8oz2l3X6NGuqSDwwmfx6iirRqPlQqKgmYCIcCZ7d6KIKL0/B3ahnpG56rVUu7LAJDKPp22l
LvFyfpG+ud/FYvKnrVEd3oXey6aaT1K7GU4mOMpH2xXbL9YHpow25E9ANHWbGy6jsmU8mNpeC9G5
7Z9PZcXubtbzZXbuFN37TtfwGzNLRkXyuGgwkGxWaphkDPq+FaBbOIrXtHf7fNLLA+pB7J2GTjEa
dvoXzToKy3fi4z2S8Ud2+UdNIpE2+AJEjWi2eWgWvHgUfMAk0O0ur0LAkjpzIPqKP8q3xdo0Lrk5
2pvZOqtyAGTyVgXn9CO9Uff6QaVgWq8OnCpYddLVyyH58OTXAre+qTNMC5aOXGiAxbmBE6WkXbBS
a9B6rJ5+B01VX6FAy3cxfK+PQr8FTBoyG9OV58eEU9RiucS2SRClqlE4T77IRnYOxrxgTH2meyJb
Z9WX/uhpXGy/dEGlSRV3ck+XafmS1I/WZr1lLsveMdx9Cl94+idlzAfwNvn2IzxMecjJICXv9VsJ
ge9JkkvwmdvRfuIDoM0TMuLnfPLOLCbtkaUdGbNOpc6KAK9EueXPoV34bLQi1jpi+rTkfFCUWu/Q
HAGZbJ4YYMCOnmounuXqHm+lWwfKTqKZ4b2FBeiMeFmBERpuJrq+nKQQOqFVA3ELQhVuS3m0rWZ0
5jBtGIui+ZrB86USbohKgRMBFXiFZxOdEf55uMtcqxb3JSFr8Gvap7L4v4IZnm/4/ANHjzlMPNp8
Xs9ya2EJNuvkvt0IZb7MbY9phDFpetwvDHlu/Wt8IGGStK9pdIt9F8xezZkc5Tn+Z4MjBiDf1kjy
4aZihXCgPwU2NtMivxwP0LxXV1XDBSA0dfAtdy6Qo4Ij+i8c5wqJSiyG6J/juoOFFN2qS7K23/jF
TIoAeNlCs7vceAVfC/U3E7E02gejcofS0Ld9Pr1ugne4mctGQz55Evm8zAZSLRq5Mfiz2JKWoM9P
VmQ1QMFNIhDWzPF8pDadNmflOLDuNwUx/h1qB1MnInfgWJv+OjhcNVVhsDlehUDBkM5qj8QUcade
6FOzeF3g0mgt/rNvwj0TdaIFwzmXOGzRXW7eouZT8nn0a2OrLge4tiHLtUyX1YMJPNpUMYHN46vy
62gpMMJ6obMG6pCmMGBOUSLjmI3WjDKmbxJyr2w+P8+jYizt1II5EV+QBFaRtEJ8nRb0OptNPz94
rzTfvQ+CKBXqWxw3+6mSIMEOSngooD9g3o820qiISOuqmJJ3lwG3IMQsN3yUfMWlqb4BAfyz65Ih
Rxy3kp2P+9F11/JBcLT0t9BywL5jJExiTeV9LDyDhpdWWosAdjfV7YaZ5VBIyS26QM606xl/gg3L
xRAFCy//9m3vz9lwkD8gVMkMPZHHZ7WdDjTWJr1iF0Y8PKfL9l3JlOxdoSbpn5OoOZ1ERd3C+Ksu
exHwXLsmAZ/P5GJu39US2OmPclefTZwBywX1a8Chztgh2bGYHdEbL4sEx2cgv92l0MVpnIe3OuMS
Z6/k+vhUebfotyJrxvbWXJOGKfjYdL/9xsZXi8iFhS0IMsYrtZtDXKTbJp1RU2TgfysY6ldj3hi4
uLok0Bdf4B59FOj+pq3JMbqsWPyg7lXM0kvg2vjFp6yF8CN7Mz8p5W5RC83AnslvMte5jWyUIwKs
yufp738cofXGkAKsHVwG9Val8MOg1nnk+4tWG/l1Cm012C+R8gaWk6Sg9oWF10vGimNXbH3VBrRi
lOrzsBhqcLQoRXgD4RF1BeACz2vPNo08xMrbadEanELyv9PrJij/QOT/ptzf3B7n2IupLUWdgthH
JOteoSPYlhiwbGzFjp6JBTe8Iw0ShZ5o1WJFqvXH8i3uFNlQXnVGkANgT41+eprzvOMW10Avr/hs
duEJ/jvQT5cCS1ku89Ky6WvKPaUcMsx9c8GlmHjrfuxX6N+gPMTgD++k3HKL5xf6p8DWkSW6J+vy
kn3e7Xo44dQ/5Db1Sw3V4t5gXx1VLYnU7aSx9gEYT/lipdkDqETzqW5QMjGWxcNGpfqWpEMcm2jS
ekkDkxfPUmeN86t2RRnmAMDqTGiKBL82zq5uZevl2NandWaK+1gjN6RUBT69ea+qTNeoHViSExd2
7lQySiPPTrJzGbdyw0eJ9x7yPW3m8MuhwbZxGtM0naz9bO2/BGRvXW1Br7zoTwKamskieaKixXKL
1IQi3/XSJGcjGGNwPycwdgvCQ+f2V9mIkM5XCwK4zp5PrZOoUFejLVMWyZVwzjvpixmfie4XNq6m
j/xH+yQrj7Q9PDlr0hl1ciq8JBTRa2cYVtR1kkWmDLvmlto3vKuNA6rEVmX8j31OeXWVnvygk1PD
wX0VdtNCu8EQ3hmlRBb7mtAk2UOGyEY87NHAuol2o1FDbHt0iFFcFnM0Y5Y97XrTH2FY2RC4/635
k+XFQAJfnjwEoRS2lohC/rWtNAXDofYWNlTEqUhV8VexRnVDLUZC9UXq7j98ZF/e6H83MsOBgXo6
bOYtiFoX8qfQ4sw4T6+0hNbdfWbM1S4o1IPxnN50GRWzcmqrcDAF/hySMzZT4bcu/WTzK9M3zm10
FRZRUgv6db19TA+uZDhDCWiA3KzJj+dRgUZZ7NOWkZ8e4Vhf53LEkB0tzIxri2/2GJmO8PD/wm68
FbRzy/BhBmA0WRNxUAcy06TEr2mRQnTn287E1SkFbuwuF+e24pdNDMSOT9k9tc5qfTzbdAn3xl/1
DkpJMdj0aCz+TfYI2fJK9Jf+OufOomPeCgdrpH4xJ4PBfNJv/IQh0WSk/jUJnbs5SkTlU8iSXUPO
CyCuf94I+Eky/vjxsZZlAftPXtBMRcOS+fU1BL6Y5n9B6aEBmWGefaPrOXkHoRm6ee738vWNPs3v
wVo00QXk+wC8a6ed0ycwTbNEJ5c5ynorsyNc3euDWfqcw4bm3tT8rkqmF2N7P61Hj7jIiFOY60wP
UvesL/cjqtOepBanGwVlYArueEFVL0vIOfItOwyPI8r2A+FPK/EHyVLozCW+Wgux2wuI2z/KS0h3
xhlHeprArlC8+mfbQB8XiiGg0rpcvLywW2rPZL/a5hd1KER9zkTKOET1eZQypyXUsH2t3pEoYiyT
KwYnwqL5GJM+bBlDG62Hl3YnfcMLdkul8DpJflK6osUXzl2JG0iHC/BxzpHxgFmaz+cNSR3FBMPN
ByHee6B1U0dCO7He4q8Z+udCsclSk/pISgUekNCTeJaGYJzBQkG9ID1/g9ncuq0EfHVDqEfpi9+P
KbmYQJLG08Toglz9rARgxTo3PuP5z1lOoF3ANzWWc+CtZXQYeG38w82+3Ae33hBq+vvXP2P5M03D
grIbERutyBPwHy/Ibk3GICaGFMaMv3fX/2PmHJLqVub+m2KBH/pVS3H1W2pJ/C8IcYQdvawOyaYR
0KeonMvVawyio+u00PCPuWGEBhKEbl/1wOQqSzGZUqD3RzJXcIZrxLAJWbSYEIsrtrnlJgubbOty
ExFlxI9F7DH2ngtLijM04Ab5QlpXeS9knViprpBul2BgoMwVdij+kDbpgssJ9ZzWBMFOZo6hbxPG
U1dQwbGih16VY/LirQXdZdBCDhObFFm14x04F6NwrXdyu+/U5U98WQADPqRoXcRJwTYqR/Z7TXpE
c99WGAfqJbo5z5ZvVnkReQfEOpfoMvi8/l5ZoEORS5if2Tb0crB9gg5cZBaPTsVGva5D82KcnSgB
CJxs41poA11PIjPzbt+WOw2bgx0AU74sqa2Fy9C5Y0A8fZlMSoD0cw2Ovj/Vc2oqKOnFzX63A00E
pTE4Gx/KObEJOvY8L+7P8XY3miBPpY8bCo0vpfXnfSjdxWqvLIEF6ZHFTCz64RgPie7edCn+fXn+
k9oDIlJIhe2nX5sfSm0E8qYo9LeFk8mnY3sUKy5bVCgRoL1KzDok2ZOHs2hgOaoG/Cee1SxsNq9T
UBUuFv8tPhNohesN2KP/KqxvSjBnrg0dM5klKf/wqXzn1Po5EaBTlYqKMmRv95lDV2MvNV1IgGQN
E+Spj+hcqwlysQdiGqwIYmvnY78/fyLqG7Lxldmg9hgwyk/Y1H3Z0hYRGmpqoj7ktDBfiNe07Wiy
L8y0uRSJCdhtz+an+6IZ63SEjMwqKAapizaTZR6gbwG9SdCTJ78hB6ySsztvJQTQqJbGhwyMQx8k
Qk7yLfZz84JQC9to7azaZonYKFGy5OWcQKou6iFnS+ftlBujuIXdw9/bhDFdiIQ4ma3gNVjPsT/C
YiLZt3/uKZvUxvVtQ7qa1rYPtAAigoT0S6I1O510dk3iy38yosx8ZxIp0wRaNnuC3A1f3jH2NV8P
FowxeZyc3FjSQlgfc6ZqFNB18tFiFihLA/xdtFaUhS9nf/AhfjJqjoqIhuUsLBO1YjNIoqGrWfKy
onl4h+94NDQNBkUJ2tGji8dFGO7OqGsQ7wICfOQWfA7J0MaVh0uj+Hg7m/E8FIpcDWwsVFB7dmTC
Qrfj5hwNARYVkAoEizxIONgyKVF9qrnIUTEau6wvmOhaUB/uPrF8TCQ1FuGChRPQqP7J2aMjKvt8
CvvXbMlkjeolXNa/5g1IvOzrPJ0/nmbWzPUxMlOpK8QzzSPYeDxXZBeEgIh0RbcOjeh4F1q6HM27
I8filhD7VTA/PSzJuQRbT7rObvpap4BVtUA6KyxzyEDa5BP2N1mErybRbhQlHGhd+b+bURJ+Ks5V
uyKVIW2BhgKUW5ZWaBz69M8Vn+6RmdoGx/PLjmZlZrwuUEZNMrLUcUBgtlSgDi5MPUukL9vc1HpE
/seFvMhOYBJQEOYLwDrak3+uNMJ/0KM7p6SkeqkRgdl6o8jOIaWC61sUBEpqHbRbJz4ouYEiNTBO
sZZ0hjQguRHH0yP47Tv76KY8prFg4gEubqCA+AiWUAOsWoykBZcPv85NWcEws0O81Jk5mBat0Go1
8+DKmsGi5CewxlxyiDEvuh9BVagszlpL3Ph73Px6BA/VTRSi8bQG/FpRo4GcCwEzF5k7xEx62C8d
cBg5FyPDqDw/iF5QSdLjcXeTbxRWbV5g4MJuw4NA9hi7W6wNZuigwVRqwDUHx8nMm/3+3q9Bb3Lz
1Haon9TUqeXheqyhzjL5cRDned53jKkxVj+z+FAiN07vaBiHl8Z++BEp6GAjBL8O6woCnkf73nCh
uw0yTgxWMyYDlnSiWpl5VlAIsCXDLv8e6BZOVmUQluIxsN7kYU/GeMvPVipp8NCXciIXwOLeVzE3
Lg0d5lkhfaGGdcNWythxde6wozEf8RJDvIIcZrWih9A8nyDFlsQXIUTNyBOe9kukuGRnhiGXAyF1
gMcQa24y5imH1/IfHHl+/n8/EeibsvJG2j87MLyVCfnCp9A7/Ek+VaEPSDIduu/6guYDQvMGtLYa
kFeZDmOghJ4U96PqNpIztEzNxO4lVHIJRUn3YsaWuigZCYxKQUO/VEIc2z8sbTSsRSlxH+vfPiP0
y5IgADdeRriJs6I+Qwv3Da/awUv4aOYW/Wz+1/6deqabVlkmguL8i1AK4uedftDnKBO5uOEW5z7A
Dp0HPw71nwQmqRlNUaTOsihvcXhCm/tES/oMLuOnFyz1UYl5YJUCTyiBuYEaoewgSxQntGg9nxTD
8WeWPRSN7raCf1Q/rxYG6DrszDxTcBiOytvmI1aGpfgDvx1mRGU4UjLnNWy26p3hrMcQAjjzj5gD
4zFk4W27kQ7CRTTcEsVV1XwZg7V5t10kCdq1ZNwUl78zQ4uz8BcYqKQ9kQ7n8tbb5nOTRVhQAakM
RV0Uz8c5KyZbnvpLUNx762oEZHqeG6ht1GIJAHgjzPB02huVPR/Re5lrD1aVJbA/scFGzGz/4SMp
KOh5Xh4UNJef1Khi149vthIQ/K1JqlnR5OgJfcA82/CHH2GiEgXpEFCKbCN9BN7s74GlGFGv24nD
mnRzZcP2ywtGcTOxhqT/Kx7J+czv/QniYUcoF3nYGL2wHWXHChE4f6lNZMNRn6SO4whGJk/hR0vw
Hr9t3hQX6tp1ic24fVxcr+h3/KEnvGZlqpgdlYq3V8V7jtSq59s5RuEYdRYL80LwqtEavXvB2OmG
JinHuAJimSx1Yv+Jehh9vcgb8d7uBYxZxU6zLCLjC0gu24gc5LwnPGPZpxK81DQabnhZ/7b7cklH
s97bh86BpUVj7dLZBlMVp5F+8xyDd+u1oEMEwOlyKOn60KLgT+sMgK6qX+f6EYVQY5e3DpgtOfir
9ApZMWlZHLFrLZ7Mv8difjbK77OqTMjL46pWdSXGoJv3Jrlgj3c0YO3pPUW7pasyYQ/DYhKO99LI
4AxegjZ9CQIxpExt9nu9AriICypM8kiJBUzo8b6T8MPp6CVZl5b8W6xitxdMwlWNe9IepGfbnEa+
9YUiGUUZbrlS70cKa8GNzTSEoQCjaio4KPQpOFOhpbzY7WR2TqVcMb9NnK7rB4i3Q/7BBAq5x2Dw
8IRZixI9EVaBJlpRJsSgq0ToL+SDnw0nWw4xlnG5w3x5WpNFQ7xfwmmpzrMzRv9o2Kfr7+qWGcZJ
0BRCY1t7cQ/Vtze8xlS/YKI8H9mXeWn9ZtsyyYqGfkO8U5HYC9kJXm1a6f7HPRgcUQaN1D7EgZVn
JM3zR+uAV0Qj8ZsGS7LMOuvY5oymR+VDlACCD1TWwTHGep+9BEzuoJJ5bXKmVWo/sMVwlWRzOHGS
tsanzxPLA5XOQ5eV3uPTpDBBj9Guv2Khgx+TZ5kBW3ao7ifNkgsJ/ShwB0zEJUBEz1ABfcarDiOt
sr9k8y2O78o07ukugNWAyI5VrkaCGUYDy3u4eDniJUrs3fn8up2448QrT9v/spzLLi0ogbHLCXe7
DN1N
`protect end_protected
