// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.0std
// ALTERA_TIMESTAMP:Wed Apr 26 13:33:40 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
izaiWYLyMPEir6565IOoVp0F+z8ra3FAKZekK7urLT67dQwlSG8siBs2ucpyxi/1
zkAQHQ2P5cpdCt72TSowet7GJ64/u9klK4uYbgXP1gIefJTgY0iuGAfSkLTcD171
+jR/B5dkbw0oV6/rc2087a57wN2SMGweSUOBbrmaU+0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 13344)
bi/yanVCEVJUqOKowGmuQwBGlG/tDGBC0UuR2auukEen9CMForyln4DW85dB9neS
QRXhKPpRVMZkigsdMfwMqC6scyTU9bH7j5nTsMRSJeA+oQyR9UpTqj5TRd4ou5S/
UEr6dYLd/H0NBCR9dq7TOQoH9WyyNBRy4yPWbPpzM+Y0FmyZT/bRzNHQHSDOJhB+
SWNHc0Gf7hC5Fzzqrd+SPo3eboYiNtNEW7NX52t3EVFGP2fEnpGESUwC8k1mpags
trwtLQy5FoXfhQ+9zYNuNyrWvuCxdt48QMhEtLjZFH/nph+vhUpCQYTr2ycf1/UF
xa7esUsL2ZbVKrctR+BzMakVniNJc+e1WgwAN/JARt+phorxXu6hRsssCbNJepsH
bSQQeA7TpK5z2opnfh2UQKLPevQS1b0JPzy0bH/356NDEN/kauy4GXGoZCMt9CH7
CT4k6EIXtkU8Xk/690N2J3hbWSeG56s/9vJZ5i63qcMpNSjVmjf4AIJ9ZGmvRf7I
zQAMW85f394qRjcgWRswP+pKTDJ7YAoHj8MUQdyBonawDzXSF7MQ0vSlIDDmmGoa
6onU5pETAZQjfz8KG7QW/S0bWycZDApwHNm7WDSYxjM22MhN5R3lcBqvutCnkhjY
880X0mGU+4LTcyXN6fYRj0o/zO8CvUZkogFilGbM3V+UptLfC5p6YXDjW/0awqhG
trkqHIK6NtNs20el+5g1ut3rnhyztu3pbHk7N+Y+vqvjKa9d//RDBQ2evs3+RZrb
dj8lr2GZXRUPzhxevg3NTCGI54tLOBQUvORz7/VTxTpXIzpP4yJSi//AZZ8OcBLN
UdQtAX57+r/MTz2VTOdcUAhyMr/GTzAjq8vjuSeGTyhN7ojp7xR5vQqVnadfzdRq
w+qCJ1Cg6GgZNSiucpL5gIGUNoY/Hm2XjTrJGNw7bO4CFwcO/4pZAGZviFO2wKTg
EmYw6cR6r/9e2N9ofkVKGLVvIWIZIkhUNnhJwBBY1lExuSM61HNH+Ikwedu+FkrK
DRyCqZ48nqGV7DrIEJ4LS9d05OmqX7YfLVmByKA7Yq+M4I4wcn+QYW4qI04jBAZU
y6X2LTL/N6Qfm2n/myIk7NucwP3DXmVjY+15RkUFqzpAl7yw5OchvwUQzr0qMhbJ
KnNaeY+BM0dn++kOulPn74+IHhVGKKpqF28OPj3yYZ2vjelACLYw7t5mBhBQ2tRL
IAmj1MC09Ynx7oYd0LFjuzZ72pSi6sfaPE0XIqncyGHA+KVrA6xJ4maijms0rSWV
XPwkWNb4fmELFEuQTQYTAZX0ACPrxT7RHIcUnkcwFSgEs4CTZ3rGMRZz0Tl7KGrh
abj0VYTYk7iDpCvQa6jU0M64qxiqZ+7TfxiDULBaHzQdqcmTmAjaRZ3q1o4a7KHe
aj2W/YoO+7pkzKEJOBekWLUAAMYgKJp9wdyxvz+wmvGyuKcVfWhN8epYNYVJDRB7
AvVmoPGehroZCxc+RsnD1COWZX60DToFwUOClyh2KOQV7oY4N6qFBnNwMDM56m10
rz4J8xoSyCkSMu4BNH1W7z8nqOBMv6LLJtRf2LICkrwu357utpN7qe45Xqv+ce+C
SoU2jDRNGo2Ya2yH9G0bSmq1e8PhXPMTEKJfo6TvJRHEqT7NeDGbzFOZBYJotF45
Ge3ZvnNkV33L+4enVvnhhk/omjwdXgszjXaeY6YrflhvBA0pL79TicGC89QLwcYc
n1BhunxAiM4x/nhR4GOblUaSUkw3web7HTyNKUAXNWaDKE1vGLsuCnmJWoay2PBI
0QHdOKRxkMzwqNSDOLjuotE32FJimoi3rVBFTJ7TSoqdZCabdVLu8q6kVL6AY6cI
AY9diXnldqcpi+nY+kUchQAWfXUer+l9Efc05KXYy1yaiWwlh1IBpM4NTJGmtoiO
157a6OBtYNNaFwF69PWle0wiwJ+qldyqpt+j9FgPx+qfuxLriwiaxg9FVxBV4Klp
8RO9YN0xU2qT/jhtfykWlyqbO3TJAVXjm0vu1F9M7aH47JN0OeKbbphoxThTeJ6w
niq208kiiRCl528UxWzV4dc3OxPCSO3ob8ADXt6jJ2IvLwyeEs+7ZQgV6byRMCDA
tW2bg0cRVlNudJbuArrDQbroH867u00gDGUPLEMxUCOGCQnlPPs6HBamql1JKTQ5
tP3DI8mCLCncZPP0MH9hB54mntlcyiZ2o0ABd02mAqlkeOTHJWj7/am6tqj1++yW
eLSgZkTqtJkKxhNvq2Q+wPisd7BNlTkWBLvHpxN8Tb9u6uuZszHoYItUfkJ199Bx
YOP9g9XjvZweOZxJFSt2rlxbso8mY+S47N7AlFoDWijW9wtB2NS5/bQ6c8L8H89V
HNympmnr8XAExAQh2sjZCGHHOA22dfHrmh0UbAarFS6Cgt3sbV+2yZObO0ZtfOIm
UfBNEf+IIU2pxsTfPHceH0w0LpXEqw1zgg8Pg23fIKqO6qMfdEqnC342dWmyu2xK
rpwat1oZ54tAU8s/DznrxodkNvJ0esVSkykk/qW0HLVYnSq8EAm9ycN0+IgrDXBU
u718IIV4npFL1WGkLisoTNPg3rIp0EnO5lTaLIduv1w+m0uzDAoupKv3QqnHxhmF
WEaw7kwAFHzozBoGzYfjd2zlqyPp9kLa/VOK6V4Q3GPoYxVaHwHpsW4uwRAGGAtW
eQ+deu+38MQwn4X6Xa5kozvMESDjyl3A34q2wmmB+6Hz2x2RfV3xvA61qXz8tX8+
OtwOsnerzJHlAiF0OwlYmIqsr+xgKcXxAiJ0k+YvQoi2WDsbGILFMn0+3Wb9HCBO
hTe0neT2E3hbPF+75mNbBsR3RZ1JeVfhelROnzAKWtyEMX/wDec5Uxirf4QIhs09
vGCHMnhtIil8xTiVjt4QMx5YAtIXWGi43rQe0sYpKWbf30UQ2vSldyu8ONi1104l
yjc32IV14fhELRbROVOrpJIqA2EU7V8sglkJhebiZre0hqD8kVSZrtJviPgfElIH
hhYp8t2xaSXwjOEVDW5Db2RZCmXI0CTItEizNqCeHpt1mAWYEyGvllqgu/CHab2F
jeyEKx5jF1arMJpeCxLqcYOlLJWICWd7rmejtxdID1W+DhS1LH7SDpCKs6IeXmjh
cU7V+v4XBRJlZBb6zXFl/hK18K/UfDRdOdVV/EicrwsgmoUQRIdJ/hQ81JOhLRiv
0FLAKYen09oh/aXQUPBhb6p3GpkJfEfQwq+fSZySd6BM/j2l1lDOmchwkOijhpxK
FDT/t4ZcVlSUPQrLQkAS/u4Cvy3FdINw+P3aQxYh35tQMD5Mp0fA/ZE7IG2e3SJO
ExJ1SRvIRLrcX4WcFOM6nY+2Yb+ETIM/lZmpG7me8XFKPn69lDe+9+dc6DGoHx43
EqfCMHt5ztBma9AQ7BYRO1Z4QMymjRx56uRuvyrtUmBRWHPtjFxibwebFkFBTLyt
KcsX9Ht64jlmxkyuxSnG8ZFiD6Pw/GcFBHDqXNfibgncAI18/rBIDm7YULYUQxjU
5lObUhPAfvHZM4s/ILHOdAUO7by0EHghjQkkmB0ByCuIXmqoexTUffjjeFI1NHfR
pZhcOq4zoWJsoQXTupHQh/sXA0JzCBSzM93YFP8twgpQJPo669ZeOLTGTZJp8l89
VvQNn4/mGCbDlDtx4DgkNSB3dXj+m7uD02QvRgKMxD/107UCJJzaiSSXOo/bm4cM
owAdhR05Y3WzEbXXNmmqj5TAmq9OBpH+unqV3HjO0gi0Y3zI9DPfpjeN8KoYBGPz
/azznU/AsT48aMe1d9ao2PrmD+OtfRL3UwFTYYMrlTWERjsHL87I/euzzgkB2jdr
GnhQ9Bk3cuZCy0XPYoPXd7RTzbCtQ3ZtShcf0oCBVgfc/laxBFCD5GJFWxV5V+kU
9YHbaXjxf49GUiyyp+KsmqyGXC0NjERmg/76QAe/J8DHS1vpuQrCWnXsY389KfcD
prUxqabix9SuDUUPiyKaGvNC3X951keBZ4ZwO5Vy+ymKh+HcDm2n387aA9YLQROW
73O4iNBJBQfQK+qGJodbOyYja3p8tnUuU3mKYaTDfx76n/0/9TYiQVlqqvQwzzsS
AyrDnpmhpW4bxVh0rjfBCrQAT6Kr9jat1CLAPBwbh+4y7isrOQr0XtLS83kzh/sz
fp3qmyiMonGcNvFvZn0z/aMpQr2VzmFdwrZ68TogBGm1nnrsDc7ty5UA94+l9lCY
Y9tAjG4Pa/Vkp+RwVTtkZ/ngb0kPrl8a2ZNjdHtUUTgVTP5xYm9b6qYGOU0ACTMS
FmXR8k8wXFeSXSRlqgNbLodyhcLLbFh4NfQgF2ODDdeUHOBECG4IBHiTH6+7NKtv
10plTJggpxkFq3JY+0zL0ivaG9zmnLWMosn0utrcKZt0D4eTpODa0POiq5jXkXGP
UvG1g5HdV1EQk4jqvZYwxk9VTFHUXzY/uDwjvi1h7suhQ6CsEgkVTz/Yodux/7KP
O/eX3fhvEGega26ueigk5CvvNe65kh6yH/5gNnlkcEOOmpmUE9KgGuWcxjDaUev2
mgy8Eg6SQxFUyIB3X230twnDdNmvg87x97XcDnTdwNNq8vB5l3MEE+kLytIzMHzD
zP71xgdp5zvYQcj+wz4CLL5TW3YX2Kn/MMpebP1TQS1R506aF2rDNBUDMl+mxutY
mN3GdASmwd6Sg5dMlS42fTBCQOa+BJyPn0Zt/jiILb2SLcfiTy/fcJjyuNRGJB5j
DX9FbM4ELld4n5vJ0ejIbgHPtyJjpfM81ifGpjaNOOkVUoX2jL6p1b2wO4hBFwO9
51Exf4R02ePujJ0VJjHcqIxl9Bezi7/NuJZFO9ihl+WI/FlYCcuFrMNXv/qEjOsh
EfB59qxD9zGZ0Ac86oWfWCWpzKT/H4emaBgJep8w68KOYtzc7NUfIVmNsRftH/iP
eVvcYvXbDNea6xi78W5pA/gXnuE93u0SX354ZJaxmFE6ZgKKbN1H8PGtO7NudCCG
BgwG01DqnPgB3x6MEDUNKsdOKdS95YcHrq19VWSSUZ50s4K2WAxw61FdG+GjDk0E
oflNMASVcgVGRecy84Um3QFTVqBOGRGFP1ZP/b90+8d3f/QhUXx2//wkHxMLCd/e
UHEwU/OvucKNdXtG4mRGDE+RS85VI2xlfl17NCzC75/HfPnw5oLYai3UXW/05Xwr
xU0lPy6dm89z3MaFTaQWwCOtT6SXlrgKpHG1XnNqry9eTObAk2VSzKXkSHxDFgcM
INIgn8Ny7Raqp03ULjPPStXVU4lkTUa9oSmwZxOXevvpv5rVuTctrO+lXJt+g3jk
X4o+Iju5D4Ydj3AiboHOZUCDLc3vsCcETpiKeJs7hSR1wX3mkmOxFSRA7yEfAi2Q
9GxAprzGkMOPAMp6A6bF8CtpUbV5qNckOxlFI9wVFfSm5ns3aSeHg4Z+hUbEX2bI
HOIyTOx6kX4SaU9yyK63SnFM5pSEAhkj3IBjs/Yg5UzJgshb+4szJQF/gAQScOPv
+4BCjZb16HO4yIYavfOU0k0Mkw3kuaSK8AdAOA7rdP+gA1tjVYHv8ZeG1PdzkA1F
uTo6BSKI/SWbLAC3/AQjckyBbrRuFIsEhXxncs4vJxl4D8xl6npIRSXly/0Eaz6Y
KiBTZQPMwh06HWWx1ucfesx87vQaqslda9ctNqG3+65rCGkDxp2KnRZY2CI3WqI+
avUkNhd7giSqeSYBIyjbG6Xs/7dq+iF5xs5ButI2ScvqZU3zdwAutPkQxJABnrV4
k+F9ISwR4QBm4wn2N6l0TbkxOGsoHs1mpgtFGO4PXnPo/5734OiuM6ARyxPVST5o
z+NdEhNkCQcGHjyYXtMflgVFtsgQAwWb0tE6dtvEqzEt6jTPwlomiax6QayYObmW
dGhhPQDwZo5NsBoWxhRGQ6L0VGBw/6KFUmu6GSRPrDcEAY9c78nXQzy/hB7acN0U
DplRDwdauBgzH74jB0Entj7vaM6nLwyvvUZzqJugGUv9DlLffEbsdP8X3Ph6gg9E
c9kn6cUoW/HKp7e5NfOjqCjzJq9g8+F9CRVCyu+hHu3AyKqFIp1d18JpwLiCit5W
W9I9dbORJ8XzX/jCghKSmuOkhWYc4lSTtJI/pHFk1DBQUG1szqJFX+8aVVQHzIqc
usHQHGF02udQhlo3lsoc+o2zZF6sAReGFEcyLImQwr0gENAHEi0bIDk+844njmpH
wDUQgYIFGrlgB956XefrEzx5yc29gCchApfTvVSDumOwe8yXanXDiXGsV0tYej8m
tpd9oMCtJ1hGcvjVF2N+PgsfAVm0BDACbi67e22nLOJqSQA8B5onJc0HkohCjzNe
RQ49ovv4ENk/OJHyZHPB5RxeZRTYKlsSWe+gQk98Td+lWGlZU4b5cEp1+VQ3boAR
JOC1/pm1AhQjEypV3sdOdnwBZZ3YeseZRiKLzaclra5kAPKEhEuhwiwIiM6B2W+H
ruZDTbEZh9bjY8q5+Tu5ZJrjvsgLvcg9XvZ0lKtg7UHzfJqE5l6CVsSYCzxB4Gca
kw02gjpuKewmxV92Khsbn7dpV1HeSrz8GApBrVvYyUEKBp3d1txaYvV+UT2J62QV
kYZq14Ae73yaXI0zb7f41o31PT+sgaFlszl49cQF8sAtuqhZxq22E1dylHekfp2P
eRzOm8rh5njGZEjYU4K5AxZhcEp6miky8sLjq+nijnfRAP3e3p2UUpGNmryPrjxT
alpsM1UuXasyAAwUquqe8Hdg97U5/52odD+bXKOgOvEK7kaGvfuSIH1mWLlLnsos
1+IxLo7A5TlVD33Rs1Q1OKntVl15GJ17ufoMO5jrO17VXz7Bd7ZoPdiXPyPX23J3
pUqIDbDAF6Nhhef55hBfn+XGBlBpql8q7sYA//k1shZ6LbYa4Gid4k9oq/WaPnAK
wCa00VN/lfn27fRb9rRdweXMSIhpW0q4cJiJtjGkPrvc3iaqOFPQWjE483IfHqf1
avu/3ZSkiuLXLDitFFA7HMliMUAkZMTcf71aaLllmxyuNe1k6x7DJ452XIMSHcj2
gD5+nufqlpDb4nClwH+Gk4hgX3RtJ5VrgQvukNlb+2pN/CAs4LXxfxJeQWoJir0D
Rs2woG1QBLGzJnwUL738zzRIFxOG1d27zEoPFEG8O0A7QvGLFZJUloAyGKCzZWMb
PUQZ9P0fkMkJEzZ/jr1IQipU3rnEQxrzi1/Y1I7LnRrujcyabztrcsYeuUZ6VBEJ
vtlrDA+rJh3hJTirSP3sydzMvsHFs52ZGOO2+FzNO34re6tLbCNx0uKlKKe1Lrvc
VAlGb7TP2/uilzL4BSoXEhNkZvg+DebpN+Gicvi5Q9hvEmJG295wEn2mj4Wicakw
T0GUVrJz4TSy4nzrsCtfWdcht4VSM9yLmIJuMxNbWZCmYo6n84Y/xaSdShfpo4Ic
QkddQgtI8TkT7ZfOH/aeEFjz9eVTxvNcfK+mgt5Yb+9G9MxW8ur9TGFsZbjmGxqZ
e7x66GariEaqDItOhZQokD2kUDQ6MTn/5B14V0uKkNe0MpFWqh1qPH+mBywpn2Qi
nqejuE59fj4SD7AlMk5+ycycK7Pr3xc+uuZ4t0BrKfU8U1+8pzSOc3+ds4fDYI6I
ILkrBw4UnNt+Pn6COlJNQsRS1ayH0LuxSTPYMLBK5vKFtk0ek0x5LndItNh2iacz
HDlLlujAJBVvLc12Tf5bRmJvo5BZndOwRK2PC60xyXl0gMt7X2Gahgei29u1exnB
XTxl5WD7ccZAsqNrJNiUCbb90BagAAtOr1CiSpGFJfizshH5iIYlvjLDoNrINlof
Q8NPfFMV11TNIkDArZ6uCm1SRdTRZV4g3MTgbyrj3QCMsNrVDz18hK95IvJ0DmJu
KJaAyOAzXT5OtvUlNz3wXjz9cOxusrOVFi224wDBib7WqGfUfO4Y23V3rSX0ir5M
aNmnhMqxapEWPfMrPu+BwkFLtgS7WL5ERV27NyhlGJWBmkFxcz7adtAY3vTmjsVN
FOkiwjqDmDq4kjDCC/gxIe8W/r6JFr8hJFJkR20+i0naRGlVYd9REM3Q0q9tII/H
iYQUKbnfuxjxULo3fC0KyJfjbApIIe0YtcbunE6uQN51OxxmaSy16r4FX6owXzen
QB7lBRVaZnPPSCepObl2pxHG2Cci7W8Y82139Xab506cP3JbjVteXoswYdMw7V7J
J44c16UU5S9Mytb5BJYBOTQwVxSkMD+Z8DasJiloMn1kd05o1N4mGW878s7Syh5h
BMgU6k5WOmDdZ7riNsqY1jjZjAIEqK6Ha52vcrxHKnUheeRL/9KVMP4znbufvuZZ
gYlQ0iFKIio4LvodhV6/RCtB5KyFSF5p/+j3w6xJvBrfeoKui8C07gP+zr4fDzyf
oGXm7FTsf70AunrhNx7Nl5qgkeEo8lQwyzqoTB2R9rAQ+XOlppdFRHSScwBARXr0
2QclL4VbM46TjPwVSrsxm+bOzO4uWyTzKwEzmao0tMUuh27mObGIkq2gWCFw+n57
f8Hqb+pDDBdIv46FhixQnLpFWTYgd1TQZpQwIrbcxj265wNaiTPGoJQHSs/PeJ8w
Z7wWGYwrP95O4Iv2TYp5RbzDIpDullGXT8UUJaf55wB+6QQ+8hxbmQw0N1TkBFT/
fDOCcuW5j8sA0W0XwrZC7TA1vEMbYZcA1NwrpjwUbdviP4WtAb13sVtoyurUyAMq
goo9f+XONinSa34+c+sb4wkmzJsE+n0sWNg4rDV6hYSgwDAKL4A67dj97TwRmBvP
yOhp4Slr+Xnm5+a7SFGqyYajH3VZGKsxOcWzdW9+NP40OyMqtwILXMbhQBvm2FIR
SIym/JTCa9Zxv3rM3VHlrROmzX/6LtAKNi++oFFvrXNuF7L6HO71l8D7WDJcT2Vk
g3hAR5/eEt1y8Py/DcCwTP94HZm8ZLqsdurTliqPqt8hNFFZE8tlfMPwKyqapsmV
IQJi/YFiVdq5WQa7z5Icv6GXFGLmYZACPplQRRHV+lG9+TD4q2BUMGgW/bMXzHXA
XXyPoeAuhY3p5m1bEIH+wAs52nGGkoDGZ01IsWg+pZLBi1Rct7JChHeFv9eD9hvw
YOlrPxxfBgcy+KYkn7+O0bHT6DsmNnt6NChN3T90e888LV+ExxY14Zq1tx3SgY+N
x2RkP/F+eCe7PVNVum1D7GubJyLLbvOib8HONywsr6kWiZpETi4lB7H3kfpaP0PX
ESfv0t8ko9nKjVf1F5vh7BUp9q3kTWoiUEHtH/TbIiAzewDtE/IuGIYTdVUpVWCN
cxuJlIOaJ+eK17X3ESs7sySoSmkj5jeGtyUxiPwh+CQbt7m8Qe6T8YONA/X2fTYf
iaPm0fIu18NQBwqmL+V9isH4503XwPmnzeGqfP5Nf2/vRuzyH+vyINLXZZUE74CN
CVE5V5rrN7otR9KAXg3k2/2CK/D75YyGtOlJCHfJXfwRWYlxvbB9a1hlAwCGPz/C
Daa/plMaljWYYaTPw4AikveNTV5OUH8fnVtB7vfCszmFdpO4FEjyfDTnC3TDo0vx
TO3SEYfRoYMbt+qOIzKvq5K//PzpFZi3gWKcaOwOCJjfVxngS20AXFlCL5dqN8yn
2AYieYseLu8V02arM3I8ubH2K00q2Y71JJuUVbYWvcEXgR++K5oP93xIph8jXrV4
WRh0vnWRDYtprepUFhHV1iqoXS9wIsEaXwhFWhyT9xBt7YfbFZyVEYWDB5KEaAyM
imXjbMQh8w/ZoKdbHM9FHS6hh0Gben0qW/NfiWeHjZoDwB9xIWM3cRkw7sus9ESn
gQ+kp9ocEe49aLLAFR6CXA40lgwev/VBZF+kpme21CEsdisYTE+XXClLi+G569cp
Fxm1LXa/WjrEJ1s7GO/QpoBJAmEaSRqqiStVR9KsYKaSrY9XSjRVxpKNYGS52zU0
XL48ohDCJOwJFFgxonbGUgd01e2tybAYE8mlSDO7GkXN01fmzw/oIVFVGW26K63P
G8CMJSQ1ct+2F/+OKTLVCMb2lpOZYBaplll+tCOCMKNqDnj+pjNWTWHiONCaKqZx
gJUWHx35BcPIYzJLNx3MCQaHP8uezqVaT0nLnCqEj7RzY+rKcX44Kgvems5hF+hX
CsKtkzCypC9OOCUnvItOzUyqI5mPpGNsWwLiASMgG0yvBIB5dQe4M9kR1KBiXk+I
VG0RlezutwSkRJMqCgJ5XGs/vqxB1Nqg3vOaCZZuasCOhrpX41zudXxBRuXW9/bJ
6QcAMk4CZ7dhpRhSuFMX4OOetK0Xtm9eGGrqmHKpqisZadxRFJUeE2j6dy2Du6gf
W5v/GWlPTPZ6076q+tRVTa9jAafTvLWXX47+ZPj2Z5Tf/lqHGGcdfdI5wsvFZKCH
lkF4i2tmdujkl01u4Fny+2yYWX7L3K1kQ3Hx3NqAnRMDRZDrRFSetl+9BvuSX377
kn0TeWWcNDrn6XxqMjagI+IozKrdMZGE3QPYQQ70P76Gt/PVsAytRzdgCcfFZwNA
brFHVh1f1ogiDWxfu6i7rdUKSAiC0DYnPFT0ym1UBdE1gSzttNpD3bRacBNGNI7C
7zJxLUpN6zzAbq53C5S+N8HdPlKrARYxRJKorGSfZj5gu+ZC7QYHKUJlDflTaW/6
fRFYLIrRuhICBz9Ua67syQ0rjEUq4f96Bk0Pj/Yc7c+gNJPg+1dVHSFbqQUYPz4u
GZl2ozHNsICOSrGb+uvMud9KiL5N9blG/gYSLIg8/tC4kYuVUt+a2WKCx9CMbWMN
zDVZ4USzeEGH8GwITmKPRQsm5YfF5uld7H3c0jeAWJftq9AqKVyeDF7skiDiudkD
2y7wKwljzjk1ka+9N+JfwoIFzQrfnaPPW2O0XGlm9zArxsAPfa+LRxvGKUT5QuIZ
jq2pdLm9Wf5lI+kKD3ET/blx0LAJFgGIFD6s0Nv76GWgIy98FxaFIzemuQl7KWBW
Z6AeY9bIIL7gpy5nWmuBkZKLWyz4vfEPsVYPUY8vCuczBQf837vvMiVDUgapQg81
Bh0WSV4dmgJ6IwonSjB8SKGcclqIpqEjtroA9iKSIBRoMLJsIFdhjo3CSjI0tMXP
0p4KPZBkU9vXFaE1I3f5OGsMwUxrBfPrysDNDVPuVQg3Ai/+Kg8s/APx5E0Z3WSC
HOsMJ5lctxJ9iKh5aDUsN6AxvedzXMV5iXwBl4qkRwMzfFBAs3/G3XwBNZldP9mX
ET8Cpuw8xmXtjB2pX3z4M5o/pRYi4dHGcKoQrZsNwKdPh2reCD+x8XJx47LWMX7k
fg1STtSRvFCafaT8vzllL11ItEpNHfTlgxPc6A82MeXVsTCzgjEu6tJaDgif1hfm
gNjDrdd92uVyUEnmMp9qHDyMbyxQnxhWhXFmeJgpCu3RAEGTTMxjsKmgLHWwtQwO
NAgqJyIRAZyjLbDXmHK6P+fk5uBN1thFSo/cRgqbsI+pG/zYVgEweSMMYEwezXdA
Zd+r1JY/709VJOVE5imYgyAf+Zwwcpy6fGUpEuwZh1bTSxX5MgnvKldQM3HKKkYb
leaBZFJSWssPXLEM8Fv0jGCfSLyybEZI+dQYlQFgzj3OuIYoGswZkGz7Og5LICwQ
nviD8ucuutCdy1BlMtCxOsDU/4yocJUA4dyhQ3foOesk2kYaS+OmYT0uuoRw8/UM
GH75GlSqCaJWPwbF91WoWNw32OahbH89CC6VtIcDaWf5D9FW7tnHTktjykx70Wei
jrkpkdfTCk4/KPuDP0V1Gy6uZCW54o+LaikX+ulyEAQolkc3j18WuK+Cs5s+oauu
xH4dUKdx+v9En6kfR0aKYgWCXh3mZgnLm5F8wEnZVefBKLR+rPGRiXwJ//N0eiNU
2TFFRy1fH8Za4M7foz6O+Coc604V+CV2X0u7FsnsI7dVdg4CSbkXmJDcFkcpA+sB
UFQ8vnQxyIMj6/Ggc2K3nVxDRe029cbupg2iNKT4cQKSonwFEfldbkF2UE2W9nG6
II/MgsPnAYhelcdR97FZjysSMNrs2rRlmma318e04l1J1qPX9HnLDfLa2YMsEMNp
KF00UjWDTh9IvR7n9vcmhXaMaTyY6wbf0E5GekOG3evlPczjwSAVrijMeD5i66qU
IPVFFyC/2ock8q4lXk9JhnqgIRBmb+pxV1X0wbZzaoYQ74z9TBqTqSgyOhgts3TV
2rX11I8E1kbGl+62fMXceJGMN7DUmoscqaSh6+gRAKUSg7rX6vmdm9L6Nt/DJewf
EG7IJ/YubgZsJov0NnoC9HXz+Xwt2wzudht2BCqD21R83Ipc4rnIBBA/m35Z8GmY
gn6LKJQv+8NLJtrFfaRYGD1pbGO7kQbJrk4kBlvj95t34MVoNm2T0qNqxLlZgQLV
qH0057Aeq1CegkfmHLJZyrox/btY64ANAZx8dTlJk4/8GiIfs2wnncwaxCyidZea
4lglt68P4qrUteyy+Q1dExOzYud9N1W8FAd8S19K+84WzVj3N+R0B6q5O5TQuYJn
nNEYPTfGOiM701e/KlAXZt7KltX+KoZ0nUPqKF4jyQt/F1fwvHLaQYAREf/1VBss
zoQCV0hr7fX/v3N80eq3oT/iboAsndFXQ8GfGWRDafD+4SFWwfOphvRm0c+sFQjA
vn2BfUGotbcxILbt86E1hSgdoFiszMaFAPINV+pMBefh+McJdv/FhCpaQpXlE5Xk
V0GgBSRtsnYm0+a+9mJUAn2cBjgARV8MHFVEs8nxtbRv+uDp7Z6Fd1TW6zoJKLRK
HhXulM/WIzIUdHcM9g2t3qgFHK/SYChO+s4Th1j08Cfo135TtRYjnxm2kw4/5Kgx
0Dt3qikTPWOX8AjfY7afTeY3ISukx+uz4OYGFM/OPCep8K+/AC4FXWmCyyAJ+21+
wxihOyp4uNJmaCD0/p7CRJTOKpYAJfaQmA6Pmr6FLmcx5brAlQWZ6VBldCLWaT2O
prM5V44F3YXBqf4JF2/VUpf1jY2mWyu7OAMGewbPL6fNrOmWALspJdoeJxeT12uS
ON1xLSP+RmziJ96Rq2sOeUge97FvYZgIi7E9hKpMWzsHRxLI3+f/UMSuHxEHTSvP
mDjLQ1c1fbayiM0dfcnuj52yEXc0RYMuhuooE7ezxOxutR9LNPVB8caRytGEBEoY
ydHQBP7joaR5Sh9g0Jyg1JPYdOwhgh6tQbq/FeHrQPDHAb6z1BTvS7LqI06HTOk7
p76WEZN/EUoq2dqTI8B2Q3wVVrFVbct7t3fml0bp9vo63Z6IruXfWqEX0G7lXRUe
ItTSSqj+5zSDJNtK11ZytnTLXHIhiE7bmYWGqCXa3YSnDJbWoqVqJEj6RQbhHENW
xeRYwzMWaiRKTGM9ZGRNlRDCNfB1UJZJ4GBeNuONzShTo9Eo4jvul1YnOhhU51+W
dXH/ToXfhCnogG9Jzu8Oftn0ep9arY4om1BVekOjZVayqyZxOj6ZKyPH4j09fI6D
xyEI4SrZHtx93fy/NUDrmUwbo8sqBvYWhRYp/IcQJozMfIriKgEZStqcNvwlp2L7
9iof+ZxjzwZqHzKEp7vMnYYX3JlJrWrQnSJt1tl/aO7rhkwWcKU3sUANSzu9lPz6
N5cDHYSMvnGhbFEb0PxQ4VPuI2bfsDzalvQGZQk60OUBbAEZIH/+nyFWopwntnQe
3TKuG0mOeLqsNdLeMFK1F2CwzDKx8mf9BxqtFOn6dPmSo9qtgAyPYvel3yudeRho
UIVUOH5yvkIc5RALtkff9sRFPPBv/QrTrlWAOHsnziPX1K/BqeomH6psT7E5Pom2
1XXJ0XKMO4O6xx0T+MovYSRygInQz0MMaFUxqJULRYLHMchWAV6LsKTCDoy9rj/j
zUZm7LlgWesR4fDmb3R0CJ2poL3CguHHJoRYhWeXuJFf6KotahFBCSzvt/mk7P/M
PwlBTXWtxMjDP9ZtBdME9Fb8d2H/a9U3Olym15Rs1VNAhmmLI9438cV5OMzBtzjX
vAueISrU67W3eWkYsF5DqYALhmDTdApdv/EGJVy7vraltPWGGuPbwjeNHeK3mGFc
p9OXXUQZAfXmtUm6SiWpMLsd7/U89ftl+Su/2Sn40PEBBgEjeHmjC74GunQZH9BP
9N9lzQi2apRQJHBS6ioUyh/Hy20VgnYU7gHIVBaOBtS4BHYIuNVG7p/9IPVPXrpP
paMPQvSX1zHtZG9DQkAoq/VCoBjh/vmcGoZPxnBuPIwCxZjMkTm6XysAgZOiAkdB
oeVH1sv22Auc4gUvy0zltDTFqHDS1+QtlEGTzsO2diHYQpVMlDO0zv2cy12lZW4t
cdQ+1lnvzT9Mb9PxtN3pEIuPii75pxzKWFiK0MCygfPB0ee2mTdJWE2xvBtWFvR9
C9n1AXvVP32qxujOQtrv9t/OBHCD+UYlKfTEBRxXKnWCZfJRk5XG2Y74PD7gJTWD
VMiPTfn1svblb1/kuAQW0Cs0rTZW1FCN205WlWnSrv4vbtzyu/35uYn0bb/38BKk
iIrSdf3OKu5w5NY5apBBXRGCe1UploCJ0KnT+D02znvT9OvDQ9KbOnA0MD4InAwc
O7UNFBy1DxSStL7baSudP5jsPOeYPjd0bWsE7eBTil1HM7X9whmp3J/zHSz6aW/7
cWccSbnq9Plq0UjfSfRT1ko+l1UAh5L7C/IbT5kevHc2nj08IHsaGHJeD8gdnrq+
E92AsRykEyYI16iSdC+DjPH6qgbmzOk4K75NZezhEfdeKyhix2VGEaQqgtvCoLvb
WPYNKLbuufLB7ACdsPIi0j0I4Wn2JErWVSdMVa80h8p+LpZjlKLuwVIx2hbZpSNL
RThub4jW6EfZOXPL3ENheFP/q5ZXij47tymWx3KM1sXuFBc+mj+JwjbXYLAYXbmT
St4e/F9o0EHHBhz8L+Yru5XZ1zUoKJKsiwmjr+68pptygUmpG94vU8X06DPHSSMT
iG8HE51CCteguw+aN3YsCoZNE8tGX5z/4VyHP2+A2qnVube/sJysFuDDLdXAzq6C
t+apq3UHnfROuDCbVM8avtFxeR4HosQEhjfTCVd/fKRSNSy70x1p3GWbPnhMiuz5
wUhEbfa0g8nykBcALkBV7JEFDzvrGtspbF8TTZdwIhIxCgCSjs2V1svlk4zAES0t
9u3miTCykvKHMWb3k2kOJghsHIBqClxkC79ZbosSZYVhJiDGw+HEE3edaOMzRHlk
zfj3fY5uiv19HC1JqxpJNXNEJrVRQ0FRQRZE4ktcy+6g7NM45D55f/AuEwfAtsqR
6kWdRs/KdLwnoyOVECiisMXBN1PtoFfw7IA062Lquovk42qJLcCPVvRnZ1nv2RLb
jI4tPGN6WQiO/mZ9bSBHFvKOA8CczySnUAHhi75kfoOTZkuVpkslHnKv2RJdp7fp
Ezf8kgp4CpTvgeZfFNln0p3L8sD85x4C+cbnfX7u/yH0e8CMn3YU6oK9KGvWPLvu
pZVvhsbNCpKw3lF0g6viXFVSO3svDLeMR3rDHMKDGO5Sk6B0QRayz4/dee40069I
bNcshqxsGURryDOCFcgBQaScyHJfHbMUuXBBS6NLsHzfLMTlpX5EaRJ9nTicN8+B
fMEp2Jn6JNklVENav3Exf6MPhrhV7L1ZLP/+y+6kwnLK7t6SUBxZg716SegezFMk
JWZ7Oq5Bj8jcYURor2KBnbv/fajk5pyfYo12v3UOc9gcni3oN3beFo44J2kq75OW
21/k2lfKKITTXWBnG6x9rwRGDwOB1WwjItarfVk843MpjV+vHadf8WEeR3dsyIbs
JOzQ2Bb8FWEXSiMiK3seUyO1wtERzC0jgZhUZgt6kpt/6KdIt4fGR7ZW2m11EssZ
7MAb+WIEHkjeTlNwv5DejGF7x++IoejybFdVRWd4fU4H26SLt7l7Q53cPbukYJfE
NMu1snjb8V7M8KkVG9nioPNgQ8xBXJKj7knU1p4axM7B+TEuDcigCAe+G5WEUoRE
8VT/N40qwrSgrz3GwxLImnnxCl5Cloq2+5yNY1+bSWLOnndaS3jM8goj6wAqUqCY
Acvp5t+bTF+ZHEOm4Sqy55TVy1poBjaYyDuq+/b+uau0poksCYmf+Qp429r/s2Oc
DQ62tdkZtuNhGMP/Y8cxUhTRHgK08KzbI42ZWloj0LyxUSq9DxcCJ+alRXUw0A+o
jBOQYuCrlWfvn3Fu7kKpyuA0k91aSjhOVqzBJ39/he+6v+XU6Gkh81oWP50mdw0H
nccR0+BWTing/3Az6S/Xhz/i9123yIpMpfKxkCcTJ0ABek7PBfZNP/jvYwyTkKAq
aCGPoskk7uw+aoQAgjuXHtMUOXMvTwp7AxIJMZZzec1hromfRTR7jE0EsmrhAUR7
KuzN4Z7WDqey/xs1HeX14264e/GcLOWX4JYaRYP+tTCN2R8c0p73urffjpEdxqnV
Ocq4ux6k8jiZ4lKDyPYlssGXYEQAHZ0xiLnzE3Vf9b3dMHflUztm9a2Mm7RaZOr2
wTsHXi5tjNZnTitue1eTPH72+2sddpCByCEPqULsU4F1+z/yIIWzL3RR4D1QvV9T
ZtJaOw//mnEaTAB2U2oaapBWA0XxCKxCxbJI25tgEJBvxtVrsbFiC77wBTH6lz3M
foiCojnjoi4XuFBnNxxnW6RIpmrRrtOYuF7zEDeSS42jmQJgiDVgc4mxYFQfXPJp
4ULta6x5WQFDHe2cr1kxLZEMAFaZfQnc2S0TkzB3hqLqccbDcuhh5Eaet4fcTYXo
89kQ9OVI8i7NbH09Dys6EGmex8KX6d1VK6EgIDDvN8+4q+P1yVXPVHxTVHXSEuje
gTMVW4Sysi3Aa1bV3YSUor/HjOmTfeBIvasXyjp/gzXpbrKiUoGwAoN7ChA33tGE
RTpWemV95Sh+Pj0YuyFu7mS6Dg3KpQF/ZDVsbq9z4L2EFXJf31jz0oj1jnwa7LBU
IMAk4EoXMPfmL8EcXhOBzPwEj9nQBKT6lloq7jKt1FoxME1Ch1U1XFd9N3dbmvNH
bBCo1vG3otL9SSRRL/yLvnwpvVc0p665FZkGZ3XNPdNqgpI6SvKo/sDMW+Ja1Lz7
sidd6q7WI8t2n+dXcpFQuAB9nIKOVocV+BmK5coRb5fqy5aNk/UH8xtKoTKGrGuE
s4hBhM1jtEgVgmwA+fXpf0Yxtjw5T8kdvxUm0C+j+dR0QTPRmD4k3194b3+9a/F5
37OPj6LRIJTDxq7iAp8f6yzqcCRPPCUiiVpy3WmLHRA9rlmDsq1/pGFgiMq4SMmn
zBg08r7v7jY8pcFLsBv9kgpZ5KfJdNIEEMiSJWS6I4Eg4BB/JT+W2T6E2Zp9xbAT
h1ohPrrzFEPkwflVBTeLiAuOcyPO/WYxO0Pbf7zn/tnwjQoGbA3jff+aOW/Iuqaj
B2KibKw8hje59LUwBZynqezulprYu7EBwB4jcNGSPmw2CZhCONZM+uWXoVQwlHM6
zTeWnCx+MZWM5Kfv51XaJKngXiwqOA9EDPZFjo+bM8DKcR+JhDLOhDAq83MulC9R
tsGuAyFjPMDYzBjp4WdGXgp/EN80LfZ7A8KRm5Rqzj74RbHW2GDUX+1fvsn4CIuA
CzeF66Ethy3qpWA2bySzVm8XXiQAYnZ9PkBT7ZOBqbTWWfbKJufgE1z5FD7n15ZI
zBiozQz/zTY4F7afJcdMrBLcUmB1jh7fDZlk5QiCKZzeJUmkuSgdAkULmsyUDvyW
cp5SnA23J5Q/NkevfG/yzy562YBOJmKl5iqq7sLPFNW1vts5V23xdFf9HJ17REiU
KNHlEDOUP7VXmr2z48DLbQLd/20YOlTXcfjyfOVoICZlIHRodbquTnjnJNg/D1ON
`pragma protect end_protected
