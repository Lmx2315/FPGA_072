// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.0std
// ALTERA_TIMESTAMP:Wed Apr 26 13:33:39 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
SeB30lz1k8NN9Sik/07KS9JjMAWIK2CvZ5Vcxv7f4CFPxpHTmc/japbOS3i1WJZz
I6/AG/j5x7FjTsf1zKNn3HYJMzwx/BWSY4AwTa9k0ZwBg3qYHaOh/rmTI7p2TozH
Hs2UBodvFDNSYTNVBUmc4BA1znxGe5NtGavPu9wp6rU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 125472)
9Y+hK2uxOdKn16he5bkQ6iT1J/FKiOe7MXj77H1CGvSgF0rLeJdnq6SmV5jqa7xp
x26EWzP/304EdD5WMD8Q8X3Hqo6zCBzjkw+xA533fdSthBrYtf+ewOqCUrva88nz
49Z1lOOkxA0IbMzzQq17Pciylk72AjV0sY+y+ZZQtkf3IoDiTGaK3sr6aYdrIh2d
s2MaVMp/V1KtTJh/CKjXn1Fhz8LYDS/DMA5pTGHsTm9gydDl0FgkBELIpq2ZKVUi
BVHxauYuGoHt46wyzGdGSjJB1BgQMoNYEHTSex3Nvm/iXZJa4R3uhH/fLuaTvFyQ
sD/70yI/iEiSdSKX8xSXV8ZCbVoEr7e5+MOS6JUB9fkXCBui1Qbf3MHuw47VGk9D
O4e1MiA0vz/s8TwMhBAeX+5z1nlesn1pkUBGE7Ag1iPXF8P3bb3EIesZhHl9kFm3
VeCJPdRJph2FCnL6IAs1Ox3bbGxictlSDEsirRfVZgnl5v1V9woaJWKTpm39MmND
otVz9V7bHRUgp0/+LYYppkphq0he4ZiYlQjz3OzxGVkToiMS/CWMLNP+IDGjfBMr
KKoOcHbEjr9yZm1xtUppxFUNV3iVe7cgPb8lpPyLh+2B8awVx1NZN+uJ2TcTRKzK
hLz7Knbjjd5pqNDZ9MbQRUBP3vZacyQkd0m+wpsX/nQsuPxlneq1i7fNl3fzhLYg
2JAaHN3tgJJLjGsGpa9ykumihrAgPg4isZpUU1u5M7Kd+HdN0LjAmu49FlTRMzO6
xQf50yA1++3npjJ8+QQgkLc58H6rZG1EDLIpoblT3UQre9bnO3oh1bS9IgwghErK
TD8cScmi1LZeV+R+WMYTh4BCvCFXe6srymz80lzdVvh82UNfCnOPGZr/Y/DWvCOm
d55l1Eq0WKdhBsrlnO2huU1kgMbaz1BTPeSDCCWnTGphSvOVe0cM3CeQ9SRQbTuz
eRVdp06SumeratbQsfOGcVDhCrqkHvVMl44+MBV/0ho0dOYYUUO3ZM2ver4unsFf
27LORKkjwL6rE3XOQPCTu9ajMOboMezvs3s2JfmYEwDuGPutLHesgHO18jpCcKpZ
6rgE6P68xeg2iHf0npO18JvFymYT7kF1Ndgc8GvglUfSYr42oDf7mrNnUna+sNTC
DC23JvC1QfiHKySzt0MYQlr2adrAmyJ+Jbw/VtHsoT4fVVNeD3efW9e8zXeskVOj
TFUxrlaJvYa9XusdXIPrNJPtVy/NdsRJxoi+XKKegJrZsh1zow6C6KoMJ8D3r8AK
H7fpmbUft3ezbZSf7uPgJWhWbm0gVAtssk7oD57EEIHEmuk59xwWUMTN7ctfFS3M
lD2a8XvHBZjgGl7nNPt8bLDvsiozBPMX8jf4RZ4H3KSDLqODoqSxe5NY8eeQuCLL
iyrU2dgAAuU09nAx3y0eZaF3XvwBdTRqeYEhJZPHdVs0tRe0bTlilE4QMLYFE6Yo
wh2E7iZrEs3WcnI2AUrD5Jbwoosd5iOFdhLT7S/ef8Oa19/UNNYEJSk3CF/HnBDK
+8FjIRTaih+6mrEa1P85FymEqvIDqTDhyNAoxdqxBBuiOJj6wVi2rL0ox/jbeYdE
76MYipR5pb6Lw5KM++bcsWltCRDBjgSuDj5L723b7D5SLwP6hmy0UpB8rSbvuTyl
0bdTe0FSgw4nH7WHOISfuJs9AtPvzBFiaOxMmtB2+xZ9/fqEXBFr6F5vundKqqxY
QUYSNOlzY+skAROgbUgKjmFsYUFdOJKrZMMZgCArLEsW+OlRcymUV1z82GJisPBe
eLRqexhtk5VqQvfgPkKbnnyHaQBn/T3xg70MyXsktfOyQImcblW3MPSKWYihbirM
rztBJA60+QwtmMUU77A0sjPxrT6Z7h/cTi5rLp6BiUUt7hP2rmv0lr2MVkp7A8Jy
BhoUuR0Vo5l/uZmddyXhNfSdRABu6qM+1K4juGhc7Yt0vfuwSFJX+vrNe98qQOSK
4x9WnUTmNEimRikMTS0HeqJhyH8ZTWKXrtn2tLdRR4ERKUn8VOhCkzcoc7d+6L4F
DQhp5+LbaNfNPZHvO83C/sbiN12bMggHFO2k4/UaROxSMMBdgkCpoguapM8i4N92
yFb8I/z0ZFmqmMveDiDMmsQnQhCTen4p4TDEyLHgYmit7E5PZ0irGG95e5PnWXyy
lLRgadzLIDweCTxSkbx+0i4co9DGJ1RLnuRO10uxTuiwdUULpG7d7ezgFsGvkBgy
iDYFKlbGwqxz2hZ/q8zX3ZW6Vg8hArcACxecKojFafo3dH9aMwmQ6iy5c9I6/cZW
zKKaY7oBvj7UtdZiP1ZMGscSx2EjZPnQupzdgR+v0AqLVdsOaba9d9IWfab/WrCk
BpATbH4hI8UCYVq64v0kfFe2BPjZOl/U07dWZbI0G59K8Po4aM9epkLCG9Zu/y1t
9EJG4rDBIoRIh+DjdhROCeBMEXzUYf2zMwt1JR3Z9MaDbYayyVFao36m4ngg+n9p
UJNx22PC3PkGDioDvFlYQvPWc6S9CH83eUEMzrL9TSZrBXVNLvn1p0BSX32ywmt6
Zpjef4WFCvxIGCrF4/6CFegvKRQzzvjssT0rUJ3qvlMdv5NkPYHKw2AiPbZJKTN9
3s99VXrf2OFOTiqyyHyBI+FicZ/LR8s7bhVlbNSa39bUOCpdcB3fYP2w9vgGHYbA
bm7HrJRqCyzk9Ns0kjwp+TaeBPMCkGT3daMSV6z+UBTsk12VcndmAra3KlZdI7IA
xR5SoVkV5j/NzStkHiVaKad08SgHZIfgb7uhL6sw6Dp4VWCXhxuet6tB0ICq/HaE
5CysUTD4YT/e/LEXJeZ8xa+FZJ/fpmozJ4vwNNebBQxxv437bx1Uj/5N6r7kURoh
kaKhPFQwUY8ONDxu9QYZ6HlnVPcVFz1lsgbPYH46yNl3O4ph6v2GxlmT9zwiop90
Nc9B+Fe06vdnkhmUcGKLtIAenmfJRU9fvn+2aEM2emP+mbXpCwi21T/FA5xvk+8W
kKMMpB5KtViEXNQdT/2kTpWRoqCYArRa1Ty5P/ykDIPieUAWaSfZfGlHoFLUhQEG
TNYTQeAz+GpcJ+QxZlc8993lwC3FIkJtPjCOmLDwPJIOlT+qosATHn4W4x6RQlMX
B0y/CI8ZboqRidJ+FBqPEk7+sx71DPFK/qeDa7njOI5FS0koVHomBHuVCA15+Kfq
BhscND1LWgyfTk3tPhmkrqzh7ENynr6lQIcNtJ3alANah+8qWTPF5yHXzfNhKb66
ssMNWxfa/uC+zafP8y/GeHnhcZGKf2YSK0uROuKGS4Sef0UeSORVHBccHFV8sfSM
q7axO5fn94rKJX1FK0rsYqO5l77qrqpHGjeqQfCSJm5PTxGGif6x7SDUWdAK20KA
FWURhVvZTHCSaFTXzUK6vFIVvE6X7JQfurlWK3lPyo0CDWKpTZyiiujGJa+eU595
vcSpzEFyBsqu73wwwKlzohUYb+GiQNKDDErs7O8m8ZWbsnI75tcOyiNVEKOGOMJR
w86HmjSNagcCLB1VQzJUq9x4hmdtL6BFvVfFBAllqSXQVmudzwt6c58TGOdiqMGD
XBI8OMJavpZ2CGw2JkTEPy8EmRLWdfsOLrIWaYvpaEnbwtLmKaJ9jhCqxBP1HLM7
/fFGB3ceUpsA68RPOfqJGUFZ3SWl/DI6+L5jJNc4pyGV0Olf8txkUV86sAHpvQDR
HKdjuK0Q0JM2qhxJtE7nofXFOTgONCn5rSmk1/1Xh/oex8I0ESykLUzYDgxN97vX
IdP9ExaGfEmGAE8AJF4mDp0mDmq8n0WwDdax0C/X/H7whBzDArl0WHWdNms/1F5R
ljrmSKP9HIIvDvudetvPIPIGq0In2VDmQ1fWo47SArMGFJnxkX1BCqin3TYUoIp0
YcY8mbDb6OpJdoPdtvW1GGx+5qra7fx7TqbqQ+s+0WLutqofoLFeqHh06RDAaCgA
OjTfHfyVpDWXQycgL30QONeMkEwr090qqN3KzOSTemb1AVvEQHDDtAeLp+gitdZ2
11SMf9Hg2XNz+fRg7B+IAGg/IvgqOAaKqpwbAo1QQkxG+rAszoCqpJxZk+dXB0EV
WdF4b6X8AU4KtVmi91+3mohtfEb28Gl3T6pIN14bVvRXiVh6LpxduNJl86q1xFwb
cI+YJFNu1o9bU2oCrxETljHCwaxu/vwH1yk0dWsmZEXfajk6H/JsX4WOpxyf1pl6
iJWOJEFs1ifDt4GjJjFdTMIsS9pX7NrUOYDl9pKNfhtt6uKEQzNleVgdOd+iLJwY
DDxhvEmnFCNVhNdp4Oo6G4SlRJm3Q6ToJAuf0WdNpk0QOWrn2UdIzWSwG0irrq/h
zKbnggWdCO8GaXD9S1U8UlV1UpHTS3NZaWHc5P2s+ywmpml+3r3Ux3vUpD3pVRp/
pVkyLFFotUnT0XiaugsoXNLHKE1VBgcXxVvn2J5pl79mveBZ3fCU0EaWazMkCz1+
0RdvAGglM6v5pRyq2rroC+oMmYayYqBEK1WlJ1WPOzyiAupGf5BUMarrsXYhu81g
KMQ1R9swgCY2zgcO4gJfFQ1Fl2PeAxKBcCUPJ988YCFrGVJ3NPKo9lhnEa5MOTjy
w8TiyTaAwdf8WD8tiqsYew1s8iPu+l46elQ2Esa/y0ae+7py8g1K+HslavcurHf5
5U4OFDggTyhFZOKCihbNf83Kobp1UDqkFOKZn4AOwFSJ6AP9q8hxFR3hvsIypa9x
MUG10/ltjDS7nLDzt1AWc6zdOn4bSRdkESBezBvD6Vvx6EfXSZRUsKRCsESnADbN
3uRUcbaC87JYOfBSCBNaFpDvO60P1zlZuguGLek0/PLF8ys7Fx2PQpRl/MBlq9ee
ozXLxvk1qsT9pkrVvKlZF+bUy/kdr4MlmJNXhU99oFhPpnYbS7m0o+O2smJ8PEmD
bJhLk/IwfWO6gIjFEO0kQKBvXTFwCxga6d5ri4cQvZRvMHI1i5nveBD9128QYZZH
WnrBG7JQebpmDWjerIsgDD3qhmIxeZ2qITjdYDfEn/mVOoEYuh3UZkSDhuQ+kcc9
eB4Jv3n/V0XjGzN3G8ypmswREmgHTVb0FSqe8cnjLe/9GhTDGbA06e6T/7STZeN1
dLcpHAINOLjnudRYoAYXyeTZPIqT2vS5jxcyLc8pkE3RSe02eER3AbndzKgMJZ69
9Nn6ltXGtMz3ExGARU6x9nSqKDnUwe7J8Y1NIgnUPcReLHKzz9q2Rw08nK1Je7Q0
1YwvlEdt2mqgx0ObhTN+jW2WzYkNWLMQQ3zHN12TM89cl1wscp45wArmJvgxZbYm
6dbYLQmS7jsejIY227CFWFAMFzPxLV69VBYLfB6iHMuBNxQiDa58cSpM2ampduft
JR2DZzu+zs3X3paEuC4sEH7fFS2iyvXGHjrfMHkgtJj9CJeZOwZcBy+2qIuG977+
DQbW89uUqfERpAnf+i53jUVUAM9UhRa4VIrivleU7U/x2tGa7ThtIuLoE/NLjFOa
hR+SnPyT02/CYLJqJsuUfsLk4IfW2d7JQJaE6+eBg93KwLcZCWOpQCvw60V9qsMS
/5KkRlCcEq98JgFNCclRAJ+pKtyKpETpDI+ETiNMjLAkzjkW8SIR90n9kaYHEfaA
7YVIJB4kyUQWWgqOXeySUMCFdCjAWAQLsVB+no8Dvxcg3Kf8nwO44jsfBHRO0vMl
85TikIORpVtsNkSUz87StUmmhbsi9ckn7VBCaVjBqrx+yJ0sESSFIib8b4/uuuWT
nWNWx+Q6mOanWQxfCif7LKrKvJyOAb1Sdl1PIjmINYYSdgTekQIJuFE6wuQGvSwa
lLRO/qJ/Kyp42rTCr14wpfM3EVRIA+uvlMfm04QFXqq2o5QrmvWU0MlG8mT/DH/0
r7Yh13tL8YPYxfXemORtps/rwgjG0Z/nhtcLCwPp1IquKs75zeVz6P69FvZpHG/G
mKDfHatqeI1uqg6rCzw0HX3Kq+HqCqcOv/zIOpW/mjERAOcTDu38TAenNCxFeHwl
Ei+eDZcFjjSNGgRAlw+t37a8nXcJL0iQeH/YQlGwLpHr1bU+Fpv6xgkL8Hmo9gLP
frTha5KBorUgU2GUq8Tr1WJgTYHgr5CyK66lvhp9F29UmRQo5ZjWQuzSgSYsGMsK
6KRDwePfcANBWtYEgLl5sV6UtUv774pKskl+dzeh6W2xYAgaa4HhvWfLZwdz1ICl
yMVx1IyY4xF6AuUbTVkcEg1OsJaf4mPS8X+R41/uGqUfJPzKglOISBMKyxqh2ZtJ
2M68yLSEfovu4p/wGpLR0D971/NrU5tqc9L8q5JNgpm5UNQfM/Nw3rCjTUO71scj
782n6sxzTs6uw9zmqNketNyMbAFrVkzBrulgcQIrqil0oWTHmj4PQmvKt0lxUueK
UvUEAA669qKobgJH1dA6bSIf4+68bTQCZP43zGZwk6sePVgGu/QVbtlroKgMyDam
+BY7E/7To7BvjtpQ3obHdJeCHRecMaldoP2XVpt3o35fIyDuJt5eKl9kNnUf4UoG
ZG6mMEdadVGfgJKV0gdi81vD1VRvnpsjOOm6/nKolAzkCWqle84aFZ7eWNZOT0gc
fNVRbBt1RNwmpyCTyx5ecb4yH1/iIibzsO7CnA2uhXe3WKrrKezFaBf8YgZ2hG2t
7FOdn08OEKxsX7KmKDEsromZ+oQg6QDlD/abphRHQmI0qYdPZ/OLYjTwaQk3T00W
R+xo3czfqTQ6oms9DnKQfCUByy27/OfVgiOHIhkX7zD8hi8ybYVw6Eqsc4Sp0Cox
g7qJd1G58JKeQBPOAw0ARCBaISX++ARq180hoy4RIXfpG/kZKpXUScQSLc4HKXUp
RCFdUAg51flFonuRzILguNoj420tC+bo4ow/WvyjyXxeAsCYRUTyLyl6OJ8Km4PD
x15kJ3jups5k0EddehQY56VzmFNGzMnsZP3jbd5cu3UpE+7n8kKcSGLyAL+c6qIw
YS8bc0Ag6HN+aUr39ddYppcTw2HJFWPsp8upVQ4lPe3zPhaTyBlOVxuJpNK8jrYV
8eFkifmjd11KngTupb7uzU3RumpWuYs8AwH4TKm4Znrk27MqeFWWRF0ESmdVkgY7
3W7Ye0YF8IWqCnSPNHoiiVqIrz3RhUQCR8Sw18gnHN4QoVv1NPnDau5TVmoLHxoQ
SRp8ALUo+jd3n42Uo/TC92FoGLOOKv32PoUV8l7eFQOoHatqrKRZ0zK2b1MlZ65r
gzIVM77/Ilkm0CyrKcIx9TESBT5bEpyktPbGuXRnSdwJHRQQmI+Lq5jKriLz+b9L
0ZqQrlk56ZjJqja2rAHY3qdV52VsMhL0ryZRydZ6apBuBM7XYfW8VxW2mVA0cKwf
q4t4CAMVeJ0qdZv0+AQFW5SWxcvTrED5lN2Nl2QbPgFaheLxWZXxp/LZyBqAoR8W
Ch5zZWlndzr9hQNIohfj/Di2Y8OBQnrcqqaPAXqBwUQxUrhTmQXAg5ikYrJ4uSa4
7/RKzwUerotwklNjezYrAPHagFAZ97/6TdtI0ajFfymkQDP6dZh05YvjzjQaYzkA
Aj9nKpdbNebdCblK/V6aIezdFoWNEu9cFI3HRkYAngj0wudQhriup8IiSihm8RQj
A1gGjoeLV+txlON7iXChq32jDVNXkK5vGLjxVnzytGFejhj1z9weT4Wt6f/FX+Cv
sVsR0przt0b5a3ecatoSDiEDKQlDtLnajX+qxyqYQIW4NrS2w4GZoF3CIKNzL7VY
F/VmDPP/7/uELQQ6j87GG0ccRtn1B+oQ9zvDmvR9V0YVFmI+mJMpcrHDJMtPvIR+
+27/rfOY3esFxnnMGdEdQ1LGab1LU9OeMsI4RF6OVRvq1A1g0fI43x1+LTUaJLIt
nMHKmPMQKWnm0SMCUMyg1IEPuDKH+7xut2mmSF2QYv7qW9qMVaV+J1HAd8t4QgI9
GGRKwJZf8BWBKlkBoYTWUh6fuBAfhQVovlGCFQ7Jy1I28vFWiCZoLujtjvZRfr06
c9w24CdReyunvXOH4o40jkYIii48hxIT8dcSK9O4pgAyW+ad0m+PMVpfSArZTnAq
yUvH5JJTQhNsOhJgUFM3D4VNOpvkWGY35a3uU/qNVDgv3SgTKeTaAAhrNKFFEIyi
T+N8AT6wClEzQhDoGraRYKnyZVKqDhpCdn9Xvz+k/BfX+6VypzFibwdywbvVoySb
TP6yEln4DTQPKu/nXniTxTMKxjJOv83Efr2xGpbIKUrtDfwKCiq2xflYaS7yPArV
qj4IUzdrSLp87zdlUAWGeClUkJ3rX3Ka9VKCaakr62uSTLfl1Ui9n2Pb/nxZiM9s
DjYcHGwmaxk6ERigeQ9NgIbZbJDwtrCqiptsQqIl3bHJoEolsQb65fsbl6HTgTDU
avfDxXeJpF5PcjfcY864VMexkASapCOMCQlp9EiJ7lOfZH0o7eWHaOu0yf5QtOJj
SwHLNlGr5EkTYvkJeJ4v4gPp5W9S8A0Jts1fAun1KYH1uj/56QBKzblt6IHV70od
6sPp8CxzpjZwyYPN0fOHLDdGLvXu44+k79EHua1FPFbIZtfd17atmgnOUhXZacai
Fp/t6Gj1dCml+alAHopjT+eZ3gCFCWnJxxLVRuiEyx05wZiJxi/PEWVZd5T9hPbd
rsTlwqp3Jhboo0Y9AfC5rt8/Cot1NliMiVUGfKLvDnWIafjC1D72Y2YEbGB6WFXt
8FIQfNLuWc6nR/REOmn68ujIRpYIifWGS2j2MMLXnq+FPaPDMKqYkkVW2i4YylkV
FbMF1KhuGNbslA1AIt8fbNMe0gCxbt+Q1CYZMOWsEECR0L55RZpV6LzaTZBq2SAR
/iM+YNON3OmurCt1IS6HHFvtOduCK1wTdqKhBQlHFZolKwm4gBnptzf+QM0dCwRQ
ELDHcKRRhXaLKiSUjG4sOn498l7LoFJHB3H6R3bFOwb3Q9IDJwNRbYo2/BohnC8y
R75/6Jg2yk7f15e2Drhd1tCUHk1Bt4qMJV35WwiFXmXpn59L+4Vg949X2dP+MwDB
BRdkmWubvVgVrQ73PYrYkvOpw/ubTl5QA/XkUSW3Bg0DrfjVjgdn28z6PRy1L1mq
wqIXXPSaEza+6dU17Cf8MuNKf+2RjGN4fY/VUOuEHrv0JKmeUAVbtlHMkufayPcx
nQ5VSoxb7XyJ9ZjM57A8U+qDVY3ychatzomoJsqzvTuLxyAWiEGb+GJAsw8gX2bQ
7ASTJwi3PNEpXsN0wVnz05spKYqPhZLWMrhaO1y6SMJKPwPic37voEseyx9RSEW/
di+rFx1v5qK1NX/Y4tzy4/4ZSffwIeukA5pTFrVDu6rN8T2O/4LFtVrE5BUm858P
U9ZlVvFScf9lohc6rg2i/2fCZUiFdK8yBeLyaIXwJ2P0adfUYXzfO+j5/Akgki5C
LwB+gtIoe3iMDKgnO3OoCfxsbxC54Lgtfg3ZWmOLQ+Pjz5aHzZcu8NM94u+UXmNi
aeMrquhs1IjbI8/wnogbrnDwGqJNNgIYsGbZ5xxtOsPxMq14icz68KReuwy/H/fl
oWuqZDN4epaQORXQQVaI21KuEX6Q8yu2Jwu2LGujXn9RHLbNichXHmesvkHiTEtw
mAbSQrrpxXdrKrhf6XMRTP9/HNhjxMNTsoIx5tgV8F7JGxQdF/28bIsi2YDQJqDz
v5FGIxBTGOQh7/QpC1/aa5jXir+FiBEp2Svj6h6VHS+aawASxuMNm9oVg1Pj7N7G
gfQ3/z/BshzLoEqzyEhLgORAx5OTr39ezDccS+DEL5r4Wr1TARsKKZYkpmbogtt3
zVSNKL2N4nOR5Rv8hwZ92YWKiIKUSJPx1jvTYThAZdxqXG+Mg72sMRigjT2ECYb3
zMqvEqpF3AabBjl/IuMk43RD1QzepdsKIwflr0jrvEnOsPlbDI6aeORGdfN811NJ
Meir7QjaPWyVGWqi9Hef5ZT4XNge+pK4EVdhBOQrVNhSqiuTAvfJK9CV5B1hdOzu
VabyWpAm2O11DdpU3G8Kw8XU/jeVr9LUDSZsRWSjd57s6wV1MsBjMM/oDNrxzfbz
euAgAexQ20lFZENozwlpEiez3yAdDY5lcKtjqoSbl2I5WNLdEaPQJ4kUm+VjAgoV
elz7ean2GPc3meRlO4z2Z0ZvRGmUlqqNuREZHI3YwEgWPOKyob9Ci/YOIK2doqXk
NL36M7g7njOF/YrCvadRWyXKoQT6U/UTZemtPXwA2OXXzVR19Vuw1Rne26oqAx3g
/ClhaWoG3pylOf8wCP670aOI+RGge3RW3GSls59JQ4PYlqhojspK60g+xnJ94/1Y
ljHs32R3TX4kcZWcfesLCsCCoYEcp0OP/CiGEeEiDzwdMOpIw4tdriY8u/NUboZ4
1ScqoabMd2Td5GgZ9nzRus3gIpNArcX0KW422YSguIrS8iSRtI2gJdR1GwYrhdz4
1UPTNjPBPghgiHY40Rt1l5zNZ3yJaFUShbSZ/MeddTJsu976lvV/5CcCUiaIJNCo
qXsr9cmAdm5AcQz5ur0rWIPzx4WjiJx5orp3Vre0jqcZa6u3jL/PBpiVd+Wvvmou
jO1L4hCVdYowJ5qyCTzwBzn1c/O2tvMUFmzSkbIgYzxdEDXvgfTdUUXWB7h4Y9Sp
wxJqk7P3XhXDjtnImrFO4JG1X3fzoVuI/EwmQWO0lYIZTPUH2yI3HmjLjtnT5Wyg
gWsAZgj7QR6JGc4z4f7GZ08SqvkFmPRShXDfXtF9vYNPZNqlqj3Cr9uyUri/c3Sp
fqntt8gMep4ntX+tPd/CRzFZtvZTNN1PG1NPQ42YuQTXKvuwycGor+B/MF6NRI7z
o5fOIWta9MWxlZkd5oGbnWab0L7LBdncM438TUC79e554AERAKaCRngcXhPsZtBS
d81T+peClgRV3mDfqVTiGPenpF8mDgg1+7M35mK17rHMqe184LDIBunK/bkgavnz
K8LU1/ATzVnTIRTS8+hKFl46/ve0gCQnvhJiVPiIW+GR6016By6C4w5tEF7HvtyI
iU5GxUdhUlWm2exIo6gwBZdIXDjz5JmlE3mX+sn/QZDHBeQJdVoVlxZr7MTQLf8w
IF+VHCW+/JUOf6Dm16DsYXrJSjlPonm1BOs3NKy3jm4Z004Xd0SxmXOHH9lq/neu
pUcTgSF3CB6XireYnTJVSDrFsBg6gvnPqiKWhmj3dHB1ND42mN31hstY1ooUGDzt
moJ4pTDF+ikBMn2UQtXtoA+54Krv1K8nF7o2ctIReQ3NAEFMtb7/f/j9eCpAZlas
rKZHxIY3+l0EbXijvjsFIGmlglEI5tbvJ5Jo2oJM1l8n7AUy1Kdl1XUIyZXFLXj/
Q2aU+hQStnwNpr/BN8R7y5G92H0LjXO1advjvGPVTAqhyyaYenzH5kFgT/AeZyds
YjrTP3/+5kCEVyXCsUen5YWUFrerivrjAeSA5XtWyddFIkz5PzxgxBw6GjCeLD2R
lm+6iWVWHE3jjOZUu2PzvGvTY/1aWvX+UtVYqydPiNV33e3Q8tuiTdhB9C0dmPrn
7io1+oJGYOL9EXkvwloxaWIQcsVbakJm2+djhkNFG8n4O0wkDBNit1DoCXZjZm1H
r9EhqB6UjVHJyHz7XnPGwztXwoZsZ1tSN6AC7vdDGdAgg9DJDJ1lqBOlZRrEuIqg
xhbkKAjqVHodat0HLyltWjQ29bWdb9UqkzHsYkZVtIWNQHPmOlC3j90T7DggUmOs
HjS1+h8fSanXbrGxSKTFyXG9vZHE7WNDMvynB9tZEMoiq1cq0LNritkNQjvzPORN
wRqGt17DvsMTbK/EMrdNt+WAzFy6zNmJr7LMniWYfgPUTJyFLe+z5MDmoo1RnThD
BlRpJLfP3i3VVhmJ10dW8G4f5JUq9Tj3KaVVHu3sGGftZqRMbqcBeO3FUWzSwTrm
rF/QTnNOrWYd9NEmnS9GQ2udjXcZ5nGJF/5RUwNGFotiwmZWemrvxWP0wLn7e1+o
byUaAiGtXaUfJ564BNpxxEBHDxUQqx6S5/hH5BExaY5rE+BVQiezeUrxrFFQkh6K
hOxyNNJh1ZlOxcLZVauSiHqHGIrcI9TaNODAXEGtQPaYPulRHGeNJM3xV/SXua9X
MVtzpZo3N6zw+jbL82mSW3PmZE2hILQcJN6AC699GD+vLLgykksFipJxIjFnt9gO
BGedZkmvq37jea7EjuoaHs70FJlHzo02/04lW1JLFJSCBe0Yr5QZz9gp1asGifCp
wWjLXACFbCCOifkmgFf5R6TWfwuChNaozo2WrXbxgv2VLuZrX6JelOnakRZ+Wwxw
bMH3T/3kRal6mAImechM3cERdr9l7f69VqSWMkOKGMfAx4sDIlcKTJEyB6SKOOUU
yLVXWfb/6nIvl/h6Uw0aNXlJFhe0Do8L6fanIpKdAh/F0EI44ALyo3bQ/QTX0H6N
eazkSxfPHCPS1BSevPF4MHX4E3j8KMhMZoQBwv9GSBJX7F5mHNA777b0YCPedvss
7L/MHmnrzbyaF7b96L5mUGnzM+jOnHYck80/IrHV9pbZWblPl1aufR6h3zzP6L6j
Eh22eQ4X1qQakIXEPraUn1y4lWh/ziZw9mTTDPJichCXdF5kh/ndrfk4KtN/4gqq
WUSJ273roVTZD6UmLM50/mOq+0ROC1RYZ9IUbD+hXppxLv3pnw0ogO9/fJGyajYp
DrHzO2Me1EkU7D9W/SeeR49Acw7RIjxXAVPCxPAdAIYXRiNcmhrQQywW85fk6pa8
/wk7lRfVvuQ6DrDGOXCDUCrx5JBIfGoqCkILKPcXchK1MKiZ5bwGngQ7lb3milQp
nmsdz0dfukldcw/qd3fY/tR8c7Udnwr+KrWq565qiWLkX0OT03OJlaeOCRy1fRe7
TEtvmj+WL2leq+Uv1fQrpCZ7RXUn0EQWlq2WifyKm4Rrm593nfK4clyeJ49gKmII
ko0drRBHJkBuf9J2B9EBNNhx7BssqA9Zoy1d4bH4RxrYzkZxMvgwDnLK8XLpJVAK
4Iz9BXJTx2q7otnHdGaV/vGCxiCN8hK/uPmUe+6fKCeRRslGpL1mUZU98KBtIV4G
RBNmnhxGL6Xa5H5PSJrYQYRAsW+uFxXVELNkQbcofDkxsq4PHlK5OKm2rB7dLS5p
JJ1iGUCkGEOK/F4O/Ouv5yEGUhy4LeFMhP+Un57QUDqDnY2jodx0Qr98oZ9030Nw
II0IgyVwavp5Ht4kGuYOUJ5Pt2V4S6X4A7NqnOXjzwGtshbdbW8Kjz36bwZ3UYre
4cNy3Np6SLx3KvlIAiuDQUc0fw7QxdV1ygCYnhgpbyn+5U4H+1kPevbR214+Qwoh
GGjWAHk/w8wIfofNzp+Kub6TNCc+kHmxYLFypqIIIddtPf5JrFlGKAihal7ANf8W
K/5TYSalrgaJSWE+eWtiVBG4vdMc5stHheaZQkYT/OAcaVWV/g9Jknlv/Skg9bNt
w/UxIRG48IL1HosRB+5nib8+D47ufJhCZHhBXp/suQVW1wdisqKllbehZAaT/HhJ
gvLAGUdPDM7BgY5Dc76HCXFhxVlYQPAYHMICOs++VrjzVxp9lPU8YCNJSUtIsed8
Lsv6piWAVR58EAhfhJSzFF6kbvrnK4Djv982WIntnR3c7HBqZwOnFw0+aoACslV/
c8LPD3vsjbUUavaYhh0aGMaopEsCBXDBykV9fcCgyBi1J07JoIpjn/ggeAIbGiLq
js4rtorkIILRw6h4Iw/EqbZtvva76tqpwdZYTat+XkWzEVRRjUYCBuYshqd+dfSw
iqJKAwEV8HcbmEcIBZ44/aK9iz/URxI5kH7H8b25QP0KsESPe7lIBpRQSnz1h+jQ
+l+SFZKK6b6WB65vQsxyDRpXDMpOLamTO6iqWSjxNOlGJGkS9r0vdACWHRHzrAe4
WGSRj95gV3vlUNQukPzOzmrTmDGwqg7XHerZq10hhzKnqmFYcPJDjgzpESu2peHm
EKp5nCmj7g0GVT5bQT10mK40ckEuwGb6BYwtN80WTbdUHHyrJwmue0g4GHgdeceu
TZn1HMUyJyDdxVCNRZp7OKkb6bTFjuxhLJRa6YU4fWdC6DbhkXCGRSHoWz0oH9wS
ng7elWo/AYYukeKNS6kO0mzlxWrLk0qBR42vlSk8ERYSqanlyno5zOCRnGemeYv2
09g+356JAtn9GUuzdQE0ud6OyTERiE2/8eqRghCCYe6fVpeVgXQ1KF3PVMaC9u3B
u+g5iGrR1edPbGgDxwfKC+xISgNFKySdgiyUtJqcZvTzFNBdKhqfb5VvEdlMDcSE
xTlPRXiNkxtpvvx5p0R7T8Zq308vzNQAj8q3RMvBA7CWyuxPwUzSw25We/ZV2l52
TSqNiFma+IKhps8inC+oDcdfDZWfB0XrHXy/vQuZVqzPZboA9Ln/Snpernc/7B8d
uC2BctGKdxzVAkz5aZCpo/Zxx/zCK8iYq4jNZI+iJb3bTc0BZ3BdntYM1M/nmKx+
+iaaAFq/4zzLrVBzmmoqWiTUTC5v5nxpRBc9AsgkP3Xw1aPqt0Lw+Kvb/eJdMgSK
3Q2tlYqdDahC0x1hzDkhblelXyPYPT08eSXbLSg67eoWVNLJXahaKw4lOrs4IAro
XmA2dIlen01ekhP7H+qoRwcj6IZ3Q+RvOYPfrhUcoorDWYfDsbEn5DlosSbwrEoB
79Zzgp8rQiBu9xskGyLDbxH17UjLCCaeuchWIeBi9SlIKwc1pKOBtl/LzJTqSNz5
RjXuF0ccNiIpVuPxYyy4JR/FxZUFxwZiGBp1Ly6koVc1w4IrKmZzd3797UF+eWhX
w5rX1kjqWMe5lxlotjY+dzzflh5h66DqcghKGvGrj+Yr/1v+tz+ladzpKDkUuOFh
9dR3AH6FxqpWyMOYYSobabTM8w3bK9lfBKLtpRWwHwvWr01YOh6owmzc2+S9C2or
NHjjhMQ9ZoGvjBU2BRbtaYfneqJDnIrED5Om4ywKPm1YPVhb64EjAj0Kxmq4I4pr
on9phQdpsxA8IISA/y+GMW7IiKGWVNYqwIEnfeHlWXflwS3CcBEITRBqCPEmYb88
HvFoDG2MrFBp/gKSp2nsf6Yj6TN0pfLwrbV3I7KQIQVuQn64Y6ZpasjOzFnlGo+O
2LMu/R4FlqtSGAw7W11Jz03qB8wQ59bKq6ajMHi3LnZYeOsakbSxrL4XllgBohir
93LISUNHLIWPBLYBlQEZ2gTbT2kPNm2I7yc00AA7thPHjnoXMWNfr4hAYSlAOkX5
5kxXvOqO/fzwYhC3urh6crM4XHMveOoUd/s5lYqldVgXdlZoN+u5/w6ekonoONT/
j6EZuGb2DlIeu/FkFS6QSfH7iVDmkfaYEgwSsEAER02yhmVLfdIOmFGRSb+HVEpv
PiPNxeYOxa56BM6xtHkgKn37llhr1zcCpx4Rjuf9S+5hM9n9MscLjcDn1WKwnLJh
0YH4a8msL85ZNCJiBpKwifUc/Hx+lT26LgtT9q8l4UlB2wU5YcIyue3sRVWynh1T
qnuIe5qih0yN4GDUnNYFVKvRAe9bdq7AJMcj6Zd6Ch4szyL44V9FXVw1/hfbc94r
erFzTPYQ0z7NHMWi2AKnuE1qG2K0L/pMQT7aUNg+Fxt5UJCKpQGenLlRHcGC99fc
dZUj9o49TL+W5oyCquVic8lm44cWVF/ML1KVK570SgNV/UKaIbv15quC92HdQZvy
6YNP9GERBkb2E+ZQ1U1G9gZVdKRevtQFGy5mGbrNBJATx7c1V+OOyoTzVPa1jtPq
V7O6jsTBtPZqejZ1oJaLjdZb8Kf3GnLlZ4je4Y9r2TU2katC+j8RgELl60Z9X7QI
iIsuX/Rp5Q2dN3agksyPJrMfVOgdhdOAZdFjUMLmEwLvg/aryom+kwvWp1Dm27es
OPr5gedPX8XICQ25ARDdPcYy8dGxW5eLLehFaAsb6zg0RDH35JOytr0EPs2YOEuu
4Ik0Jnhp1ZRvX/R2Fw7ACSzaCPwQvqos1chAAjkjUXW306J06uVRBl/RuUDYI++b
ArbZkQa32nRcx5W39J6d2Cv77O5lmctrqyQsZ+dexSKNn5VCeOGbXHZr52IXhP8h
8rrCkdVTKszLo7lZ+dISWjI4+4MC2yJ+9vVmYkddA/PTluMvvs30XJJZ9VRIG8BW
qDfr7Z8dEHVR1rO7QRh0f5PIF+3uCNljXDvLLpel3IOBphKmw9/uGHFedkVe6MzW
SUSdqf83XHTX/WnHM0AMdaTybDjLLsMmrEKFXg62dm6xpBl3MKP/uX453ppfU3xT
T58nVv5dMVXy/NypCOyrXBUU5+b3DjaC/gKhYxxSg//IT6dSMWi0Mz0Il0ZaYYdY
qd7upRBzHzwwNSDQlTFXoFl0JzBlSZ3ZPLA3LmavWVeshw/OD06UedfX5LU0np3y
CuJ2Ah7k7+Yak3nDDMhtCNELKhAKNpdv2GyQWkwMC3SlGJN2/lK2NhwErMEovkq1
LxFoYnbcYawIYNChGhtQvJyDAoPnH4lv4x185tbKw8aW3QbqZrcfsqf+dNvOXcG4
/q1B2gLUnzqNZ7J4OiAESouxcVE+MEDzr9ZoeFU8VfeeX1RciEvv+LsxCF1qw29C
Cp8Glq4Sn3uT8a6ASWhoHNkSuf071IMYsiCtKwCBOW5KPDln4fvnqeG+6BPKBeAq
+mXGeCCOX+UpxljiqYcMFCGziYByTznjLVtl7+dsMraTCxsptvsDcK9LuGHocm1D
basAnX1qwwAPC6T9Tbev+zh0V+SeWJ5FxLmm7dcejPkoI2qmml6KVwZXAR0ACUTx
lHERwFKFYUWMkp7qipuBqPjX3eg5BRkbNPTKq3IualPC7DrR3diX8TqXnPEnhuqk
w6rbkmaQ8kceHLhso9BCQdZ6bvHfhs9jDmdiSP1I1ZZMFx/pWUCcIzrKHwmXWXcK
E4zJI1lyzI81F9fKV56XKmvFV5VnQC91OiF3rXI3JSvVjV7wkQg1MYCNwKQJ6Sb9
y5ruZFVGApzdUNnd8QBDh2rDQz7gr/e79bnEoKPwCxVsKQKpyAxx3l63xWCwVgEp
U3gUp7v1cRqw0OPiBQ6WlQxrofpMJ2TdAGv/XVN+L4XOeXTjia2xond5HhnjXHFN
qLwrhKOB/CZmuIG7rc/hDP5Yx/I0ac8pYaCCNQlD5NBbKCvIaiLtkG2yDAL4jRLZ
uy/AevjWlc2uaGtmqQ4Ogp8PATq28hXRyWG5vdc3naxgQyMjxTNHXaLgpBec9wPZ
e44xhGsX2BvlNhbyCc9krqmRi3XX8gr4bXlhwhjE1kYot8XmSL9z42+ZukS8eApN
9ErY4A6g8+fmooM5wN20msqfFPnr+57bHQ5CvZPFgXhn7AY1hLPExfpnm9faSNqZ
XQHR9z192pB0EWVwOqwjNOaj93tscl7sldZmaJ7wNYBX2tgYzJ9Ar1Zy8R0q7CNu
2qgP+MTX+n1fEqFa8IY4AOJqajogJ+iXkL1UkplSFdip4LALuZWzcaYx++SV5drc
8Wx5+KNHbMoyPlU/ERn8NdR3z8W3p78ja2eHFL4J2zR0kSzTHpD04hVAm6Nu0fGq
d0uzS+HA1HYSF7Ezonw8DcyKiSOkSRPlvUYsooboRMImvJPkoWJf+lQ733PjqxIn
OQzpUKfrs7yJ/u+eo6BkQ8Z/Ms2AH3OAjTQakugmlGtK33gZp2JZdeeBdC+JswfX
aFbevWdc13NjLgOjLOC+eqVK+ld5dkmnDDUmbzWPR4gXPfeDN/d10uPGYW/f7wHZ
rmkDq5qTzKG9uM0kTuiOiAW/fqwEHK39kuIG5oZ6VwYI4cnXo29K8EJOLs6CkFcp
KNx7DCrazCfQToIw0plYJ0rQuJJbdvX7q4SCwEf8vrsQHgaueN5nD4IAMc5tt9vi
/WX0BnfoRIOqjVlfEq+WF5KmIJE5M6d5TbWGRb/MoWOPfFIs7Oy/+9SuYydJObrE
+6Vf42q79CQaIjUWpCaTnP+bLT369b1wWse4hmlSdD4a2o4ry34z52eMP+Ld1wnt
FsfVYK0AK6sqdVBTSeeEYV/e1V3E96OOuSLadmMByIYMg0Pap2R9Es4NP+Ot9cmX
z6CnAhUN4y+nfwx6gXC8ccrGH/Sk8Prz2kKsEGaDYFqi5kcyxBhSo67xkGG1sBzJ
LVIZefS/gFdW+OQCg8ny7CeM4F7QKA3rnAwfaP3iN4EUCS9qyoO6RKPl4gtKd+pW
5S2j57gPHn9yWq4dCkQ65Jgvl7iPGIZWH0W2+8oc6carEDHdBtmoYzHUfJ5QDVEa
IfsBIyqXvS3QqFQRZY0paAV9bTrFhcHh26fyVqH/LiodEb0/tYm8iY/YteWmSlkv
Lm8NzGZAcZ81ADqieLxa8Gsp9ZpkALRsFcroxXSu/fCDnF1mPZQ+/SvsuKkAWAWX
M3uZ1SbfaqVU1aqqFZ/JZPItQEDc/csayEObRs+ZMQ8w3BKUw+J0VVDvPP41/jKU
FhwjBmsVsYYB7FOjPPQVo/b2kFDiXvaE7ZbbAAE+wi9JEuj++rSkwgNGFc+i65zC
kjq2WXy3ttHFPreBXZRGfAC+5sHR1T7CEuiPYrcHpJi/ogOP+hL94SCKME37RXH6
r1kJGzxmoRw+BQ2MA/5V2RctKZFMiqBeF/DMrtJkZuSYPqk7sfvWQTNVJOY1E6Op
VA5hbg9ODGAcLfsMUK1GsRRN0CAtdTjCiuaras0AgQOEdl1uGk8yIEFN+CD2rjMs
L+cPkpMxvm6gikWdENMXUPt2FDKj/jVlK5wcVhC+BEUDUERVjYeZsl7lRKY3k4f2
A9sZgMfjzMx5QovoHmZgaQjLgijhWTgJGiUzNeRNq0iy84XbB1/iKHWKsohR+7oK
QLTrZ73DL5FYhNg2Tx6Yu9s2wXLIO8nPy0IfLbRbSRbNWma7v9eOZQX1ykkcpBAU
6j5WlNu7IEyZ3Rcya3xxgHpQAFxtFsi0Yd6B8vJ2GLWkf1jsj+Rp3GvzOr1hSEcc
b7wtEQpTYtVBirI/zofjwdxOTORPK2foPI2B9jhAVW18Brdqy2XGijkE9tY0N+00
kd/EaFzFm2RkwtK4gFH7I+nVbKg7tC4vrXIfDQP40h+JwsyPPVCzGP1XJK8/yRLJ
KKFi8ClVkUW2+TTGgUlUq5a6Z+DVmahqAvjYXBXDbU80PShqvEZ/Ij0I9256OVsl
oeJBafGCFm/sXjB3qgq1LK8SVIdUR79jHcFbc4k2u7C+qvntkYTpPSBuFBtio9Kv
yxPPNXNE9MZfdLVGlWY6gcvhVT31G714gbGB0DKpoAZM1NSVGRjSJa+TaFWZ+KLu
SHl84q4Fp5g1EKbQGc44zdoTMGHWDgXQF8YWFzA4Ocs9LRrp9sqhGpTtimKxXcgh
fpVSSso3DXEFW7wqBk3HdXFlNcRDpCvBF22TvJLlgt0BoS5rmeTSyIOnAQUgGfGC
RZiTOSE0G3uez2ZDJir8EHgWaaqirYPJecyDzZE9/GueoNIzxGHsYeOLhZmHBntl
zDMSUU1M+H74876dyCHO8Y/PNRdZLJpvu91Kb7cuklJxUUx9ZsqFdMwZaD7KyP+n
0pDHzVr6TqV2+tg9YtvMTAtemLyBljHc05r41TrtotmFFTXo6cK9gb0oUp+78Cwt
LJqkf8oGzUrIf0Ql8jc7N7rf9cAk0eapfpqm1/Z2toLOoZRv2NtlXXeK717oMoT6
7BgPx4CmPQc6yevbKqA0xtqePzFGLdFid82LQILjcpkco3Ml6T/RjX5ljUcd0503
hloZybnbRSD95hsda7UxiZnpcf92R9cf5KmGq6M4MRqceXkB1XdrksMXW3VDaVfL
FmpjCYL+gqAzfqIitzvISVdr06egueViddRPv4DM4ULKULrA8YEDJrEkE9gW1I1B
tgGKdhIteV8cTwG8jQukaNz5dHr1MzKrCEMWmkGxThCdZkXffVnCL0cKSOE6fqxD
QRrwvOHoEoItC0CqlAxDiZvtODgwnhe7RGgdqlvnED6Awd5Q96rp3iKC3qslTwnN
bqmT+HjEEkzbhbKuigRyZDcFIeambuER1sn7HHLyf7vDlJya4C8e2IWKFiSynQ3/
SghspkqTCgD/Um60rNgXVWETwStjM8f377mF5A/mzuxMfEFVtC4pRO9M6looc1h6
k/LKkMxhI/bb6iedkaF/pv7cUaWZaw/Pg6mZbQs+maf+5ATMu/nRugSOeuCjVuwB
W+OPBkt9MnamI3S9cxAMb3g1H8MNNvuAFiN+d39XXIyTlcDi/5dLc8Oq57QqmEfv
hhHyuzsaKGVgowF9RMw3k2BVKRduSsKx1dnaIj2FjeoGnOtK7iVyPudLASU7WxJn
Ufv5RaaNuJV6boNITvguxBaYbfCq+qGsj9w+fxOIXcNT100KUcoZDBhnRTVie7fh
Qke/YclxhQNF2P9oaBUDnYtIB1P9mt30cabO0aHJFGkqp+YscFpZB7qLU/7m3ExO
VweMc2uM15ed3vDMgiXX7TWvmK2WYNtGmrPRFnm4xTfLM29NgDNZW7Qynzj59KRB
I2Dnl9a5fzUhM2p72FfOuUbO04JM0vgIba85lcALhxt6/9B46g+mBJoCkpmqEazD
EDUSlFHP/j3NEEWjfJ3tAHOrhmTPU+suW8VA37Liw9N09mSQ7E9jptMoSwM4khaf
nH4UeJ0k6ywA90jgyKpqOIoz1yH0n92bMxsQrcew2z/sfpI48zah3gqQytRC0oA0
oGJmwabRmhprbD3ELV1s/j2nsIt316ktqnF8vU6ZnrWCR/MnU1UTPwzCwl4+87ua
OHvbpenfjcz2Rd/zKERnLJpWMAmQ/d/lijJG6f4vqfh7a+47s9zPYsqF79x6WBxM
SQVjAdXPVoogvDLLMDGJsOIe3uhGPOf7NdGp1iDsULruh9mBHPVXAUg9aTO+j9ch
ENW0F1ZO6LDuKqXAuLeqTnfo7z5pd/v7sTErqIM0XIDPX+bGcjFdyNKTJ1rKwqJw
V/OpFDwPEYZLA9URk58vGBj96rVWaJBPuCmLoleOQSyMXOWw5uUx+uYHUwZaY84+
2WMoZUBwnor8qPcBZQna1c5whZGKr25N8/7muM6YkceXlje7ikPJqkzeH4Rd7coU
dSRKjAxeHanAHCKA4fMOMfGGOyhIt26WJoKIyEXJJ5J0KPgMlHL27JXjVpGNQ0wj
QT/mv5cOh3lGx9RLcU0ij6n0VlUt/Za+uxOHO5V7Iwe8prWXpxPf2EK6okwRrda4
vMXaevka4lgmITFHoXyPoRa7EP4pi+OBEIySTEBYLmAu3100+B2uJxzRyg1VYXEl
1CvSzk9v8aJJOG6wTyup/o25c/flXDNipxsmR+mX/5JMhCEmEwZRbLypWxE4jWEi
b17GfON80iI78mZHjEWFhkvo0IKyMNb8HWDQJVy8m/ZJYeVQ08mLIFe+AhCZG7NB
GI3ZL/v9qPJy1yi4cKdrMN75KIQuvd5DoCXsbnvoSMYq1lu9V6osa+WcICwRvinr
94IqzPmDZKYRimGnmHDyhyzZ+urJKcQmaeVzkT6YSwR9EyYhKkbElbU8ZQGKDPw3
18WHXNVz8PdgzdcwTVK7AcG99uvCvdlXmokGS7KWHdQwm+OZOaXv74MEMZpSGGYy
EIoql8XzWr4DaXGhYG7590rsO3X1dFKsIMXPtrmlQh/nAuOi2nkbxWtPIT1yMv2Q
cemQbLFua6Btp/Nv3CBd1mWhub7pYZMJ8e+mOt3X9yGsXbNbE94oHTx5nlX7b4iD
zPOleS4I65LLmpbDZhCX/Oa22KgstuFlevFsUamT2vnR2hElUcaSjI93Go7AnMhX
aRrDUyv7oAfwTfurjldZ7MbFYtoVeQ2GDdUNYiqruCGGUefRPGZp1WX93yElKmSr
olqsWdcGVfafw/aj/52WYl7Qeb0zY+sHBxT5MGpRRczykPOV4YOMGBueDDSncNBa
Q3FWjguVOlzag/2o9keXfzooUiS5C2hPxkCtG8wV20sN548MQxPVgt7Zh2LcRsFm
+wcWo5TfoGQUUPkEpZYZblj7o1qvVkLpK5ISR21TpZGRJc8sGYTtq9ZT2FIw0pWe
bg1GyvPZqpS6bWZA93rwDNpCxM3jaARq8xqVKTzmjL3Zoy+Pu80VRvRO9tzkkWeF
IDSHd/cohknEoQu43TcXqquxjYMNgNgWhJJygzAsA1Ol+MbtsfO8rWlq9qOAl5Cz
63wyHx2Y/fJT0Q7gXw5bxrrB4JQAdoU8GAGZ7fLme+5tgCIqT0tZQVa2eHQzyvYy
2l14NasrsGiq/KZjZ+/mUTpXttJu6wGB+Hc0+ZfYFwHrOh1qpTOOxG6fWzKxIKyu
ffF4zd7vdeJ72+BAa7lkCLTW25+erphQnBMq7QlPTGnYIrFsjYZ9DcEZvx2KNuuT
2KLf+grbrvxgqaPGnxP44/cTW50OOlGn4EDbhxoCviWiNo17dt1sDiM7f7QIK+lV
b45B/1CqXGTIECKVoOZG7ZQCJB040jo/5QkdLq8pBOwQCVf0dn1pLPqiu9+wtEvx
XuntRbXuQguTKv67FpONoDTQSZUbG7yCnqTWf4XxhRW+rVSvH0JdfDHI4o4L8hc6
lApXeWGy5bQ3UKVHPABY7QuD+yjRJTbEvFDzcvWy6sPcGfXko81YiVoyF80TaN1E
uEondKt64rYFZzZFRUpWd6HuqMWqvTEcszuiinfndkviHMIEP5mWmmg5vGFUfCzu
PNDwomk6ZTr0U3buoAPEFwRbTLnOcBaU4JOw9RnXcGfvpzw+9v6Qibt0kQlW9LWE
FHPF2uTYN5/2+maN43UZRoRWzjr6IBxlJPk0izIb5TXwWLJZxF2p1enOlfe89STE
Iu9IBaRKuJ9MqjqZV+Vzi5JY6SIXd5YZj6ACGy+2BxwIj60DyzRlcgnJoxNAbTtX
u5YXT5/bFdgcPcOIedyxdIt8oT2cKxx5m1SXaJLAHe1HpfDg/ocDUyYAzdOMlomp
7H8G7C6xaJHRjesitgtsd1ejJm6XDBUCuT7NRwL/udlSGR3UGImkasczyPKn7onw
bK4n33oI51SJXtXPYE1DJAm3DFJ0ptqKzIXSKH8uGyPaPxnjs/N+vTXs0on1U+QI
lCuwekGVQ/NjQgoatTyo4VTo9FbeNuLgX4Lu12JkpHkjyERuGGSNvEtHBn3j5yv9
xw+55qJaFqW96k6pKyLxLIim1Pmn4TtUqWn4g33IcQGOFhdNfFEyRTK6E/tb2+ED
qm95kVzWPCKirMCKLv08hLjAlySbFh0gFkuPqab+t4zmisc9ab6oFxfkgkCCsDzl
D+kqxlLvdb9VJPVu75LdEdf/b/7dl3r2NK4uTcWipQzB4aMsBABXBiXtMtRsHhiX
NS5YzCEHhWfw+A/WEZn4+pCl4vZHhewUhkOiVOVzuC45IPzEJZ9qyIUBioYUrBL3
0olG7kHy3ihRqDrAGFpVrTyyuMFvw5B70htwQyTS+G8bnF5cX09Bn/xQBqeyeOF6
bVL2G8wK1y24JNMlacITzNbba62+c1AV15oi92lFtaLl8xfDLGl+iiKdF4sxpT9X
94vL2xx6LB67PGMTY62z4QMzYmuNhiWQWasJTAx6Va2t/Z8iYQbN2YT5n9Fawyqz
E4BqySsGPzrIECkY6Y+sJEKo8NYBdUUhLIkq6kwHlcCsQQ2R0LbnKaKhkBhI7T1/
i9dGwGVpBdx8vEojLvnMSqcn+9ZKhuEBcPfdWNMsla7Hmn0vNppyZxcUWPJQbAmB
G+nFiZujkWWbLzuXcg0kjio+dVpOnB0aPLizdGhCwpfEzWDlaSkG2qpKwY2k13Mv
OOMp7Ebwed7+ddAlrDJoOgcK7aqmbv2zgtpZFCkj5pfVRlbGT7sfK2bDtI6BELsF
P2k7RPQ8gtIWxx8hDUujljQ4/xVBcSbm0+HVHgx8MUjWaSiXW9niV2CyLzYX1t+g
jazC7iP40HGUixjLoPhEvZpvnfWDwvRJWqPYKdSkkbnQ/C0hPFwDH8kKDQ9dPDMc
/U8+KylR42pd6roKAuX11BqrYQrP7K1TVKTPHaWMqLjEUEFEhjnEl8i8PwGyCUrU
VhX9JqusGwaTuNow+Zq8ffTurfGJwRx/hqQoNjnci0c3A5paA95OpyZFc0p1XuCb
ocGI3BgqS4pZQp/SJXdcaj5S8awYJDNE3X+GXIy+2p8iPaMUhVZHnU9bnCT+Zcy+
tbm5oDY7DC6SrKbZYz9R/m9RF5q+AFIOpjsPskBqXsyqmNCcGEewZMBPjZ0mxEz/
mJNfAcp4Dub9+C0zJr1gbHYrZrf8oz5A5Lm6Bn7VWPF7O7Q5TVvth7Wg9N1jUHDT
bsBO50gXZMSF6w2x1giSd3o1GDo1YsxmAtYi6OLHFlM9O0XL42zjmM8KUoggc8xu
Bi1APF8CDdLaAIgploBpyk/Hk9lD6G+unn3dg2Z5k0cW231OzsCXutBV83rtJCde
g+RJkzywFGiy7Cnmr6VMDEMDmr907DFCMXrD3RgkxIbeHuS4GjubKEp5YPRttd+M
ayhozUpZTdm8/0oNi+jKoKY7YoHP6qS6XUuvBj5d8P7s8ASUg4xoONImx+PEsrbr
jF03n7Zfe+OdPALulXer9QU9sVKlNNORJIguZ7HNPRI+KtP8VKRwbQNjrUaOUUXY
WR2jRQ5ZArBi3VGpr1RTQTe5TzQ7GM/XHNh47aT1WlbYYiAzhiJbS2w0QgxKt+gN
p4iWS8R5HX8Q4VoduMpU/av05gZKv1a8yBRIUIPCPCsz07QBzQq9M9th2nw2N0HC
FNS/nSFTh4Y+/69pNNdiYtrcJnx6W1IwBwNhrjMg+NpR0i64436qVAqpKIJPzMTt
+9vtj2XHdCfvj+ze3bNB4xxhMH5LhKnBpvn7mR8ikjF39+64m4zDEGxkQJBhr8ZU
LYLyG4BmE8Rqy09s+SQ0HN/vjLLah9ojrpAIKZKnSxbo/nvdRyHQ7qk7XmbBm+4+
LkP/W6N0fljEOONT1f2burVO2tyY/hEwzK+uvjnyNmPF39uor0Q8ALJaQgjntjgN
LqFoxy7MfOc5FqUJpYKey5xRg6ki2iyV2IYlIdu88r91qDuDqP1RKNHnugeR0U1o
NHTDMUFzV+tVniK6OZbzpP8tU5d7UaoArdOkfVNid7otffEjpVv8xp3NFysjlqXo
AAj9eRQDvoxj3trkNnAUvVEN2zib4gkkFw0FZnY3hgsjMa/9aHNggdJJT5H7x9/i
GSL4/UUDbvLBTr1pgBfSa7x3m/AvxzB+7qEkFBDEIbwd2Ipo89wEcNYzOVg3BoFK
4b/bfgJwPZrca4R74zUcOUPdZWnjbEHHetwk0mV3ebixPcHdqTCG6PPUccElAXBJ
KzYvoqpCf3EVEzrm9YxNkK0xyqK10kre5+w7Fw8OKMnu7BgiFQpAlUYZOMLW6pws
RpxBXQlFWLZIMmB/n3XBB1qG4lfaOa4a9xUR4eGz0XkmgvHHgSY0dSXniFRFtnEo
NDeo5Ch9oR4EkOKHB693mnpILH0xftb7dWmHM8fBlhPMgNr+pod4KwDBTIOv9j5o
nyiq9cdFAqsC83CnvAskLFLwijQcaWrDuL4l2/JS0N+8hsNHCl4JTZ1+aPLFqt3W
4rnhwCp3bhXDbYr+G+mSS2K85dApn+mWRSVpNLGIITxLQ1eDvD5VRWGjZGCYZFd7
Rbw4XeKVaR9+6/BXQjXaX9NlbNNY/niliDHhEvSdxY3ymxkbbjWtMgwpiCucVLvA
MiPvuLcGgc+sKKsrboLLrNu0PfaELdT1vKgMXhijgXk95K8i0kKjfoupH3Jk0K5f
7fmDhVbVRrVlWV/Cf2cd5VXGRIJjCVLZiBRwYNImViKjgn45aqk6VdSHNVNb22Jz
w2ZRshRYwymkRDo6WU9/qfbMUWyKLMbA8EuZbdijG2QRL5cGqXsOCy7TKc8c3irj
olF5w8dVpmZQjFwg8j9aU/t1eOlLveY5SpgiV65Ilc4mSpQUAJDSWdL/KDPAZ/d7
+FL3cYNdt5jCUTPEDEysb8WnrwTrBOKEm8jyfc46aHpxjhdnWeXlKkFl058M2Vsj
Z4Dd9RmCVGKLbBCDKE3Bvbn3+NMXv50g8tteBigl19brhOPZEr83t3+HOvCdEdTv
JuFdfcujqJMg9lDOdhoWhh8rn0udXts5wXWvBY0CCivZmSgznpm/KSMW64hr9bGi
Rx0w23F1zN03pI+ov8ccw2mj1VY1E2s5IFNCVK+MhPTPVZJb/gpiTI1K/eOvaZad
u1sfJ7t1S+kustFrjjbbpMorjagJ71VNKJK644NxeJnXId13mB04fAk9wHeX00bg
VtNccwQjqvjyiyoc8QMPXmxz2D5AhBwrLuPFFrSwWrbG1cjwLQKJN0df3HhSGm0r
NMSXEjb+/lBZUztBeM3suj4ay1aJ/Iiavi5kgC6LA9JOPky3v+5gD2+fYrFh1JOc
sOFoNzZK83sjKvnbQ1Yyv6Rb/isJCO86iq0iS48e7v3sV4J/gVj2t+kI6DNE/gQ8
6h2mpHTyr4TPLZnDvAW36Qi/E3qDegvXK/Ga+b2AOmeRqG5AgjKzUfK/VV25aqCl
LA6k9vU7kqPVxLlWWwRu2hHfCNtVSRiTq0NitBx9c6WnDRpTQjSHZQtAMCaMoIFq
2DqQdw2oYzC9+Q6uOfof+ycTQ5UOJO1cs/yEp+H7lo+jQaQP/r0/iIDbqgY5HAYB
yaOwJPwIvaNOJAwHBqqAM6o76KEUEBmeDjM/D/l4ohFb4g8cw4iGWOE+/m++ush5
vril+iXgRAT6yb773c8P/2VdborNgjNKEY/XcqHsUoKbxHj92qyQm7mzY+9DP8Cv
B55auCop4GDzb3br23HN3PSePURMIEMs93WWsPV3geMMdw9KpAxz6pGR9papFhys
OznjASiHu7YsYZZbEW5tKRl8T+I6UVtS590qQpBm3Bqr331UlffpMNYgK93ahCTS
XTA/sE/A8PIOycE9zzENwnSKFfR/uBLzETPJlWlEt9WVoWgGbYYRq6CJjqNKjPo1
suFdWy/BdEf5huEjNxxPXPQ2UyfGpFP/1KElBT9Z4Zyv/K5oB9h2imngki1IyRmb
G0j8wiqeIzPVIygaSGxfcqzLxzjDt0Fw6GRbxQBXAV9Y00WQEeiVaPUdlZQuWrjS
Ow3qrqcV+9nj3B12Jv0O1vArZEXSSK7WHBTy2WiGl09is9cf/y+bfu8Zeezr+mG2
gzZAP0ZKIUHSbNMAw9hLwucRloVN1jQx/gXro7IHcXOmkAQEjIykVMZ2fe6vYR0n
//zvUQT+eVsSmlMNZDuLOHIOCnQDGfN5LZz/VTJUark0cbpKol3cjAMwNL+9Xwy6
3+YRpJhvA971P57RQbzCTBliv9hEiq2gAr+UZGxWvogtaHWE7K84qOCbFHGPo756
L3ovoekxzyxtJD140uWlCpx0Z/mUfJnVSJ/6o36kJmBjMso/75zdwoeGURK2az75
lZ2GmOyrkPGU+Pza/Lad//FsOBxQCpAlWZBdyIX9oV6hiVWzI+VZMNN/tZ70vK0V
JJ/A+/UYMaJF1RTf3dliOuSRS0LKbM1tqlg9oEht2M/MHxpU9CcupFROfU6NL/wn
oj/Jcv7y86HMHBe2LRbtxeYu/PJNPDSHhUVM8XUtX8G3LfBvj2OkDA+n6k4dOB1O
s5SC2Y6ldJmGa1H9j36aMA3yoERXk/5B1QhQFRo+vBXK1e9+HDlPmreE7jKAo4/m
3Ys4P5769+X2r23FvZOdXJmEzCFxIuL4IWnd34thYiwQ2vdu8I4pwjnPic8RrXIY
HDnJhmcrjVaqlxd7NbYaORHm6J5udc3SLE6zm5cW1+idOOfNIbopCOx5rFC+X5PF
U7lLJRt1XCDiPpTLjYAXxQ7/pxgSIPeQKQxkheVRTLjf6C6yjFBEOv19Po1+eaAV
QzQJ74QaFqlwsyuEvtjsp7BWq34XAE+npfIUUHEWcpIgyI/XLTdIsf2i/rbsAO5i
F2uQyQVBfLNS664TffgfDapw0ticGV97Vyc/84i9b2Msog0TyoW9S09w/cA3NvQP
zWFs3GASxr4KBtsCpdV3Q34di7phAjUBLQsmV3jIV45EGa8H6shnH3Mqs78CxlsP
LfAzm2bMY3gQCc52rA7aNer3J5kNZsFb1lvbIZYFTKMLhl/5FEIRkhzQ+gUkjtwM
qLY6hCUFOj5hYhLFCK4aJ8x9ufl2N3VH+vk5Vhsxcuee0tdUtA0LM3HTpriFgDOX
Svy2pSSHnQ5GSqaAz9SfNgI9KoaU8O7o6yIlFvUjvsWiXdrNrgyRRpjEK9qL1qr2
1cm2ATZ4f9Sbz32pNKaFR48pPnGVPCmv7Z9AFAyJQ83p/VnkDuY8IQ8WKc92fvv9
SXls5H995G074ue6+jEZQHMN7NxVJNBV7JNUj6p8pLAoU9bRuI2ArcGMrBlFNOGt
2OmXSex6H+YbLFnpMjfKKtsA1KuaVYxTi19DQPbSwMiTBVp6ZKezuuhJEfFXvuTZ
RZplaCKAePLJgi0nNviJdLJoAtF/lnQ8qs2xqfNuPrWgrAI4NZ8PI6c+J7j4MU42
Zy2I/qG8bKmLBtKmWG7pgiu43tvrBQXmRyRxOq01cES/jmacHfrBKO4JKXlqzCHD
TPWi+RPd2Moaq/DOMXiLk6hwoPEU7381yiMbXRJXk2w8jvDLTznYFM7vdcUxvzwX
FoJ0WTzMgldkBFSOekXuqVg2fBrhtw1fvDAcCsE/2VvAE/zhc52Pc+J2iHYp6cYu
vQPZbAY/b7xJAoXvsMcvm2U+IcWhZCF+Cikxb+CIeKq2rW4w4Z7hjJhjkU+CXEX9
/cDKNQhIhctuvMRbBmIXW69G12LEi9m0ZcZB1nSCPRVq4iHHo8Gzr4wsgJu2W34g
UASYEpVrwMseN7fgq5l/ytU7ZhCs3+puG2h6XNCcU4oZPZEns3tluc7Ku7xyDxpJ
DzUe/5wEOIvWV5RwKhy0cN/dHOoqtmumO7FTRmp6olpCbuDrJrqUzDbItG24/kqf
0R5TQfEGfTelhCBZO0Y1zZYif7kBtN1BobK8xbjc+iiphXYZohMX5kz/hsP2/aO7
V+ykPVNAZvIiTEdDwqUwG/rANsPT72jeWKul3wfzOvS82px12j+Rcf1ZkHt7WE5a
eD46vRXJ2DMFWJr8UdGn1fVWh2UbIhK+4hArpavvmPLW/SQ/52XmO2lqKUt5raK6
hUEzYKHz7jJt6JHewM12nb3Ey8SI7RG7uCNKq3G6Y2MpxWo4eayT1ke16g8hI2Hw
22E+1P4zWo5CSCEJtraMcjJWEZpbzLasV3XB4JPsawHf3TMH765L+/BGmkuboihY
j8FqSMvWKes0iSvV7OrZeD/b6hU2pQJkADmIKHoUt6TtdCIEuqhN7FWV34ST2KcN
RZXH5Mm/Are3Rc+5FPiLLv8XZMyTt85VrgmOKHR5xkb+4yqlzvFVFMeocrJI3K9+
EqEgGzHJSC0871g++RhNg+KYlvPjYp+Pg+5MOp2oBb3c65irMSow1qmtynPtUXA7
3R6+2CiLoIrAq7kd42zJHtrKd35AeDNmAvQO8yapm8fkZ3MbjmScCweVXEZbfd52
tuNzFcnSmxRLNrSjaQSVTugAyytag8ZylowQCGwLFlaOWZew41xBgVWXBjj7D9ky
U6u55gaewtL0y7O/Wc5Vr9DCI/0C5+WC1aZ5l4w6CEjbBB5Otj0Aqf4MMLB92civ
DrsS7JcZ5G0HtoGGt1H4qMILxUT/ow33M6fnzc22W8X63JvHMJyTBI0roqOCRgUD
9YCjK8kobo2pt5wSu3vCQiovkVef96JgYGKmFnk2Wjy4aEhcb9ZBzINUoyFsjxBL
XVGQC5cUdLQgilFvSC0BoZtBPaFaO+YFGIXNhMoxdwB1AOpcTw4mB5R86JFLlVyv
Jsfy+yPnggZU37PUelma9JCW1/Xz9+d5ICHq0qSvVPS8KZGIITuevCjIf0ao0JcU
bXAI+LEpECkZCin8sC8JC2wB1twTr7dK1OP2qmp+90XwogmH08Yh8lz6clmkQ8uW
Jp/rcoFHtLLsX/olI0csX4I7nQtRTecooF2QPjjkcu4sbPy6fTw5r845m2tgbal2
H6v3uw1n7TUcTcawdmTQj/fZOAVcjupe/2eHE879r+AocpK5ZlGBIciF/VF7Ikxb
pn/X6MTyDuGKS638+PMysrgYbbdTgR0IMbv1sCKoc+wM+gPI+Fwer24grd6PTgN0
j7m46bnzfQRdyNVAgd7DZjxfMsdRiEpLBWX/IP6P8LqN+p/l3eeXKEVXYgild5qc
I+VFyQVM/HSK4pS3sdnDGLE5sOENpnQhD1P8t99TS451PcyZt3jaa/3QsRbtJt+I
TXrl+F4LMmldSLijwBXtSqnrs/RlstSRBCxBEOCMInGEbKpHRClVn6qpyp58wnq0
B9f6KTPteFRvkn7A+zm3Pxf3FSjthyLV80kPGYVJH03yuwQYgeFcdbp0nr/O0q6o
4dArMuGNxHIovQL9g82Bs25IE69l57cB2XO4x+m/NRQZh/tjUGx5H8XWLuDdmOkp
TrT+Xgo4tUVVQKnFbb+MdBsinp27Tp2mJsks5QQZNwZ+rpMAHLmYpsHfNTSyWMGh
B1smdVRccdcuItJaGMQQfnBp1Zw48Dlg/TePG02z0gWMTWAjf8102+1wayG2/HOY
D0GPMF8WDvPONCpixbOBjpUY64vmHpvmJWCzIt2rAVUriZmajemI4niXidUU4iET
uxWLoaSsNISvQ5UGlEEVd/7vKs4UjrqSERh7FCGBtf+oab26r35H9zN2QZK4pgtV
FIR+Gv9/BRsPMn7+DazWmbqF6ZauJc05sWjo1rNHrYNQJqBbW/93J01nemzYQN+y
hDyXphElXMcXT4Ex8vk6fB9vG6lvclsfSpJUAg19ZxKS47wYskztokEujmQD0rVX
XlehdlhnkwGvLPI3SPAVnk/UjFsU+94O+P/XkHtyPbvZlhrqe99LCcGQ4rUAx04/
VODXxkS01eyF/0jZq7oSHW3tLYORd3mxR+epdeb5hnbDBtHiG0rzORZaBciYnxPI
fZdHaHQvNsYIoPEYKokXvCk9rLCkA/PRsfGNFSM7kWJQoXfcXXct544JoOjaWC72
dTg2Sa3aKe14R9IZ61qVZDMpQdPj/UaDJAKzIw62EO/oJz+nJl6oQYXrk1NArgWu
bZ21Si/AY1skDCfHBc/6p4xDgGpG9Md7hmOLjxDN4K/vbAEoS11mNurqeOWSmhBA
+ATWZVj2jt56QHLYzRzlNoDD9yz3uz0fi1YIfxGt81C9H+6Scz0C+J6+3XLICbRL
fzkLc0fSGxfwXpT7HiBWQG9K5qyJVoLgx94jk+cTRVGuv3UkNBJONSYvpSRmiXk+
3buTGzRrEBFM3HpzbmDvM/v+9umDIjd00L8WVDrLTDA/ca1qG0v2bgd6oG3Acnue
0P7OTI7RIHyxpqPn+1Y1dyno+NPnHgMIFZwBriZFI8T8vZBH7LTZe7A8wmxlmmo2
PNlBH6079IEUGYlQ2RzbtMvcjTPXVjX2/2/3QXz/g1n1fn97Fur6qXlAIqF5NRpS
gnS1Z6ZCuYd62I80NStzR4QQI9QvM7u5iUBDiRvLE2iSdembBohe79AoYSRdp6NP
TmFivXYZIlB7qtDn7OWCp88q/L5FlrMDoZBxYLUpgLCk0SFCp+ABwCDADyJe7XTH
MpFrYxcKALvtYg+gqahRr+AE8i3mpHMZOODmXzPzZBcWzzfS0PUTP10FlVUXR3xe
4mqjbtUh9tE9vXfVw+RFEWYmEbLYntKYDMG1Sws4BxeHTnjkUVAgMicxNqqFA1TE
WY3UjVGhSPU1EupH7/t90yOixufSrkoQN0QFdFbUq8lKPuvcfM/YVHido/skYSwD
1b1pT485VFXjzP15rDPf1EWO7rHRsNbeKwxjOJaNo3RKJ1wG3gMjhrTVMIyU33mO
Coco/w+8X3Dn4sEKKY+F4M88r7c7QPU/JjGl9CMBvwCAGh26TPfthOyFhxt3Xw1P
ueXXAA6mRgdU8/wmkL3qvZHTOf01LjcbDhdb1aIoWfF32slQtrAgpcdtPh+38mCy
44liTaSIC2hktZQUz3jKl2cjhZCq8MJpx0ZY7mKCTG78CrvhPqUXfYr9qqCK58Ue
y2AOUz+Ac+/jubwZdeVlRH7xkhxt0g1OT2XT4OhTbl5H72GzAgrtmOstUOehPN5l
yWHRn/t8Xov0S4tjw235JD6rar8YPQcH5HJQWTVu0LqFr6tlInq3AMj0aY5AXBcE
LKOcV0pgYG2WTA7dkJF/2IELb7p88i1bNG3a8mrMhJ7Fjw2uWA2u9wPY42gQnbTW
IN8CPvKBBx7w5IfxvaGUdPs8nkT3Pwt41yHLtQg2HGIwNnggyGQW/ixfiH3htxpc
NTk2+EkZz0NAKLRjqqIswTlUu7eS+w5j2zPHakgYdkBxvrYy7ys9WoWxxpjn33qz
ICWuxLr4x26V6j8MnyvMKQruJ/9F3YLtFUFYLazViuqzBQ/AcQDDECbLjjZoV9g9
5E0624HHwCsMLS4k4YjJ9R0RV3IAYFcjotRn57OZLncpQrdZMflDPf2TulAPnlJQ
uZL2xw9S0vHtzkL1SPWn7MWOW5KYkEUoWGUwNMGsqNf9wIq9EFtvhr6jZC9ci7Qe
sjJK+RnQ5GlqqTLd+7k+Fk8FeivXdp4mWx1PWtMeZz/PNQs5qE3OkYQzAP5ejGp2
swiQEzNxa5FNYcVC66hER+VmEb9j0HXC9pYd9SC6BhoRCejjmlDGSFEQihvn05Vi
xo9EGD4fDtVfXLdQskOTYStpNjvoMGUCAYr4JXH1Nr4g+EpKNScH4qnwWfYgVwhd
JefJJExvmbP0byBYqV9tvkWad0Ff0d+/5ef7Q8KEqOecQR4lvSpa7+amBrmaDc4S
pdK5Vaavd6noFQxVN/hJ9mpcVYDoafrlwyI3LHC7WAVeaO+BRxO1nRKxwjOVhDff
uFH4vFqyrVjpva1/MJIs2DYGFR4MOLrr+BBih63BbXi9BelswiDPg8OSz2lqRKvR
pAI3E98KCudFfJBh9F/S4yPqb0QEaTH+iPN6CGiOzleBYbDCb/MBYtG7QwWnDUWg
47YSiJprg0RQtauu67fn1IRK/C8JU+IvfsUGJmrQ/mtjui4Ea7HiYF3H2SWmhryE
DeXsRCEGEgaYpk6cX5sEIPk3EUwZaJ0ZrJXeeSy3ry+kXdkuKhTnBYmopZcksMkf
hBHbNfq/r2QeGn+lBsSi6U+DZNs7gIrHvcUv3ACt5V8jAA/cgyg7T6iZjii6ujMN
AsYR7FmLRNZVy+H3B89EZJNQ76g72sRr99Cbh2iX9Q0y5VNFtu9WhixGbDtmyWD5
DIYv0r0uYQjQfkOQYQ30IREyE5MaOHSsAF7U9sXs997FG80FDAstjuMrbXqAw8c+
LIzmsTTsjIZ75PIWPv3pbylQzsGC1IHMJ5W3vlUjs4MfHRs+PvF/gZ+5yR0W7LfJ
rP+6EpGW016n4/PJG5jCD/q1WFDSqOER9bYFN2qX8ca+T0T1Z8mdZYYhXsnxESSB
mUCyxIBdNBY4NReX/oS9HQhEyHlhPfB9npGd9h5opy58114AI8E5RPG8OZfRU06R
ITRz04xaArcQkdh+A/B0rqkYtdYyFs27rHezLmxW3+bXeGhAloWa5r6dPCX0BZKm
/TqC4XkIevnZ22n5SkGfMr/mDf4c8P1X939ew80StGgM0Ygs73IQXYYHW8XrSNSd
amd1aGT0842ilM9FZJ6zMIiSDvMey/XezAvzNMMkQUusi+Sx0oqFu28Xv+sOwzKu
Mwa6BPaJMJaV4Qc72qUGhAKChg/ryTt/p2SNa4W4OsIt1UKFeZRr3tV3yCOQXfu8
ICI6+MKzMwUkp2t3YGvNXt8J71ZbnedfHE4fXi9//v6TnPVKVzTyKrBHK3/F4bMI
VMzY3XMGpw5+gUYHvHgz5oSK3oPeiMq9FFgYqZe3/l9XlOk4Eo99W4hT7XprnCS9
418kJR/TtAbBgZTx06GGpF+RD6CxYxKlGjL+3tWUAhCsDZ3iC5WWIVhoEKigtlS6
hX/ukMGeZBbhi86X2tfZoKCcqpclP5OVP8dGxWEkFj8YcvA0BBM4fmKdCBLY9NGd
lFA2tGkSFDqh7X+XmYV9VWG6Rnkw0y/VQE8lzEM6km4B5kNai56ndILwvW/BGb8G
cf0ftemEexlObcmUPArX2/HTRdDbSp1g3evvsCdxcXvK6HNNOWjrnZjm3TELszmu
Iaq+5qV6sFM3qAf3O59jwgU6YRtdUGGxSjyb8/YqSnLP9Tdb36J4IOw5eWqkr2Pb
rPpgThrV1Dbn1m8gh9cy9mQMRWyIvckb8M1D1EJELVZDhx+aHMXc/WvniS/9mSBT
g2XoW1GldMHXU/MCEb580Q1C+cTkckgmUDX7qPpSJxY/CdrBMj2o7xMnEF56UU5x
LkdiKQ2y9Y0hQ7uuNDQY0vRF1LAEdqRUCh2ENedKZiNCozqF8Qn56/LUMyu4Vbgf
3f5lsvsbI5ceDMDqI2vf7swTDicybMp54Rp9sRCWrvNbjddlU5n1KVhf6mcUeaYi
yLM2ErPC+Tvf0eaSXRONM7KNHAaJzuUHUS7/yegVMCqIbeWGzoV3lyqALkOTurAU
11n6sMiIOQ1eok30dvi8oAuzzkAWjGPlkoPicF33dFBUTVDQVw2ETUb7445V6yHZ
7nszMIr/LESsjN5i4Y4xqfMQ46KSywc5J6TjuDJZ9FS1jOIN+zsEjVNlhJTrPygY
QG/DKYKujGCL/jqehWZ0Y1ycn4mUPSMz7oYx7+7SIgrkuMpUv/UTdQGQswMmpP4S
KWMp6hQdj4rEi3bOG29d3SZBQYwur8H6G+CCoSfsIOwL6Lry7ZwCVUTbI9B3SAYy
dKEN6ztiU07iAVhnA4nRd3EXBwYyBX+IM4uYSRDHpDcuQR09CncVfqw7btYkoHDA
1QcEflHI8s6BaWBqU8e/fAJHYO64jpY6U0YMvGBXm9B00NATR7fjaE6VYunGOvYd
elXBfL/QRGsr5Y65TESPEJnWt+5dDbArFtTheth5ci7f60hZI0UDQVP2GDHYTaNW
bx24sBz5+Qt/9eSeiSnRslhrrAKn6AR5ZqC1f1a0SHkTVo5+XUZ1WWyM73/hc/NJ
ZTu6/b0hEPltRCw6ltt5hUQdfIdIWPThovU0gqC2P6mCQIdvsQwlAK0yKayCAXw/
8uPBCFAmnskApDSf+BhO3flVb6qeZGPWk4CwyDDMNd4gS5k/qwbYosnqy6LjxumZ
nwGswkM4GmCp+JgYE6Ti1LPWmo3bKZYThxopvID3kvWirA0YzFw6nvgtKNnmqVYZ
scEuYgZXUKdrdQzkme6FD6eDjx8IXq9jsigN/ra3qnOdXs8qfwDOcrMl+2ikt7CC
uTMFlle33HT8GrbPh6frnymBo9368EZR3kvSJE7PNxbLIBjNJz27daIPJ2dRCShw
y0W7kFRZonTYwwD4WpdlbH9MuIb80ah5Y19N4hhKuvroph1UYn9qiHAD7t8DxAg/
fxFmHuVEhcZBkjb9W/tAKxBqDKdhyO7Z/M+vZgwzOiZy0Khq6KwOWQlzdXkS2RJJ
MfxVweC8YwJA222ecpPLqxXGfP1tYyGZhCHF+99ziSK3D35Gs7KuoPtAvGeoeSxk
cH+XC+oyiRthH/ylWpFwFMnpUkx5z5DPwDNiMCeKI8EnSUri++JuUqcPhSOLdyEb
ESdWuMw08hSJVe2JDabsBAJ6q5/eHABVoybzAsrar4nSdheuLjYAKU9do/gFtwXZ
Ep4nPH0Uxb7OTbV+dTSTsYFR8s0HFBpCVUJUgdQ+Y70pEoXEzs1FWkSQH7ryykb5
F7+NfTeBoQIeGrbznrOvvdxnJRuVZlxXzKThkKasZvaI1OGrAamX6tpj3Iv8WNUj
P32k9HYfhrJHDonKnvp2HTbZvoUoxG+iECuVIr9beoBlr12AMggScynsw21640u3
EERBA0KRo4mCJN4DUkRVyTVEo2IUmvqpAQzzv/BA3YiMR34Hl6Wyt5JfSFrJY0pS
CZXYTyfPhBD83yKMH5BvoeYvVUZKRcKNEIU/B8il8zWLKdv11DdqAq8kqa3qNaOx
HQltma6lRgTzx2zAtw5M8HskGN/xpTcai6zzNVXFIZ6D/xHOiqYjOys5I6i7OPrq
71SJGJZnmb3wRI0b2HmJf1zNw4lIA+Y0wj0NGeGnBMRLRVl+bhKnY36myrzaZlqN
irj89Uwg0yDurL47wevv5fEobdFJaYHz8S+NcGxw+DMF3YTxmKEQShtfSeG7YKUU
zsn72Vyzl0rdKNT7yLfRzTflo0X95NW+TpX6yQAeCm0V+gFCqqdo6HdLqKwMUnPj
APK1UzU/iFgkNCCSOvHNU6MGcc/NW5mWurbunLLrwI5zjtb8/g89VCibFO3NSu9i
xWLQpIMDxVxoi7lDGjpL+owxV8Wn9C3Fh8yBSbRnxM95Uerf65uWQS/x5qCetblD
9XtQflmh2AXIDkfkYx10bMgTbkZI+B46irKfEGSzU4LaALynO8m8GnZz5hi41mnS
SE+51cnK3FggiigYHw8sFElhGi71EsVplXeElKwVtElWLng7048/eYFaZDZhXW3k
L/1D11WfoaX6McPW9hP/HZTEyOe08t2qTW9sYuHEKRsT2V79/VEj237kJXKtmBP8
nKUS93k4Tppx8BtpaKcwXc+/n4AD1Uzgh0MYlMOQEzblcTDJrnDnB6LoG9UomqqE
xjAQjg5ylyUER81oxcO3meAp3jxg0eQyW7wahMzKkBtUf0U6D7oWCaEMCy8p6VSM
y24L4929Pa6OGo6zB1V2y58lN0Z7aQtpxHw1WqL7iZXRJOM9yziUmo4e6PmZAmha
O6mvX7iwiUyOMe54BxlPRjjUCIxTjzlhVrZLU2nYFBZbt6XE+N7wgm5ACJllsAK7
ZQt7qxLEro+lFwt3PK6mv1517EDHB2BOwBTUDPiqgEI5og8MHCaq43rrhK4XwJWr
YH6P3RwpyNR4BVQUzNoyGSlP19fIYl+lP/847I8tu1DL8YF7ddCR4BziljwvAVPw
gibkn+0pNBPM92Q+lDmsFxZebN/uQ4MgMytsz147coLpFDAIsLQaSqIwXLHJEiwb
pu4c+s1jrYQSrgT6MBqLd8QcoXpFUneaeVBvJE35V7yCl/DQWMLvKFaiO1YkI++m
VVab7erwxdpZMRAaFFUXW5ol2NTqalTKdlixuSKBn+qogJIdn9zdWzVvsHwYXloU
i8wYCPZQL2kQKgxvZRC1P6ae1GRPW5PKDI0vleZopZL3xe8B0ZZMHm13j0RM30cp
zqg52xsHKRPQnZRe4B6+dlkgw/NU/0V/gFKm/eynUj+cw5fGtv7uvncp0oIzkbnb
ul6hgSak+2EGMHkbG+WUhV28nxyq/+dIjl/7pQdarrrANZS+F/s2On/vrxGYqwpg
LWWrVe4dI2SndjH55qfuDJ2p93dIUMCeVJ1CSNS21/dOJ35qu+9Ps6D+eEfNd0Fm
mBxT7y2dL8nh44K58AimIPF6bFaadeLr2FzzgYYnVOFC//C5cGtlf9QgLHH+G8Ig
xss3dGCRb84U/O/lrMyFOyy3Aj2R+b4YiBw3326vQMWqaXDyx2NHuVLiamY+m1bO
oAhrTlL7XZYds5qVqpAg7laXwKKxOgQC+OY3FWsHPPoLEeb71r2bDjo1xOHfJ06a
n4ZMyoMD0ncz+lbix6OGyVVK1k/APkGL/rRH5QxjXqHw/8TPaLbCONQPqy79KMl0
R2qG8twvvo0HA2v0tNAPpRhtkRtlzcvF3FQa78rD8c4Yq5Uh8MvwDlFgLUtMfefk
/z8sfuvtsDu5sS7+UcMMTuldDD/MWEXAQz2LxJ3ylSUZtK11SHGFo/0kNSSeOwIf
qVHG6eAL7SOphcthqZHxRBuWiM+eHLFLrUJJL/gerI0L7hsOVVY5o1nTdiXWjj3e
66F2Wwhav4PXmNK7jsNRlVovpy2JpammwWCdCW664C+LxtC2gELC75m+pWXbQckC
yX9Opwu4XeOl2qAgM1kdURb4ZO55nDEEg4GS42vWUePb+QbDnGAf/fvdwQAd3orV
dsCpTfGQQP+wnPfTWQXV0V94yjD9AQeiCcOCuv1vRtlXfsQUVPr670rV8/5MxK4v
tvWAs4fHZp3jxGVaRXvFaR7JI/5gwCuTm8VMvjqo8/69RwPmeOUxGDnb4UKrPxoq
lL9gsoHQ1ZhjJfgX2FQKKL/+Rc0qsbvPVPOzdd5fq5es1zjZFjmwa/uNEfrc9+Xw
nghpdYkqv9ndN4EulRO/kEI7Iq9HktGa8dXaPazTVkVOy/QKor1++dcUI/VtR/Xw
13bPjdgVwQLyv2CLPPfBraTUmdVNqRVGg1dWUvC+JXW4+/jtZrk4Er2ug729w9+y
80YeGfCWUe3XyFV/hxTBGnHEPKjY9t1hOiugrY+Csdi+A2bcVP8X/OlWU01CRWW5
rHzU6MMsAIOnmyKgolmapehzEAzjQ3+6+UWu0K6YgJpyFqD2SZikwd24rR+FSoh8
LrLDeesph0oYwUSOiXG6yIGyA/fxTVoiqs9DYY6LB9oRAYUUF2XzJBF9FSUbr8kg
MowTN7NuBo7u5onN2DJ46gpb49cLrpAw7hfPrUJnmuf18Qh7wL8lMniZpF1UwFeI
jmuB3KkvgqG18pBeqpxQuO6P+KhYdu8Ri226ZYbTaKQqM3EAskWgy/jxy4qbcGrR
4oLqs/Iwsg9QDfMbfIxy2HZH2/uzXChpB8bZTf2JLnlR23KDLZKKqNZy4PXTsHgf
vN85xdWMp8J42OJCnbI7Y/5t+hokT8d4GEu/314O3lhNTKOViGNOqujA05COoIkH
CL4DQ6MHsa+NBj/GzPmA4c0pRqTIvpeK2SLcXRSvCzAjn0iEUKjf8YcR3PJw0cIv
/9D1gnJp3OMBL+b9GjgVhidfxrTrg9vPQpDtNYLUbY0EqHoe6bmat9dDEjKpzV3H
cbo08AxaUH5r77U1uliLN+9X+sNkl37m9DW7G8pXVHafey3HLpl7l2OQrQDaPAAF
TitCdvQ5zLibpzN1DRWMFjF9J210P+235OxLj/Iep6YhoGYGIta6yupMZW11x0cH
sX2gtwGB9fhGCfx7/aVQxjiIGqgcpUe0ebYjFX520oqtZ4Y8TgGfgB61vcv+dN4M
dSGQ0UxWSSzrZTBocvG3ioOZZ45rd11dceEhnyCJjWw+Ni9pJKbgE8d0KLqYKCZu
n5L9tfZtus/rejPikT4pChRQeLu+CkUG5Em8KE3IqQvcU3cjkz7EJgggOqD8rceN
q6nCEr2VKd7GaXA2MMPcpXIClIm6ZIcDBF+7KqLY+Ql3zuzozLs2LdDQK6A4xIT/
KZTgoX3UvzQQnbZHql5HcCIN4dqEAHrLK02sOUiDj4feN3OJ9bKTKZ14iWhyO8Y5
gDJ+Kc/IMRiJlNrje01FUk2NtGeLwkN1OYQSQMeyoVMwOaIioDo4eEGv0zLxEwj/
Ud7LYUYmAzzh5DL5F5eBGopU1h1XE3v4rQGeIfnemfh/7TiGLoxnXZly4yuN4kQk
oZvmKlmJHAN6y8CAAuG5P4INzD8bb1GbErC5b5F6qjfiq08pgoMI2StC2nGyRZOi
Buma01bjxDav348QVgQLGFDjsjVX/LK+naDAALWRHCJ28cX0RrUTDUXeaRRStK1g
FGVMKbWITod/lPS50CEK8anb+pM/zsp5xs0sfHlmjZI0KhsOTrAcl+aKuiV/oHA0
WTlG37b3bxOldxfhXCHTvap29vv5ll436mMld6i7mSoz0zbyPkX2Hpzps2LutfdJ
eORqbaZproXPE2PVV46XAPPvL4CgsYvc2uDsMzjkLZOzDFgR+1TB976jPubbZGCy
qFQXYdOxZ8MZIMwfskWlJY5rNEX89WHFkVjakhBGIA6veZ4GuN6AfDzYaXL4TJhj
EuFqIBCOxX0WZMCV+r5x74Q0F70zkCHkmIuJoLhnaUWilLBzdgfCFXR+vi/+Zpr3
tna+dFrowoQNJysj2BGFF+fvZO4risOlPTI9CMKKVCdQz4a9fSkuyGoBgAWwQwzC
D7gf/lZlpwxtvbSg9dDx7H6+5WZQ9wDRCBU4++hLlKQEFXrAqYUa1bYyWPIMKRWH
Xcb7o83U4EjrthHAu2g/dGHEMARLlhiywkmm/jXJUXCrbGz71pEb6ClZxa4O8Uzj
mHyuLORlZBvqUyn8fFIHtK41rtkecbtdr9MsVgO0XCe+S76ZgSrn+3+nMDHKLJPB
MWZKaLIfxk0PMUpWlcVQcgvmPYvUmCBg/E8F4totpJ0VxqEL5ioNZdMazWh+xSHC
Q8m0LiTHoNtWnvqAix9vP6xoKDJZef5A7EKVPOvlc8KqGYepTEuG8ajt5EqD2N5i
OqYKRhhfyu+V/p/9MTGuKcIxijoR6eTHtE/51zBlvg7vo7IqRjfJQfHPwlYUROYL
7u/JzWLfeXywPTFYLsxOCEesGoN95G9XwEuS3mgeio2/fqL08+BgJoHjO403ucgT
DduqOh5RN6SbMmvitBsFQnSWs8kr6QfN87FjzvrSCzjHvz2T+kxqWsmXpAxFDxuo
+orRs7KwnMdTf7bbS6vbGdjkCYKm1VKlFTj3CfvtNhh4XlpQ8+Zck2AFb5+HsK5U
ltWXqBu1nyCVWpNz0wtNCmtdPcAGP3i14KGV5G2LmxvwiL2EVrOd6WOaFfOBRz3U
O/GcgfSxpYTXY/ByM0x0Z45tncZOd5sajaz92WZ/Ze3s0b3RkMJMFLqjZijUzYdB
GAA0j58R6t2VKW8AzvB+A37T6yFuRzkT7JYimKjWE+KpwCq6EyyEd37dnNZvRtlW
gkZ72Csu+tOpdycle4cQGzeQJTg7eeqIh9HlRi7leu94PvMIx1ZjiAX/uHO7nrIq
E2eCviNmOkNWO0BptZjw2oNeMmep63ETKVYwDgI8ZqryqVJeCtSYuCBOKQ9s1LPQ
wrXJ47NoaeeaPc+EbyNpAS8diVjuVgSYwrZAOqVSQ7sobWJN+rgJRoGqDziQHMtz
BFiOwYIsrTgtT7UZbiEXXtopssPrMhZIQMP1zYv77hOsF2e7hy8XQLvwezeb9mAb
+QH61L3HCVLnoyZgMrFTOOqzotUj+2ChDWxrgWiXkjHEGywXYONmknfeyo5D8Mgx
UIzTZM36Go41sDHS7Lc+zPaLi4wyHEQzke7ZECFAjp2Gc6qzauDURucpyff9787p
MlSYdX/tTH944iEQzI7/Tqnq9sEAJHu0obLqkEExZbMRVDDxDmo07fV2LuyeE6sS
JiBEa4bHk9H4qebwvGYj1MofXCpUZhDuzJCy9LkGfBiiiKZk5wVnHFOSssgwyARi
26iWCR9j5tyu1dRylMt/sVU0Zv4sAVVHFRgyYSr3fmITj5L17DqJrZuL2zkeflU7
QtWFMCKnumNNRwquZyha7z1Pp4eF8v+HeW0cK/e9rlG04Z7qc10CBEBXO5NB+7Cc
RoNv4D/Hl36urHhEzJ+9zYzm2awz7Qwy3niXUb4SnL9PRM/63fj3+IvbxxrQzpYG
pOvPOLgczv19ie4dMdsFTUJtuqttiiyL9wCHyGxMGbRruI9dW6OKBJob4V0Ldxf2
GBbVtEgBq3fHrDMP1IpfGp4RToqbwBuGmPF60645iJKahs9p0B0WauD/8nldqM0Y
k05G+0XKKznG+C59dTEXGBgFBnMudaJ2mtXiyBOaZXrMLVaE0BpD7QPtR/G5O8wX
7V5YaeuO70ecGhM3bttQqzIHfpjeNgN0QokQSf05jQa/hdoZ2oxnXvqqQmkr7BQw
l3c6+CioOSc/CG4xhaAfOSjFxRiEWVErochSRn2a2vISFb2DBsXDBzXe+y84MZLW
4lR2AneEnsddAxeAdRq/sr736dZots+dG35loFyuDm7rW2TE2HyXXStF7L7/6C2I
Q3RMbPtT7cSU9HugYh3YolcrBlsTb0PPoz+us9lQZviCAjyuDh+//tVxrNh1FcmW
jvYG6xzRHLN4S2hKCQaaColJA9onH6I0zfKAWEDhsPAn4r87ehQ6KgnJb2GItmb3
2kd21dtq+snKOXfazedmeHKxgb0ua2jpJGYG+x1Jc+ugIfmXLImVkk4vuYYQNnNA
B647TTOOe9GG18taqcmuhvWD20Vvkq8PCKrU/34yJrjwQDd0pe3TlXS+HDfKZvMK
tpbAQ192jIBe5TTRd0XIRZkrNL/j8ivRcNMBGlXg4x1a3eU8FEOELvhd0yLRlHQz
s+oqydwyu9k/lcesfzaqjLrTEl3omH7KMZZNdF1Tzn9AXMiaR/Wo7rSTwD+5OGho
cOjeTmeer8yM5GcyOM370xnRHOoAdT1GelrtrPg2iHqFr+F+Sw7RluON1wD+tizw
jA7jYReJkkhZuLBp5Ne5w5CyfF/Lzkd/RmUntzdzqA0qW02KJIjH2LwC0d3V5uKv
+KFhUPI4kHddIzbb7rp4gVxU0D6VjkJTyX9zBlarV+V81PW7bvx9dYPI4XAv08D8
rTWAq9W+ib3zPfRiWWSqpoN9sXMrjZDR28WTZt/AAAbm53XM5BbqFXGSY5Olx7ri
tV9HuHyxDEt2T8K9DLNFLadJo4m015NkPm4YKeLbtqgp2xPsDhW4yKIOBdqslw7Y
7uW4d2bh6D1jgMfYD1T4WMMtMBgQIh6UtcDSC4iBuYVVFYnboyl0r33GCvMRdbIM
nnVb6mD0bFMc3sPNRoIfLCvMCwZQPzevy/EG3TQDymOguLY/DhDG1ojgxmOesThw
O+oRo282rRbbzB7l8rntJb9N2vgCsVMbQ1uNUW/FyK1e9CAIguN7PKvs/lWJ0Jwf
scV3oma/W40n4e0502+ZQjovkRPg7x5G3ti8YVgMdrPW7zg2XLo3scsS6cPo2cAg
uU9nQzm3DlQpw2EcBNsOtbR28Wzl+yP01mkt2r1XPFL6eS/wvXiafKPQ2Edu4uR5
u5RZC58ARN2/rLQU9L9KDOFz1mbO0NJLpEgAqwrho1ScvExcEP6OZkz5d+EZkPjt
mBMNadNzZ1MVXRinYxptD4HWWnwk8yGLF6/Zv1ZhphVwNI1AAuC8gWZhr180D/9I
h/JkV3p22eS734jmFyIg1sLYauPiegcOHbZ+Jmn5/fZd2jfJAq5QggFiV65HkvYx
79zoyg3Fw1x/EDDLYRwmrq7oZK+cFxSJjNUajBogNihzhMLhQ0pO0tYx+Y8LACHy
LuNas3+RsKxX2qnoSdF/4qve3fp1mFR33O3+EWvlg1o7LIWVJtmSFshvauHZHJMj
4/+OWrBkzeM6uUKs/AH0WA8bXiqcRATGB7jMbj7QS6YQVJoUwgHPWR1OiqGyuBWN
b56GqrEoeNyAPxIfFfwyy7/3WXvUrVgoDAnUmnFZD+z3fCdTq/sJvVYjifQRUKrT
5oE/zcGVSA4Y+yNsumbqBDwGNKkg8Z2t7k1Ef2u8fiaKLcpZ5P9LGygXnZYPPT4j
qPOiKdR1Dfow2Uz4hwsWv0I7zQkR12/llVQDCKpEmvuxESIeBfTIPfPglvo+CI8z
w0zoYfchwYZlktDWmw4PjObf7dRuZPH9tPelDUu96+G1v4tKXvcotcJ1kwLawDd+
VFBx+7HmgV3Z/GhjrCHWJY0ACdEpokNpgZaGCobAck4AbKzSheTO2DYGNnBeWBIc
lmc/xb7QBC9iAw5gPj0YXo0enf2Bhq6s0S8G4XBLFVT7MTggQmK5ISsQNS9TFZ0e
haPbdtYApt11WBeH/oNrDqFWav4N+B/di5ENBlzBlFHo2+436xSeKmrnvQfZC5AE
/o8FD/Rd5l1lgbhsCTRvrjnfrmPI1u54ru+VYqB+nxm+aH5gUCP6enU+1ReDzquV
KyIimiHydwona4HjGTxk/ZuEVFtjz79aSfMLaW4txXXINkmh1Xn56Fz3tnYgei9p
Vo/SrD+hF5RUHku2mjeD+z9Ubaq6UDa7ugzfcYNATY/Xm7P3kTagUT+ctWIocWpG
RAN3knRlY3HLLqbFwOGWF39ulNEUbeYkXTaLGACtaLzOEWWNB406geLgMHq7cUb6
udaBZSHvRei1YVig7majvFuh8J+WxmGYb+eYfRRLQ/fQrAeCqyxMD9YO+fiQaxu9
gihVF/sP7WyPBIkJWWuOlsyucc/GKNyc2uIqteTjPC2838HkYUuRP2Qdj7SRwx/n
SPl2t/91eK7KQ802xYHfGEPYr4/KafXTqmdChFV1SNRe/4t+AUAsAPj9hO5mC7cl
LLqVf++V8MI734YMQttflksq95hjP10JskhZi2LrtCPiYyluD17HuToS7nnN/pMB
QcJ2DVFGjpTL2QW5LVcTL4sOcIBD0FmaXZZI8RVablIcaWVzy+p5cSlmhpXrxzE1
dAWLT8TJhbmagcn29Wx2ybhNG/dnOiEN7FQxM53FCa2mQhwaCbGAcLxeh9QvYOkT
FttIScJEwoIXS386KtD4V/Ru7mvCl/m1dXD7Df4+ULa6RZfijLLcbN+Rr7JVWHRo
/7ENb4XYNGqx9W6Nj3MpCb11gvX8irhXvgR7wWhhj0K3kpdS03C97yKtFfQbn6yQ
th5Y8g80B842HMe/L1o0oQmkP9bMjRIu3RW1n2sVPuhp2kprEj/AOSe5NYFswjK+
aohDPTz81oUlSaDMmab6viRwY6EeIWf7X2LGmhAs9CVUFOLZGNHldFTYAiqBaemB
fD+pNkiJZHOfT9QSOJF91n63dTg4kWLr+9pVjc9Nl9Kxx6+Z/0vS6qVGilI1VT2n
EFqN5pUNMnpU3DhOldbDYlwe82DJXR19/W2sWwkym9oPfWyJB3T9xYs/XljUCeHX
+WaOVS/6N5Q4uJGwDcsySwEBJfSYjlvr1zrSBiVrSXJb0Fio0bmY+UU6kinpnVU/
zMwk+T+k7n9rVY4juuKPKnfr7FyuZCwOYg6iov++qbanTFAlTnQtCHOSQdbpaanC
l0Jkg5qwPn2DgmmjxWGnmNHPl25snVXVBFWmzTQIZKmmiTAUaGLseBk8QaNwFKsG
vb5EqnRHQhj9Vl4Sac1wP036oxQHFjUscJIPrkmv+Iq8daIULOyaicZhX64ieDQk
bDE9YyK3/CwGo6+r9PjJcxqOf3blvjgDbF4ap/Sud8TxqXgWz4FbugY84G2vG0rT
Om4Rr/zX6iJpRxDumFi2V4to9Ib73BTcVm/koDccyfBbtPAMw4GVR/uVrYYsfTMW
zmnkJWFlUsCVBl2wOs/PabnvdDNnn4U0BlAwPAs4B8LLTtMm9+aPPDu9XR8AO7JI
IzZVwkprtSUX6Jrl2SfpYp8qfrJY3jH0yHUIcWi0Mzm8weVWSTT8+EAnt0xMxLyX
UnCKxXpcfJCqADhIJ1kstVaClmOluifzlXA6grmd0QyvMhg/w1ffZVrJUEgw6/VR
yX8WjPSbDgn55W3uGSJXBo9Jf+LNrl262BCUMP28gK9Z+KbXDJLPbb2bU9yYGtgG
9ydrhhSSzK7VNkPCYf/E8nDvDG5X6ojTJ1qnlrrpr4bVp630pTku7k+XiK4FtPPt
SqoF0AMriJNQemE+v6oGKq8lFrEUqRW6kBaEPELbvWiKGBdouFkpF69yYxBOUd3E
3kFKLDVV33d27yhAk8r3Tt1P+WNRZFkDg89kGNpXWIPD6evtGJYcMEtsNdKWmxCj
Vt1GHmB2ODMrGJ4NcVTCtgXxKcYlT1+3MjLev0bxOiQsJXzbLB1a43NGwPg4m6DL
phkQ0CqA9lP0B6JmVsV/bqSEeUFfmpbad5MkfPDcwYbTsrgJnU0mFMdwdKrWB4P9
1ZFA8BKDhSNDxIEzuU+cFV5WGVu8tUo+uqOjJL5Al4CDfBbDGuWSZuQphSwOZcVP
3KXsCyjkuyvOOmoGwtoG7570O7T49zWv61Og8sVN2ieuRHxbaTIxVTorjzenEJlk
izmx9/QJKAy6l0Pp1YBrpMq+ty7STDXzKA+u2AI1MGqExDBMfwIT1dnrOE9YtlZg
OhEH0iWeOm5A6n4xYsqctlIZRENOfIRMNlc/9avhTM82BUtoM20veeV7VSHUPiYy
PTJefpQicBamX5ypdOKXltJ1IlkIJ/fnqWZkkGlZyl4VkBeEpuC5G3gVvAcqiD9M
k2yMTx+qxVeusSBzh+OyZgsQQP78ZFpJ1BAa1dZxuIlY6D5k+xohyHF3q2KLi9RF
I05+T/cY5YLwjqKlwFZ1GS+nlzwzvLK1zesKLzmYkWcbEfBZ0y+LxU9A3Ds1UuV+
dwix7DUWcg0KPx1rp2wDSf8QXsyYbkRKYdIyadjX0qhHv+NHh5+8R3Zf5RKfxEaw
xH6gLHlMD/UnIsp0jRXhU+fsaXoVm4uAIPSeMoVys2aQs1EPmN5c5FQyLZvdXNu3
9eOWnu6I/vA0I91nW6BEnd11V/NgaaMi3Zft0n3ao/suKicQu/FbpJmVBsgcUVqO
ZdrEt6rQEVbk2Yr+nPmt6ZV301/NNzrLES7GZCZLVWI3FiPRlvAgCR1/HkjehyLj
kQXYoSm95v61q9jqEPxp9VI0dDKnEiKbOvGhxD7tjQw4OeOOm0DGQq/RvYhiFzWg
F7oevhiPAJ6o7sBtAEnEj4Z73nWjIYA4lm0UC/FnMnwL8ljaNTCFshmudFmLW5oL
cmjxX2RyV9arYne/CZG0BzGv12ZarXT+Xx6eRUwIIYS9UW15QhEQ6RMduXqEVwG3
hjY7bgCIkZut1fnedg4BlSWw6h+F9n9lZilb7PYOqZvbsyIQGyqIfGwsMR84ilSf
r+wNGQcaiY2AotRhwIr7815U8XosfBJ7/UrAE4RMxq1WxQlRihEkJONjsglEXpRY
BmEg0e7mAkSWpEkYnw60TrhyXaCOP5ZUrLAoX5kHmUtQ/LaeRKJq6erIGydsLNAx
4xy4F3bVflnHfFlxkXLjSTTQ0qbAJqbTVpOQt0d1TNDRO7qDie44bmOs00NxrEXi
GMQlExDTglDeJuoUvsD3iy0qFZEQodwHsm5n+iZyiX9ECl9x0mBB6CBw0zBUW38/
TH9Y23eaG1CP/OyzyMziEuIzXsY3NQ+laqJyMWLA6m29ivooK16NPqXq4uGW2NDW
URvCbqqjR84JhsaiNxtAYLwcD5tMLmwRqNq0UsD6thkz1hV+MT3jjzrmZppgxdBg
cpkALG25RlejnsHwbyTJGx2Ud7cc9RrOdiZp6vw+ih58AdhDRTtiYlnjyml8WrA3
r1t+J9UZvhTgUh+smRc9VY5tXEu9mWdS3nbaFpXBUh2lCWkGvNc2mwt6Q8NWWYzq
KRHnBysp32ExnvQcgwsatgTEplH5UaXIg/Pnt2TXtOXZc7Fh7fIIfDbeCdcb0B+G
k0SgWMjd1KzAk4QbOUq9bPwZMk3eSom8yIrYNYFbvjSRt0mkFGOa30XH8DYTpL9H
v5Ob2uG9uS0yRmMR2Iv3c04J3CT0OKwwYfBc4IV95QiAJyCk/+x6DJZnZl8xRnt5
Kolbp6ZMKouPfajJa0lL9Csocua3hnPejQidH6OhDPpz9IJ0uwr3dEVZr+A0ZY2L
lZGhIy5Yn8LpgjvH+0VaaMpJBaQnEEYryF+UpHp3DG5FzMu6im8Xx/BNe5Z5kOYl
50/5NWf6x2rOcjWzWYasnnLusB5UKJErdVj4S55LkReaig7sKguXQIwoMeS/LalI
8RRF++syITFyHencv95IBopIug5O38Byx8qexGOIQ3mRchYXULDkjaReZCEJRP4T
hFXPoXs1hj4L91zJP1tbkanX3/zPVNGFCKCa/w0g611fMX2cddBeudJdCQCd+OLn
/iLr1QZp67HOi573fp/tYFgbUpLKsZPPOXzuwif7bTUdzC/QHfr7iC6wT63uaYjZ
npM8woZUtVLFh8by7U58Enpa7jkyQr2Qag+w3kj0qMHGITGidIu/MSurlo93WxsZ
ch7Nm27iv6fAYywmEPocUktm3Q5k8m/G/KtTtKUKnbpi5l6mDIP94XtV82kxMy5j
Vfh6xUW7YbeNib4FizadT2ADZ8pD0kuLf9hmoYmjpj7RjfK/8aAHqiz2qvYrRL7b
jj6jZ8tbXtsGp6JRTFWmGodkQED63JwVbxHPj66/i71Pwm6vE1sPDXZsIcsQZN7j
MBic4nmZzmdlXl5Ky0ZmIIspu44Mr8TR53Bgkixrx+PoTCLMulg7dER5ZhEvn2HI
rGATpSxy8bw2DZqB0gCuxRHUCIFDGmVFzuN2P6ksl1L7lv9GqhgWqbe+jCeGms2k
WJ6RZixN9ucUpoVUWsJwinrRnfQN/+yAMRl9se+EmAsKsbipgjbK6fde1yQju3Xx
Pjbtv8vkioBcxUJ1bXe23fxl/DgwVtnvxRY871MlUFRXFaPEZUUt5DCihcANv1sW
bWrAIGmMeYkYMM0EQXVbbe1JoWTGDdr8NTCZYi8D2GF7EDalCSR+5JGh3QjIdhjp
VRqBSVWHXsqsc8c/XAqPwE3VMBgPtlI8g5KNMaKvyPt8WuTk3Mg8qJdWVoMMIvZH
ixhQJb/zssPG01+5v8AMeps3v05iv4ob5Bm4B5AsIgXWqC2+Lnj3BMfmAoD/pjua
2F8adv7tO37UPcErry0XTlUdeDbHkqxUshzC8XYFH9IDW2CNKowGNscwlzREzxVX
mw0vdKB2WSRzqmxki+Rd50a5P/Mk6MIwiJkTV7ws7sNYq8KSD7xluJKJ0crDhUek
1gFZfU1lcMT0lT196WARnUOjZE7S6qdbtp20el1HMZ4QoiDxQLYqDBbV3sQcZJXS
XtPuYECgtGuKFNfVEx3e9Emoqoj7GFSCWRoEko5cfPwnjf9pzVjy3YpY2K7VThkc
JDUJGS2s+b8reEvDjuTGi4DJhzskcqVlTyWPSIPl88bzotQIsRGCn9lG5Bj04zF+
ybYVO87jUtWvOUzrtnPzAXZxtqwbYv3T9WqjV7PmqWfGwa5k9ZADXCQvZvfCv9K0
w5rhkZwD++o/pclR3CHG9Fp7mJvJKYXPElLQgJaSe/ASw+tiHc1itKIuscKXEZvZ
wEEdOKwjEKH7+roV/UtRLKNxAH1kAeIF/sv49yiImd4SLREIe8clmirU0oMvvWRb
LDDa2NkBdsUYFNICsxgTVXC+/NLFfT1z1GTmIxGMXsWF/ov9qEYGtkKZe6t8RGL5
FI1rtAi8CGf/vPlm+bDmbrU1dMsH5nJCwzM7uWAOmGg2gr2gmENi/+2T/K6JbEOm
85j5l47j0mpC5B/OnVUnZqYBP8YBq7+oJ/aDpK5Z+3Fc76cBleIiSO8c24CH9wfO
YUfPGXRH3BwzD240hXhAP5lz+lmyEo2TaTKjezXp7qYTxUXEjj0TxaTfNf6znAe1
q59fPRoUoQJYt01o/0TI7ps3ONBCewKc1HvPdSh+5s7gTAhCSEQYsn0gfv7c/C1f
EGuxGNvqxjscysnlXVaZIRlSdj5CyO9G8yGxXUMj8QzUQjwIEnSR0q6cUm1hogAi
1P7hoLzA8xasY9Zj3qGayIx1if69cSEhm8+BWwrkttWUwVylHmxVb5kVCdutKYgP
BjxdsdDQrkdplK7RNI6QGMoq1ElAeWM3JjFBkGGgNm6beDKncQBLJ0puL8c0xCJA
gZuO7YEwTnO4kmmkNulHqu/J4JF3IDvbUPusP/JeTYiG6+0/kCS+6Pf4sbTwdo/s
CgZ6TTOPMVUAsD1rAwKj2JAMc5Pe/JqXBpt1kQvFfALqd7KU7NLWpOiGUnK+snWq
miIaY2W6RmEMb8/jv9PRCaM+8x1rMqnlGinJ4RAmEz2t3mTvK1psbWT5RPwvx5Rq
3TSAl36kIq/atJsvCNovaYMf5VmiMeYHT5JHxnC2Yu04xl9oPZt4xhN+IPOFKsq8
JmpqVwRsT0+eXxOZtNRujbE/e0BqXWf8TccPatLnr5RhkqLjM61bmSb+T5Ph1xbI
CmuvT3+OPKVPYmoZMkTSmu9qWqAabblpO13Qj4u5/sF8CFO4VC09yCTdSJ9ZAbGE
fDFyUqF9/xM04MD0Q0+j9cIF+/ohQrNeM3gAu8SKeB5PVkxp0O32ET/gid5XU0cq
k+83j4OeMG5XTCOsFYpuKrhlTgwBraoU0EPko+3Mg0KOEnhFatMNSJqMXxUEbRBV
ICneNZ3ZvN9pmxYruCZvAGevajJq7XScWpPNmgk4cHkOFjCwedcnU5EQJu/PqaQU
FCCiGdCvVpO1MYZEIZ406S1PHAXlE+06mRP/D9wE+4F6NIq77qtRL+/tqUljdcI+
JmxZVpGzvytVeoQ/HEH7a36mTPnx8BAMkxD0nfCB/FHlky65tKIVtRMyBTA5AiPG
2N4XgPBixBOe66BynFEfFrGaXyqnRPXsZ9Ocz0CZJMiu1de86YEJychG5bqMWeoF
Iq+MqtU33HVQbkkASVFAF1VtZN9hTP7c4PYbWa+EDufEfXwHr46StxPSasmiNuno
Eh4xR8Pk/DlrelpUAyKvXoq2d3I8xBtVkA6Z98krAvNlswoZfR7PT9EuxcNBZzNJ
HRM5j/h699deIk+8FdUXxidQ7rPRkHLrVxjjo2pNWfaeUxt76zyOxqeKldAeXK9V
YOOg/AKYnAaLCrOwpuIEUwd5gtHaqoeffG/RlkkLl1r8kuCPgsIr2iNCpEAlrK+U
76MafUeanw0xnLwrVmQ52d2Vy5Ic1aZE2lSW54HpkTXpTQLuMq0aEg0xKajNunKH
INz7WteKIYvtAaLsy2G3xtHHgvVhVOuB7gbFAHRWigXu3uybbmJ9D9d+sMj42SYf
hTGD9PA8aV+epdofMPQ4OA1197DhW5hleSfQ9FWOIRRQdNdYMJu0Myi/XMwGGO81
9NkMq8yqQhsZa9hmQSQypSOVLp6HFh+uYhlVBSc4fqz1uHJ8OuxeCb9WAtlbYt9N
KRRbesIyKSXTB/qyS18l7WApyEHNKrHudI6/ZQkuJytyzu1NqGZ53ukaYZ0SXxsx
BDgI+O6QgiRvMOzW1Z6+M1SYDrSsJvanuimbGcXm2PD28a2nBSe4Qxnsw82Rg1Bv
XNxs4826EPR9yk256jUVXvMxBZNlMpfBViBrIAb3ug3VY24BvUui+sAK+Q0Zkqc2
HIdkwzueg6mtrO/MeInYixG4E5/+UwLD+aw7le+RCKMPWjEZZfsS/HEYMr4qFtzC
azYIqXcSCgwOqHbWY9WkPBC1Bc1N31e3roPKtybQcHBlQ60BStrIZuPZZJABzkNO
4eTbrBGZHplvyHNpciX29GyperrRdn4w8w8vfc3BD/chxR9OS5dyCRaDMeqAteEE
ULBW0eddWiA7svhRkiGr/+75RV04E68CTn4AQsl3P0amPBAWew4upqOF4Xk7VOgj
pG/kZqBRhR9hNp4kLSYaTdtx4OxPNFgIcKT4xD3fVv2XhOvMX0rhMg2SbP8cI1ZZ
sHxX8tizMjqvAyW0ztgpht7FB/CFpFVOYINe1BL8D5LsrZz3tlT39NwU5iB+pUiK
sMqU7rBzlkK7xVIPnRyDpDB0X3gXF6uGR4FAgVO+n2kHM8CXKL44MZh1CepVoCKd
dTN9gSDHA78c6P1YooqYerhhkrP78RkqjxRPkYUGp+v9IVmwrTA7UNu4ZIZT3M/H
2LO/mj5LIrMrwhv3cR2DCaRXvJhdokAAtGFzY7WR5L/8IP6k28HK+B0+k8kJvRoU
ZuuB810cT1d/U5uz/IBYWRfsIhFVp/zLAYwtFu4QrUGNDlMGF69huo/0Iuh85btd
CUMw2CAyIGd5mpLfZg7P8FkPEk0xVnUVghPw+3AkIx0nJJtVNYbX3eJKoYhxVu8K
db50ZnpKspXQVTQ/BCDlk0Tt3skfk49K8+E8K2KZEW+HfIZBVNAZKxpYptvsxNIg
Wc62mxm27SDykgIk/KSE3WdGoQhk0LD6CybdE76o7Tm3Armx8uTbCCD+ukwj03rF
AbjtHvF3WVMkThjB1kkGZo7CK4MABx0nxXvnLquzDgzamhE/k+mX7MzadpNc+UaI
yH9K7rrS4wlL2JN9a3I66n+I+75R52A2E+INNyy5dn01Ep066Td+rn0rSpVaCCKx
jxjjwpcrMPQsU9XUfq8IoLi78vQoQMFvl9M+OAGO5S+xOHiQPjKt22nxY8GZ9jRm
NuiRIfhD5sZMNcFPNUT0itivswSM8i81VkInF4ZhJUzGfHRZM7pp+Dky6i0OutXt
qAN+FC0MVov/38Jt5tfJESTN+bSuIwYg8NERW4r3VKS29iQzgdJwAliHJmutzMOt
KUXEKMz/0O4kGkV8PHO9DLb3jLYO41cti3icIogK/BXr53RGvBfBMszNARm3kh+2
NbI8Kk1KA688OVgJUUkyCzFd2OO6emUhGMpmnoDpo//LN3mCvt9GmOyninWzg6xR
KQM9fa4TITzC/jk5XGv1X+TiwM20Unjy7PvlxRcw5z67qWu2/RzycO9owQ4+1K2Y
Oj0l4MaSGWOkM4K2hUd7SyBPMh/KgJNBSIFxWdFHZWm3n3sWxuE4wUQSc6ZBovHa
6mjxPXQebbxUDjRRqYtspc8IZMZurkRdNoW3pdTbD7GSaxvJSdqPqjvEgzR0CDRo
zOFm3O4BXMNen2CX+CxKwlsqTjLjf5Bi8szx1r9uz3VUXcr19pU8gZXQfD+mZKdR
pti2/tMfLZQwQWLluoC8HTMmpXt/Ue9AJ7fZ6MfL0cFvAglmudFJNVwiB+XvZZ6H
1cZqJ7OM34qbh4NomkQ/fvd6+gsK5ygJgPCcW5tPDaxGQsN4DpcekGwhkrhH0Aer
iQYnKmjVubZBSy75LLmAllKlKkoSOt37xcUnCPy3f4E44cWt5IiN8DBf+nXEjkXp
UF+EQg8RkVesStJpSy9GiQyNaoK72jBelp94bvfiUpDlenSYQ3MqhtnvZZhjwhko
qbB7MKdcsMPf2Ef/AVaUCc2gjF10YBu49DAtdWsRBdY1wJOeZTPpou+cJ2lOHnL/
0QKfvYzvb5Cn+vjPR37x8DIgiGGszqQdy2M6N7JsbmuN3RjCubrsEr5epAwbo65N
rKMhhR3huDaAfNVaVWzrT/FaFpVq4mmV8c+xPABJUnWbPpL9Ay+xDDAdMzdF5ksW
8r1nGFFL8yp9ZxDlmdV0IRBdrhLdraBNHomMdGvEphHjfurjIPOusqa/wYvLyz9G
naJaqiKiyxuTgnhWUPlpuCTJ8jl1q07VA3GD7JyWg8v4Td8TiPa6Jagtqmk18HDK
glR3Rarq/KFMDMBCofWHwTZOoD2IJfpBjG7qRS9aSunerpHR1KEjh9GGE2YxEQNY
68UnEnLIQut5+q0CjlecqeMtc4rk8v4KEWIpMlAitaxuE9UjhiPpsyUH0pEbWXwO
oRcNkVntGw0a87J5j0Y4meYFWmDZae0E4PL50rIeqC4aI6s5WptuAHkm8LqCBixe
9dNab2nztv97nC8cLfKX9lWIoyODGJIHQKXLZdpZUACjhEK7EyCGTm0La2eiPWxQ
HxEyHA4nNrqAHcWGuY1sfN/rbUNnIRDDJ29Lv4GhAN2NTKDV9bmmixUsMduwbL0N
hW/LlTdTaOnCqRqARko8FU6oKF/Rnbu8lAd+Y7/9vsPQDRCLnsqPZmJcFQTNqiYQ
b/FpC8hOi3/rVZ4pHouNuXcu/hwSNp2bR/mlQTAvbBlFOgof08ICgFpZEUD7BZgA
YjhEnPl+9h2GOhKclP4S/8lsd5MFub/Th57XpMLneaqT0NWPJ44Vp1f9v0P+dtbN
6+uMqsp1/2BiTFMUxMe5esFHr+b0q7h9PUAEvJ/CLYJxJPqwn3XWCTT+hqfsLrIr
b8f2qRmL1sKPeB2dH+Zw+YCs2gxVyN0gf7+8hqOXA0GBKMdfGENNzPx82GROH8bv
eP6dPfQrqQRW1IaGhkcfLFhxirhQZ7MMo3F1eEPW77aDI0QjKEff8MB4IRue2O9k
t+DBN0luMAc3ChfcEFU+a6nfA8UOjexi/wCZeC1FEJuzWfXz8JC3sUK5Ozlxg1/F
X+jB0knG2psE2RnhLZCwCeYlAQ92d2DbFxzTc8hPwDSgve+p6sEE9cBu9y30UvuG
WttYdj4qOz/fnd25ZXxEuoyRujStR2ktan6UT5PYFnCW2ZdTK0MBKw43GQ0+YCjo
1BrfmW+kG8/ct44pmnDN/+20LtufePUutHAgWjIR8aLV9hbCxMKZt4Iwz2PyAqKc
1UZ6kfo3Ogg/8u7JxonSLNxRAAYdtH+VpaM/CpU9B+sn8031bPy9tkb3oyU7ermG
T3vaD27C3iQH8A7I92N3Zi9AGwyEuq9ouw789IXHRKQFuPdesdP3CTvdh99vhy5Z
x7LxeMn17AfYlXbKBtuu8Gl6aqvci76feL5DzejhywuihPpNwArJyAxv6nxk0nVn
z3OEIFx681DgfiXx95GHSjgCdo5M/s3hOqs6l22JGjQrVc12eRdYFpUGgQcfz6xQ
GzDQl0uLyRIRFdzeFtU/xy1frKCQITX0Esbjg2+sAq7hn4PI3p+MM6csykxNgdQp
ZcH4GHzvQYwR59i10sQjPZbwPKTM7LNpPU81ChL012ITQIUU+L3iMlM7u8uOHar3
GC9jfx34LxbrH+tP61li5QNOGjhrVymfwGMCX3swFyzcvy8rtps+SBdmYfD326ZD
WD0YQ5GCLJ2Vr/JCiFPSp1EnUzckoGUdD6WEDRTNaAwfz482E94lvZm5Ms2Pk1W/
n0EHX1a9mq0trhN98jzSz7aRTORv+Qg9KYM+yC2S5IlB8gUsAQru0T3rKKaztMyC
Jn6bXKU72AqOQcAgXJ9NE7HCoEMpTpD2+PA2UhckmMe/PQYu9Inq4WWGkxozpKIg
+DncCVxZcIkr+2JthEgz/SNv72vylcObhWrGfY6QHO+SJV47jPCUtrUKOUd466lh
SPEFC3aEiuw5m84M4/xm0ZysUBaOE9k874jLnAVTPOnei94dLbhj4OZepdrDLI6k
8xw/W+612xzuX6NXgPdOl42boqWGC6xsYHzfcEGOKQ+51CgVUEUVziJ90vntMaRV
GtFUslXI23t4NX7SEnr8vskjpck4vUCbAcG8LZAZDGOMlbAze6LRu9+Z7ON2OMx6
V+HhC1WxuFyQUc3HRe93SL0ojvWEKICoaWWtInIF1GLbT2R3YcZcV5vwSLVCHV1s
fKOuVPCTiufW/OJwqjFk47zby0J9Z8sQgNeM+57n9ZsmigNYsAAn0AoFo66ACvKp
fcEwba9lpZNDdQR7OCP4Wyjkd22xTaTGEJ8lbHewSjssh8WfxyoiglrT7jiA6Ic0
aNTr7qtRo4AK4NPezWQKM2j4PkjSB85iiPcEc2IRQWu1e+apPCZ8yDIQ5CXsEwFt
WPGBSpKJwhSWziyGMhYfqoFJ/8r/GqgXdMWSs5vKuKYnPdsDfu8v2Rk/wEGS6HWx
uWKhJPmfzwZ69J6Dgnrzg/Uh2o3tFhDD4wfts+XtiQfj4LPJcFqbuIcLJTQBezcy
GNoe1JqLS9kxeu4E/JrU5i4F+cBKO81+MJISY3y9vJlB4rh56+kY2zmIDlys2Xgr
Jg++P6GXBmMt5hbZCyVWWHjMiO+YDkYoxx3wm7XYj3LkkEj6WaVX6K3BLOVNrPND
9zrMpgxdH00AOqpttsINA1JikA84Aq8kwHXTVuQGBUtqd8f8xajRMWifNGKja+Nd
Pb4y2udM/mll3jqMIAUNaV7xzDbABp5WlBmfvbAI1cPN0QDZBdSJb7ubQNDS0Afe
WsYDszPcWk2zko74bJyqORvwI8YwGyme6d2CkB0kwXVYorS3pj1UnsaIurDrd7RP
U7pvajN0O1ORAVfHrrhCk8x5T9qctSlGFR7zhh8n4EUP3ikjGfAU0leL6f4SCjrY
6sgrPsmXr3N7EFIy0Tl917EseS2wsOpfUtBhDpYoC0r8Gm8k2KBddn7N2dKy6QZF
Z2DCAOYq9tuaWByWIu2lwiVkA8ATJnqbFdw3a7nCb7FWPLKyx+5jHKBdywxBbO6k
AwHIUVzt8FdZuaX4rc270t01lhU9KHtdNbz6EpJPLD1fmQ9Pr/Jq1vT7HguiTXxL
IU+mF6wsafhDUolAL8YCKBrAHb+NSiakWVdjHaSIJduTWY/yS7vyKHul3i9aU3Lt
VUQYLbUlU0h32Wh8x1zCy2/M5rLO9dGhroUE7tth6vFmaYNJrhAHyrBtKbJUZ54x
GcvOHzdyFgZueWdvZXrRRdmXK/GJgMrJmmpX6QBExNqzf4jV7BWZfnnv9CM2gx2v
uAQS6Y9IDHYejCw+dMymp4goW8rTo6xHFpdzQ5aEQG0lGJEJ9dyt9bed7c2K9AHx
BCVPCeBPX/0AFECONxFUQBpcp4wOLGXh1/FalGjTxsJ3njTQdMlkCcoUSBrmavOw
rp9rNSWoDJxLZjVOHuwdBgG6HEhZ+7MZD+Ny8uEXxrnsIRkiEGhnG3Iu+Kyz4/0W
wCYZdJy4TWgnqiBWqlji6ZXngyv9dMjVMQlkhAGmmheyft+iUKfzsoDWgqvB/98H
xi/VmsnK/fppxF7xDyQJ0/TLBAjQIuoY1Iqb8DgFWUBJKl6nBtTLavbfVQuU9m71
iIGcm1EETo6FioLLM5+SZ/noSqkgdkPt+vx0P56GZayQYkJi1QqoA4R0IKN6wBta
Mo5aMOaNjpperDnBBLvdKY7ijB5I/AQhkTpAqbHP5exO0EWbQdZCBuyt9oUhUGhz
d3iR5tSjhKBPNM/4jjYV9AlId+Bp74IBqZOB3tOxMmazz5GqUNh7dPt0OkqSVPWe
OlYw0xKQxm9pP6RsrRZYCEJbIWsVO/VS+Ry8TzzrjiW1Ko6z0xZbbfgvxrYAjj64
4hOT0Whk4Z9ccTLDkwtTQuszMp5QuA6kQYB3ne4iM8VSw2C2LALp42QfpbytzXnD
zraUDOOONK7hGpqvHSFc0TdQtwaY1ivTWf2fSoHYGBCPz5JfOnjDAStOPK3n1AuH
E3/eB7X9LmJZdSHbJx8HbQa0DnP5bJHGHiz3McaAEqE4j9eiv6obJNJA6Wgr3OJ9
0jmc91NWoZJzwy5hpZ/SV3q6e0epdTczkf+4z26Rj/wWe+hyJ+O+nXTQdlRtevXu
jXMXjgUAqvggvpqUAvq/NFRdlg6l5UWCGompVSdYDghhSVqILkEmMFZ2k0pWjj4Y
srv8wv4sAqhtPou8uyKdhJtnA1hwVmqB/15698p50CQwY4bhVNzjWNa1umnN1Y4o
CtQ26SSgH0dSWcfuxOsVozRCALN9eX7kLLsPejzz63soYLXSBHzTA9O4ZNeYHEt+
eacAu2EYfzJ8OrhKvXXCoMUjTvpIkcJN+bOWNZdR/CaKx5vyU5WB+7ODBN4snFyp
uz8r5qGpamgghk9dKzsJFzZkM5tG+wm+7IC4OYtueRs/mwXCuk+BdsTm+DsLsjgH
OBMhOHL1B9jAAWhPXvSwxjuleUS4oGRg5c3Z+laoBUNCoOxpDTGIg5o+49c2HEQ1
AuORaJGNuf9if+nLsFZLxrF//USb1qnewp48fscWaYCyuTZCvERleAPkWjknjifP
3kG+dJCctYHVtqa++lh9HglTiZRCNZv/4AHVwO3IoJ8iZO1FdK1O/BZbmaUHHHWg
y3kw0yyNEDvlJlbX1uykHjikOAnCtMWjpMUMsuObcFYM1zfnaG9pX1MLfdz3RHWU
OPwzuo7Hp8iR1BlUW3fAH7fYrv3Zt9W1GN2Q1kHOvF0a24GQixzpeovvuRUamhlK
gYn7fbfTImOpnfRDATI2FEHR5dQ1ddWz4RGUv8y+4UNUzTMxHWxdnNpKz8FNraVz
niJ3n08rysWNNPUYNICxvFFQeJqOO34nJAqj1rQNBn3yR/Lc6BSXa6xF4sXMbak8
GonkzZv6r6WrN6t+lobqxCZ05rB5hqwo2EYk2lXUNIQts4o6A8SGSgjQZpdFZkrc
TP/TRYEtspTWDwdUAuMNsZhfKU0lkT/uZtMbm5JAw6sJq6b1Xz3ZJQ1eEsbjadBf
9yh4bHPwVoLtl53SXEW+0M0+hsVTuJPZW68kisHgPRdzLH9wdYS+b27DOxoaeGuJ
frYbeoTLbWClCY4O4GOqtNXsSqUup+iIZ597MULQmy5F/xKy4jLpkfUa7P3hbdQP
OvJwsObbfVQNOE45/gjgKNwcH0A0JUwHmrRvgyFKb2qU4QUB1IwRVtawa0Ht7G04
prmkt4aA3Qkc11QsbZUaRsJx3/nEfqYLAuLaviw/6VlPFFs9A8z+G44miX1WFng/
6K7mMokpR8MHW2CPE4JK4y8Ieo01jAA71UQmfsN9yWhi7225vTvQ3ugLgVYSSLSo
QguCl1kvqRLuMjAiquuiZNy3fRx1nhyHDGWcPbfB+jFH831qNyr3ebM/Pu5VZbcx
jQ1XO1op9SqqmFlOecskujvHEJwFLUcPynDwY3ro4dqtJ+asudsVn7pjXbFEYWX1
NOf1rxa+ngDTXuGOGaJSjrvum19dvfdW2hx4B6GGwUTRmOkA9r694anA/ZiEGYmD
/jZOufhJm4IJO+9yZMUcyMRrTbgztXz3Hw51bxgJc0g9Lav4B3NNYqACOXlYw3ll
pK/wSqoaMvIN4rB5hvzx/ti7iH+Ux31kSCDGfT4R0q92yTPU5oTMCmnVfx+5GdCe
IhlGeRMgfriC/RiN6BiY/oVwHIzv7AtFsaW/KUoChaHFK/hao53WoMA/ThcPDt4S
L3P55zGbmX9LSPK2W8po5k3PbDRtpas7hjZN8dmWf06ZKpe7TcJMxu32NTIN71MO
fq5d2+2lVA4vpcJOSYZvUqXzHRv84FhnPooxPA0H9oAvxD9Xl4p1fUmuLCwxZbXU
GYB82397PwQxDmFHtWS4HfUbtIZpAoE9S0e5UMMSuVsluiKK06B7UmMz0dtzHkEX
Ot0sDXhILWCpaUkvnsEt72lN5JlACbT6cBVpPSbYNU5vgcA6PA1J1ZsOpU2/KQsL
ypjO3Ej6uSeyBM0nO64ufHUUmGAhuvGNNyz0HA4EghC4WlFldrrwRMHGnF1fghh4
nrV58QUJu/xetm7NeBO2wwkGcbMUvLAad/FJu/t7v+p1DHjFyPOhaffteIQKNPmG
onrde8nGB8l4fRSy/tHwJH2k029BxIxe4b0YTuJSRhSO4p6en/b7lAvUeTJd0UsO
6k6VU/vXzXr2ri+cPMw/TBO5gycd/ebbbxutQfwICgKbkuaRZ8DAS75rq0X2nj6l
1TJInKfaGELtzksmN01tTv1+6NszkPDEDgwiUU/y21NgryXJFLPe1yKVhx3eKRHu
+4p12PFf8RGWkgVUGGWmsaYMg6AzpUyxyfSsJ46E/3xFR/IKAx+FeCY5VuUOyBZ7
pg4KstecnQRb6+PiS/hjNIl02K/WZZMc/tcCgwXkQjFi33iYdlrR0b/q0T2giVOB
JSR4dkCk/+QY/3Rnw9IoDpeSm3C0j3NOcVMml9yoByhPCncdMiNRe/1gJkMacmO0
/ONSfDw7oX1+i3uTQu+PEJI4tT909boNEOYbwLCPL78CL90aoLAjb+JxkfHk9hpu
u9gV+wtKly3YAdMuQqpRBGIQnMflh20RKNJEEWX9XmcnHuRLlS5gVuK2sTABQYRT
3ExoFRN0nMdUg5j52s8HoPr5TBQo6D793SHFJgy/Y0wMZCTEVGslEpvNDs71GeO1
f4Mt5/Z1YWZScCJr3/fO+kJEMSLWv/ig5gWMfXNhB5Xr9GLER+ZTbYWZPq1XY0Sm
iFLkxpyqT5O6m+4mYL1nbHFLt2IDaOPnV3vITk+6iThF5JJqcdfjMRitoUC/MVbs
lOuQ/TbdyVyou89LzIR+r7a1DX1To7L2MM2BBqD4g8PyRVEn5enVqVDMupobkkSf
0gi/KoKat/WszAmoKryfS5DfZ0jB5yKmwI+5hcliSbOgxm0MgXjV9RbshmIz7gLa
LFvRkbi2OYAglzl/eSnO05IDEmpqV6fTsr0kBnpkJumKhMbrr6qt7baVDQx+Z7md
iBG8jlbupEcAjMLw6EQsNaTtSqL1ksuBkn+q9eRYwYIByFP6AoIAxUg6DWo51ms+
Ccgex3A8PggzxTP/NW5BzDnODg8vR2UhAABDeGYOly7XagkC6OI/GZBlgxtF9WZR
ItIHvxtFcLim5ixl7zsmB3cF6Wo3mylAy9F+MNymxzXf5ul90V85AccZbiKJq/22
zYpztaGtSAWX+hPfMi4LVXiwwAmxpe8VCAk+CwIHCXyFDMSPTYwn6azKKuZsoQ5c
hpFck4sGR1TgTOYIEaEefQmpnXYJlJEDlcOn6xzwP7q3MgDXsKQ3X2EJqlTilx6d
jDoSThSgsA3aKTMfjVspl4wPcM04M18HEVTMmzjZyjjX+snOBmId+5cedmJVXvSp
klQbKVatDAcpmorT9PfcuP3OVLBoeTSydHzGLaebwwwTYqdCQF29w+VQtoCGElF1
0zlsm/qhraeiBigaFL3rHZOMY1YsYRbAesUJZrqae5pbzPC3kfMCQWy+m8VJ0qIb
gTtpAnunEK0MI3zDwO6zemReKo29nbgfloc0SruyyraexybJJ5+73gxWaGs1YdWL
RZfpX/rZchxTx3/4J0SHdprT/P9nklszf8wjnjiPN+7G3XFL3lZJvGc0dbURp1xv
Ci9vdqgw7eJvzsOUcSO8HhA7Ez41371XFvLfbUbsbYLQsLHGSlw0LaJgv90GsYTg
G4ePhKCAAu4olqqQA5E0prFIu0ngPEGsWHq3jrENdPhL/DFb+WaCFk/6oWuc7AQT
tpO1/cCVB9r5Y8+zQI2BrNLwYxWRGeVzR+T7CBvMcQn4SkqpewEqs+zrkOYaqc0p
KNsqJuHSDT3GMOh47c2xnq8HZmn+sTlZWEGo/LTP+sIh4dQX13wUNz8iIoF5PnD5
V7ouZ/+QlQFaudJwFjCfFKnV8CkIEkcWKMX0gqhKGdFilJCVHA/OFiOwtETllHFT
ft/xwLOHUgC0cZPR5PMTSfooMSgdH1e6d7CX1zfgj250sqEFQ0aPkqiWgz/g7dK+
NpgxvcN2lZEyisfYPADTZ6vHZR0vzBWA8CowIqBksutk5zfqMIveE57xQRfpPY66
O7dVQ5N69cO3gAqhtLSbZzKUP5SOgINq7sMM1UE5qBkxyrqICLKQVXNpRGR4Iqt9
TR8hm4EvyJLu3IfzDPfW2nKrGwaSuJEbyRxcKs99tCRmd9ohvt4GWaqGixIKebqY
9WjoyA0EEyGqvdGfvl5CsJ7tK3BeSrNLDgAUmDZhGoe8r/moUGwC+eMS6LDaONgm
Yia1M4EMJryfFUDGqA41uX1CDtiQ/ZDosyjsiguZn6P+6exzojuZlLcmZg61OA8h
bNTMrBC3J8oxcAyb7tgWJrcnfomCdirAVcu+qhD3UhIuUhi6p+ozEoX2mPOdv5YG
lEMUVuX48MrbRScgGlir9Gy/TznQR7TzRI/3EvIF2Fu/V8zMr0jiF9Qe9yOBG7GF
R6fE6ytfHPr+RJaV4yzFZz7k/om5bLlrHmNngj+AL8267rXX00SUN1ZaF15NbBUA
xnQopIaSX1Inczw8/OdYLdJbFix8iiaklcDFcwycRzl+ei7QkxTeFvJ9TmSp87R/
xwBs37TnbaHyU0/Lhrsva/i/E6+3W+aVAAz1KmgjVjt5wnCCQymE4etReZwbTC2m
yO7JWUafTPjZWsq6uaJ4Yp2mkTNPIyfnb5jEdrtB4z4LYfdUfis3/VWNhblMigRj
JVxjQQ/0yZLL/IJCctwUt1H3iR4weS+d7NBDWtxuv9+bWjy6f9oQsXc4XZAIS5yy
eKiSV6aNcZYC0LRj2UCHcTrW5Xqbi8x3B1eZTUMJ308WGJaoCVkt0sG7PyS3dCIm
s/zg2N5Gh06MBRxsX3RHOE9+dhadtBaaf7gy2o8YLWjhynT0pnO4bfDyX4FEcjvA
tBothadz8AHME04smhfgo16ZWJi2E17OCNODoatvqZH0JCpvWWVAwMEZeWKXFNqE
nCPZh/0WcECbeLD916gtr6z0CKOCmvwjDOk4kwe3mpGsk6/rrJxALRsJmIlz6gjX
0++3vFZEfOgcc5UGBYZoCfhAk11r2o7fJjjEgNU9CdIH37RR4AxzjxJvyke0YlSs
HSnM5IOwrzst9kAEOZ6V8dlxKhbstzlpzWI2IKQpCNvY2D4nhM3JqBqnwz1A30PG
k7BE1L+PYCS7kQx0ZjVNMH1VHism/jGL7EZ8Td6G/ql+9s7pIUXjBIyf4mD1MNXO
HuL79LInkpkarCZkQYoXD/0eqFU3XZSKddkcEdean0sPQwuWEXDUQLKqUSfhrOfB
hWFvcLHbslm62xafh1X+qMvQG63P5LUHAYp7Yk4loBKkaU53HRvQFxSWQ+XTn2A7
64Q4jCVj51bCSlQ4TGoLI3urWnnCi0qzvGT0M+HKT78oYhFU8FHqPE9PQmL1PfcU
+UnFuDRgFMXIIPngltvNDiEuX84+QO80ipTwY8XiwM2+XZ7mTxCPbjOpL4716TM+
y7ObDGdc/kHCqQYzZVck/bylbcvY7N+1EYL05lCp8FnZrpAe8tTBubSmKPcnKjyH
QvWsXvKZc0LsWEtIbgXclJl0ufIpr/SeEPfNsuZK023YpKshTnybFchsQsTi+/LH
xy3ydNZ604IbQeBK4IticyEfYeTPm1EyWXOUq+1bkfWg8NKIISLYIa50s4iHIxuz
Ghd9GVmyHlaCwS1Yjyj68bVVc0gM6Vo0xJWmOc/ylkd9osELeDwvwOnVWptW3zED
TFmMIjWeWCoiIG2FBj3pX6MEKNqxErds5q5T2VYHxkeLfL2cQTMngbouDxS7zl4C
X0up7kRGxv6PDUnvEEvEuX9ed19Zoi9bLlSW+fbFPh34a4hG77zQZg4cVy7zagYK
aZK3eJZ8kxjNrn6DZGUCh1XysAvJOT1kA1Vm6u51/VrF0yxbEzrn/QmW4QsGbVQX
A1e+3LDMtm7zS484giPH0AiPTwaJ+oXpDl2emocENVim+Dng/o3XrQVm+V9Jv55d
jogwZhnN8zSNMYyKMz5SrRvkdNDM5IQgUg2eE/mN0bJBpOXY3rJJjdeyOAjEyceK
ybgBzcu3lBv0xC4lE8QU2meI6q8u8YYWgZ23239rdVKtPEAdeT4omginZuICEJwY
EvM6JrByhNeTVtVEiyoEcXmoKfPmu57v1XjrCjxxq6asF4ezWETdtsYHdeI16wSH
6CYCL6ezlLy+vp6Cpo7xlBvWQRzlxa44pAB0tAbTMVP87OSPmFv/eWt0UjX1SnXq
CF7Hp9kdmO/LqRDUysZ4SuvTXGymiJqTUjUC6yUvA3FyfZzDbr2IivuLB03Tulbk
bc8QLOVkAw1kG7ExhDQZjH3IRJdulCmGLIIAkib0ck2lA9FUW87Zqr8coCdpjZFW
gCTw8WBvQwEZZ4LdvtXR+RS0AbrWAgsR+lgBviyMQUKRG6vptaUOuU/ZV1Xusb9Z
2o9daNDndfhjXZO7KgyS+o3ZF/MkgU/+m4mYreISe7rTC/KuOxLLpfK0m48zYyAC
Ltg4RL8CGflqcwH+S5khxYkODDUnMranjXQ3bVO12Tp6hLHzCCTqo/H6UKZjPMGF
csZjR3gvxQlJSbDvveL3LXKxFnXNC+iFkOUfCZlVnp1lUFMW2fnNouuvFezYDW3H
oTcZYizvCCLljiUnPSU4wfXTFMI6e+G3USjRsux/OixQJJfLdtguQ3FjY0G9sts0
lO2G6v2+7Ug87hc1IEJKIHN+4gaHDtcGHaknGVAEPsdC+RC46rmPesShMuUsxAEJ
5h0A9nkngH3++ujDJ0ybu+hyXFZrD/V/Yswe+wm0wlgMoelEOgQWCZVNhpCFMQS/
wYI5dck2zXmh8N0sACMnVatUFB7oi2nQt04vBleUADjKyi8tYJo4nS714NDwlHxq
rNgKGvj9RFcdduAArU4AdJoN8axOPSYroTeKnhlyuxh6/Amv8pPDDwFnvpRCwrCV
U1rkS6OteY7/sCBo7F5YyylZTDJhiwcBfw9E+U3NoA0CIWaooAP6hcFoTTZFaWHC
Qm/F9pe7AZV+xF9XBkEl7QAD/YRxcuxokB6IUbvPEkSbLsQcQDuS3BKqtlM74WBK
HR8OCDlPde4ZopvBYsw3EH+Tr4haRZ5u8hJuf0zAIHxvLZo5istw2dDHuww4BecU
r//HeBPocPuT8A0rmpuHttppFQuJcY56wRpUJ1/D54zr7yiMwa1WVbf1mnr3gWf0
qxBzxc+puDBiWtGuhFkbDmqnrnLymDeOUs0VAST0bHk6Eb5eLTL2DUXSWI94z2ub
fGRDPyYAOqIpt0xRmi8Z8sNN2XEvpB8LD+pB11iD4DDJjX3FAmF1KGz6gkajg9Zk
qI9pJzwjc2PE+xXTP/qrADyl5oqbrzWC1ozT99rP6wP2tRcFCBuSp7x9CEHSpPln
BpNd5XOw966B3RLQBs1FtZ/nXfMIKW4W94d0OJJkgup0McJ8XPVpe78eu+fSza5/
eB5OXrxb80eUqeCTCfioUZSCgUnmKNvcSNtqwTcKGqQYaQTtxPyifVraszFSeCmM
3Ob4Y2oCkgztdynorYloCLlzDgIqkvhmD80HINlpSG+MuykdeHHuqzkOGbM/14gS
vPpzstOFrqOyI2GWPMyb54qXjcbnfRwTRqjneKnJOIhDespqdTjudkXZju8ULivp
PjxW9s5/xdtmuLe3AJ/5tJE+GoI6wx6tgnUStZu2chXCS8Rpw0yCOQYpBMl7nQjY
z1ujjY3z7UUoVoDHQNZeJ3C6taH/B3ZCgFmrJD1QaczX3P9ufXDl+XMTl6PAMrft
ex5Bq9gcS6/U58wY3Ro6O1zEKbc3B8WVsHeyz1LAEHY97UxCY7Dl9/WzS7ELXy4D
yUT6CMMZWhn27pyCzvVItHcZnxRCx9HNX8GfdSGM0sVxt8MNcArvQLhpdFbBlK2N
HZSqH/oYICe9X6ERuRrAwDl2S970tbeXa8tSCGBiB3qyQ7yK1uXTckN8AqnjOTym
Lm13LCKIBfndqdvPyw2k0iDAPsKg2K2ZbD5kh0FsXCs/QwzzqzaRF7KSnP5zpqEp
B25lKBWMe6q0gu0qam9reBPSb97fBWIIhRzHPIHFiXqqBdlB1fO8hHbLlmdVd/Ad
nvCcGmuhTAKqc+HgDduJeSdi3V5h+pn19IEBleAkj4yjj13Chmx3MaT2/gAzSR0d
X+i5jubAJk3NgTIWwR/arQdvhfRjb5KAloq8wYACzHvz7/oKFRE3MFnEpi36yxUP
ZhXH87W8mM+7AdASEyhvfVQB46sRDc6lNiH1FHfbZg3uUVq2eytTM+u/Oyl6LENc
Ig4RcaBfBAgrQZnKWm7nyA3qui4kiEorolVUvVKnkhKY33xwtFPGYQVVtzJ9yIo+
bJUNzabBr8+/ry4JqPUNoBMzr8NUSexT6nSwZz+kau1sxapl2PlHOf8rvlGTBhBN
L9F7B6jbkez8FNae2CjnXLBjAnygqsf6rV+6L7QRHGcV2EvkbpqlRutqZ3yJufk4
AHRuxAF3Tpyln4Zf33N1XxlzlvMpUZVACeJcrTNeoDb4+pHcK0ZcjE8u6FOI+Vti
8Pv3xr8J2c+GkGt6s3IE4rG5Eh3YHUdvMFwBL2OSWdc5vYKttGutIsChjLAx2QK+
sHGIQ3b7xTR5Ai4qCrHo7OPEGR6+AH/y7Dy2IIcMZm3jpF18c9C9xhIT6i/4FvZm
Uox3Rc3PGCnmgM5BokA/CMemE2WdbZXL2ABocqqntwiHC8mfR9U2ISeNQkvPk1XD
YwVUbrdhAQjL4kByK6VNMPamkz38BZCpNTcQzA8s8Kxhm90EWPllgvNOjwcT5MuN
j3qfsv6DX5hwjVpUn8Fz+1sXGXJTEIGIEg3trYOR0VddriyWAtDh6oGsm0bwecou
XIbhl69+a8Nt0rB1ypxZ/ZsUbOis44yn1ksAa4/DHZzFmrP9oxmqXd/ULId45Jjk
DNkK/bMJ9JuB7CyQ5LPWaOGWAJlVk2u541G4fq8xjHmt1ELPTZwm9EgJXNob9mwr
puvUzdbW5xJ64ufBtrXqbfuvRBdC7LXqf/aARvSmSLg4CmA+shk3Usv9lwebrn7Z
z0DA1qy+Cw1THMAE/du/8dyH3TAII6jsMxe302cdZyS1iaN1UHZqWp5SL4n5rtaF
QtKCXc0D/3qrHUNkBwGQFuwu/cSwtrLoeaAW38Dg4GujJHbdDkQcjThSedEio/aD
5rZVWVyDkVjbGIeE87pvqAnNIdCqQK4BYpuh+1hBNJmFhBtMIP+XtRP/igAU8RME
sNCKWoD/qM1G7pX0Z7OFMSrCu9KJTjQ1u5+z6YF5LOGb0yrwpwGJmmPUxZg7q5CW
fxQlIfUl11np73In11g7aaipDXLUrO8hJmQhBjQxHYsZ0seoLeb2Vge7fJWsmV5D
l6j6r8rq5YLCrBqhuNGpaeoZTh8AxK0Da6AWUJCm3LKBQ+iOSWH7IRuxsQP7R+H0
w1yVUO1rekQXJ8Y260PXqpYo7+8EXV8OySeXhFxtwc+v+WfmyrnXnsAH7SCm/kaK
tl4Me6Q2YXxWYB4sUMemTJphd7sKuY/cxL7syD1cRt+eIdhHVMsoe0qL8H52lSX6
yQ+m3ShbA4uDhxfdzBW6KasofVLcdeKBaNROuGnMibJqlb1Bu3gNnlo3p12ZaJqe
SuVPwV+de4XQujkWWvDXGIyflzS2xJQWqlere+Jt9l4dLHacPhD2BKMeMQNr80qx
FBIbI1QxLribj1GMjJ+eHTX9mP3i3I3dFir0FDnZky+kiaLs04K3/jKwyxvnmHVv
QZ0k5fSes1a5w1KsQUMBoA/nTJvQCofd0V8wUC1eSGEJKTALEpWxhpXOOPb+6OG8
NCCZu3TWEbQgAuynrqizwMCOCPTZ7sYNNJOCSlsy04f3VgXjdps04Z9qq4gqskbj
UKK2zTIhn9TSjoHdzl9BdOXaQ2YYkgvU3nfu7nNjExWpa0NQFUQ84S7L+eTrHJAC
ra2byUaieIo8PRpKoUzJBoqgB6BNcNyw/KYSkYW8D0b0e9hkp2vSsS0tr6zumaMg
4sFNmN6ovjq6WR3bhafMgVvYOZnir7wRg8AJZqtJ6p7vTU5f3b7kIDW1k1IqsjMU
lf2pQCNDbkNeaziZN3hHsBINgzBxHk4jwQSeyEe3B/edx7A5a//pQAUzgbyHEdTm
WBqNDOIAQDwnZvA5mgB8hNIhHT1dm/ggV4B+sTh86mWXtCvvt6B6RZNZ+VM5zbvI
Tb2Sl+aBsx+cD2I6j81i0WoAzfQkoE4YZKV4PN9lqFNnn5hob8ZIlKh09oghrIXT
1sPn5QfdJDiZTofoMSZolSFN/sJcYtRYrwOZWwfbCOyEDoXwYCALXHD6vj4/aS7o
uLQDh+8zae+qQmbeqL5aqiZt+J2sBPq9IF7sMANrojo4eDfdEqaCE2zwunDe0sYY
Qyz0cENuxg05N2GACS0KtVTWQrH6huoeianoMNeBKcmWcAOHSo+Mio/oISaBM1kt
MxDLx1pNSqOEEvtDtCGwl3K6jpCgEzwYbdX9V4BPWAT08cJo6boC9aLJULN2BawC
anTTd6w9bjNCx2XW2ty4pzUxoTtqd0Ou85e9Ae6S+XcuY4G/61TBwDkCvhjLmqVs
HMwYekXd03dBxztsrmH6nYzWs7Q21Gd78Ld44zr5jpHh16e/gdrGHOzxhaVCHlhe
/tiH02uqFvOY6rjkwWqG7HlDqiDxWl0T4nxPBxn7KcfhkZRLP61LaaMS5YkmFCme
yE4GROVvOypvYwNFYyy1lXzJcYB9MxOQapeWlk/OOa2z2HEmW7bDZJW0gHyETtUw
ytP31IPh+QiEAyydHFEGBBPlRh8IPeK4KGyXdlQxHvCXDxd2UTpxxhG74+ghQi3P
IOImBxGIFZapAqYIwdG7Y8n7ZiT9h7GZ3ADRxmK97/CzA+FAEJf17hIuvy/F2Fjr
lKcwR2soMJn0B70WtOR6NfoCULNwPiQPvfkM6Q1IuC9iJUgXqASElYC/no6l/5cM
VQFILEf/qxeCv6kMCEsfH84+nwC/52p0q0Grt3rESh4gbfgRJk9ddCrZBiz4xd8H
sMjctXIoTuKe7yDp3Qi1KLO7hZSEbET2Qpuq0QLPuGNL3Cc2DR58TjJ+0S6rwpyf
/QY58AUSFFBhz2I11urpnl2F4hSGfq6MS3FJZBqQm8qnt197cG09PPd021bVIM5N
WdYFOvfjT9pLR1hiY7BYKiywBFtJWeFW3j9FG39dr+eHB9ryAT59lgwl2aRppHHz
OjMG25t1JfbGNew3AUF9mftQKOhm6+2lEWxRRG8PZk8l1jLlRrg0vC+rZc0F+Njt
zR6hjpHtZI119n84mve0nrGR+hp9cnxdzxQ6ENJEurbFxr3rEZiPTIYX343agTNX
KjQuRZk13FMO6m57FRfYGWkHosFPPNvgrzqBGQ8G1DOEL6vM7J2RG7nBQK0c4hOX
MLlor3OtuouMqKYsROqkWOoFegtUQZIUNdn3WM/L69SW6AGQM3x5GWbolQ8O0nLQ
neWLMbEShhIMoamXQM/YV04ohqx7RGPkT0K9tKmH34Kd5SlEQ+tcpSI35UdZaWwf
hAtf5D/rgngw1PeCu0X9qc2saSRgpX7A8XN4g7Xu7VZxBL9l2i7wjE5mUfXEeLH5
uOYV8AhMnuz+43sq/N1qjLft6LaTea+/1z4EuuPG7lIGXQK8zUiG5YMbfGZUC1Li
6HduLOX3Ts4QeX4flVxgP+WZ75v8LQj7rhAP/UdncLV06RW6vx8ld0RAYSKxIwRb
VfMH4HSqLZm7i1iukIlu48EV5XCmQ/Ket10x/AUuh0L8Ujz1QD6TAeHEg7XtrH5A
ibHrEpUvVKklPXrFV5xoAt9O74tlS0h1tQyPC+d6Qk3KbwW2aCzqlRUxtkX7pxZN
9vEYg3TRBxwZv+G6QZvusi04NGako8Xqlrq79jjNQzcDWgM80k/R8DyGUmgKxNAV
Nhj5Ss/NoC6JVtvhpw0OE7NFgV2SSmcY1CvAvokqedM5HXUsO5+UMyhu+oRLi944
rapg55Obnrwwpt2gouatMvxqYJuZs5LE1Fk4+LzjHjLZX6094jasDQyPhBTMbEB7
yMeW2kqreUSsn6hjGEZOQ2ioL+InV5zkJzW47tPFwHMv154SMWrTp14yJTzraOyP
Eaii75t6voVcaUamzTVG80TYw84mK84Xj6MC1Onul9xLUcGdiM79v0cxKbnBsL0V
tbCDavcMMDMDr4Lhw4V+mPSRDqNSjzyHFDhBpcVaWBZP6MEK1Q8d+zGIOgfKd64Y
kQrrMyxPEgXEE20FF4pLqUeMJQK1i44DwzgXIqf0bxOw01JSlGUOu6Y5BYHWAV45
7nr6DOjgL86UdvGU1SAV6aaaaDjgokQQFAJkmQx/bjmv1xvzElGbKTo9/uKGRzDr
Toa3O+WShmONr44sRkMsbTT3DpQznpyoqf5UETndpPMQC75/UZf0cVbzaQbgccQb
AqB+WJFbid4mGNwkDSdtQos5aABVQQQSQiCS9hjLCx99qeH7rO9o+1sKtmoARrij
/qa9kCPtdHYdeEBCsJ8IkUW7/dIJzNMjdJ1ooGBg3hVY1pDKy0V3bRXUNvoWJ11/
rjoJhdT1fNAfptkfXtRGeJH1E60+NgTrVxeGUApNPlmg61C3l/9kJ/ULqzNVVLyr
TajSA47TMtgphWGo64jbbaKIvL5Vq5ezmEUj4VzgV1dy464nq0ALwmN9yuZ+0f7T
lfB8CAv9QrMaVu9lBI1GbEmByNirPClDt7jOvzP3H1SEGPcdJKSdkx0a1wH2jBdg
gXAXzrE/l1pz7EebYp+2vHCFa2mtP4aHXfQZDhvqKEcq3afEUKFOdDTiZbJjSQ2j
GWTedEdArE+z2+2HK0IvzDY92fez5YXWyXANxc0vpWvTm5cemRvz7xHUg1PAzROS
Iga05RZerBZIFIxBss8KZ6M5ma+YnycT/ClzWDGaHZiRlw2FmHaEQiW8ztNsUbDp
HTJI2/eL9bf6/OfC1j5OLzBFSJQrVmQlHnqZtMybFswkeVlXAZzk/RhEyxvsXKzC
kBZZ97fPZrt+Tz8AJ/mLKRkpLyhxShx4ZF2TvMfLXnYeCzVjuXpLIhk6rMcjwEpq
Z+brqouXOjnBktSN7GsYTUW2CQC08b8R6O1X2kAAvxCwKuVP+TCkBqK2aiX4IbwC
7zc9VVimZb2P1LVOqGy334nShcIF0qBynwqANrtIw89DM4o6nlNVK1B1ENyWuRxW
e7GukDHwAfadwwWfWQjrUvE5/V+i0tZT5z9xAjy+7dko1BBQxnYAlUIVPihhcnuG
6+Y5qhQ+kdNzxDvfL9fS0X8oL33JS6lybywG9sDH+N7/N0EJcjFhn6QmhA2Gj11+
r91F8XHprvqM0LJqBcHiaK/8QBA7oXPs882uZS1ybU0hfH2JbSFrcYWuJHrE69vy
iZMYZ/jhYik4ZSEcilQRmLv61EG7slBAlgG5/kWWAiptqBBUzwmtCc24K0BU+lFQ
jDmOYNgAmpX7SeHoPoyBubDPTagDB7ijk1U8QywABJrm5BuC4aNRyD11wG0FNNjd
4za8fg4VDwdw1HeHPMe9lhpzwKu2CdkN2D17fmDpGkFLxSvz49mITDwOlg0C0BvG
e7ZE0lxNOGG7GJ8EKT8aa1XHV+Ln0egAGRpibRYKbZmIIC6ecw+DkjbEFMH9w7bH
i0Cu+7rdRR8P0JoiYZ41ed28t1egr6WyVt7Lze1DXDqDbzAYVpq8uC9R3ptLICNT
OW1XZdVdGx5to6nJqKGFAl4geFTfrlzJH8PznPGGHp2zqKEgTXnFEDQH4ccSFWCX
Bc0QAxIPfvOaNb9+TtVLKznNBP9oWfeloL648uyo7uoj2KyyA3iS461rak1zNar2
VsnIIKoh3xC9YyPxaolyVPUfhSiVfOSgJt6k1BLA0/+G18/9G06r7dMFIf0k80BA
6cXElesfiTzljLOnbejSwO6uCCHzEpx/5MBQSx4do5zml5ZUF2wnV/CyCmS3+J05
P5wk8o7B4NcUd34/lVDINSwkMQ8IPRIKilu3DC5CwXFLTQlmZFMJHICQaQy1IQjW
sIEXdzP4BulOvV+F7MLux+Y6/YU3vTTht4+o2D3UJYD6LkkHCb2M2uDvycUBl8So
OOQnTSop0mUkbJNeDgq0oI2IWWHII6D/kDzUWAu0sq3IrIwoToj5P2kfPOrIU5ir
kXQqnbyMMTgiNdaPLcdKkx1y78T6UHBmml2Cup6wwe541j+Oun+j4vCBOFHEtogu
T5taSSvSPmQS0BuwPsDmSWuu/UurJwLR+/SYCUnTeGAMecWIan+z+1ehlak9jydo
5Y94RxxoLjj1pFuzyvyf4/DYR+F9FXLGwDM9N/jLv9jvpTvrEmCTtnEDpyvbZvlS
NkBKIHJkXMwotZiJhiUZstgC71SOV4Gbv9Dp9cerht2e64gWa7fgMEpUj/+nITEK
ZLDU7Nljv932OvkPfH7QUVQAN5aCOS8O/TS0vpT+j3JKtEpL0ap6qK1LDtZbvEgM
/QsFICg6HJjD+cbzTWQzyGyd2ytLCZ3OgJ8t6sIOk7iwLA+KPXrP/dDtXA3zuxBe
7yrKhHfy0ylc86sL0aLIeKnD9omL6vdWJOpOG62GRA6lpPrGCZs7MXz8S5lm3XhV
EhzJ1DilW0g6at1BFMPqfzWeYMKyOaVnxnwwYzkLVBEG+y3vL66ZVzcvW4cSPM5n
CRTJwH+2id8+Qw4szpdIaIgXBVfhB9J8GhQHMb9SMzGK20XvFxiyq3C+hg/J4Aau
17XXqg/OCZRfiODN5RGgjfko71zb+jnscTVvUAgkMyG7WKR3GsyK7ACMVFOFvzI+
kC/WUvfRZlCV90+poxa8DJAf8ut886nIc70auo+wLFl60HbB0vv/A4cAVCobH5GP
mvrhpOhbvhJout4uqjhQQTKg29aomJ/hB4WtkvjYieonMby/TUO0xtowl6Mu5yYR
9XVv+kz47VaXlDmptghX+TuKFsTmtYyzQAh2HKnmgUrh0PxRu/kxW0D76rJUnJJp
MVBsJ+lu79dk58ig7vOxFxHuMvfmxZ7rTovj/3uThYZVNxJsu00wv6AfDc7yPZSs
DJovIJMuyd8N1XTybGpldWSKRmVFEnkHQf5jim67TI4Zp2HaoQ2E2CoNX+tBaD2P
+n7h4w7Si3MWBRv3nifJ9mvcG9gHbpx8tmbE+XBxRG4mKLzB8WxeET0eQD48Fakm
g/UggHWWpqszCzHy5GHcTc2voY6O2NQ9d3AytBJDO16RaXvi6XvVg2Y4ZcZQ58le
nHczS4U/NV7uG3TImX3ZBjvU//1kV3ciE0tbn9xCGuL6fs4lrLV7PD1AgPtU5c0a
qpndUEuLel+cLcWrXo5px+wFHz2iK9e39elu1muXlmmscaTr2Jd6Ax77/vmm03yK
3jFCL9KWiaMzzn8dT9USc5pdj9DpJBm0UM3dYTni/q8E+F+EoFOAJ6eBlKD8vqVp
ubD3h059KReY7vlm/VV2zl/VSeT9C4hzlPp4QBTf0IzE4w5l8hBYgmYKyWICsxV+
YeIiIsYm4uD4Hp8UBCJoGv2El/fQwRvpyvF7M1NEqeWysUPlQndUbx4m12PRiUCW
Dy/Cih/MGzPFNpnsyxncWPZG4tGFfyXOOaqp/YgoKR5LkxF10ca6bjby/ym/G53Y
SZzT3x4IPCNaqt+5ec59xLttyGT83IsefgAcpqXO73DvRNDHKzUO8pTT/HU9UbCh
tK6iZub7raN8jcaCfGLOGsCl8F/Yvti5vH4RyUDrW2kr/AXlFY/xRkwsuM/mIkbL
cqOmijtQrmn1ZX+UmvMiBPyqr1Q18zIlu4/3BU+qPiJjtW2EJUgWDW7UDJ3NLIzw
w5XgdPTjKs3X9Iyv8H7a+zaY1RFUu4EXBnxD9AAJ/Hnz0mJDVBeyG0gmay9iOhLd
7Zhh7zBI4gYF5acdTkg5chteIuD+BLYk3od4OCm8uCL60akE9Iu8VYiWsrgrnLyx
0vyFBKeihE8aUKooOEjObiv+giQCYzetA6OApJFlmxhFgw5COzF1i8kWjFPRf4Wj
c/1YY77RhPQoaDiQa2yKB8AH1IAz9vReWcZc+R3flJT5dHZsjwDzKsK8csRVDBBO
0TL9/FOX5z8a42kzhdRC5yL/6qpdL6WkLmqZaNEHlNnqRJAecbukakrTQrR2IhtW
2DeCgGxQNZrZwuCAN0xM4s2QXR4Qr14oZ+sK4gV0XJaHJtBW2BDy8MM/pOj7SY3B
MlQuFrOwOg3Az+o0OYHdK1mLanR+tJgU4TFGLb6lA3HI33BQf98t0C+y+vwn0k3D
k0H3HtW9hSiIxtpfB05snRR+V8WgYSHTRtj2wQMvkcIyuTocSUu0bj7WTbOnU0kt
qCurDe25te+A9xt/97KmnZ/FhUyxnCupHAnrvYSLYiF9CqlTxxhURmOlC4phwsJO
cfZ15UlusuW2n15wVz7ZDOkcvcPiCwdoDXBNj4VQPYsnES4tu+uKW9adt37qUUz+
KwBf7om8Zv64uvbj1p7SJX/cH0OGTqREvgEIKHVW0JWQuZMWFwsDdClLifgHQErG
Q0pPfsthdhbFeL+yArPCVM/FhLeA6P4HbV1Q+grVV1iqnJWYs4OWQ57/tud0tR8s
gaJKZ92KiOYnnnK4IBYKTs6sJRI83gQjKOW6dIWg3rU8e1UC+n29LRNfH2m0lepA
7WrZ+10ttmGj7KL/0C5EOwSLT799rBX5t6Rr2E7XtdnQQxXscRm5eypAdUpRmjdX
d/rE6A7Q7T84Ebrdm/jL3lr6Fb+sSEZFBu6Ig2N4wafpTiK3f4CPu6i12BpJPXDy
w6Ihc9et+0Vqa2A9+4+Poxd7ZQ05gyX2IxjaVG15uVx0QUSfdYoarM714yPxSBxw
80lflIKzh1OMps+ARH/D77d68avLWiKFLJwdWVNDi+7jUOqZJeDoGrJw7iTFXXs9
P3iUReNfFIfrtpauAF6wSYjTxMJS4PWU8Q2gQn0TTOF9IK7bqa621h38Ap/t7SSd
IWLH55ukuM/ReEqdiOkg+Y8JJAOVrHEdysFPigKQlBdiZhSe+sSNr2XMwvDnVNb8
2BdvjgJ2LPE6rvW4u31O4Ykf2TeBEXAT0+BTlmb4TbtviE6R9meT68B7/QjXqP4I
S5Wlic9g1QOK4bx9hGYwL48PhwFQE69PZtG5bTM0Sn9ohC9uzC/o3cqa/bm7CAag
AXhCalfRtdeWYEro6TFlmbhSkgTmluswg9VIWvA+bntpKlEaxa4X+RdHi9bMYqjP
UObgZkR7guJccTR3+tFgpUaiSTE2gTV6VGP2iby9WRSGEuQoM4SMA396eoGkq+1i
nupMR3QcCEUMhmDRor35vjaSS2GO+/3DDfxzYUXl847cJhs1UjKu+5RMg0RJSuoK
7CJxzgWxidU6jvNMduGdLyLTKCenXX/67kul2lvZWfKeaSxR90ERAY9nZJ9HXZ6p
R7fgBxjCnuKXtUp5b4ii0hl+k3IZzKJUAV+pZoUZMVZH9QWgV59bBHoMOhfzaliJ
cod3a782YZ2zrbIth7DiElWiXVLgCvVHcO1VNd9LDwjVA+1/lGfmuPtXBGSl7sMH
MlCFCyacGO/f6z0hi+2Jne17OEoRvlTAEYZd1MHTgpRFKcHzPNg2xbFEDQQUzcSN
XOrATSCdtvHTetkgNrlMplZ/sF4JDtdXKZKofCiOXtIhKgmTQUjsvC7idBuHcZVc
4MtIAZGIQaT33UdoWKCNpExZ8CdzgJH5QHevgadejT4PHdwQiivFlvxKE/U0UOsI
Uz0pltc1PVLMDCTp16ly2HAwOcFP8+krSCTW0iBqAaUROky+8issfle92Ui6Ztlx
deOURckblghtHaGkADXny7f8LhiR1mxvAjg0heZ+r3R41BPVXY4SmOv/H1n3LYZA
Ew8a+ZVavAZaWzLT9Mq8YL4wwgyv1TRk778XfvmjY8fkqLPofoZHY7hSFutWzMvG
CTgNxuNMFuADV2k4ojqAj9q71fcI0Qwivuf0gti3z9MXSYzAd3UlJUO3fbUbcHe9
P8IhLdxokR5EwUfcLZvmI3g9E6KUnpEolrk6L63mZQIY8S8l6bFw55dSC/lu87c9
plEDrhSzSAkiDVx0eIFxep4IdChP5m4l4JQaDlbXLG8w25+IEUMAlaIqVcBY8k68
+u4HnLk1UIAwzFTtyQ1Wk8D+P3ajlX0aDE7QrChxSw1SYqD0Vo5KZT1GAx9YYivB
7DfnBumyTRLdDQ9PlV9ELc4XCNpYCnisW1eebt/RwFwsUEVIz0IneoOobFS5oXqB
AYgRQNb6eubWuNLr6w2XtGRKigZuQ3bh3idUk6FbZ6lyW4ZYzz6ui7UKBjfmnMc8
vVKJdxxCUnbOY+BtBDQ/wAzYBp8OPQpSGYztclu+PKRe0vzjIEt/op6wd/9JzIaz
fSHWrdQA8Kw+a7g7V10wwW38ZhCceJ7uX8j+GXaXGMBtPk4tInspVGcZrOOZYZ3A
OjkHc5u2O6u8uzWsaAWzB987V+NgxtbzH05oI+wpmWmXkyg0vdmDst9ZyLCoywPL
HaRkzcgR/gVYTwhoWswyvjT/OeMn9mQZ7KhWnDjccGlpGopZwXgXls7dtYGw95LH
nZTuS+DaNZrCRa4JjlkMa2jBPLXOTXPsEzR1Xk2cEfEbKN/lgyAiYp6Y99gqcUnC
27FlPb5xxR0YyIuM9S6wdsg6TjuDiQx2CQQrCXPbVIx69vYh2VJY0SFv8GWQYmZn
vbXF+lv9k0iPdae0XOZ+VlsqDH86k7mOvpZQyqsYgvebwHU2B8vewaOrSQLuJvac
8vgStjTY+aPlZDRs62dgkPhfCdQ1f5diQdziTYSszsE2ttpv8zT/PNgQ3jnqvYNA
YR39V0q5A2jaiGPLV4oGxeVAtodIIVQe10JcXJxULi/m2vS2OnMBq1yeG7eWMSz/
yruDU7D7x3FNdW8/AISeEn+PlcycKMvSPMSnZkJqoKrdM4ZoPGE/8YMaLSD5Rra9
XpXvbwSqimGwEGWnw0iOWPf8qS2DtAiXkqyNNW6vOXDLgMNsFgwr3tJNkcMIBG19
CxuCJa5nDF1swPV0HYby4GuJFfFvKchWLbRBc5dSLRn17W5HqSDuqhQ3JVV2X4Nu
gfI375WMofT95uIM8Gv+vYreelcO2sF/TKCUnJOWm9Eo+TfL4MZvQ6h9g5FIpZ5M
vACOyvfNGQvCNNSWoxGoLexLO646r2CUg9LyS3k7C+L5xfDDtrbt230l8CC3f2PN
aVdT4UoqBuZJHGTRg/WwHTLuylZL5K6UbXzL0dVhF82vx4mtpTju4vlBth8yXJIO
4wtkLDNi+D69CRgdBvaMVOrQlSp8WM/+2ReZYSV1U79QwEJgAMFvL77xV6YEBaUT
pvfVWhqbJ4pHeD3/b1rkZFeDJlpH9UNlHCCcRfxejnPsH+k3g/9TZTvIJ/REmVR8
/vmYbIDW+XYCupdkrJeaztOsE1LLSfihUk2JqaS5jbItw0jEMYgToTv/JvHKxqZZ
JqZj+wgfY1d6PTC4/ybPoTdiBNQYckirRluFDDnDU4pe7Ky9yWfryFjMhthsbIa5
x4IbfV4NAyrCMRNAjGe83e9cVlWvLmPagv0lC4crTkcdo4oOS14ucMrZkDrRHBFv
6c8xKuBV6jx1srOqvtAsZOWMiCgy0dvFKlyK2Nv/gzWSq12uQ1R+M7AP4eWuJCLb
SkH3C4ef59PNtE7UG3+ApG7rmfPijqkh4EG29BWul0s+V9pC6kJS4ZUQI4cC1pzo
ANBfjQDJkVMmKdkDV8zBG+CL+9x8YeLa0zT34l3jd7cX2ThGe5MnLZpIeZJVidgV
NsQyNQCx7hq8Mbja0n843LE5KwQkY5Z1y5UAmnxzNn/yA62ofBUegimGXHoaqusd
7VqPUR4LhCWI36yowXo4/GUO11GbX9fY8T3DkPwsqSZSy6wyflpYRFWtH6vsBigj
aDpj5tMzQqkjCxW6QvVvSTX5VPYfhE93/PG6fXzritG7cv6hc2BQP8fA9+cnaVyY
Swc9Zps/z74qk5M8ZzBNdZLs6lKkqgB//GG3pCLLXk5OKy+oUPGxwu3QDXLWN4ch
1FikRZvCAcFKzyQW18ozd4daNeZQhxb16abrc7T94kkWa3FHxzWSJdYJ1uzCiEkF
2Sm+wcB11u5DqXvESWJ0VJVHLZBamxYsyTKh61/zbIrQHSfyTDrE/XNwyFEBd3xX
yzDPO+G9Pc75Jk4zySfmKVF4kDp5oqQJs3GYUWYxP1+ukS/k5/5uUuavjNoTU1FX
KVOXbXhE0+1mHaCidm6+hdbwmOkMs005y3IgyArHCcRmUEhuYGw53D1QDMY6QfzP
8VeMv7pEBfOO/t1+UA2suGqmCCU+/jsCzH5qvJ1KBRcIWsx8mXkYoJzf3KlHXFjt
9+JuOoxni+cKUbxlnm7/IdSrGfSkRoRnhxMshi3GEj33iR6P5GxFyS0OhwM+0OWq
k1EUEJ87iEUubI7jojuF0gq98IzJ2dE73zbszNFM5lsXSl29OBCM68xry2eBNq3N
vPvKEMU7ZEdKP9m2/4eUIiN+HZ8YVUptc57VqeKeRZ3cAKt3xyjytkFrpB8VXEUA
xlOJlDlWO/wiKA2KHK7nvhG7rIsH4vjsWjQW96AvBhrDNEPMT9BQru93BxsqbeDb
9QQ3z5v94i7EbqTnBCvaiqbUxqLk9oRjDRC7iX2KwxuwysSJZaismV2psSBDuLuG
nJx8I08EAidYDioQ25iDBqBW0IDqlDvIALAUMDrwW0RAsecR8Y0ynINg+ONvB2HL
CuLRPcU20Z0DqcoFugSjkQTe1byHxYS94qwv7M57DckYrn0XTUeOXjTr5nq+XnAn
pPbKXFfzugB78Rx42dHniyNMjn8iUYW1weZxX/9QRwNLiEjx0rCl5pUgL2wpHN1w
AhMSFcISZKX5fU+KVlSDbGnZR7gCLo4pl7l5lpnx1YialHIOdUZM7nq2NfMR+54R
uouSnRpNAxKnuzpkKTZdL4AQ9ML8QGFtNsAvwe+Q3WBvnDunnKJPN6ICbwxWb2y+
5Z7x6QLfXwVj79/lFIB46jrplA+bY2xcs9Xh1WBngCOrT7NdrZtcqXgHg4WbBKgN
y9RDIjw9zWncZa2WR53Q8ctGRBMpmg1agniw7+4Xd/ZelNQsYgO8C8mZrxU0AD75
LrRn0BXEGRTApvVxu0WkRvPqsqvoIIhvf1E7E0tngaMESO+7I7yk/66gFBois7tg
JO/nyMleqXE9fjmP0GMdiedFBWbPGT1MDw43QIudAAGEN2DUymdp7cavek3D3hq2
G+nA5Sue+p0yLvuscNwY1Hd+hXz6eaK0sr1W2i3Ah+vVsuMCW7V0oLKWZ2Uyju35
JX8qB/OAyvzhsdzQ+q7zWUMf+WN6bbfGrfy+FHeg9vTHCHp6oZeUSveWg4y8i8Lw
NvkrwW/llSLw2HyB8cdrIcR7/OcA1cD0GLeitIq2AADsgGMGZi05a+HpBJxegjra
r8qN8JB9493iTtibnq1A4khjWqxAgw7mZN7z0rM1AhcSZZCi65vRx/qGhM/VTXDZ
Mn4+3080DlJErz7/P8cdwWrkRwHapMxwJr/HKKac9QxoNFGXd9wV/wRsNg0YEW73
J//JIw6ELH8rYE5qHqGHhVVyz6AHw5C/sLVMI77IzVH1MJqLU0UaN6+TwNS/OHp1
SG6pvEnAu5mC5LHPb9gXscRbj2YU9dsWPestyxD1YyzXtS29JGz3NTO3IFw6lI7S
W5QwUhXwushvxKMTQEyj3ks8kanTFkmWpwiiT0duUvya413GMNthTdklgIvCH6SM
GolGgqGbMUTR8+C73mYTtiBEcbHPGYOI3L81BmIDBzWxkH/t4s0VOVliwmtOhKLd
uKgRGjogQBVe0CWQJA6iwCKAeUhMt2NjyM8BUwonIEbOwTldrx5h7Ce8ds1EBO5+
rrImErp+tV6E/uZUlopPNurIr7+V+43F+CDrlBjIGfm+dA6KMU80KAaT8MqnEjDJ
sV32M0PbQJvpI+6JrY5/U8IUBo3yd44b2gn8krUKkErRXY9joQieAH6T7vY7jT0i
qMKrOMnrW3q9mf+V9mFHPvnJfwBE1JKQNz56q8wiOX8pQYnyL0aWfAffzEcWxP2T
uvBDHod7+wfe44tA8ZVbZ2m9U3H6SN+zlpcCJzzaWIHZlkR+pXwueRABwBX8Kfpn
VMVPRZKhvPch2t5GA5pgzTwiEq/9lAf8VVvDi/TPoQd6Zc2L382Raxsi/E3lPXpu
X23bdtGZdHqaoYFUIxGNO3IupzRmYF0aTMACdZfLbz890HzZbRjN2arQr1bGp1MQ
22E7/g5vngLP7ofSHROzHrqfJnlTMWjCJQ0Tl/bt6pwN9aQBfWUSSN24ImAUNY34
mvtIRS7SfYo5dIYF0AF5HaCwnF7DVinWfwaksdKyAVYL6+YaKn6S/prmyZfwOOZq
kkUqmnyGNy3eZQGhNR5oUtW05+G7mDmzI3QvIhrY4bWe8d260ZUKDrhA6+J4t5/2
lkMeXdOtj7ygdkGLqdfl22HKvj8fFSMBEp0lZHGisDUx/KYm8dsQSDfplqrZHHxa
421/M6RwgCzh+mjdlgMa1dZB6Oz7Q9CiYbyutslmJaP4wbLcVhez+12o2rLYmeSV
v0u+DIKEDxqc6EsjBtZ3B+1shQwZra2g96pkmfOctLl0CZbYoOiy3NpXaujHQNwy
fsNHXwwSGf8D0KYd+8JMnLXLaGy/rfEpdZCpcuFHYKGuKzGY2OJFM2Xtgqs+ft6c
K4ClqrUv53Y05xe0oQmAzA8y4X14rLiOQw1AQBC7mJRUvsyUpG6FNDHeBmEcQyZ8
9osYtwPBwQd+9SrK/AqfHVf3eek2nYPsDfFHHAxSIFZuyCS61/kIffMr+R6Ssxt7
7R0LzOfvGT+rCUCGo3nxZ5e8L44K7l9tcM40OtWObSdJRxjFp2vm9KJOoCvrU6/o
qR1MJ1sTj+DEtpW6CTsQbBtSecWt6nZ50GA0SsH+pcRp35j4T4rLqY8IvjwhvIq5
kjg+K0lTbq2eGRivO3v4TlX9iP3kHaRoJVnccxVqAjNHpUkJ4UOYrYnfgLWtkR4E
+Gy5albU5zkh3DryPZ9Iie8YhDAlIIfswAAXzx/INL4Vo6R7XNcc/WhgazrtW7p5
LEB6+9LRMRdbgK/Pwzy2/cDQTHg0cZ8UGmAeRM/hBZzzRYKx8gDdUIdw+TDROEAd
rUDXogwYB6M4mF9Im+wxRpy1UPbnZOx0/Z9RzkYmtSdmOw+lOguPPcU+XOdLUN17
D++Xue1RzsHpOQVwOmr+FhYXirTd6F49aaJ8JBOqFyFdOlGyDpYuU94fCNL9vYGD
MUpAgH4v/i9U1WlB3Xq38tzSvQYTq8GBMqZlX18gVXuyXfdYlI4UnjC7T/F7MqGM
ANXTq+7v8V4dF2XCq6zS4bfrjboDLHop+a4Rb+2Tqq04Fpu3gBhxdJ+pNrJ/1TRn
c6Prq7zT9/zqwnvyp/tUJXZL1M2JYx+IA64d07YC2Sst+/nSqtt4NViIEVliaSGi
pWO7EmlrsF/cK7nhFriSL9Bt/H8p/+E9Ozdti98yZw+Nmq7h/We+nrFZOK+LRMKx
mEtQCP6WQAVuc9M8Ne4j+5AGFuJY0lqtvlJkCRzLrwYNPrc22MN2TiRYl7xJROP6
XWYpKXhkmnAEgnAl8GGMRPViV5Nftt9wXY4HVp4iBYdisDmdHIx3JD/RCLxh/cmq
Hw9UZGDCibJwDYhpi1dVJKFkzAYDWvMOZ4ruFEhuFaBUYSHcnsIwUcPNmFib54Yb
PFmhLcmuCzcUrIO7MnaOB66SCKb+tYjNV/1aE8QDb08EtlvzqNxbWN9FXjTFZaty
OSPk4FzmDbpvyFq4h4NXYYHwqYwxbhelQT+j5z4C8NU3t5XJABjlDZfNTKy25B5g
1ZjJDd4eFJiW3F21VFrhm4e9D++wjM2QanQY9Kp0gc9NkSUkl8LxxS0PwatirWEY
vdnAwVqFGd2Zqn8xfD4Jf0SdObN+bDqFiLykK4JqV2Uw4PP8MsTSIj32nPkfU0sd
cjyW0Ys8RwZa2jM/K28z8smDH+fRtwV1F/3O2EQmUJ12kBJmMUbEjSyTa+mUErj4
zgi2bbUCKgkC+Ts8PA9hUWCfeRDCaVadDh/nMwS5QE5Zn2JQ2bbY8cXpNlRw40NG
qWstMLjfF3B1T00OMCGTHGtVrjKVEH0OPKGSwVavlEUIPmmRFzBNahlHoJPP//X9
GNYZtlj49y06Ss7NmF12e05CVZVc/4mTPBYfFlDY2pmR/tFTONEl+ILhcfm3c6IK
5rchFlqWBryVkw+gg1fj+S7aOGsrjimZdLPv7eVtyr6gKs2SVcDEIe/2qNXRf/3h
cd/Rk1ECYrqO5OAPIm9+Qb3Wig9LxFgvK89d9XImzP0WN2Fa6rjnhUSt/0zdRv7C
cgkI9EnjvMGY+p9aqsGB7mOKeuB6N85dtO61WFasycorJKZnSm45dPOhxbIyGPWl
YTH9BPG5tqJDi0XVSMlfTiINm6Z6vi9IWuvoEBA59zwlbKoLzKG0THQyYfKhQmlP
Qz+0gxoD5YAMEHD858JQbCKJ5zNQ0Q0kBvd0AWG2N/50x/c4y60ukHLH0ExUwSb2
RhUgtWJgEjT+6Z5qC+iLfgrgkSSdIVxp1taa0uKdgk7hxtW2qLaO8LCjTRkOzox8
UGlbeii/x2WzuE+L7oGfsTcfrFp/imuqQdiDW8j8mw15iOtAVxOPBuxp158pg0Dq
F22HSX7dElDw15hGJz7ODG7J7otrn0+/ffkwVMrY8QkTdZW4DKT46v95cwvq5Hv+
zGicl0nuwxtz6jF+E/xpRm8IoAYE/ybLfO/Xi2HFVM3P6uslGA2YPf/jUg0Noe3h
95tBEIHNRRVfBf9A9/IrzWKwsdFMfxIKAS3GlxLJDldWhoJg1GHVTJaegjCWEGEr
mV39MEejSc4t0yTmtgzd0RfJw8lZZWNSQeBovOYk3sBdgKL/Rhvzn8CUvvsZFJRC
eQv0osloRmyEXYl1Cxmfj5JiDZxlIlG+avmc7aLAwYPqwhoQh8GR1CoWZebIXH7P
2mfTD7aZqy2TV4DE0NTSTsggkLNZISlwm4ZZ+mDG8hrlgb20GXX6kUkZgbGDYZMf
gCnhLm9x/Rio+GvuJsSxg6KVmhygHLzDHuMPHFTUj8oTvCuZEIxXGcIs8+NW9yqE
6HHaHm+XYJseB/VPYh0IjBvO3pW+q6AGzSsmM6POcjpe6xtunp+qq3D8FP4g5gck
fvAnjFlU8CI8HGEKo6TQ4DrK6216tXSIcNpNLTsF7ddFa1GPYNal3h1/DB3Px3Bp
XWFsqLsF0OCc/yqjKmJNiG1imDZams/X89bi8ycvcOrEAj5UDCqkvEdUZVtVhXER
lSi1b6R9u6doHzz4LsJUxPEKEwR3P4NrAHGYNeUWaMLH2vs7IZx74LdLGbgA3HRh
HuNEAbIvsomwLDE+Tx5vzdqOBD2C+lZBdbMsvGSRaFGtCxugxCzcZ5G0tSAo4j76
YQ10vjWLL/C0Iao+V6Yijzrtply+2/vg5mnw+b2odBATQ4FkXoL2b114sGxVDhQy
FU2obnExh4n+wz0OmaDvR/EORF2drQVsQWPerWTBzb3iwAP85vpWUBdQfHQ8NHXS
o3v6WMQq7hWnQ8ba/z7aNzyODv3HxFH2efhQnm2hF0OB+yFd1DGqjOUdN/Ct9UkX
AVlHUbY/ufeMIsLoht8X7kIEQOS0zxM/prgZljvmYkg0c8aVDUBhoeLayo+OS0DL
puxoheFR3ynOXibFdWPcbSfIz0dI5cZvXtd2UGAPjPnUOTezuzvCMmYzR0KVcqW6
Jnc7//iRq4oLEc3fBtH+Tg8CNKg/rtjiNKPKVAwYTx4ig9Uru4Qdf3WgY6rUO51Q
tAt3IgWcS02JRHDYjexhQ/S7fWQS8I0RPfvVw2JtwLse9fcFa6T4ZBI1M2EAUDje
qkqTOd9Qjkjeg5axJzq1S7T0NH8tRaP2nqobivGGN0vRcclf8NS6OmZbTaVAChrB
1VCRca8L8KLAHdQEICxwNWUP/VImSjy7zhc471uxg0OnfTnIh9l2HJqv7cM6p91y
CzU0HuQXRG+x6/WsIhU8EI+xpkvGorMo6Hr+yLcz9B11UyyUdspR/0mlLaGHKjQG
E8wv+BfWK3SXkCvLRWwyTZL/6hV0Iqp4va+b0VYSYFqKC2ZZV3QEUJJ0HjY7KQoU
vb9aSVC3cDpE3okgTd5AT/ouf907CFHewmResHeKhN5sDXQehkGY2OuwQmujXpYQ
PaYZ144pXeTvNL+b5Ev1rt/1sWQ8AZA/rrHQH/tHhTp3/zPy3htGSgRWysZeaBdS
4igrtEQIfmPpKVCF2YhhtiiqU0+9s3JVI/M6GKm9TW6xt1zO1eP2jTDzYbK3NEs7
ySedeGufN0/W+TnOtxbeKIb2QgGEC3BvSz4+WKdSQRMQFe9IoZIJhlAFA925oVLk
KQnzZGUF2rF5nytGCeAu51PM5KO0npdmjwrpECDuok6ayEzgYc5+l+vbQW483VkH
0ACY5yKuweqUw3LuCLogFY4HBEJUz19/DSsSl2FUPYuRE2lMoOe9ZnHnjYfdFfb4
S4mh6Yf3WfqwDyFqIUwA4KsJ1hq6W7F6T5gevKkZ1v8+JJJnUAjuc0F5n7FjYk4A
gp6mhgzdjcwt67ABeF7Xh8ruaBS/etmyb977HsyqdUBpnhgFdDaI3EFkyo3R/I6w
RYw9kHh/XLfjnSwRm8CfGJ7xnZxi8lF/eQMn1Eo5Qk6mboP2ilgBxX0Y1VHStKoG
AOzu9ZNO0dqp1LqWmKMhWtYkVIj24cfVanit0FgMjtG/DRm5tjByTxEdjSIABpfs
DWDk/Nv2LKIYuvye0z0WETGdquZUHwqywLFLY3e7PPMNd2h3PPAOq8H/a2ZpGvgm
LxdNte8H+QKIxoojS2ThWe0CaFg6J5Bx5EKe7jAi8b3Ukvp3UKeYiTrBaNLKTXRy
HTcirkAW5RjgDZd50Pe/DSFwhnS5Vtw6hqbPfWZy+jXmySX5jUtYG3w43K3XHFPz
6BAcIuQCGX6DEHZApJ6sOdwfZEdm9TYTwtqbsW4YvjLf+BcvdujFYMb3PphruTn7
AWU90oO2zDUgMCNhRFpHYd+kDrGlDtmcY0u7dTeCIt7UVDdnkEtbiunoVsCEk8YT
/UszesJ2g/pRiyIe9s3NBrKueu8D7uunCZNyrKH7AKzluf+TLRU8SJh5y7ukYrlN
9ddjUYnJ/GCcXLN1UpuQSSbXZUhfE5LGQOI0NCZ9QbQaQ28gRYE0I2Mx3pllYGvP
NhptFyZc/5mvpcD4Owo6colix8esgnKDuAFoBsJ8korU7Q/RgLPaMwDyXSPJOCyc
VDrWGfwRvuWhThmm/sgnxfXgXgUnCWZQ6Vq+XplB0vm8HC3uMxWceM10Xe61sm2W
44CGqh8MXOEvaAtbC3uJzYsCI7R0ccqZhWcO1kjlrwxfLJfDlQ9De6ZvmuFoHw2B
0P0qs86RdAoPXok+8soze1jdasf+rexe4+NmFeZR+AOrZTcHJchviumVDFDKO1Cb
1aADlRrm7bm3SewiYXHs1NR1Ialu6sWJHg4t455JIxuiH2rzYkvaEkGoVG/eQGbz
6No2vocHoOmIzw9Cnejof05gEzAgh1fgBWnCn0sFe/JLrUUoeZLhr76vnmfdN2sZ
grf265Nu4dofGDJnJ4yzahGKj+jxC+QtHomtcnw6LDkxCTTcg7W+UKdZKKGThFVI
s604Y5TbZIWdNe8IVmg2MrkfB/v2c9lVpzMC6qL79OquDGfW1oF5x2TSlsvkxLlJ
RGzteB39Og6XAXmvg1cfo9pXtnIFkBFrEy9Wdh25+XOzDj5CBkdYZhbkdY9MWFb/
ehpiRjXVEejsnwYoBI5OX4w7X867pwMyJbTNtAo984mA4ByGp92R0CSOTTUZbTk8
DQwfXn9Zot0RSx+Kr3irIOCy0lrIF4AB2LRutctrgnC/ZMYTjzDR54TGQrVdZlk7
MjUDoOrzWy4ofrvA1cl8irc+LFlksBPtsjoIm0h0fanDurfwRcSsgNu53mvd4Q8C
ODkQ3AvXy9hr1kGEHMRsL8B6V/IvxEWSNt2vzbx6VFpJbQ/bQzYNAgMqOGhhmrS1
Q4EVKagjWWP0Llg81XcnsL+uCxJ/K3A8h+txPV7AYcpz7KrJnQ7oAxcbcQCreQbL
VB6YNElcwwwepGzrz4VhIjjzKlsjxUvzEa0lRA6VYRccv8joKXG0We9vShg+3Osc
YQNh54ikm74pQnRPv9h44YJSDd7tDtV0ZkWZSwK1o6heBVgnA59pGpclfxuhJTVi
21IbzHfdrsAo3w4//evqHmxEMeROltozZhICAOsNgEjNSKNqyl9dJNvoFkj0neWE
Xj2vFh9BKkCXlB/omtSbd2TkMJE1jQRn80q/wVZwEf7x4guoGfMTkpBFllDm6YKq
Y6gXGDrzOyTW8blMybVAyJs+H0Na87KylbSnrWER8BHmpPqRc/aivKro0bvDG5dm
PbWwdJkVsGDMOtoA4H1LH7WVRxlPEP/oSwBwOSngDX9pBzMWGJCi74QohP7fc9K1
KEE1IoC5EV/sy2aq6UhEx4NbPYnm/nRW0KIwQv8E5otVAQ2koMe6rNMbEpqtNsDw
XFKZmzrZOzc0oRcZGd14oYbpcGDCPO97GSzzZf9+2LDFPb34quBdjSLJ8IzVd3b2
YYadZex8bbnRb0pxXraQ2/dLZyuAH+V7vgts/x40YJ7wCqVMaQaL77/v4MCuDk6g
2eS1SLK4esAuAczNZ+1z02bRnC24NJu1hH32BiWTC3+/N0PcJNbO1LLLeNNkxdvz
RUhrOkG2JX6MwEkY3vBLOzLzqnhTDoaA4K1ct+orajZUSS0c7rfAvRalcKtELxX0
1axwGQ4l7QWA6BCG/43rOGtpi0+6JdRdCOqfxqkNC0XTzERMpcPPLzMsYTspHg0B
cNKNJfecvC4YAAdkWtS0NCoZp/KFBa312Ox14O5/U9uUcyixhvgViaQcaDZpBabS
NY4y+i/GE8FiOOcufeRB8eNPV5+hZv6DiLBFTOmvd7g4cZBURQ3AoKmNEc4jprgE
RqGWl+rYfU0QbJwlfK5A5U6hYfVG4w4mBscYMskEkd89UnPjk5CqodbLOx9piVZ/
+S8ihmC8omoQYhNQpEVOkQVx81RbqHz22+2Uf13XHYj70hWElXRvgW++WWzORlRV
p7GFspu2LAUVaOge9wya4/rGZ30fFF8t9oQTjQTCYHzFR8Rkd6VV3gk5/LcELv0u
f5+wqEmX5+9xYUuBsNz6sNx91sq+dQC26iB+tOb/V9DFwlcepSXtb+fQRv4SIP4L
vgfIpKoXOfdyq1zKx4ioB+Y5EiuC7E4g5tZvNae6LZBtQffKW29faoxS3ANx7IPW
h2K3zg8NfvIOvVEKUFjCiIOXRj9VVRMdyvRTnfQsdEzWJ/zEXJGVV8olasSFoRZl
cJjfcPDU1QMNPC5JnJsKVShnkXZLqBDW0Ln/qWGA9Ygczi5ypqui1drimbNK6QFZ
unjx0MhAf+9Bvu+vXs6ZXKXvtuiAckxRkSDnlgyGiWfbZIiGkhdOGOyAliWpB8Tr
2z5/OX5WVZUwfWsnWD13GMalKrjAgiMqICSCrmcwRATrhOrv2vDHs+6oLkBy2iTl
TI2XMHskBAux7LsS0azDdkOEd0YibUUpiz6Kuj5HzMuIIrWOnuicwtjJpvwJFui2
drGGTi0olZnh6oBnkbFlUimkABJvkPPIyKDmLfBsfDsNFU/NaR5EH5Mra8jJpVWd
vFUCybaxXGryViti+Xg3/KZ0avVLeSCOJnc7z9AYdv5ccMIzy5lyKkd/YLWt5BhO
gR7VWeyND9m1wjEQmNE2PXaI7DLvoqqBIdok0ZwSYkXY01Kuc7xR1tDdjam/xekq
RcVh01ywHET/Xk7jIWyZyi5fYOAq1ttLqF8/ENdNukYMoAcC3PNydu84Lc6ZZLUH
zNnn4AQv8++uICpcZ3i20YlXrMKK4P7kSTxTf9KK5SaiU2WNy86TdOtpZV8jGYEh
aQ64Z56UVFWuqQUEXzytuKNvrxzbhAFIMQJtI9fnIkv8K/MbVlT7wkEGuLXsxaPr
QDLUZzb20I86U5vMGfgct6AVDlqWHpcXy5lyvE2I1iMcymeHH3vcFwlRIRNHVTWj
Aw97jqKnQkvYuFLJYViSwAVhNQEU94bXs26XcPVaCucSaN6SmTF5d+YGxpt1tu+c
Rhan4Vs1+ATl+A5oouAVS7I4QyBfu4eGPLADY1n0D/MtNAaQTfM274QkDq2wZSox
fpgbWS3Sk/f8psPGpdCIWGpcgMyL08gyBwxJQcVMBCIBU7SoKe8NUOnPez8n8sMS
jD+jwhrrOjmMc2cm5wAC93sgG7cmwAi5PgmA79YPuOwfbB2WstzjR1JXJlyP1zdJ
hoJluFihD9u/izGr8EzfT6CMOhRzPUdmiZckxcMKWgXi27oz+d/l2T1JBmGcxpUT
xZKmIX1zxZMOAqNXS0QmCNH8YoS/B5yrMgP+FJSK/pX3AlLrSvGhKng6nz2vsrfm
RaNqNRSumFfteuVlEX3hipjVvQLRu0++pTqdzUwUHf+jlHyboutq+WP8jUZUk1wD
G13ULjfqOR22OU/HQR1taD4GURpcpSb5mIcGCxXFprJi2aciGh5ABrTs1aYjB91X
/EzM7Hn3P0+h6A4x9JARD5I86XCExcFe1lHiee0rbCvRyzx1jIIaMqgiC9WGWB11
1BjuBlpwJml5UJP4xWkjkyYe21fpdRh/0X8JpNTdDGDtX4+xGtGEX7OlsDWskY1+
CZ81nq5guxOJC/gYThmY5RuolK0Qod6gVc6Pu9LnymbPOuq/YgShaCov0HtACHoE
RFRhBmOspLTeoa3lycfTtXWl/VWEMuUXSjZLer82SIp2+W6REqxg9H0/+7YzG30s
jqlL7hHKy46OxUVw7uc4csW0wkhlXA/PmRvxxl9DEJVMX/jrQbduueddGGGh+SUK
B4FnunLzcY2IBP5ea3XOlteCewgX/sb36P2n1M36HjFcZJstjPL37dZdySZAdtBM
f9zjDfUE86iV/hD8WQgwc+EoM8TfMVKWsqKso3RTRE/hY5Tzl1OfR1wDvtBwVEA8
UpR85lchm3frX261AW/vQ0qtQmtj26prCtTyAqdZ3NSlc979Pu7kh0sCHp2+n7cr
wx0tL2kFTQAlH8vzvFkpd+jU3qya+bmmwSDPg6rBkwMDC9rrhL7po+6s4vSvruXs
jL0XISYX+ZoHxskSFtvIptqJbZ5dsDSdEXtuS6jK65YTvjnnHAHfjpsOBhKUPFzb
nj1k2eLXhNP/ODuzHBeTZ7uhiSwlgT7EejBTf++mUYbI3CRtebuon2b573Pa3K6o
FWo4Tm0HTsha3ulLSWjOk20hf6vRdZH9wzKK/LhUOf1qYIXfNQLtERXV29ftSfQk
T2vXkc6sGwOIOuOP9G9uPQxbuCDcUKtmsQSPWNsDl9BhFkaos/ysq0Wpo+2xbHJD
Wdrq/ujEfCBlQs1Mw3NvSphrXYgaPABy+Yx6X8t/St3EJQpLhyqPIsvfFsw3RLIm
1fxS7i6jLCv9Hw1eAe0Aqzbd2oBM3Dilpr6fbeyvBAN+Xwza0hLq9GSzGxCfvbHS
/BORK26lTE3/KCe1pJMBozmRZXFCZgg0Zx5MYdWKW+/9dThmdc/pK0onDsIs9w81
17VbPUzEthsRORltaz27RzKqsFuKIonDOfja0qWRTSmC66ur4iSai4EAzAvmJAo3
jy5poekbQfgXFV5hHbzYZ+jUeFcRzRi7pqpDieDNT0FrwZpPwk2LqncofM4xDnEB
wmK1czUqM1ycu0608QxQMRi4O3mKMzsPJ0tyjLwj4ZYOfETYIaGH9/akLTzc9rcY
iP+ofooJZssf1m3y+aG7Q59GA8ncSKTkZPMd3OwYFL7XjMhAqeN4AFbLG8WxBWCQ
5+bL+EJZfq9O0Cudin/irLezpkcF6nBUe1n763m+yuFBGjD2Qs9PjFcRrUaEc5nA
GmKvYFHIhF6/JQSLIH41P0mopnTGKHRHtJGc5SMyi/xDURqtdybrw0vzkLf9JGq2
R6UtVlyOPkPqFz2nDKHrvb8rylhWQIxoxTjvg2/fFUCK0prQWEQ55itHRkTkGMsI
A12vQWXDhwfJgKz9B+aC36qWdvoYvZTNExQgC81xJWfpgBgL+rg7Wi5RU8bis3lR
FTHqC3EngWi8zDpYeGtdu8nDRCIra5phAnJcIEdN2E4nXnCgANrLOCLgHMy35Eji
rw39viMOwddVjuMrSG1WzloK57wuSD3fPJEkbnqZb9uL2BWUNWbieNcuxWxAGmo3
MNTkie/FD1mahD7wdJ7uN61dd/rg9pNFCbBedmPZI/fSXeCihTGBxiBIAdlSDK8o
x3SElgyor8Fev2iKlPqlbBuHxPFSjXw5qytbvlqWz26UoynMOUegwbla//4ZlxGI
n/x3zHBiYCx6YVY8zBJ+Ga0iBvbPkYCchhty92n89NEEVEag48WfS3GouEaHyihB
CuZsc4BE2fvHufLjzTew5f/euFYHFTz3jvxQgbzXYEnSTAcpVaHuycwrZidvZhNS
JSGWh4BebaUKnQ2jcpuu5LJ5JWmbVR9uzCx5R9tHFXE+GeJXXoG1eAjcVX8+iPpP
JaPB077oNXDpbIdqwdSXwZ4oQUj9kT/bzcpixlXZEgtaeUXjJXnDtZhXjm2SslDE
hk7NkDiqRadMMNqaV+IAbLtzHBatBmUNQgX8h+oIBiqIvP/Yf39ba645bS/tJeIu
TcQhnAHwrjCNYuUD2S8EzJZ8YTVM/fDNH8Wiid5q0MJf5RMCMbxs3/83k6nr8HMP
yfaEspMDMTwdZI6/kdEGjZOLyqKPL59eST2eg3YT3pOcERfSI30+erNwAlO9LEPG
q0NzjLokhUhGHlLfcUrRVUkzb+YlIGcNNX+lezJESfy1BfMXiJLw/Ex3Ovz0bevx
F5OXU/HEVWKFNQR7jx7f/+mQV5ulwo2mI8Q2VHD6xmtZmj7JxV3egt3OCgAQ3uIR
jfsWvHxLKoGuDvEWQOCxkiL7wFmZUZ1UN/jYTnPumOfj9hb/Ql2V+tC7jIzyWG/W
XchXl8JDzyxOj5RI1MwqtxPg6RJkh9tKXbQ6LsWzUaATQ4rscGtuHzc3zCvi7AUK
xfMhxTBPNY3rlrXLsmbD1eJ5aTzLboYhLEHOaSad4AKP4lO7M+L80/jFPo/Tq+hZ
DRpLy7Y7ZzVcHhtDp6PnN4x6BzkDlZhwpczaKe9snwI37NOci6UNHthqwDSBg1JE
L2uSVoCEHUuaDlN6h1wXSMGcBGNCU9P7Zxri6qgS63dmNmVy1UrgnWF4QCLB/mIX
6200vqDUMBfSJ/Ho+oaMUq+3IWEzK17FsMSXm5V/oxBVMGDOrOkUQvzPrkjWMf19
uo5/fiDoJD5M8itlh04UC5qFlsifJZT6JvnTz08d3M4/5iLGwUVzGAhFSf8kLMN5
L6JCC/O2g8T7ZYVG3An6XehUm1OjBGglDE/481uaNgMqsxoq/32ei3i2hvPngFFQ
yImz3SQQKcyUAWNCBEdaroIxAeK4y6IVpFo0BWwdH6TihZ0ORm3/Ysm8abRaP2ZH
g70egGEvSD454vpKkiV85qx3KZePZpeF4b4engQlA8hNFdDm+Sp58XkMeWRthYXG
zlIOAqt6ouFYgznZeBe/cBCiFxOvbjMkx0yhVgB85NjrDq9xiQx6ZtnE50RV6dq/
QO0kUDp3bYHV+nlCwUM843K10Wku5nnsZXNeJkKPJpr1usmrqOby9aU3QeZYqtsb
gEdjv4wBMlo+mOME4u5ftzbhkanMMmVV1emhCC0Zz69+lHulpNbURIbCezQfNcHD
WrGpAJK8Orl8rpuRiwljPFfWmfJ395pMzmAUtU9GVaNSXgfZ7OqjZHftfMD8jKLW
2aymtnxf3XPjwwcE/pzfsT7O8/F+G848XvLfk9wp/mqbrcdUthbq0nJAuxSYwNmI
WuZC14spKikuEXE1cAUwFQ9ZujBEyC3K2121Ris187SsLXwJVKcQZXWny/7eIUuL
KrhriUjSZd0SkGmCnVRzKJ04UmJ8GVD2c4mWVqCJ23AyiwOmlZzRM5yfQLWd2Hnc
qiBmFn41FwKWONL6ehGV4dZ1CjUcBw7M/HF2Z61SuG30MQ50Ggn5bWxTjsirN7o+
1r7bHbQy12PvFeT/81ZP5znSfRy38xEXr7t13UlJ2+gT1mNZW+xtuQvcDCcwVgeO
w0ADFSYXehl5B2LGGxrMFabRKrArsjJBAZcZFTFuGglyr0UDTfIb8kqMhLAA1SvW
KH7aVSbA8LNQXBr63bl1u5MD1hiRKLVyYLb91y+BXuInED8nvGXV6hptwz6G+agw
67mFTFmGT2hEsz0VBgSC1m+MB29GnxPHEaHlf/WqR+WN+rnmnuAywHlp/7zPBFks
nDzQOPQ16l6LbnKmy5fH7SHWJNOFwwvUPL9PRaU5P190+yvBj1Yd8izzXoae05kC
cSwUrQAx9ijpjPbB+F/x/QGCnGfPu+1mY1ir1C47wvNhrQ20PV28sg2n+MpSSkGL
dw09uUgSBan3mLZzZVXlqOxd/zLILP4tH+31G3SlxZJm6AdbRL+alXfCkz6wIbT7
xEcBybe8JhxnLpswi4gDAAaUrJDJQQz4y5mUCQ37/RRMpmqPLqB4ruiNyGWrHrHj
5eIEah/rEBPXuIV9Y9/RLpSCLA28SpuGF5RT2JKkRbyKPNKUIhSfONnr5Nvvm3nU
byFWvP4IcAlfdIx35n7PVG14TZk+kkcR7obwvcUnyf3LO5BkU9C3T2rDIHigocTp
N9lKKxbqPmX0o9sll/twpZoPmjBQYYlBsm3v6yAFJ5HWBZrlmvJhXtImk0W1H8TY
JgL6LZahBU88ti5+1YCM0Lp/+sRNKluMXKijylO+Dx37eEC0f5jUvyBA8oIyrUWm
hzvTD3tHqOpwsc1YNqkFXRjrLJakwnqBLAkiTvkgTxbwctngxuRLppusS0ErUzxd
uMO77kWKU4VBD40xnQc3eEvK+5qlWhAmnkb4NGRamo70iXrv5ixkQDUVWyKIYO9d
H3HMggxhdRyKO1jr8ooarxRGJfBiEpyy0BC/LXQ+jK1U0pRNG/KlBpGn018fbB+2
QZwZeBq88V/PFh2IsDvUytuRrwJhghM7ocT3Q5gLnvZNBjJMcTILAhiY5jH0N2f9
0l+Tb/e+ERmoFOe9zWKr6WXGO7awrjelIUIBAnu/cQHKGZlZiMO0BJzVpKzKXQ4V
mzS5dF0HFs8S/ZSznDxmkqCxcD41Pmge9JUrrm7RnAiVBwi1nUquLzoQtQclsbyd
Sdzng4KWzLroEhdqcHiO0qyncFDqfwk3Bb7lEASNg87vKBaoNSSKzvEmPmFzkD8T
wQpf5nkJTBdu6Ug1c/Bdusy3ud0Uz1QXLkFkOdOXfczjxk0rTqFje9gjtW7SRxJp
kU/BJSPO0NOTij/bu6YFAd0BSEmLCvNjD7nEmxoBurN2ln2TRAx9DzPMdp9du7ir
PavfaRxD/8XKPz8EnpoqfAzCkQUCHleT4snzoRk1KjuYogRy/RVmrJuEMArhpC/U
xrof7FZayuLISXm9yqaZHy7fk33j65+VgQu1hs7hsFfRME0kZbk/ncuW62LAuzsW
cNAMsL36iI6nJNE+7VnKb2oU84HTJEFXg7nya4x+KpiF9j9i1g+xhBXSeqPQlTVh
QNaYUcKNoychS4RCWMOvXsdjmKejGbg2Gu+SjObvBRXRBlV6+xPbQYrflf5uaSFI
0qQH82HzPcAgPWGqG1FdSdDNjrg6lCYuP2VZbQ0olwEz/MdMwcHakPJB5Mrmgc9R
m68QhCFHKv3E8E0a1ostVz4I2grXaBy7fSnKvl9aN0CCQOHRfLTb1tLIn97OZ9jP
ZfcvlAC751PK6YkqBnKM9w+BtoX0yvs+TygxPDQ0AhI0Vanpyb7Dl3o/qgcmKEkH
iuD6ChFTWJanYrmULvQAB+qooSQXdD1scZ2934m7/112tz0YvqrZT7KpBfWz78kL
SCBxYrUOa0/gYmcnjgENCTauUY8g/5x0crMEnw7qc2rH7y5WJX+jZ2BxQRYLyGB8
T8S5Ep1gFtapsScfFMogXaYipObuNy/kQZofzTyocnx7WXKfwWue5+Bx+v/Adp0w
HMmFkKXTb2ZuSsWI0EVMrZTjQyXcX6evBV5DGkNnGFGsPxXHGaO14a5HS0OFceDy
ztsfoXByp2NwG+ldZWx9IFyJxY59Z0HpuoWSaEfExxVhQuCmukXcyvnnjlrsuCDO
5TRy7XpFfHp874al/nVrOS0Cw6GrGKT8odtEjHfqpIal8MRj8UeFX+AzDPLfQH0G
0eYUIJjILRSDJy9J8IZH1KRvK+Mp2cuw/RPI4fmmMIJ8yRWmVh7KW4BjmHb/V2Cs
BNyrhuwcuPP13nNRxV33DNhjAtR3yWtAmz9214GyzHqRevTv6+2PIpX107gUS5cZ
o8AYe049nwfBpJTyS8sbtQuF9pX9FwNp++3sXFzBCGvOyghWcUa191fPzsU1hI12
lspF08wRxRcQ2MReDT++92FITWDRc2QHCxI5XhtNX8M7MltgGcvmIg4i57Cg5drg
squ+dIlyXLRXnYfbAMUZoHCw7xmMeDwlXQT9oBMIQZ0mA48ceiBRnfnrByItlqqA
8Dwu1dDIt5jI9cfDbTStFv4DBGM+VlWxQ8ajvO4cxkNTg+2HYmOgCTYZhcSdRDkv
9+IkzUigxsqB+1qVd6rE2Jsx300OMzXmMGLAtOpATw/ZgYU81DwGZ5SPfmDjpH9r
As1VdxBO76aU5h8pMqOzfbesjHZkrMsEQEr0hKU0ee0Ebru0OFuBh865GdWIuHqL
C8kcV5gnoKokhim297Ah96MSVsrxenYbGibIhVyg92kZ/fRTRKpYORYKHZolKAqn
RAQ4oGExlio0jLRsqiLpRRYR4RO/mE3GiHfEivZGqmElMCIMrQoOGooZ9Zp80E4t
fcajF0JFNuwjKX48wxzVnjlji0sO2g2szegI34Y6OYkfDsyGIqsBpWTFFkmGGSTy
B4fMEM/Va28p5mVh5ZJ0bDZrqWfwXCOga/7jhBlMNbYbPPgEYzpNM7Fcim0qaRYk
XjO4dD21N2nGJUmS+tMQc4h8VayacPd1ud3cTL2/1DOwXOYYZQnsDlG8KCTOdVYG
lVkiPXqjrM5Xc8mPHXSWyOmFV+ogjW6Jr9iaZ+z5JxYE12Y7yCFlzgnUvaIAXzUX
emen8jlizEjzFLuSVxYcndQ3X0fqx1OrVgeW5icApJYV1zwxczlWzg9fqAqmEomi
Ysv+Ox9MjD5C9FgsXQxd3zrqVjOUtySsQMDaiT2GDqgH+Ug8DbxOqGiPw/hoSbng
yxno+M0y7saEz1QDx7nFu24FNt/YTJsVwBWw/xJBRdH/6MQXPgMI92VGm64PKa6N
tFi6/f4vWXmByW/CeECaK8vPkbnen5mwjj4NbIcwL8CPtglxHMOQoluuyIkjfn6r
KH62oh069kirDS8ATtxryhfepPc3g3Az57+DR3dqZKbJhiMfOLJeK2Y3o7uxEZop
7vxMJMZjMxkW/EZn89c2BjVkA1beQVnnoWUjIofHgvUaHvhak3+MCYtATpuFt0PC
gsz3jMq8iz6Jg0zUCQEzcZ2epI6ciiOZwanbdbZpsKfxU6N9OEefjQs09edd2M31
mgRyFUnM5yPEXWIp+qYrJug30TkYDzvEC0i0MH2q0nbK1E+lGhI35mtFgPDFC8QZ
HcuwQxtE9iwT+I6e6/5IKql4kRz0TNI89bNfiHkGd3Iie3/Giz2byWPrRSJpoRI2
InZ2z9qa2tgRb7iv6xVjNouKoTFzkr1+dkjfOLiO+uh5VfgX/RVWOLQHjCJ5rgj3
b/UHQQq+zlb8S49UwdbVS6tLU7hmAPWmoDbyQAVF3plTAxrUfcr533B1qLiz9U7F
ndKtyFvEi3x9vn+xf1eWU7c1Xb3jpVFr05yEOSE5Z+t4qesUaj0rkrxrCG4Uiu7t
AzLZQfELohNTtHk9hFu5yyO9GhXlruFtNMuIFKze8CLL+8RxSgqhMRSJcm5I/MV0
udSM7xk+kVChhGY9QsuS/ughvkFlCUwFCTEEBkLP5tgBgqmDn5jbAEJ8HPjFLodG
WhfCR5+CC+dTSi8JDqeZ8zXDg20SoaVl5Vhq4lumun4UTYRT7ssKDI7TBCFMmnrb
y0QBd7nSpq+FeWKwQH0T78JgNQKbNh6oYXR9gRUS+tCgaH7CAlZfUNqSJuOYY8Ko
vh1Qy0O+nva5rD9C9Sybvd1zbkI3l9pg5pq3niKbng3GaDyjI4MHyxZlETcNqslS
ZkMYATB9P0ZiySdBF3S68H2uSzd24LVKLAIHu/jDpI9rEFzkkhJWIJYCPztKZTuj
VFUZ6uWchWoSzb+HsiYO2G6oA6wmiqPa2+9W5dvOiLeQJ4lJJpTi9is40ujlFiL4
tDN4Fkv2zrUHcyLtf40tEIayK6fpx/y2YuOf31LP9bx5CTiAjxA1sLHnHks+GJGH
m2WXui4tTDDeefiV1P+HhZ0Vs4EQmRPeu2IdEWO4vFG3AS3il+1c1pSJ9y7apfjH
PvUrnGVKezrQahX9kOpojxtba6B+/bpIs0iA9W/RcD8JSqrXvQNkck7ZnMLSOSXH
pSjvo/XDtmAXWoyn08LZmPHkjJP2MIYf0b16WHSmbPxh67mrIbOcuCRybw8BqZON
tltdCWkGqncDSSpV6+t9J3T5rtNPCnDCr61O4x97YJy8s2TWuwWCNSLuDXYHbeHC
4LxOLeS9cTxu6+AgJ3pEOuPuNbtOr/ingSUY00j3Oopr1K7Il5gy08CQRM/TxZVQ
49XRPwzJTJ8rgYRA9lj/JxgStp/5/H5xjfUZvv033Cv4a6jDakcxQsGawpWcXjik
pMht5Ez9oqfke7vBf8DXe9vWHK8rhUZe7ZmSesc/wnqWxu5i+LtXp7H2ZcCLF44x
zZBVzStNis7cilqVz3HVgqxjY6pIZwHopKwSbN5cevvJNXbyTk2IouAAfg0joxNS
HFvuw6ocYaubv199agOnBhiiHEN7TyQJkgWBQLgpa64fOYiRKGNCPpKS9yxg98I+
K2gfya7TfKRs4JQQ/pQ9Si32D860xcb6VxIrMmAXEKHTNTWrP3ZxUpVu4pslbhJd
uE2MeXw+DzHzpPiFfPRn2VaHMxKMLit63yANtem4LhjtoOUSPVbNUo0xchjVZ1x3
r3LqOXEVom8AdCKsza80x1BvjMrnzlJNee/461+5JTZ5TMovWTSpYM2hutK0Ovte
6TEspLVrecoe5o8LNcU55Kn/TnFAcZa4RJ9mNV0tBp+uE6EZSLo3wNVaiJQxZMRr
azkyvYpVHO/jkXm13/1J3SzhDtJRlKjoxdUzSbaj8aIh3LJuu7lqQVi9NvJFDBDd
aNjYUVf963sP7CKmOdVkiXgd0CbAkFYrA+DZ5UNZJLcV5rktBpxheRoedTbQ5JU4
zJ9lF+be3Vg6RP6BsLpMaj2mFlhmMD2oW9iKbYQaYrkJLK6fBLo18s56rQSDZq8C
WY9N7aPcVxX+/Y8Ewbex/SZTfWdhSdGnfXRh2DGx0y8UYMxl6u9DWHnPeOnX54hC
2Q6CwgSVVG+OIULNtOgpadYTwN8t26NA2/S2PC13ePv0cQitasgtMOGbTwp1ZFjY
kzOPTzKv7E0CvmW2qze3eseiYPS5SjSLNpLrxBudX+Kn+7hvxf8m1GPJTWNbV11I
5zZmGmF435tgZcj5XnpfNu7C0czdOl9KNhAaxZYk9321zOfiJGnS2F+hbYlDkK2a
j9J6qcoghPUHDCeFapShioF8Fylvqg5eV2LY+nc/THDPW4TFPfnj4F8JiMe+4mDg
dBQIF7nMRSLojMiU6DNRK9uDNrwkWf2BNvBmwxBXx1lW3JBPatdbcqyGLDNMGmF3
unv0EJq3GDDSkCTzQMM42Ps3ZyxJrCE3TE4pGAWOdSvIVjOZ5jtJRMdgoquOK+51
V2IYTup1cm4mBfo961PsH/NtuvBgiOmGZedy6qE/O2bQ8WEoIXGd99/ywzhqoaG/
c9v0BwEELTrlVdx2aQ35kJrQSRdafvPkS8zrks0RsfawC5Ox/c/ekCJwaYtheYNG
WSCKq+PUsLntwvCDr5wcU6QjsljTgfnHjsa/UF3WNekIluF4zb9KQlLGBpZHv//9
L7P1TAdagWc5F7VdAe22iUGA9kUPge7qHVU4cIl3prhhbUemvehIDTO+wdB1blTJ
BCqoISDibM1MTUV47xu11vdBY3BOvPfgjzZZxW83X+aK1TBW4nvC6vEJ8O06QL46
7yPF78KkZKNcuBEJbxkL7+orKo9WZtbuDENlSJbrVf6LjWvOpaAv3ta/BN4t477k
CmE4ZkIKAXyeMQPlCAa2aMX9u8TkaK/rKjpxuhIyabvaNBkhVehGNYzTbNa8F5dx
A6ls8nt+oWo/5pS1hN+wpq3hXypw5qU8ccYNiSQh1vmc/1rx0EyMgutpggA5+iMN
7wuYLXolAQXRXPMeLmInC6ZZ/+mPNeWQIB3NPmaw/tTF0g9x/MCLv5F6jqj3v+um
DHcBHNyPy+uGrqK3Xxd6S6JDEPt+KZjItUkbf4kFSYqT3ThwivShQzZCRjQ+sBfm
l0hiJiAGYF7/OUH9J4xdhn90yrRtn7a+VWiYotlvOEGRY8A/vKvIu1630K1pK5zh
bjmXhfQh0BC/mRhk/GKNKgfNjJ1m3p7dhBVHTXwoq3b4TRXM8DWaGecAiJsPRWg5
8QeI/6R9sSULdPeY8ysFBhXQKo455MWsTW0Od3oTSHL7t+mbSLLiog8IoBXIybTo
yoVHro1nKCfkDJcXqBW0Y2HQj5avovhtmTidM4e2VddMr3gxKO3VIGNhmZ+GPKv7
Ayw/YbEtetkpyFbih116SASRQ7REOZTM0NmwLcd+W4wnUEk7Zfb088VRUi3CDiXN
QWeGim7h+JujsZ7q8/Ds2+hgStYiRN2jd8XQCya8apdwDmCCIzupup8GWxPfue+V
VQHnfodPVKVUmNtL278fKMFilIt6jpisuleyaGSrt/qBAmh1sx+03qRYl0jOyB6s
HVJ4bqKWdO/Ucntrd1YQ71+V41dBdDNZDqAaQ5JecmZ2lpksjjvR2VGZKds2TN4G
+gHQqAoRmZcvuGuaf9AflsigsZS5J/yjgMi4F5a54WumKkfg9VQbwUMlGNH345Af
/Lv4ND+QeZvjBhx6mr8WBPowP3zoDZ8Fa4hC73QV/NQqfWiX/jPQ09a0lDCPFiOu
Ay3XeoF85pgP7H1i5jVnKaaz8RaMvgWOIYbZJZPSZqHmYSQDPjIipHOYX0DyPnK2
Efsc5WtHK5wKzF6Av2bTLBGu86yhWxKLrBuXkEVt7FlxoKNfimPCY9lzsHagfJxu
phRGPzOY//pMEnA9IqAOC81gN+7WqdOOALv8nCsHzHaXB6Q4C34JSv0tLXxZi6Br
JrFCeNveYhIdqB1mHiVU6rsYVblnHvVzZTVYgBsVmWH9trjkxq6GVHebGWWPQr1Z
aqYdeHu/WqdyAB+eXMO47GoJpjWZkSkw/F+S1F0qxyHbddVm3Cyo4jCInRzTvNMs
47j+TrwiyI6IFEW52wQzpqpMd0x1Vy0p0okM8NMEDL7z84ZkwdgCiQnDgmBKiRhm
5CNHN6dR7/ZFWlPkYwYhlfgm0T1ppygWggZxnt881oybV3PcahxqIbLeWcjYWz7e
EABE/FRgWuTkqAbhWH3S8EafpfBuDjF5pmzzVSR1qvfUKFPUEc2Gwu8LYBpREYTi
ALTjCkx527VdPvrl0AQRLmrQxHHnYDihR7DT9k/9cnfiyBBjuxJa+1iYg/N0zlSH
+nujDMatImUBSfVW3z+rarXF6ISP/oNgDuYkhoO2zw2BiKGj9DnLYh7IgvBSXfVp
h2F/850opVIPvUZypUuBcVLOL50AnH3tj3MVebPEyrOFnZoo17bQhllVesZ7YIQp
KCSluFLujgtp6JjcOYEKhrWBJrPBsfMC5nTzqUX6fFPQbQUeYpSVA+I/WXaA6JGf
YbMfppYdQuSVY+Vfi5XNv6NlyPGs9esTBNoj6HrVqZ/BKMYFbiY3IrGc5po0wgJP
qnzMk3TpODX8DZA0LCVdd9ONdIsIKQ4ZRJWUkQYaPpKAgqsZyKeQhwGA5ssH3g2H
4LSjprbf6Bnj/vWxScwmIQHO/thIn2anV8PNfGDGgCqkVIdWQ9y4erLYOETMOH+C
Bz4UHoVtb25dFgBabJziFVwbjrEEC7/8p3fjv69LxWS9TbDJSRcV3zasSeNuYuop
n+k3gBiIonTbGyoYJkQXcqq0eUNZsWeTsMG5pjfNViNuGNuYB9mT7YBX73e/5QPE
ZjH48AMOa/0CVIK663nbAipQ02GImFFfHsX9cZ9TQ5MvpwEBlXmojb2IxAfzPLDv
q5GanhNnZIjzx+uXvKfIeYguxppICvJvhsRGyPEf9LTINzXymDAY4fU8Ur/sDiC+
oq+0EXB2v+ZBBLjiqGWyHY4lMWQSJM6ZxM4CTHrIy+vAG8VP9f+Gc4QxqZpdplJb
cROpq249PoedQLcHyhwByzht/U7sSLgRT8/ACGq5r8ghw8CR7H/9QBqeZKG5THdL
VTRwGpBlgJC5N6FTGsvVPH4jZZd6qDWTalwA5oTHlCkq1qog6/wcs3/atqO0aTDf
PiEtpa4+aZvsVG1z8H6YFyQO1iv0gJPoZTxewItjf2UACUGfjexe73gQcFk8bl8Q
nazW5iNW5gwGnGYxx8zyItyKP0VgI+IOwkUD6NI7iYVfbOaOT1PcKmCPdyZvwf3/
nR5/X50/HYrdP0geAcE9tmgt9IjgFBUUnTT6xF4IaWP+w20r690G7++FgsG5UeNr
UA3pDnLlWdoMPKPb4XxEEDlXdyUoz4Ib5hF8a0bWk7Zu6bGyHKhmD5RqENhxYs2k
QOjbs0AQm7BWgCbSn//8tmm3P9x/9koelIisw5z687yx66PfD5UpjwazyPpCpttZ
hCgL4c87vI56XvvNkdMbLMDv78Em0q+SgjuucQfpbSLabQY1Ar7D9xayLm0aYjpG
yBhWTd0u31IuzFnM3HDSlTkyT6CUfXbgQlHyB83co5GuaUguNLxMZq1cgN+ZDDvk
44fYBt03bi/2tdhECOJSvRbmNvHScZ8XXKn0vw3bG3EWbotsh58u0FvKLe0YvTrC
6fiSD6fHzlOAyg3apf94XG086uK4zPXtgtBS2cEed3qFs4eTdnkzYr6COpCtyJwH
2CAkBaUn6rEjVcQZ/jbPGdZ248oN+wyz983kPRJzKDiu9Kod1KvgRBDlE6PMuegP
+S3rInMAyeGrq8udf+sd5FD7fH6N0zX25n1A4BlrCgTLQdDWgU0E+9NgwBr+7b8I
+TmUGjLSllhcriaA/A7B9+pXR+bTgXPs/Q6CF/7Hd0DucaWyYHwTG7zV3BUjFBxf
u8Pvd4Nii+qM6fmrBFN8VTyrVSFqT+Hz1Lrfe/Jn+W2DcKF7iK21Hwdi0bQAHXLB
r6nmPiEWkM09X+/e49gh7SBU/hDMniIJLBRU+NuecpLR9ndmWeIVzyae8uft9x/9
d79l05Boj4o/MJjKHwLCQhnaH01f4PZxiSXSzJ+vS3V76Fk6Zyhy6ZDw1tYLAKKX
kRudyYUpjn+IkjsIvxYzyZE70+gsbkdNUw1xUyOls0JoznOOcYWrJLIuYQv2GeRj
wkAu4eJipiO+msgs7BIXjn9EWY51hzcHIagvMOdSM9VgJELTRi0+tnwWRQSXX7L1
XQit5bHnHbQUty1l+B6dWoxuELG1OuqQnsLoOZpoT6qI7cw3HVqsKzfUbCaETA1i
wODDLG5JDEAVklsrCH8TvGLucIXkiHBws7/UsuXyMFbsQ5KPLdHBnVXf7XCPG9gP
d785eqmLVceliHJx2inBJQZwHaFKUwipIOKGODf5rIt6reE3WH1CTHJnwE7JpyVV
OzI+KikjL5TVOfTToUhnU1+9zTrPSE1ZLFnKiSS0Ob5n7TZoI8m2UGCrIhAvzj9B
OTH/1FZ9YN240EyU75c+spMM3MYmzQWdeYjYUfUa1nunQs8MERtI0t8w6dnNsncX
fAmKRT9mlrJYKND+m/2Bo8tm3Ho+sywVdBhbF6FQb2WW1ITg2v0//6XddoAJPkY/
+MYbWBxv/zgB6Af0EpbzIcnQL6OOjBDdA2mIjEryQi3SjYQWunCNidRc8y0egcFu
XfwuI1rDPPkJYGLs5UteScxsZPJN+dvDDSSza8n+O14M87RnhFAX5zbdxd9uRrRv
7OoWTaT5F/o2ELoj9TS9+nKH7eNOuvnXtW2PXWp9DtiRLx8Bmi6Wbu3qQX6F3WmT
GRxoxK2KgQkV4B9CUwL/h4A4RMz2V2hNktr0TPCR+2B87xx4shYIkmhH4IPC/+yL
RwS0rR4bLtc5nj7adO20HLTeuSmuoDD0hU9QluB/himpQ6vmBGi8Crv5b3Qs3+DG
E8IXCN668riDp5D4xWDjlU2JpMg1s+fLmpMW8ijnHUEWvdQywZViGOlsP+TiUkyq
nlEcSfqYPxxI6hZtA/rUOCxiNaj3nfn2ADXLjkGuaBbd86YGJGyh1uzmlBoxanK5
FH6x/mblVIExy26S+V6j4tUfvVl7se19EJCNOBPDAHD4nSUtllyTYFvfsrg2XQwJ
KReS2cwA2HRj5X6LyD5Fav1hw/Pryuuk8MNDeTQ85kWr6GZqGDGa0dfPLK+igFvn
BcGp7Gdh/spAgyh8hZvYmmWuBdeOu+ReX+i6RJfUL8K0QuLTN6OUr1In3Zek9ZRm
DvTT36zCFD1Yc72vk1g3dYBy5odEZbjI3du9+bLnYvqd885c52zAyncNMHIxp7dN
roFrrsbBF56RHRCF3behhGRkSjsXERpKaRmfXzftmAxxyuyuFNplkHjerfMHANz2
qfdLkIYb8y2ED9B71AYxfHZa+GEP3AcIP0FomtRxjAXkQkdCoN3YraO6KHjWNqfL
g5Tn1mpWJMIcgwdAcuA3/5US5tEZR8EXz4a2FRWGA9ks4InD94s7ZfXNxJsBT40z
kP9jqFAWXrj+8s2fwaoL+xuq4N7wdmN3P/T4kpn85wCYAgi9zuGuld4ruC1jARtl
N46XIcqN7fb67X4MjowZJ4PQLAAHMjqDd5PmrUz6vuxe3diZD63VT9NWzhtx6fb0
vWbrW4E8OgOcL/AoMHhfHnhiDhyrgGCqw6HescWj1OdgrMW10famjLZebPMOvdY0
i4y53pmqN6OxaoNfDF0ymiUH3qijoBbqki5lzxOsdyl3dhmEJ6ltzPD7T2fo8+l1
s+lwR0apmofZHWVoJIrPz21iO0xe6GlAsAnHo70r08f0bTiy/581V4VqckOD+7Y8
8yFY8+DqtOmBAKU40p0KGq1HPVg/w42C0egkWf5nQjB/nGNwrGxNN00khd2VG7se
KgyYtnI9K21Q60jrUboEKnQd1vghQAi0w3M9uOOAZ6QGcC0ZuNQNThQR6KSk6L3n
qSSox9iAiKAC7lESnjpEhInp/7jaa1bVcBmDH0atHGYw3tQ/+Rx5ngQXhXxsd/cE
/9nI7T88x5rHX3c+1vYBe6CP0tE1J5IIvXxLQqyK7+XVhlkUG7r8lChV0mRVLQTa
Fr7m+MmROeMaLmO1fAm/RohOI8ffF6uKo1SUFlIiIuYoa8iqoDWQKkP6xLBYZTb/
ZDZNq6iKqWK79GNO6vkaavYjzg7iTZN0wUL3sBxQOyojwRIl+1XZkPNP3XOFbyZZ
aqGVXeAAPXyY/0a/ejybMbfjNNFMzo36QJQ238qGjvDfjv1d47Tfuvgbvm8UfIrM
/xbJqPbk7RN+Ei+f/lkQl3kCOatfVD1coGMRrKu3UrhC/Gc9sJPJ/axTXUTOd1EU
ICUO1Bbw3KDDEhQwd+xQFQofSuJMW52TtOewzcZbfGnjpN/HQm7ddrcJMWibxDuT
owpPnpOChwWXkalf/T7L7BDO3KLDXgn49ffhX0tHNTjY9mMUdU5bgc2UGlRUVv8a
bmcoVnfQASaaf7FeJKWwSpfUvZADpzrJHJL/OnYvZyuzFhOLainVewkQ9kJu6U/8
0OvqDgVNmTQ4s7exYWAWL4AIWHV/3JPq1RvhTapr9ib10Qd/xcy7knE8J65Qk7If
Qhgk6IYjG72qxU2/h98889PyExvD96n0z5f6jiAr8o1rhIcvJIEav0TnJuY8Qykn
GLPdTKkgodqY4FrOxNOVqk3IO4eHvUmzuHggv6pYAnk/DkvNROcznIiV6+wr6pyh
y5ysmsWpSQ5Z5l/R/pWPRi2ungQAQ1VN42abqAffDXnOheUZZiwFZ7i6oFDCId+M
t6g7jcba0yqAcLoHBZko69QzQKCPE2GkOzYEhjVrw37PnZIw0vFBMXMW8QSfH7IT
+S1f3FJaMGIOlNJZ+VQ6nCxthX5pl26xHPypVaCutgAmvsl8Jn1nwc/9JuCSFjOQ
QW/07YjhXIqJjZXkVLVmlz+S0VnASgaJIIzSwmPK7B4d8d87yD4tMxftNt8bhMsT
4p1e0jBOhpyxo2LCVwhXu3HLzlhbllpbqBqq6Yib5pNaqpaU6W3L+wQjLrkcXsU2
2emY2mtlYif2nPbbknUPdTdTECCJssg+POVmuwwQDQq5YlqNBK1n/iDSypXkpTQR
tGcwcY7K830ixLOPou5ZrpGw8ySPLxryHUrMvfk8dTldbEBWc3gl8A22At4ze6Dj
SFhqbxshgio6+iHH41dBinPfJP70DzcZnbctG1JNqyU1BKYj008xXBb+Sx+1n7DW
5ku4yt30ElQRVsYGov971B6q1GsdWxx/BFYPLbVt+zgcFyhPnDR3nqLHrOjI9l9F
yHqxT1dDgb2XtuQ+MPxbHOTLjyRx/R/59Tg4TN0QJqCIWEYgE4TVzYn0ouA2Qrg+
TAyrDtjOFqvTOAM+IH7rMh7MighcvFurNORtnqx4gbZV8ZIVwgioEB6LJRPHVfsB
hxUyqZT2tn+cCUBGGO2DgAi2tGalidVAsasOZUnV7VvCVpbpo4ijNfFP0qQYe2tI
y0kDfwW9jQzZVCyogT58UJlgRu+IMH+X3ngmK7jNRGucFoivniPFdBvk4UayH6Bx
D5rw7/6TMBjpQckRQRydmBmtta1LNA2Nd22yO3R0Vg99hNxSMOVWOcsPMROUZFOs
9yPbiCFDtBlulj4paw0jzrWQ/XyPbIEXUQT7LlIq27dfXoWv7S90e8DYp2wBZ0Oy
EbVssttgKoAqldY3G7PH3C7jTiuQF+sUMqvD4JJNltU/dSbQ6HDuY+gmofTGFBTz
IIW4qy7aCO0Q5lOsLsOBr+KbsCbkSTNioeVABUnKp1D+nJLmeNhy5LKuejDs4Q/E
TiyPP/X6h1zfKV6J1GrmkjO5dVjBScgYS/DEt86XFedCo3LwLnM7m3S9fmJpqUZX
kz7Kd2PPT4uR8elxiaWxjqZMKDKtzcv9sS7Y1tokbCUK2AHqFwka20Li+PCHtQ0a
zB9n+dT2CKBOVXNOjXUHPPr/M32ayT+qQB4YkepF4nQKzEPZwatffgXz1TJu3Vqb
74Z0bSEphME+PXCFtSzR9eZY+m7GO2E2phD0mEaluiITOlvy+T3878D6terQl8iy
BsB0YgZx6cHdto2reV17qEwkOuZFQXYEtdR1rEaQX0k2DPmiGCiOR5mtKhoh+9XU
pKkwD27G4E/7G6J2JmVEeWM9kPIVbddKAOva4k7bU0Y03OQxNIbXiiTN6/3jVp/3
9dUYNy1R4f4SnRAvBVflyISqNUHiOu4cFVzq6DxG72PPGlhl2NF2w7u9jBsuAfwq
h4e19Ie0Zo6bBiwGCTgyi+MOjR5W+oogWKOHG3I8TiHNTe+EJLm74AXRIWaByIXO
TYt6su2fGtytqMQ7ns2hvfkroW2YZ1yNRrU1U3cWKWZbtsOtDSyd3pS/UQlfvRZF
KyPy5BxjHbuh5hhv6sbNJGPeVkxgpnblOzjvOrNAvCgDGQBUn90YgDL+pbExtGO6
GJu+VrO1ojTMM3wQwyKlSHIxg9qSyOJoQjDEDjxbnCGq04JxjC7RwdWdWxCUk06q
tjhPxhINgIifev6wX38TpFHLCrUswX7HMCV4/+s1Z0qmXT1pOfr9KYmSa1bezPek
93affhcXKxl72149tQCiQSanGv6xfAC309dUPnT/ZzJrfux4KIJBZJo72KWyCzkB
mIJIpKKl851FT2bYGKand1yACG8dCZlx1ulQjfltFekNWxkwQzd+5RczW1bai3OB
UM1iRYOSFywqn1xWwfGeMYUOeNchJ+jOArquBq8IYYDf25JRe5CTp+kcj6+Loo0y
8PeER+9rsVfo4U+HE2AWVJ0eAVloBvuIt0WF6cY3pf3ErdW8k2LfY+obGRIeuBZY
lKJMOXn8vMUd+UoSS0mw7K/9/KNV7ULi6/nmjJFxIOE6zEbTw7sLDlze7MG2Mo9s
2l9MsAYf+Qd7Miucia5vzIgBsyUFE2OZbEtGtgbH/4yqDXrbIee+VYV8m++nwuVw
0Yh8y7JDPkUPHBxn4bdR8NQHSyj/k+/Q9AXVULeRz5HYEt/e6Hv+rIVvOOOg9upA
1k+lHw8gqa/KsFvKFlt5LRffWEmV0sJ1fa73mbqz2YoyJETImPiAVAxiYwHYW27N
7mrhl2o8NvWunxbBtlkv8Vv+HezcJEJwWpdlNPfBmNCK+qC+SjN3JDh/rtqFsVRR
iy48cNRRFLcYYFXOtMmlZNAK5vgQz2ECnsTI/4aDaYMpkpaLAnAmOD3AR5eVDAll
5cAB6X0+WPHuCGZkyHnt5vbAblMLbO3DYSVoV3W5SmXzaaHM1XYQT/+iQovCkttN
FRjd/65TbaAVUuBDKHGn7yTLvQZCt63fxOyRdGXRHeyonzEhKeTeJbhPTddmu4+1
vuiy5lKmAcyp8ggxiinUD4pNoVPfLXpnw+gEJiCK1YvsSu5rUsU6TtNCZHLIl23e
S8nOTFLzoUQiBgwdtOlcl0XhwG5zWc+4oN96LPDCFOnvwRPZnoV3HkKBTEoHebya
1r13YI5WAouYIyxanN7tBZt4rLtLHRmf7sE85iUejC4FW9d4/LYmYxuDhY5Ya6fg
yPz4Nm/Lh6WYRP7gadBc7/+rq1DRKHpfrGtpF3vuxfQWGEL5Qg8clRWNymqCOgZ2
qJQEy6KD3JU6ZrFL/atldXMddKo080XbMGBEb/fSfNF9EaBadPdr4fpaHd2EkLkg
fXRwACk2WVzfyHOudMJ+WXd6thJ3YhF55QxUfyi+u7VWAETTgDt86e6z4cSzCGRE
4iVwbfzoAxdQi3nfDk6TDawOnE/6J46Dlp7Tcw0MbRoVC4Xea+8ieSEeylDjCF1o
KurhvpoGgHsRv4o1TAvp/V6+g1MQKDpfQtKQbf/Cjon4VgSuWC6+/cAB4SHHpdjt
aDuyE/Lr9qwwHQFR0njo7cx5pUlrpgXQd2TasoYrYl6l2wcCir3aCOkwnUhIm0ko
5P2ajkMntl2mi/y/3palzLP+B9Ok4ZBjIx2PjmSX0UC5zlYkL2Nq/pgRF5zSAjRv
0uisk7lS5KpxRyBLjkyPo37gM6aqVHy5rHkxWshHXGUpZeWolUcTAaakev0T6Jfa
D9kk4oXqVGFPhVjDTjX82OHwqIBbAjGmlHfX9G2AjWgr6RZ+iU9qjr0gjF4HwS68
XrmHMiEdsdTpHdxCJV2Q3hbTuly0gYhMx9Z5f/BOr6lxSeRmTa7UJrya7OSCR4Rr
Cob80xeevmyNhJaXDbNDga+SI6QmH4JLyQIM+MP0p50sG1MGIj0PmN/nDAzPAzsN
QcJD9nzPbolTif6MRJrwSkzH9wgFVvUrrLdQ423wP/G0eg+diFjWGx2n9kSvO5mc
S9CdNg+3bNQoclmYBGiCl7ArIlLgsI0/gL2mzuneD3lvhSdvuaH195VtJA2Dn7Su
4GsxbzP+JT8Jj3wil0u+uLjoeyQTBgJaQ9fzK8hy02gYTFDJHX3x7hszCVlqX7fP
Cr24SEG2StkRHTZNSuvuvpJy//2BCY8DaB5veP/q8v6DybwmMWBLf2Byas83QHbv
vXRjD527VcXxMceGjIxNAou34SvVE9RQ3/Ssj/mHuEnozslKMjIbkXmxLRdutUPz
u2shMOX9Hx+C02+46HoLK05i16de9a5MyM7m2afRts/KrLZslKGL8O4AJNwheEMk
6jZEPzZppjPLpdvt4NRTwarKJ/rgQCMmcdvnp186NMPbij2CkVK0F1Bp0jrrsWzx
pTG4NwOH0b7B1EmckGJPbvCTB06hJMlo4iyhAWLNKCXr5TEvk7hMUSo60usWLF7X
/Er9ywyRcxqUrTP9I5R8gYRJpRkQxM6EHYxG+oHLhxof5uLuv6HUQpUGxHqzB+/a
FkjomAbdU9f1uvTQeNgKu024Xs69tyAwaO+3H1H7JqYTx8CscscSTsIz8TLAkg55
IzvSPOmY8RGudQtpEvzNiRJW17RgYl6MkA8uXVrYQtw6R6sc3zUnylta4oaW8uFn
Pewm/pz06MmtJYEBPoy/4zQYN5akzuS8M5MDU+L79n4Kn4tT1aig2mGRQVPU7FCu
xpBdfcBqcGVh0E9WDoHe/lIsZKy946sA1/bT7RbNP4daBAlkAYJzDq6L7aXKTboO
45UlsCOqXz4s2WQgm6ktVX3o9b8zRuba3EzcvM9cXB52btLz659RIJa3Jc7JXX+q
FIIDzZ0D5lnT5OooRD/OnwToQ9CeKv5QRDCUm+6raRov0m7i5xoJ8u61CZTGTPGd
yvh/hXdeulQbW9NEJiIcv0OUdW9cmI9Wjq4G8uj7393cbHICj6Dqa4mSLloIj9O5
ryVbRmdHtXwN08/Q4QjDCNRTcakMAwsSDDkoOwDlXy5gy6Thz7apqQG7mng4bKRF
6BBovnxI63WJ62QS7z07eOlzvkrZOISOd5T4pRW739x/OxAecoG4h4cNk3Ygcgtm
MEXB7CKbygKsYErBX4gcihBgBcoehPFHzSyHG3ysMlWeCLUawE4FOwBKX3bqj1u8
HN9tzHaEPDhlkQhgYVDvIJg00Zf7/xxNjsCPMYnjtcXVYtSMoDT6q40PWdRlsF12
XnCMilis+zZX1V5bPXFytQtysTzKwDQZ0Uie8CqBHtmJG1um//4z8zaewnygQt33
jQ2WJ+NRdOMzJ35HgxtuT5YJHRIsTbRbJmTtWcDsR+To1nFu8Uraxwkz3mA++yfv
6OpN35dR7N/+bM/IUgUSYYExUE3GXXXlLrTNVzAIpPt7KG3NlGS8Utq7XMXQjK1z
5dlsZRcut0wH3fNBEJuG5CZleJLQpSNaWuAY3OD6abQZvgOZor6MtJ485dW+gemE
cUIt4hve145tZFNcKA6wY3k7FVtNF6n5vT3j4no2AtrY1LE8aqd/e31QqNyHdKu3
NzwpOiCZQAI7LbR5sq5v3lWzz2BdZc+Hj6zDNIw43t8aVsM7xbcTGyCzTQJUq1dD
NJkKqfWcPLRzi33Lf+SLQbL8Goh1WLLuxU55oK/GWOu4JYuKJp36l/cmC5FH3+1M
KprulA0Mc6Itx+CljUMXvjgLFYxGZpScAGCSl63cxC8s14+76BFFRPsX1s0rC0qN
1AKcx/6CTQ2ETYlBkRlJz8jZfXCznEfuvUf303LmlINnVQZkd/JwL8O1MfxyHGMt
YVCbgVVcsy/Cks7maJ+5a1uFQgu6x3OAqOJusdcb4DGeyJSrALXfXcXnXHWTbybC
lAM4FZfFQPzH6jHUDsHw3WQz/pgdIAWJJX0SEQc4RR/z6PPYXNUL25E3Rw18M4Of
2jPCbX2zb0jijsBNyCKMuYPUhIitjKbHkaP5ljeMp7yyr5stJH5Ns4+qtPbrN6Nm
v3jRseFs4RHPBLIGca3lDeJ5jOqRiI4EIXUnnC8Jp/1/JkalUNiFRxbSO+wXvilN
7tlHzhuJlj0MCsOu9FO3pacQFUYOuWpD3mF+UFTp4iQKK+LUnKVGUgknUfiCtYPZ
RDfIG/B1m4GtYnLjb7yE1FUCRodbUdcMVUv0AA7zMcktGo1qrlsHbn+YGZzWuFl/
CkOb0LTnfYub+oYQhPH7pBrt3FvZd5xw2bjmNXEQdzuec585io7q33wkQ1HShel1
tIWIJRKVgNztHU94R/xpfiJyqOqGnKXo8NPY3i5ZFzIqgyDqk/sNrzXqsy4986iq
XRM0JdEF1GieDn9vIw0anxaS/Ue4vV1WTPONuC0LD8oAmEUTWEfTWbc6SQhPEVnf
CsVdPKBRy8fIpBN8qeYipER/ebNK0UTP50XcRhZL0pwgNAcLh++Fw0DSiYYQSw0W
KoAhbScrdVQHvo0gnCSZyW/Os9+8O8qrM7FOoQ+ZntuHX0PsOl6Xn1GL6Ait+fzv
uj6D1RlA6G6HcJ6/TPHPT8PJ1koD23au2mlINZ2NkshGYt9AQYdWZy5yGzEFvaSe
V7HjRZVnmRwcql69Q0mW36xcW3vfAlinped0QhZUQXYnhkaRlpu2TKioIjLBNg+f
iDroTc62trwcVW98VnwOc3wno3RcuWOuyhkzX1ox9yIMvO/l6V1QxSovqYGEYv9J
nNwiJa2O+5Q/2Cd1vkE0WJuLU49jlRAxDgt5TNh9HLa3k09xPSuA8y833cSnU421
UlHB3JeM2wCLtMzdyKVsNEmaEUaRzNkIVEJydEP6bS9MUISaQEIy9n45/XjBV/wc
zzcfDNjkCsblHuEUW9yrbZwylMvH5XrnkhcP/Tl0Djn+GQGWyxqq6F/wuvqxuRNE
KHTKYRKfazDTniSqaNx+w+sgDeSAiWNQLzknlB7OAnwt/yeQABGymYNDRM2UqXeI
ZxgXbbFVj+CUiUvdq2NyAtC4zsAo6WLKre9VNlC7O5x1r+uwMr0FaK8oLbKI8ZvE
NQaRspBuq2NSJpX98v5TnRJP12FrEnTRC2SxhYGh8iLznA3vFlvZUKIzFYfn+qlt
NK4pEhKjyZg6yvefrbu7OSZvUArkWPbrs3/z811tpT6mY63iv2AikM0JiWQsq/oc
KNk7H6ZZ8KaBzGTFUYmy6rc9yO9Y/2Nstg0boike6I/1ZqcXnnkueOolQUVxrPU5
V7HqJ6Qd4qVcbFhGXXUdAWyKTldgNfgjzyt9IlZUGSgziHeCUo3aRF1TQJuvnMJz
987BMA7HjuWmk+jnCytoZZmaTRbQMBsq8yvlSA6v4wfchZlWPlm15S8bHQTo8gF8
OnqL81mdoDUfVgilLXLqeL/le9wPFmo6n3qgWnniCPL/Yat4pCOWm/kqZ/I3DNrV
tIkqr/LmXj4q5QPPCTVF+ndGMYSnIrO0xmhV0sNhN7F0f5iaR6ISEVN7BqRC1fWS
ISgCnk9n6kI7awEFeNH+jOgP+KhcA92tafT2UHzjBEu6ri4ei8Aa7Tc582adlYvD
RqG5RvzErzoTwf6UnmvaX8XsSdV4XgAZvD/zBvFogerw9iQ0bgDjk4R+DWqLYeJn
Lw33QlMGV+KQMrWbNTaMUz0VK0otpE6hucIYVy7r3/2Us0hhUL7A8epDj6RSWXdu
jJN6pZRgYhsVl4noLDs9zUqe7x+dKXaQMtP+Nj/Udcc7bEQmJHX9wWmBwId7bFWv
Q6qM6CXvW4OgJQwk2nL+wyRNaPtOzW4XUTzejGhTXBlCgD/oaqzWnMnqIUjXPydB
mos3+QM0g9V2o97NqhTx1H0kvPdzaLpGKgsb0xJDLudEZYIaEBdBRpwY66g4c4dx
PHO3MuF19EFP5fTwLbRakOz6tUtBUpnrLf1quR33zNqKp2FGACdCBEpvkID0BGNF
sfoVJLj8buAAindzdZUD0KMBrsz6ug3JIU89VU43l7yfAxsRrwFaaZC+9nEp9Kkz
IsQQ6f6cn1XCngCSWByu9YkNdoCVEE+Hz+KQO1BOlqK3alHHpd3D5JhX3d1B+ss0
RFAYwqSCue69HDsCky7+s7EiA29P/tPENK0EgbPw6Cs9t+l1InPvzl/yr9JSB89j
DFuEe9IoAavnGy/X3wL58CGHG7cWgDQ2VCWSzDiB58z9DUVDrJ38jAaSTAI4zRuL
mm/DzeCyXFudbvV1Wt0/R1CZG9ADTl+bNT0006Zsm0xD29MApe07Zni03fanyRgY
JCbm/2gZqiqpqtSlWB0Cps20SZjXRW6HTDu2mA2OvXsJBSG6GyEdZNVnpLZw6tU5
A8pCT6KpB8mCLFgtoI52HHkwqK6XnYyOD7oQDnER4S8XDP2pqb+dfSLca6behQYl
C8vdIP4Y4nxwuM1pZ78m5R2ZjW/SWWh6uN5bpNuuOJGbrfAQmQKoywpQZyWHUnpI
c0JXhkhGBD5YVZZd/ejZ2lTR80gs/X5uH/oD1zZUP8l9ICo+GgWE+ncY2r6Ra7IX
VJ/IPcrxmX8zhEj7CeznfS4zlXPpYeSj156QJYX/mfj+ShghfAL+8h9gm+Lj5D5N
/3/TOtRMfk1z0IrlKjTqEFVyefWENZZsxaZJ6cBNnelgs1cL568FIWphDbqT7Yd1
xYsL0ti3D6IXSdBaVcIVYVPTwcLVA5i4/6YDxbPlHpdZ+MIanSy7IQpNUEyENPJb
MlwxcaCJ2PYw4C0rLDmid2L6OFA8KTnE33z6kXwE+eYCSmrLpan1YyAE2a30poTu
bqvo1HhFOBftjjZQXs8i6jIQ9kfTW8t7eoSnzSHqODOd2/KuFY94zso5mpSyKB4A
XJhYUSLuXXK1SCHIZ+Z+Kn6OXVIP6krTEfzyzV4rVp3aYUcOKoCRqnnQTkcYtZXv
0GM56vzW0tw3xa5PA/tyvtd1kZZez8xzzE9I49WSlPdbdY0o27RF5ip675HlkGH8
hb9ipdX4cxfRpNm3WR+zlwMagDsxG7/n8HRWRl0v0IRRurX8J1i0hz8FLLuItkgV
4Ex7+YvsOK+ZGvKU/XPpQdVwVGnoP50gA8hmwUAJ2zI+bvNfT05gfj5oAahU1l4G
SjYe4W3Q+J4/jU477GL+h5EXMlRUU7f+r7RygOwjA9VOJT0DVwx4ZtBMRAES5MMD
lI0tUBkMjmvMn6qJm6Nlv2+hu6xd8g616fwVQHoPnLc5ROqXzFWIdgDNkP1XDCLB
IzORvRfdJ+m4w43kNip8NykpgzLt0c2ErmdyNxmUdaa3QC0HcBJVAdUQtykMa2lX
YjM6QlzEoXqm8YwysNDgCUcxVvuOiOTKsw2DDGo80GbEPVMtq7PN8wizGIdy0pk9
wUHJlRjatBcbf88Wfk1DPmvjUW1jDJ87VU5ABw+xUKse3g32qmvF4idBfnNlQOLN
/PdimJmZP+XJ3T0f+tzrURMIdHS5Xgo5TS39q9WNqB9FYbmlp07phOYlKGqQoQBk
D4oVDTG05VE7TyVSsfw3baFjl2PXwu2nKPBh44IDLj/xC6tsJsxzuTx8LD+Ts65A
QAFRf1MCurflfMiDEHzNzV0Z2TDa6hOV/NI6RPVoQvH5w8lv1rn7GDsoWqCB33D3
IiXI3Z2cChMlv6rqMVL8g6OOmXxjJguf86T1/UCjvthH1aOJX5OkQazO3YgrCu4m
aSctvbwQ6RaKbYrxdfpj8MpIkzc8QMBywYR9LKGpzjBgNH9PelBD/X0cty8RKRnE
PUxVkgUOBV2pM40xndRcMaLKnL36ZkjlYOuKQk6K2HyPBtCnV1D5z7G/wTlplmt+
G09E6eOST6x0/G7YstzhoB1qTIJ0crGLR6AL57wzaBNbxnOHBGWlak9Tgwq2asxx
84jRnfPU2ZSj2xoAq0RgmM1JB5fbMHnuxgIo4jHXqs8DB79yVn2yxMFszG3IDtMJ
fJVXY/kMQzbIdgt9u8avUzaZQ9dyMWar4uEHAfyKqKjan6US/ItiBoCrgC453ebs
VpRoZ0oB4EElXEkRtz5Axx8igGe3TDwgV7/bHWn+tW3PnH6w3J4Njv3tiipbC8mv
Zj0C3rNhi7zTEcRoI8VRNQJ75hN2WR1eeFu3W8aW0jCq2NpZNkQ6Sw8e8fOphf6w
mRlSrPsJlilKuBDuvBmhNMCugBCOgSLgXl84r6qQPnlEGpLBSwjZTGB5U7r7nOO8
msN5CrkeA2vD4ug5BCtFyssuYHLnyAgZk5AWx9cSs/zpxj7qlIKwilaEl8pR41a1
OB3iraOoQ4tS21iOo1gS/e1I1IiUKv7CDfNeNEAkGZCrHYDa1ij2hwFCljFnnqNj
yOjSvmHholfm3lAKoDskhLk5pCUGV1xgWajZlfMs4YAgMNz3SZ+RrWznXPUgucBf
d50RUDBCeUnfKYmkGaB9wiIqD7cg3FrjOvPehvHWgFe7G1T2wKpgbM7WRCnIPdjD
wESUOrDKpo7E3sfUDpd7yvQGC2GKF8zyicAYUmhGc8YvHp8+XyC5nrZCMV8ep2U1
lvFzTRcw1RL39Ui8fKsgS+4XPIT4DveDcY1Kaqn+LFrYc7E1m0nQkB0YwvdjJCv+
DnKAG2xH45XZm1kHXKYdcKkrr2X0m8HMHNykfe9QTGX0fv4ej7igmJB8Hek18GA7
3pEOPYWG1WIxRK9zjnXNv6uNJxDZtyDFh7WT3m9SDfl31rg4iRKFx9/9tf/fh60p
aQW3Tx1KznoHtWxMXU6PSJMqqlTsvtvimS+o2RQ29Lyx9EFDdoqsaEEwZY8wgEGb
iw4qlIQlwouMtWNiTGDOdLeo3wH6+tthWchaG6yXfeCMm+YH/pOIWjCYdjBCGAow
v5qv34opwP5kg5iLe4rIhmL+fjXyE1208tw7iXfOI0Od9wkKhULa5Nj+FrA9ABgF
nak6igBdmQmtH3QMEU1mteV7GzijGkOcSgHbiPc5bbgE4Suuu1+9UU862KJW6W0X
3fk9sYHpnj1Xf9ClERNjqi6/y9pXCQ2HturOIELSOCqaKjGoBR25XKhAs5txS9Ri
kvPcQtkeEXTHCTk+usMbFLWgpbaDaY+0DOwXMmzKuy+GVY0jk0QveUMO19QPHEyx
4G8duEwRevOuFqeau7+e8P6nVWZUEpm/umwlFUh89hU0e50eRhNNVtphou5U2NgL
dAXVqUrHsOxsbZVZFDZ/UPafmioa6//ORuREynE7zuygbepKP18FNh1EUOKkMh6v
XT3rHiyEwe10rcA/e5O5J8L5D8FutcfFvQkjsOFY7eYoXG4PS1R87d1dJWQZ+eH2
KT0bokmTEU4zs5fcwU2vwEahrGj7DLYG6rqyWUKAP4ZnkITFstOKy0LMmXru5fda
uWqsrF+kp9mBWF/PcVFSMsxrLdeE/QtlsR9YKoNrTYfXnuArFhP1KTTDpWejheI3
ahBfqNGL12F2+lP2a/KzdhuHXAej5SHbONPRvMImb/jDJOVcefemxQNH7a1q6g9B
lnznfvls83cfe0PWyZOJ7ap4LE3ceKTj7ifhyZKhkf5h/rHEjkE4CQBtfdviT7Mc
BWAWUxVr371/KpN+bC69QJ3SEFYSnicczE9W80IKJB/TN04JYzK5vlJyfDUUlHzS
0daQ4DduI/fXL1nhny8NwBCIRWKm51L439Ln9mF6Eb60HGhc4izw9by5YnqM6KBV
XXI++91sXKYojzlvn+RgXKiYKIgDCm/62cKlWFcQTTOBIQMPI0jqRqiAjvN3ZEv1
x/tPeuqWnHCMYsDZB0+tFa9kfiPcHtmFyYys7p+Yy8RYFuZt7nQ4TmHYLeFwSEcP
ZYO1DgZHhAPOR45dxIqINAAb9Ct3W2S4hzBi/Ph03V8W0jjzJmCEKeu9SP+qwhF9
Osesh4MBPkvmPtqnMY4E3jZuC+a0DgmUevJgQ1O+5SqPICuKJ5JtI+PdrIzYjgQ2
vN0cdjLAri3evA+a9kONxj4ZV7i/6bbiKJuWgvta8j63Krcnr7Qy/Ha5FTHKUWib
G/TjjYB0KzbtmVgd04ZNOk/xw5SOWfOwJAF6C3YzRGUhTNL/CwvPB3xyvBvxWhHL
y/5e6vvQQMJiMxvgzXuOMUzloK4KvuO3tI/kmqQP9zUKNgqbq8RJCS2BT7s09pZh
wP/S74GWXwdXsyXVTlVaP7OefUfAg284mnF5Gq5qgLY5S33zOfAiSlCtZFkRb+gL
Ej4gbWp/iWeTSWrrVDb8Y8nN8MV6cN6Q5b4TkJK41RbqgLkDBFD5PAzfLRhcrE9N
GYg9SNczqhwQvKb1FYvaRNuOSwz1rMkbGHaGGRVF0+cC9xZF3fUwteTgFi9RV4YU
y0LYhtqhCE1U7ZPi6qpX+MWDcoWt0d2lCtEXrdHSuuvqzSPluv9cEIszlMcxZKme
nxLTbvDVAMUfLviml5m/Eg+tqy49ihfHp9ZCY+GkKE1im+tdoscsiHuo5bbnkoej
K40lPQ5a+Igsx43gIHQlpeYW5GPaYbFC9aZ0KRHp6q7hrJ2X9qkGHNtJK+mOfcZE
Txz2Gx/+lfwdQi7a9AUBfUASvHO0LWnh2dNSSuGy09wDQsGlI1Q6yT++9Z2aPHJU
HvWocCRDaJT/sQ21xpCWEQbfln0cPSOLzusgE+6YfYWObOD2bOqHcf1ZxvTPS6Tj
umLkN9uxZjU/Lo85nk+uyVrdJrOOKM0BBl3z5L3v4sKOPIm79pco0+eSsTrlR6yr
ZcVKAgwgU+gRdlUiBA6JFbDKkN9RY4y+L+9jv1apAmu0ug1ria29LHnuRf/WivQr
suaEdmdhC4VzQsAPUaGsF0AbgpiwmVETtPy8wil59jrQReF+fnXOT63Wpp8oK78T
GX6w+7jJy3p7RkPQ3hfXif1L1g+yF3u0RQ/+peDINL9Qsx1DdTd1I44899ARp3jl
XT/Q2V0a3YIleq/kUF2f9jrh7CI56hM3e6TSIWsXNQaOOiQaZIkGsf0RJCBI9gr/
8eEa0UxS4sQreqp4rMgCM4TwdcP+IXZ5Kxqqa6KfvkLtyexWhTp/KLcT9226VK/2
i0CKd9aQj1u0fH4hmF2jAzaPRWrAZDoIpPlD7Wfm2egyJj5AAd/9M1dzZr5H8SYG
5VtZIwePVLn15XYKVXiokJfLuQlbcrwSRoKO/ZP/aF6kAXZAdweiXAVUZCJ7rimr
RKB/jClDIoU+OMo7W/BTaWINFi9lbVNGK60qTouHaBVBKek/rER8cFpmLuWo/DJH
WOg+DMjHlxFAeMAQa9G1RuvryJLwyyqDOnIxp9tmeCx76QJbzCx08KyUIqYFfnBu
YaPDjBculML0mVpD7GifGWy4b+kqf+d0I6x4kEGCFKX6vhOLe+/W1gUVkKPUi9Hr
q1k3xJoHpMskN4K00FzpQQV/8Uhx3Q4IJiZ9O4HMoVBz6HfOPjjgyaua45ELSD90
l5CWJFSXHduJ3zjYUGkEMfd7+/ediOvhr9736EUaVLh3leBut3i9rPRc/RAsbvgD
wEneNDDKHVr1Dw9Ao3bHws2w/eGApBgnCuy3iWRSnDfa1pyKBas3ky55OyETTygt
BkmPcg2m3CbFteQQmxnuWMzUlxQZz0p1Q6/lM0HlaLtOSiP2AC/VHUgCmMnURV2b
K7qf0+J54jAaqFn8HKJqVwVaCoOab4A8oJWMmiMKvvfOhR0WXt4v/xANHE3lxNiI
hiOr6OvjIwQ1SCDWKOtKWFv1jE0UJAPQX5oDXRnyaEg+LNkZXQCVVHjaXjAHLgwL
pVCjjkkmQtcpfuLQ1jqOI9WVOZTQUC5IIoldE19VciL+CLCzHotziu+/TjLyU8iU
7Z8zSz9wPbX5UmorCT24VaEy8BFI4lmOeqwxvxHEy74AcfxC2tu1VPAlFxndqqBz
0qKmJKaGRtAaFS0cDM0p8723jJp80voAA/G/rSI03rGYHMLyJABsB9OrUCzT/d3Q
2G6blKCcQXL5xEI0Yvgjc++5syLufqE5GjeQUn27NI2VelsRAAxyM7XYRldVVdEL
QBS0g0s8reIFQJ4Hd7JIEoVC8wnbUU98Rc0wcaTHKwUbH/AG9b5Dq1gPxs0qn/Wq
3vFV4V+l9TK/NTUxCxRNMg4br5We6ljIoT0G1WpmDC27mwOvMlgqWxmoT+kb7o1O
z0ABeIBoI/gHOzsY1bajEjRsTVVDz5Ikniy0DN5Iw0MXmN3nekFe8tiTXhcoBDau
nizg3EdJhfQC7ku5/UFV/oY6BxWYr5eNLMZdIFRWPOeD6J9xvqHStJEfDlKDhiEH
skKxggC0skZ2JzdiJSh2UNP5nnTVS5aE5+3hDIDYAF7UuQ7tz64ehXRot+9pvKR5
IC2O6sG1caFhYuCua4zJ2D+8uL5fg7+BSobP/Ei5JG44tAD2WwQuWAWQAD6f5AU/
SO8vNehyDD/02dhVwQrplAHQdaXUrAOUGmZ6PZfSN1Q11Ji6uFfSXo91p6tCjzkW
C/ftxS+pu6Dm9gg/bfDi0feyZmuzjYLnbXAirYVitQY+FXrvTz/Yfyy77kWpXI97
gfhUQVtDkP0UDvhoOU1s457wj+1jkDK5D3ltiWrHnPl4JbwVgwvJezhHQuB+SEqQ
5phmfNCZdyJR76hRQn8QvMwSiEnVr2eS+oNL2wZyrI3i7RxdK2SQgLNJYzVYMgM6
TZfSmrnIt/GskvQoHxX6SyN9+WjWe2MYnZfh5H1Mscyv6IGut3k9qRGubfVfblXT
a/dwOU5B5DXMBsicwRBOzrK/fT+U/WRxi39B0Gc1WyHedNBZRBuI+uEDWCWDNqTP
34dgRwFkjcFPA1lntSAuA0xEFKoj5TjL75oDQJYlRua5WTBWVLiBS31OjeeYVa1/
CjXHgNTKh8KYrZMYvGhwJVXa3bu6MK/bZW2+s0yqlGFvhwl6fRbVva31FCnvNhpi
acW/U/sKndgO+3vumO6kJ7MCWK1PbFPGw4rE9QtV52LAFm/KpfxHs4Kx9PJGHcBu
PXtQo3IkrZ/u4nr/CPlEqsgbbO4qs41nmYAf6tiHmv4IqrvtX7/SVxuXhtK4gfu9
n8bEGPLzc6xsRnR3cWm+bXIXzhOkImhsu0DhIm2mUMKCyqNwWSW1r5AV7tBtVRtn
fYUi4UuoBoyo94ZToyo82GlRyKI+OTMJ4XpzAMkPcRw3KXVkpVhPhj2Q0uDW65y+
9f9tRnzdAHEzADl1Sx4xPt/bgKRiOCElr3XQF9hMcrfClnXwPa2QPNgi9tGmFYCk
wNh/mglHYQ8EcbXkzcEQkdVdu9cFXXvdWahFB7MTRdbJK+VqdaUXpb4RZSvTfETM
X4TBaXn5lHEhg5xi7he6MSRNUwarM7RpmNPxPTVDu3DgsPkLGiaetzzfQrQKl759
Vq5epPvht2ZtaEP5qivaQFjnXrhE+p48qZJQIjeOsQR3HMsi+HWY7nNHoZMEbSQs
Psuoe2N7tUeE6fGLEzZKmNytNonJpD08wjJna8Nbeu77ITse8GRDA3WBl71H3u0M
auOgGoDsosw8PZZpT4fpAWOYogajeIxwJXzZ98BP3aqSYZe8D12RY43UQkSO+dqE
FeznSLbxxjsXxXefTIzrLVKJCyLEmpS4n1H/tfm0Ux0eKEkQZ3YqYw+AJOufjMgJ
wnSikMhdowMUS8wt+WO1iTYkEAhwJO8U0Es+fwbInvAA3UNnl+m8vHZIgo93cRRc
KBnNYJZ2LNFTLQxMD1wkoj4L+tf4kU2DTtiJPe3aM25JZtAlcdX7SV4s+e45eQH+
kihXzCByzKzg2+QrZ8KnzpzPPxmluOpOYKpUQTSus97z5JcDRnUqBQpspgz1T/8G
Nv84p0Ajymujr7ix4l2v8iM+N3KIG7eQGwZheS4+ifn43AAQyjwU5EwOSRZaPV8y
XUYUb+3mBANLEmEDjWHQgu6J5RRNCGSpdG1QyYrWfdOP5pwGfoZG94WwLe0MFHsV
5NSEQOMS4L/foVjmXlDiqjHsxCEExLDhO1dp8mWrhLVZSej6ajMbji2aZz2+F48b
/9PzqHm3/kU7I3FsmjB2XxpRe56Jd/4YvisbHN7hOub/cDE16CniIRQzzSu7xojf
WaY5fV/l5nQ0oiw4MSwCQrj6FEOzpDst6sb2YpMFQZAG0yKe25xh4oQaKtxx4h57
rUHfDFRuTrUMaDm8cFwmqhlXJYydKecBGlWj1uv5m/2JT1iptkUrrCGzIJFc5IxT
q6bL2dd5D+LMGne2kVsymzLyeGID9y5HIZz33ZULWKD0WoqoDe5caUyoxKrf9vCj
siC796Zzvg0VkJhnZl5Q0374G+7jWzlv4KFZPlx0Kd6SwKnxnJONfoVs0ktGmWdA
WhiBBU3HHauEQNETg77ZGfroF4QY9jh1QbxVg/v/CJI6sCWX5nJ5HNGw6ShVPQzw
pU1Iu5Pflpg2BXYmLBxVbXaMrZMNx3VmsL1WFoJyVEip3HJX3kFyEh5jgfexQq+s
xRKq8w6ScFcJ0GhRheDpQbxFi63heA09qKaXdaiZbIoEQUax17pHywUKt0UjNHPw
pWDEU6C7hn/BZEcfEFHTwISzg+ddSKed28KnRI57Z/Q16ORcRrNQqeUz2e/5I+7n
oju+k8fKSufv6xsx9GU8R0C8us/pS5I7V2hABy4tE7C3rIImsRHGKSD+N6oeb/9G
rJewTyRU+8X/JHHOmQhcXuWAXCPlVXlxC4J/2hFUmZDAuK0pjra+QJls8BRwR03j
SiLdP5qI2TYv0XmbEWoWZQ8086DxJFw/Woy8SxJQdOZoKdBrPd6lyvJdN1LemxHl
lsJpTIZ7qy4kyy54nPHhwyGTh1DkHdEAyX4+z0/cKrcDeBQgKWa/5VbuOmSX6VeS
+aBcSwMaOx8MJt6SOGMbDwhZ5zWGqsl0cj1IxanZ61M/AquJVeBb9tSjP0wKyGfa
NfGyw8HWjIN0yk2M8WteN1kIkkvwXAIFTayz3XuWn5gcheWzPvmXteic0mHd4z3V
Dmg5B8BygZqPSNwWn3fYLre0AhHMn+x0ZjpfpP4Y3ApDWkmwR3D56NmiQHgQ0fQ6
3j1fRKE6Mcj+jjG9MVTbEA7iLVnsYN9tUBKKy4nyQwO7wE2rfcEF87EIrUwZFB59
C+/vQ10e0CXp9ZTfbJ9dwwr7owXWSGM3Qvq2Zyh5BRTRkmKCdhXCua0Qvth73gDl
sa5KPrMfqEQCDSVEgB+edLxCO6GHU4a/XHIhnVb357P7DE57W+wLjKs0Wcd2WXRg
uAtT7atWlm5d7irXKepYkmLtLesbOSxFPqquzdKyEfgIUiwxb2lMb48Q/cMSkd6y
zwsLdsVgCYwcqp6zHf7oDtd/IOU4jVBtl3E2j9zB/nZEfHQSiXG8fky+UBuryGU2
VdEChqCw9nUSGVjAt4t8PwUedSgVw7tOy46cH1I40kD6BflD70OnjQGI5oASxnVd
bzQp+zd2VVkzipyGMn0cZlgVtwkvSD5Vp2KsP9kxsdogR2AA1qF3EYIUHzzi7lj9
osILgWVKrv4n+ezo9ej5N1HrGacioaGmDaFYpMzyIn56ZiV+hBeRGKwHOW1TdG6y
cuTJuUGzI8bHOwGVDvkz3hxjs+GJxdvz4vx2QyjBtSmg7P9+5FERdoDS0EUU2r/p
2Vr0cRNj7/6LfFXTDEKeitJVzH1k5nnRQvakWsNUlfeAiHGAXSJGZQht5xTcH7Hm
WXv3/0TuyBi8vzbt6SDY0fBraN9ZV2Cm7mij1ouF5ALPXswhsRWNkFOc4/rQeb9u
EJnt7vch4B/qFs9dhiV7NReOgV2CTzx4jFBypgQiVcaG7PxXg2EYpBRipIKuB4sX
o5cr2eLfUnB+NWdYPvbBA2UecQjM06wXs+GUgr6h+0NTw7THLeQJxHddd+52Im/A
sfv6hRiblLr2qLXWlvusIWLhvPKFpy3t/Gx5EyAENT3+v0kmy9lU3WtBEasIByRF
Dysw7BuFSKfIuaJx8KLqmJ4OTwPLkC9MiQpBeAVISXBGQwCzmoibLneUmv/qF7py
6spastR/nI4MfvIVT7LpxHmtKUeHSVuE9f1VF/VimEt/OGBaY4/STo37KoIblGJN
9u6f3rvUKbT6qvWmnEwKwx8GlJ7VMFktR5uNt6HMl0rMAbsiebHbVewtuvMVY+lC
o4SuWHDfgnoEpYDOZuHWqbUwfni3tu4RJfa3KAQX2OL5SHkWSQhz/HRl4UV7Q5JX
7ZhmN/RcmOKJX6traggeWjky+fcgzP/5UAtz1mt31CUVjW26z1EPe1xdPGv9uZeO
/5aPyJKItB5Zrykz5EEb7fcLQuntR9CXknIgGn3squd2OqIid/4ZoXh2d44eg5Py
JknUuOP13x2MzGDK0cHrCFOofnv+pQMwhRmzGsNtiu0M23/ScEiGvDS0Z+qK9liM
nfDOD4KD1arLMxVkpFAwm3iZrhS34cwiAXq5cdTv0UcDs5py1CbxxS8LLRCXMyhD
gfM1N3nNShYSArWW79e7IJQ3wDGcdq2iikb3c8PJi9wltbzxhYnS7d53Tjezcw88
iTJ90C2BpjcEV7sUYjLLbWk3Z7Axwjyri/nuOIceHAUXmgtSnIT6LqLgIOGZFroW
vwgAmL0/Jie9HYLAf2tV9t5d6NgPFWgreN/UEU1v1oJMJ6Jve1uXIiQoU3sij5lT
c/vURruTMps3hemCPR7CRMEsV/sE3CX0VybglMyZ776tX4Z6aXWENnfSjjA49xir
qupyYr8dF2lEQjo/m4nO4GOqXrGiab46r+Ap4QT4n/ikMxXetuPJss/hrfkQ+N6G
//snXruJLlsTAfYwQYWla4gJuK5yOLKQGzXSFIY99HUIrOC6hRvtUd6TdUFcoXmk
ehY0akTNvhUkD1j50vJq8aW5Wl4vwY05+UTPvMFf5NEGqdwagmEIktNvoK/7Znhw
iGUsnFUrGVnqehxbaCZfoQEOjjyxeeuUBpy5x8s5tLiS/Xntfj0qoAkCfKjkM9g0
4lBTwRyK8QEwYGqgxGmfUYRX9owr23dIsHtm6G+LCSUhQrYXF6SQ708b6FLwaq5r
cRNenLnd2GCXWj3RZ+bYpO1aU2q20bxbIChAbuF3OdlQWXzi525TVCEm+KiBTr/O
XGlrZI6rTeYdbw1ksFAwZ1lbBAsvEdiNBRmnfVB6mcz0VW8e/7I/hRGvAOxflYpK
6FnwmsdSz27h1lLUe5s0SklRFaWZr6/A3hkBGgQ6IWAKZcBl/mTOmZTN9do9EzNB
fceG2wmFAshIFm7ZirQTnUgwyWM6VVXtVLYd8d5Mg8S9PrOCRDcee7d2atkoX0sQ
jNCgf9Ohh1neYltsX9JmHR53GpKQQF2KbrGqf1+5o6tBf8heyN7Ky0E/5YqLlWa7
f0D/EKOxi7T/SsbiErPROefRzGDXy43+FeA+O66YKxQ8PNXPsqMfGZ4+lhiIHZZC
M0jwxylU4KB4NQQVt0L4TvOyigE0w69Bn9As5aixuuH4DPAW/UEsarQH4ucF5iR3
X46Vb06VhI9xAmwHf+bAY5ieB6Wduh18I2/bag4OOwYVG6hJ6D2uBjRMLsKxXMQo
Rcvc01ipkDWAFO/9+Vp4jPvNWLDeEwDrmmDfu4L/Do2jatQ+f7KvKYIQF0gYRILd
dVp2yJMGYSvLU/0fvuXi9civstHpAISd/IAaZ1hCIJR265ww3z3UD+n0F9bN9lD5
IU00bzHejcHmFe4ynoRiaA/5t6rRhAo/Tidj3iZc5IAtbvASNtXcwJpbH25K6Kun
fvDazsM+nMqwB+sqIhVndgxtz1PBiVl9vzpJbkrPbA8bVXyYwbd6aZgxHmtu0aiA
4N2BeUYrI+B6tu9hXDQUFPWCTl/Wy0i8juMulFAU3ogP5HICfVRruhf+LgG3AMmm
uuzOhye++mcomXbD0zhiK0rvmkavudJboUoEOQfOWHtpR0aCF9gff8tXQIKs0dFo
qi17A/iKBAGhEXPq+VuMjeZqd0v6ZGkphoVYTbBZg268F24fBYS/Wlnz35cc1x+4
Er0zhXs4qLYkcT8JqTBgud4jGzne9lHIn5U+YRAV8usw5kQvUbxBdYZkpAzoddm3
lDcmJWGPslihV3670flGBn7bf79mlcIHRYW+IJfNYN27bUY4fDeX/yCvdE38T1qC
nhK0bIolHVcYh3YNqIYH+e6XtralTU0RwaJGVl25WqTE23YiDthCLy4Txt4DVyyw
uff7LA4U//3+K5LZXhvYPDdF0JrBgJgfpg/+r6So+UNpZoVS1N461PW5ihxRXk2f
9xE9RtBmf0Rv+ViM1szk1aKiN3JZxJdqeOYzC1zidf0sTJcSSLN7BrdjicL5u/OV
EovjWiQziq4X6/oelQHzGxA2URf0vItSkwX2VyYMSit0m8pKNVtzd0KZYBEyYujL
Bj6gTyMLhjTVv61JE0J/bLEQiMS7FFeNxWtzAUlXVkSkXI4gdoI8ePpDf9ZfVV9I
bImJqMN3FQsI64nlFKfImok4Qiuc4cAcqcQ3GecH74S7gMG8GAgZF09aG3ho7P1F
pjHjIWjBiwsHBZEtyKD08vBXnXtP026sZ0pZ8/z9Kt2LCo0ZIQHckTSUQlwyM3Gh
5TQ+8S5rc44xny2pmE8gorAJtQTVSrkyxBKngJM5DkNclIzhz/qvAizP5z4lTwVE
PVtlO0X21pZwDfx33j5a1DiQ0dPV/nOJAZk48yvllC7eHB+nX5R44kUWaq1bOxDw
F5pXwx78ekz998qxJqdEyXnWcNK0Y0g5ickdQxBcyIin09N6q/6iLg/P/ktNgYGU
kJY6/rIIDQKDK9PFom81Q/nZ6fHVwbyKskCclsJhGxZ1QG+nz54xEq/gvsxN9Cjj
UVmYPk6W6vkRVcpMahXpy0rPyqxklxO4NVKAVe7KSAFoFtN+/3iwyc+gC3Omp6cj
5rv0YSRNNDGeil0wDX5H/nwIJT7CJ/4avqqFtW+YHOTISR6hyqZYRun/m3XKYNs+
ukAnpwCKiaKWeNEG3HJX6HF98KPx/7sCd9U0qAwpu6sAT72X93gDxdZz8kNYH5yd
2l42ndMHtwHduiHx52NlrSJMTynoCZd1CfTABx+fLaqRCL562ZdnLtEZaPdqbkY/
nClLtFazHwt8Knvs9hHSf6R+SZ4kONLh5nSAJ87RYlXtjx2aFR1RdkB9Uv3Loo17
EHOfjFVUi5DZlha8z1JR4pOURs0frp51kpp75JRvArFB5Sz+eMKPb+WO85WmNFLF
mR+7BLVOLFm+kSE3TZiMuJReYEfDhn+/6b0UfmUFHKzlBQJsRr9u2Tz51g/Va0O6
SQ/ERkTie0dynnX6Hh3ZwHWbmyXCwbymh8xYDuoF/8wNvBBDVW6DDN4IZNooExa4
boUbfKN0ODjb80JBnF0mpagJ/Q1Bx98m7ctItlG3jB0ga00I/SfPLw0Y6RlvnwKu
n0OMDbH0q8BmlgmBYKtMbotcojAT04Lp85cftYaG1a2myTHtyTgwJ3TyNdmcLdRC
hwJCogRORd/p+1t5r5ywkYxrfOJEh/5uwq+iYaR1lwPCXWFhjU1oauaLJq9CCAh6
alAxu2oihgr6b6tJwrMAU3zZfNY23jyyp2m47t9yrtvUMUzv7sdK0szYz3OoAgW5
T27LbRroq1tVBX+5ILoxyBAdLYSa2xBKSsk21+XJRern8uoYfmDsuuE8rjMMqDYv
EwXYop8wH2nHizBdir2QfQZRW0te/3i1f3f4T5Eodgsket+DSIEcKnLy2nyKV3Jj
EL2gOcvMq3GwyDPfzx9uEcTdFYRAmLcxpdZC9TDc7DeFprzwsY6A67LN6OpFGtRc
J2oPqoKPMjPLlgL31I2V6O03DkBqJapUDLNb6IoqIDIKYjlLI5a1qDgkF16rtWpE
2vv+rkT7Zsw0yaF9hd8lhDfLWaosG0oSYv6QpftVHVXndng8KGRwuQOzz7ESQCQ/
1+T9/mdlSKGENHDqzo1XxctHR/N5rt5ut+QQbvka3Ov4/sIr9Kp8EcpAGH5rE+/y
xu/ZmrUggzH8SLEX1Nzobs4J1s+0EVvQAbM4LAKtpueNzeiFIkCcDRatcmDM01sQ
mznerPYqYPDgrBmaeBMSleOy7swWjW7z7c2Az68CYVU4OK5wGZYlbqWoLTAYrDPO
3v4o8OD9M8t9aAhGSiD1JJIlP2gVLSi/ouqPFawvcg7zallfBD9O8Du3wOGJdthl
cFx668sRgEWFhW9sKGxl4T2Mzpw42VNWA9uLTHH+nz8nXqs2332Syk1aB4PXiABr
0BghUHhEoQ6HBbS9PenSPJiFGs7ctT84KOq0JvEze1VNIyvDke4YqWoJX1XhAYil
Akn53HfKLqcD3SBBOjdAHjUKGsxF9bZfFXCWrmtcNoFZ9g+8iNGjUUgEfWIgVPmK
dXs0TEepuivzsnVhj4Ha0RKxwgLx+AVBTJQB89pAJZ423gTn7TzG+SaBMdvUIu/S
mreXHatUudj1Ksis/PNuRNusPUpIEKQW3dJtrWtHzbOQiY0NykBcgs8z/YXr68uk
hzPbeWh/Kd9I5BUD3ZwvD+SG9qBQCvlSbOtFrf53E8Njltdfy0pV9/4D0GxGLbme
U4b4kokQ/3In2fOKepW7ZuBrcJ/bqp18fHCwaLr/edBqX0x54JCdMx/1LKHtPDIx
ifK/Hp6/nYtRBhbK73zB3qMFNUT6fN5x75gTYEIokSVorznfUITWrZARie3cxXq9
Gf/MvGMAmewMg0T8nsyy9SkoW2obNTBsx1KIGKI74+j4rhwjY0dFf41fYIDjuA0n
EhajPuqn03GgIrkkSWbvsuvrhuMXKLFqR/yPDykE/tPDrecJN+Lk/tDbgfj5C68V
cdx2obRa2iRCoEJKpFE7m6p++TFwzukm2fh8pY4Ab7CYlgCy2Ah5C1+okTLNksOS
V0oAilrxPIXFd7yOvpvrUGoreErrpXP4PbpfQVmTsXFTwaMi461mWY9XBcUiDvDZ
j0Q/QlYKLFXtY4GPd1ir2SZ5jtZfhct0mPXVgkqMiChxInv6CthhyN9Oh1rPTbgw
b2n67LVTl2cn5cHQN8Dp95QPxyyoEPbzT6CjuXZ3kRiqGO8SYeAeAsllw9p294yb
8An8ONPOeWsHd5u689OKiZeuMYjoEVu/T0nDK+QiaOfHt0aK9g9aWOWYlXf9vn3j
A4W0dJxNM8sDgKR4ixUMGS0BGxxoCPPBDqHvMn1hV5R1xIOeyiNgZ8W4YOce0Qdh
xhpxzms+KOJRTtMLIE/3VxhGpvrBLYhcuqdCQOyTZtEWnZFeW2Z60WW8/MQHNfLD
Lpq+UntBHYRn2/fuver+hRRrxsNAqfhNg2Ah2H5EWHGcIw6y5PiMVEpJR8OBzMCZ
IkJU/CK5GDNT/iBh3n0qqqmhPPOB9O4Sr1uBjGmGGoJhO2aOLTgLPR+qi0vl/qWb
HhaF1HZodPjgE/A8Vfw47uMrN4zymipS9eqIVl2mm9z8wBcdGlOGYJ30z5rEWr3u
mpI82jZ2SFQqb9GOIuyklEN+KlmLanryUSRdAor75gBtuMFV6aaWab2nHS+pP0s1
HcwKTqW61EvyPiR6OsY7P2JZAX2A99D5hxfkq89wxZP2Udne2OhXZLw6MHZJA3bq
/ppHZQh8NCNGnuRlsiEBy2LfAelrqjubrWEbnUrrq/MooZRGClgOwo6e2rt0mcfK
tUt5oALjYbTbGQ5qu0EWnKJumUShweASb0HVweDiclegY81J9mIwhpU3tPXLzxUN
sB53QmEP7O1pPzph72nvB2DeDKFki6YGk8+bTFYm5yNrTIScp2E1mcyE2F0AsCKW
MbDFE5/cA9tx0l/YoBaEzDcJN4QvGAhIE/9UJKhOqLEFGzNEC2Yap94gZNjcCVEa
t0JuvwotKEX/4qK0SjWTXc8u7SS8WApi6TQ76vnhPBT0MSzKJKTM7Vmpxzx0aVPC
k221oSMR5uME9zH5lNh20Z50Zpj+bDtkjDt/LLd8wN9yLKle19jUMH9ytYYSV9mu
K6zCJQtx5hO/eKmYVQ79pdloOtnJCSoEKRjINtRl8Hoc4ivsWt9y6VkRfeOa0/WZ
+xLvjLfneDchRmy80ZRQb2tJLeyNt6r4CzzNFQIrMiwjwMmgpRaqMd4jMcBCiFTE
Aa6xGEgOYL/6QKVa9DBvLBYj7CFpOyJoRTZxbxMV2TxPKxbq+kq9CtD1dOLbKizK
4yrtjqngTe3Wd27+vizjywDO5bI9WCUfT7N0zzreqdaFUVXK1dBh728i7dBx8HTZ
C+WKQvpCrtZ7RKsK4BIiaOJ/iiYYRBxCWUnHurKzDBaZlRpOZxXIVFFqbspKeZXX
ROND/7Ln8XtHQuYdRuIEYxz8iDcf57p+uuIzfkFm7ZmYuQwF1Bh7iK7ey+pmvtnd
Hd1r4XDr8qV6WpsBocrarQcCHhxiWN57f077OU2A8nhVzncaAuetGzzHI9WapAKW
7+LkSi2k9MCRH/czbZSGxhT6KD5pCLPlrFY5cTrAdPFPySP1Dq8qZ8bdRdL5MWi6
WaN+EKAcBvZtupz5ohQJZ2jeLsDPc4q6+Z8G3goDwBVBpKMuV1/BDMvXPvA5j0/L
xDmZWrtQOH0gsJ6EyexBgosRiMTyzde4lJfamQdPn76h16OG7B1Eikt81MMsghmF
0Kg1CuhtgmtPTMDq1yYiCeWfU22onN230uvOzkjdadDCEgppiBaBhfqfhf8IIV/6
5dL61hn0atCou2QDpJoL6K4kLuGDVGBmxFD2EHzC0gfk2sgY5+DgDDeymb3kHakS
EmjcSBHY9wiKeK3gb8G26qAZus0hGVYVJwL1nEUPNxIe7zcaVBdjgYQ/DtTHLGxX
AqwXGl/5iL4psZk2uKbaa86Q9tWBv+Hi2jPcDt2VC9L0zQNlLVVh+/BjDaPKs9nx
v4Iw0LeEAaRJtJd4PkGT8S54YVgCrJsQrMXpt4Cj3rBjfiVU9sAQjVUTNMO9UHs5
48gtpDEqd/GadjtjJvUgQCP+4j5GQ0NSwa2n6DMsC/Y8nE+LUftDs6St4gDUMgFv
sD1iuPGYb0R9ywx0xwlWPKCvWV/qNKi+qr8SkHSwwYyOdjvGAfeOX/H6VoDmiGym
h1x3zn6YqlkArnR5XDNNJ6VKMMki3k9+qzw9dha3zPhcxaJZXwfqJxOI0Ppr3T1k
UBPU0OR01QYYgMSjDYc9BBqLgljI4EK3LV9kThMsVJ9CKfnX3EEeCVcJKkB+s0uZ
dQE/GgtLHM8UxYJ8vuqZeQhO4+8VIKR/4V9qXnHEK4yuoYb9X0jgdq59GVQ720ZM
O8aL3hY9mQ31DbBVq+Gh537d14tj9uGKECON75ZWPoi/bXarJzH8fg3sHeq7ekfK
8ZH3EbbGtR7riIndl97VN6TmAfzQuzVSmLrsRUwyI+Tsf6WCYlUv4fuz/7duDOcx
dl99FEaUHfegu44q4I7Q4+/ND2r6kueJaLQu8fGESbmGp0/wSy+TUUPgx64d0HdW
AJ3X71srn7VUiHO6b6pJixoeHYCp/hJRzbjwbW5jH27NNY7pQgwEULCd9rc1VfMV
PIm++vEyVbZbCBoBgV2SQkrQDfEQSgUHSVduGmNUWGB0aGHCHQ6zkRE5p4E5nBIa
YuWe4W5R9Hbc4i69RKDMOt3N2WvA/lM3gfohCHKMId59rJgWawwzOz3PvgIEFGLN
sZve3a6oJ4cFeRJ9lpgFsUVL4PNAAFQ3eA0wAgQhVhSpNVd+PvvpEciKs4LIhroj
DQJv6u/AqRcKlI5WNH0ou9ai7tqfAykXb9CdFL1BDv01xBM3DaZ3eg7MAZyEpAnK
d+GtamHirWUK1ani/thNt+GnNYjRjFuhiJ7SDd1PWf9m7NCq9A3cpCK3bn80n+mP
Ht2w357Bhzwr+80JcofYaWX7fYxV1XlcZC+n07JIYLF0QvP/RYl4NP3CXA0NAnpD
Lajf+/Lcd8jifD3Eu2I1DwRlF1bYUETLl+REFLp0GPXMoRL8K/vCqClKIc03H+fy
Rl4+zlKegGQM+U4myQwZwPWmO6k+oEN2q4pPcYlXuqnxjmfgjDivtenhpeN/h8G8
Kf1mvBa5yma0KE1pJR4b2bkvyhx3q5UQo8EwthW4Nz4cpvD4JkSI2TFvUgHRkD9k
dNVDM/t7F31uth6qbyTKOjKhGHDan4yvuYPwQdgqpujcdSVkoADu5i9awsVnMA7n
8FWe5yC6Tb1gMLrICI2gWu2KR+UQq68lPlfdos6Rv2eo87sVuO3hfkeFvf2bYq8H
vOAhMDl/K825y3bfS6RkocutVT3ziCza3P3M7tMSQTPOtqvkq9egRea9n6PGVwpK
Z4vk1le/V9ToMV9lnNnbCo64GFG+pnLkjTGZIb0SImubeMgi4xt0+Dc2JmP0lHQB
6m7IN2fxA9/eQuN+ltvfLUGXjjNQYdXNJ3KqNNUMX+7rrcp08c74AGcz+RetwvT3
bbIEYskW0fOFitSmHbZwtZYmvhLD1OEoAhHAi4QKk8W4r6stpFVymrRGGGTJI3Z8
F4sDz9g9/VDCcPigihDx6xgNW2qwrg6o7hMsQFILeHsl1g4MEZ2zzmTa+SKKsihi
SKMipdmywHFExD1hoHe5JgsdIAe6GTD59VrhK7verChHgfFPmLZtebEv7zsxb3yE
2+qaeKW01pGNvB5zJfdRJJ83catHbdJJe0wR56L8qmAohnVaOL2TM4f8V54kJIGy
UzbxoCJL7W292YEdewsW7PUineLdxOOCUNbzVe9qTEPPzT1bg3X0x2viD5nUNYL4
05o61f/NGwGTb0H7rVA6uEDIitV6FgXiw7Q1vQBVa2w8fzpuCTgT+nCghS+uEv4p
jAo2Edn9rHAJHmr5WiJzZWIMLxO2WKoVmd2icSO9aV8ouLzR1JlFhI+wQOreRy+X
ZWmUcdFYL60zfucRlb7WDLf9xpJ03gr22yJObLHGhw7E04wITj+bEwa2z3pZTPFL
bHJnA0SREaqcyncKd8Qi9Zqnc6JtjApX8f3bKx5rGpwMrh5u9HuL1iNX+L6NrfY4
yzHBBXzy6kfgzOjTKPz8MdznEDXkdiSRrWAD33Ni5Trtx9X1G6f3+SYI+XLQdyvL
lx7cgJI9hCKWAmkCVixlPCZqc5p0P3f/bdQt8OxkX0tEKKyqWIlkj/BfPUyOo3w4
vf51p2WPTcfTXc/OPkF+/qDky9JDJIMSCvkPs/yp2ZMHvXLQG+urw1RyTo+nX/sJ
SlqrUnUcg0wS8lENZz1WoUHYJ+hLWjX7Cgcmas91k/R6R+K4w405ktwFBbtzq3Ta
+G3Dk1eWU8CqXyRcpFbaQlBntzM85ybVuCLmX7TVYolW5QvhIzmevxs3oDrGdBvb
RcOh5iZtDbmi2eUNB00TXLTDTHvcmOfxlxYRWJKSA52cMEC4BS58dWtlbKgsXMBc
o71WB4iy548AoKM0+OxA4DpByFg+OC4ww/VKIwtNX4Mo3E6enO/4E51D/PnDj8cM
Ie9GehRbIa0eSVSnJXu6Gz7juNWCaDmIT9ZETZTDgKNfxnVsOdKgQfOLqH/sBiPK
5UhAWUi9kM6k32zKAFU9UH7SCxHTTVr0FPsv6GsAaZj0EbMczovQ1DY/UUt5p+0B
M8XTyD3a/qXNEX1c/8mUGZFuB2qpYpWYJY+7HAq6fn2h/34TIJ9wfE+dKfulzHZE
t4eddAjeWpDB0PgWBcJLYJ4O0UFgazbOTynaLgxWhAOZoi6sA/VbzStIuxxZZTyw
RpQ9axZJ4uazKX+Qsz0uSY5yZP1BbiyxSM1+t9CUBrHheg0uTuCtr9wPEI0zIhNE
cEH/7svIzdP+gJxmJxqKlu1WH5GTKz5G2wlfkAdRZoQtUSWX/Q33qWdST9UySLuP
lVjpKz5qexunJhA61BhHTCPLCHXKecSmmPS/HSq64zR3TuACr3nB31KQ2ldkou8f
XpPgioOzYoe/iF1f11ZljKqg5wKtEI9DVzkKdZcaCwZLGZfdOdKDeOOHcip4xr5h
Bb+FTNVvSnaIOTvX6ShixouXCNIy5iYrefuKot897BoAqkwfOlHeNFZvgPJ8/hzD
TLwIdeodrYGFobe0BYxo1IIp42DHD5jgTVwMJu6okFPA+erukp873Spp0fGxx8E+
wl0c4StuUoUtRiZzjp5bdCujdosLdQEPzFxqJg6drExCjaziILDrGS0H6hJmYRZc
3iR3xYXW4j+Hramv2pZ7+AkQnqfcmzq9urRkGZ50LtXYDv2gqc6rlq9vPhsM4s+i
rWfilH0nI4FA0mHqKb+dFj/25VxpS6zbyoxzO5MNXB9yGZYmpf1bhPmR/5WM2HxN
3Xv/6DLbq5zjhCOa4g+3rROm0bBCgS8ppnF5gkjgy3os+ZiBUY0LRTFa5hxZymw3
t9OEVDJBbPF0TbQE+ty0GdWxLBONtSj7leQKoGH2h3Xe+BKpny4d07/Rxrf3ku7V
uaNTqDu4ecaq8YYJ6jA2P0oQ6JrPFvGYjqv7wGwS+8qlIM2TDRy0tCIkuI2pZNHS
aG7iivmM3sYg4tAuV0SfoOkHQFOQRmOWqQNt2L5P4qusnUJNI2aBKFFzvjT79OtS
hhpLnGVn5sh+V3DclOgDZLfYepkM/RTPfzV6T2FBZ/nXYp0dVuZWAylmzUQAJgDX
3lUCvWipLs87oFI4S5LNRI5IR82Ya/dgGHT/3VpRwf7/yY+eKj35yIk2cfO6ssWh
vxGvthi1BSME4XXgUwXuPTzSOOlYIDtrXio+PbNxBMFuyERmx7L+Z4iKJxbgSlPJ
yvPKXwKczLUQBwrscU+WGT3zlItfX59ZgnsslwShoECY4RsYVKTpEYuKwYTLEG7l
hAuV86KWxa6CK8QMQqlrPfC1E5D3XYm34QzqhifW6LvxKwDPF04SRyC5WCmN0j6l
2qymGnO3mCjOM2KtBKW56Rrs84JpZGl3ROIpd/CzLtaDy9QTUmC0FgEQUF/ZVQ/H
EPOWyEJtK6WidFOeAXJvWYigErFTK0gumPXKRmLbVkNZBxkKyPxz2gEpk8iiQ7sg
QBct3gO46sC07d0rKXAwUHSNoTg0ZxpvWqhst6EHCQB1wFLSeFpWmtBFGf3vf7s7
uMPb2SFUTJkgrtPK0a8GrJpD5hv0WM/LB0l6PrIdJIP/52qIdJT0HYkhUw9MGXvm
iuMRnFNmzJe6zXO+qgoexcclOZW+1BuE5xWKuM+LBJjmma7BUd19M9L7gAR4GAiL
ZTJ0KNHwfh79oTTgd5Xyi9vkaaZNM6xLInXxsCu0Sq5O+VZFUpSy0uUFXxaeQqcH
rkBIL7zuT8BAyjmcoeRBovLy3BVT0dCU9glpV7dVD0NKvOGX/MlgDMGPzP/WWecx
lNVBD35ZG5iywrq2xQxRv/bcXSO3/f0c79lvnPFEKTIe1oh/YOjjK3jhcjfZFY84
pg3h23H2jsU3+rAXy0o4TLq2FKy7LuOA57fCGidOukHy3OIDkM2CAcjBSwlOiovA
Hlfz2IvRiKiMz9crvcbuMIcURzc+RNV25/G06LvSEm9qZ1Lx05JQo6wgJZKmwrvb
tUoXZimjoJ9dNmd9i7VjV6O4hWzKyAW5Gu4jzC7DwmAP7ICsa9cPpWo4QSUJtIzK
TVhQq6uGO3s2gh3n4gCg5kL6xl9H2RDQFArkI4dIfAgmiX48XTA69gc6EHL6gFJB
PiYYxCqm7B99rrHHURZWavLWT1ABkU8UH7z5CsW6gTvuhMGJWGZLGc3o1fhi3VGf
bGfw1iBMBUvcMppKivFe7pEfnSux7evw0ID1huKVwSHxAeS3utFtwi1Nz+1HpvGp
39c/UUsQ22bzNyYIEeuEYq0QhgTb5bDpAFSOo53T4yMpLMJ4zbpIhxtmz/2TjlGH
EIkaQfixqVxIJOcuK3Pz7OJ50NValQ6oKcGa0PtE1i/7bMheSd0FLv+tMf0TTKrZ
zmKRU9aOyG2bnGPqcW1255NX6DpR+IFxUR/AYcHAH/70PnFNDOTRQffSqhELhRi5
IvFQiSqE1Zi0BPSTeGwE/b5kg2yaD3nH5icUtvHj926JKVCn6uG4hQUfdQRUK3BR
KlVjBzkhqhc33KDRoLGtgb0tdeeIrk80D52IfK2OFEt5MfiEASiFuPHJQsbSW9VJ
N99WkYZmMlZ0eQYRLq1ptRXNuY81i1VYVVDifd8Sj3WIAPwyMdCtZJScbZFo4zs3
f2Pvf6VQc673Tr1cumiqM/Mpb81mTinHLVGkGf5nmY8blG/my488vzEC1tpM0OY7
9ruikM1Un3VcbnSXRfn4GXXbIdR4sd+mpsMFEZO0mseujEXWr53bUMql9fluw2yX
mmb/QAjhIeyaY0q6s3wUvGVSZnsx73dR0PNq0pE/QxM9ONyyVXI2xBR66ePcZ5iL
3soD5J6tm0vtjuCwIATc57/Kkznu26/kHJ4UkSS+DwVyw+Fu4+fJq0Q6/DhBaOq5
z7hzAywjpIoye0sMQtvfWi0yiPLSCVq+EJro+nkDVtUkAlB/RgLYidxQq1zgl87L
bo319e079Rt8pb8gQMUcTr94R/SdlLvy8z+XzEtgUxTVKbXf+oB3xo3U38+Xb1pj
R2etarjgfY6SbGbzkI2I+kGsmvsMDKgQ6oeIj6qN/UQC6A8YBs7y6fq87HM2EJmT
+ahwD4IlsUl1jS3bGO3bUeN1qrETgHs3UqkvFpLHXY6Oeo89TUDXSKdKqrWo0GFs
1t3lnYAePZ+8O728aOuVcBO/tu2KZ/mv5BMuKAC5/49on8b+gdua+h9d7qlJ8S6F
6MgXWm86WpijnQzc5xBLJvy9h9MpM52v1sEWMU2ZcJqAgNUET82AHM3ZTES2Ced1
2BAaYl0GWcTa2MoXGd55xTtaTzVzSOaDzQ5+7Coah/TsGiPRul9yQp8cPdaht2gC
FZs72XrFdyxViKzm916t15dBfl3jROx6zzyiUylBWUJPr9mEMYV0gsGBH1apix0W
9AmzNj+rEDw6Zu8VQDiEttrvsYLr/wj151yZr+Jk5btw0SkNonbt4ZpsCGyaunNH
yoPg/KzMi/1Ggp418a/Nosb/QaYgEyOU0m4WF4sy6GVbcXU8/WpH5DSrvy8Tgm49
S2jSg4pzywh/Fk8alHUR2V+FP5dOHytyApriawnIN0YZbNPc68CscXVoURh7WI73
q0n5Z9DWgzKNiasS2uHgJHDODea0yJxGnGIa8GbCI8LYQrx6RlbmePjccQNNwdE0
GrzdGIU3EsFJZpYe5mwnSlKkLRl7WkIsNAqWG3w5+FA84eZAAJOwwoubxGNct7Db
eJ/b1dFbwRzG79CfMntQAB6e4rClw6UgsV7D/x0SmF0wAgQ6Onjsm0oh81jwY69K
gnq/sXnv8hOF3IL46K4IeMCzE8Q6cjnRWpOp3fMN+fhqkJTy8q7N1ZMPgXADwCYV
HefuKguUASifF7gP7pIjhxK2CAORgZjXPcUGYPvLiLcr4XWbvTWqmuTPuF4gJVZA
w5HcCHLYsUM59eOY1WrvVW2gIEQd9vzsYHZw5Ft5JIyra9UcSDMVliPwEsDCQcua
H/9IFWaHBTsmS6dL9kHNWIsoMEBBGvgmrsri6cUpTq4wZff2N+d603BPGzK5Z+rs
YOFEapocuxXw5kijyjhqkQH2NG+vxM3h4JaZwoCop8Sc8XBvOQZw2uNiHro1ML2w
7S8IGicVvUDRIQ74HiURDhOMFuD4ydOb4ApgxJL4Gzkv7hv7hOzMooq7Jze/KBXl
ABD163Oh5cq8F7c4o2xA2CqLkr9cmhNdyHUfxsIK79+IIpRkKRKm63w1B97OaYno
e3uHQFSzEmZHUAr2yZvPvhQHNxPJzRifSP2d+UFpDHTiVQJRMlO7UNTKJ69zwYNx
LYf2akfSdvEv29iCcBoRtlCvthMKAkFADEB1WkV1+5ccNEtvEZaZ+zqr7akbT/WM
XHbL5rpZQtsaG0rtnCGFVivkQHouIHdfwagsrsma3UkNPdYnq/xl2HSES/uDRDHC
ieg1fIbfjY3DdFVQbr4t0RRin8UVBJ9pBoL3rG0ZQzh7A673cQn/d9N2j11RdSHL
62b2Plj6AqDyTqYmCLU5gZT4pso9UhBQm4gIjNKEfsP8xI281HvIe0lf2y+TfyTL
wZPTjZUiMPwLcEgvQlJpPjQiYUTAuZORucj+peQ1vqcNq7tbcEkVsfAVUyuMOf4a
3yJbNyZYD1Qb7qzrs9Qxhg8flb5j10Gn9DLyrjPKSwgaLbhzbJzVn2XBKMpcVPUG
QUS+777T8IGzpRqS/yK+zmY/AKCdnPDUje/a3CSehDgURP47MgRiVAGPojG+tgRQ
c5gjUKXhpUWfPCDE+cZWQDHzx4QTtJG6M68a12txtgHJel7phtMRzar4Pn2agisu
qbKgZvXNlcV6m3V5B6sz5AT/4vmCNBsQUcwbmKPP+pt1SN6HDMPH1jLCwRjIDK60
Ox4P7H1qS4bd2l8JqfgR+Br9ldFJx4DMi1KwUNJ2UL02mQV27e5f8fYH7WYSft1/
MIQ/epL45y5SI4MN1t5oOWYz07K+rzLLubdhPyU+fdpk2SbGIZ2DEcefoHcIuVbO
v3ZHnvDtWaUQ9SWCSFy0kqelZ8AeDQsJ66NMdxostmL6R9Y4ChHH95gdj0xdGedM
+pddLV8a0lHe9n4D8++CrDS5eNgvPUEM+U7yFo4Nf8mtAA700seTn0OmqxqoMMA1
fxxpLZEoft5zvhMdT5eTDGKjxf2m1E4V61DHCHlxZcrGHy3yub8iRacJofww+k7P
bDBDBm8do6oD+MKvprOAl490HK8Pu0gTYfS1mMNx+wbszuSaVVs4Ccwb3KpDr6Zh
g7dpRl+NYYp36m6WhjkFJbAGhUGv+yhwNwHM9uJPaYJjgOyR1PBonQJdCFogdHKy
e4ynP5oY56ZBuh6xhk2zZbfV4fF8xFnfyUDYIQGHotMuHojJoVRk139CyuIGdp3e
EZSWyKJIfbw+a6WKWtAvAg4AHoWMts1FPKrmSTyTLPLMrBEE4PwpBYUESWWh+jmE
3n+I2ujnDe4M67b+iI+BKqDhnslGthnvpboB44mBKLRUcARQZfSLH6LgwplCDwgf
eXmrCFDcNFM4/qDGYfz08QcF/DHyXxDrZUKg6aUkJUm3m2oHieaPe9DpmzVUPDzT
yklxk+KmnUJMTAgI5yngZaGS2dIoHvkEBn11Rw9Y6ZgsoLqTpp4qJyykGFvjojcl
NNsqCKIitFd5yZWKjUZsjXdNtlX5CxWRXvXdBPtzx3OprtasXO0Fw6bgmsSUxK6x
h8xicUAICW7vqvh16/wfwwePRj5UCEzbn2ticM5lbLdoX1blzODQfav/dVsC3NxG
GEM6b4eDMKTqxiBoz7Yp4zXs8GysykdxjO7xSuB7leOEROXa4NCTSQ6KYTLQgi9N
0JW57UayXeZdnYRBxEIAwXLGIhJAGDrE5j1Nqn6r4uzbGOjWStrpfwMCMBK73iV0
v/c1KWKxpEb/WoPE/gwuG0s5BdNKJhDcnjG/77kkZ+8OE+GatXzS0wMhcTf+1wAi
K15qn86Y7aKSgSCBW6wt6sfXYk61l8ZebprHg20o3k03nkI2iCeqh/oTwW90CQqX
g3dxoZwOC3TAKG10Ow13e2JKt0EuaIylhTI5nSBZkWQ7okpJvJl2WQ9qzB4LUEja
pLwNQvYbkq/d1To2M1cKv/Gd/zanFyQehf3xHJ5SXIgIzbVdbWyYRBx7goAPQxFC
iEpkAtRXy2Hj2JOB9SAItV5Na7scwck+PTiBqDhuTDvtxVVGQWI5PzcOyQa7bYGT
hPLbhR34/GhxTFaZ+KPy/Igti25ofRz9ivQl8MQd0ydTfLkqd1iQvjcp5w6Cp9Pt
jyc/xLp89djqW2UM0hnQfrUlW7JlutXxBwN34mcZZeNTNrCJ/jTjf3lrhPwqxa4Z
vcPr4PHQAdrCnZzgrZ7WR1orlCrWPegfH6xOiOC28Lz/1c/RUwQ7lxZPK0t91zBq
WNHwdzMmlxRaVCbsP9nS7iP6QGa1+IKP+DnrrawIyEGAcbUxPJH7e55jpd//J4H9
eO3RqUnYywDWXd6qFJjgpKfOmevNwjVLfYDqU6F0mAMQiNBPXoPbD/ghvRN5ScBG
b2WkZDGSW070qdCskEsXPJonWQqZJHqAJXDP4CFhs5UA2cKcnihf921AVJsAdxCt
CkgapZtSB2ETCoanhdXUPP67SfgcsxJ3jUz5XP804fAtrZDl1CBUguZ8Kk6971UF
bD3Lr2pfWvaqBZAhAwCkW8ou6ZY4BAe0UlLQWtYBLia9UKA1o9ijXcvd90Si0nJD
/GQnlKZiuuUSXP4zp+3lBRM6WD1ix1nrUzOJGZNHJpys2YQD/ItKHSRxrhmPnS+O
TjaPyckUWULaR3kbX0mR4rapFwsLP9kBLC1JHbLs4buyOLTnMXdqj3u3ecZbx9P0
iH2MqEP9oSZloPauoYx084fYigWbeI7SM07yhDzgxQ9C6N/SmtZD7kl+l34RKWFS
hcjGaFVt/DAHsmzviUlIbFpFFdrmVlLTZliDsM94URaK8xZJvurHJDWh+Dlm9X9F
MLPwQViKbwUrLgKpUzp9uahNisTF7qe16dxkEAgIKJkypdBAory6OoYEGPQZ5rYN
PFqZH4xiOFhkZ6oe67lsRXS/Nv6//ygBhltfxkhKxvm+kvLkfvsSUZW7Wj0AvYwl
uup9PMs4atByVXSvXMLCx6oOpEjxQJyW/EPdxISb/JpIlS07+JNIQefCdlzjJlk2
bQrmxEi9EvGjYG3sndtr+YCHApzwOWS0tZMgw7u3ak/UcXe/isWAfvmufJNbCSw1
wty3LUH/4chCruQOC/adavx5HPPPW+oKl4qsWBzufgCReTN6tj4d4LOmlYm+yM56
FoJmySgQxAru1eaXHd7x+jEbG1N/gid6/C5RlUhW5/C747ogR6McAiu+nvU30lcE
HBJbMVgkIQ5SjjQvdT3thWbMdajwU/JWnKAllvoL3MD7RPiJDcPvxcPJy7yacogZ
yGApJMq2P3nhGcFnej5MgqNqhr1UXSIEw7qznz4kajAmRiTIoVttCXtMPQmx2Bii
gCHoKcltSFhEi8fyR4M7/ucw9dD2VcL9CWgxB42BrhgdUfaMIfkj9iUexeVPOHhL
uVc8gl0IBBVZcLT1A0n9y6GGK0hr9439SQ0GD83wwUTrYjoXgQSj6tWX4KmwGMVE
tLqqv/ilpD2MDOCu8yn4sr9apkOwEyPPMPqEXCKllMqmZFvGfpgsvZd8N+GsMLXj
8dd2mQrJmm3jTWlFe1674YlFcYiWS9b3HTjy3f9PedM1gBuONbctGGKkf0s5ASNj
3oXgFLhjmZ415bVpEelV7E64mw6r10blqfKzFLBucKLNMVeudS35mvsUjMVuf2MD
gJkSTBu2TBMmPuMJcT6CGiERaIgxKqvYVZ3NvzBCTqnqyBJq6I/sMayZLjtnlmV8
sJVSRvi2f0KMhkuHTjMN91V6zEL7on+9OesQ+ie3ACg4gfS1y1ZLTW3EPo/ibefL
ZOHddt5BJP3EfSWv2FAQM5cd56GakLl0Jz3trZiYrhvgff1vx8nS4CYta9h60pQh
RMqLw9IYpQNFO1/iLpK+sWY//NbaggH/fqyfp501D50+gqZID7QbhUPVXNQjgPP6
Cq4+9CBnyLhtw1EoHXafwOVGbgki096FKfG+OnM89fvbrFkDEa1/yrhu5ybRoAwW
Drp8WDu3F9MJZvBwEAG4Y70dDOUC87HdbdBmqx66lqLtaz2wy5foojAIZRxiUhOs
bVGSPVsSeFb17HBHkENUv+Yi8HGu1jIOqplAeI1p5vTZo3SUHWpNMK6SZmMrQORU
zoMWDty/p23zYSHmj5/KXwRqBlhlbY+ZVsQ5P64ADBLId6TFI0NBbVSOiQui0kr2
GLT/vRoGTZp1kg2b7HBNn82tBJ+7FrOIXooBRih3u0TGiCtmhzggmIremupyWwd2
b7lWVYXyw4ZObKziTChCBA81I23xhkZVTe7ixG5nW7Gtc1celvhLiA3D2m5zLscM
KoOAWJ6jTDEwb8LejKgKFpZbBGWS58Xll19HDXZYgPTg3LaIsejlkkxInGU/G+Ii
dlfwjKn39H3lHR2b4MDBOVVjQlJVL61SrPyFlOsiBFbEgqEEIu9V0PucpwoG5Us3
vuXlQ0YC+Vw83IlNDkvfL9RA7GPPTok9YA8bM8xxWJuKAOX8S10Hyk12soqAGzzT
TpLhWwBQkqLk+n1coG4Uh2JInzCXSusLvvPri8An0M+kpCw0h7DtATeGet16CzLD
DngIuHxR5D9BynNbdU06rWFVy0Y3Rl4rfZvVh/UIfoLf/UOzKcVR/Oow236AFpcU
BdspOidQHgJOgi4/1ooCHpjHXSRW2h27P5LgJ2FqLhIcTGKuPtpfnO36/pCg6gGh
tZ7JF0RPP65rMUVgC4bkB7SuhWLRinmrEcK0ZxGPhZDlCUPeRVhjKJPjBQB83CKP
cBdr46ql+JipdA9YzFOsKjms/DFZ9Yq4zWuMDlmSvKWzOqBjaW9es2nTkYZIx07D
sKYraDHELQPxaSNzstpYkqmmgMB1QBt00MGD8HbTMCDGHixDdbL9AEa4ivX+LMM9
8rl7zFhyQOqIUR/t+mnrgBicVwojiogPua0Nz3clGzP4LO+w5UbGL3YFUeeqKTCa
3I/GRQ4l12NCo6SF+Xu7oojc6UUa12pSOrmVRY9FCwL11iQvoN7nkNQv3Hj7pf68
XaYgprMtVUO6u4IpnmNb0dPiIZVS92+nzICDfSh98oemPoOB1/oCxXXEXvW0nvrh
tFI57+TL7MnuNNi9LdiHxpfZNq0WSrJB1JGq2A/dHGruKRRo8hhhYWk5ypwuSJgD
xCFOTJgqTeAilqzyzvn3twgcycEytm7MYqvW4p7jaUXiCLfgcduD9Uu3VI7sewRP
kvePUpisYiFCp8EdUVyuOxHchybJid5IqMkuANktoo9VQULMMsukrJDzwGrTZRwI
vwYu/cvVA1I21oT8UwaDL4jQ0nGTy3eThUla0k3IdxVr3tZFGaE19fgkgxttgQ8p
0svoXHuLMeeuZJZ+dSw9SVrDxpdXYW947N1VdQkVjshyW5DCcNEnvqFdSe4dksah
LhVQeZELwhM8xV0HQujFMrrYoMZD3191vGG5kEI7OGT673YO1QbYLLUJcy7n9CqC
29T+JGeoBVuT4Jwe1YiTBKK/Bt1qnYAMv+EEP4J93/0YaKTCNRoXBkUjkdmm2V8w
uB+kgFBR2tet/z1H+MQEwkGp1SrxhI18F+iPQLYCETZhUk17YsIeYCH39qIh8k3s
Fzv9w0LYTd+b3vCr1lGOmEfdXtPm7ogCfjMUABEIUWUjsnAX/nTnqLWxvfwsAjSX
DmCznsWTpvvnDYJeS69KAFQuNOKdWNtkprTKpsobXf+wUexqBO1tzjaV7sWwDCUJ
xFtGrADzG0XOtxMJNT81QVsUgSTyAazdJa2t9QtPNXbCEOkfT5Odh3pX49DA1b3J
eag4D90jq6RLVCTo6rebqJhF6sm6L0tLdCHs0qendlqs5Q63tdV+u6KYD03WzBvG
9u3aqBUMd5gFub4HPzRqlHtBMbumbea23QL6qFDqufjC2MeVxXT2+BWmsOvt6wng
wpUw3Tq3LBs0MORhIkAy0AOvVS9nXbMeOGfJMCI1MHsor6QVEsyrUrQiEYaY9Hfd
Zpdo1F1RacFaAybJmOhnrV60R3/ErF/Xau61Zbn9iGH36OwF+hdk+TcPhiPt/dQH
Uhu8R5rl4rJYW+ncNW7brKNesGluiS+SjO/9XMp4cKFDnM2bGsTlqsYTuUyS3h9V
bXFQ0jRoFnc1+x4LkeH/JZn+l6cnbSQ6FUZVxJGwFpHzQyDFYVEjqGyjn7B8O84m
f5tJu9h8X2F4v7LaXP7FTkLMOluCF9V+VCjmNaC9xIB+PWabyeqZCIXOmKdT43km
gjWGSYsXl0lfDqCcsJRTGjSQNLb2CqmCbO+VW9FsgpLkKh5ImxavmfI0dI7M+G8T
ffYPYEPr/kj2JadVVkBcOvagmkK4k5YazZ8vfRMWuMSgc810LDa4r2jeNTCztKTe
X3BrHgmgk1rLM39ISwF1Ag3xH50sRowEPxnTIHmQgQKoD3/9SL7L+ClYSwsBPOdV
wM1x7Fh/2YyVri7rVv74WEGYppC+i6SM2/ipwCxw26sK0WUE1IkPgAnj/5G+BYHQ
WU/bB6/DVKl1b/x0dQVVExmUGNiQLYzpIFEhbkC9vPD9jPdgqVLUyjgy55iGjPAT
1VzsE9oApYAc+HUfTRETvSvnxmFL9WGTg0EMuRXbqbisk79h44aB2h5v5m2terrK
9Ta6VU368bJYX1GjOOyDH0xcxSSmpz6K1CgAvcPCGKF3hB9f+aE7plGzhXfTFse3
R7FD/VuobCBQ8K9qyDLStReEmSykAyn2D64xF/AHLkxVy6ar3d4KKwcGVqkUWSKZ
HZaFpgXI9RWvwMEE/6K63h3qvtaRWeG47TyTT8EaZrg1Ujz4/AglNafmLYV+HoQe
SqDhnz3atg/Y0gcYrcSwS1R6+ivGJdG44wG/82IAp9fJpjlrkVLh4540Kl2zcqyG
Ux3b3xgs/Goc3vBJaP8PJJ4wGHYmxVMmQdHKBgaGSHPIdItLO4Becp1f8+5KcGxH
cJooY2yLqkWdRM+ehF4hA6+iNfkSl+aeDiRAOWI/TPZRjcsVJ1W4zz5mDhUP+mcH
6rNDhBHQtFdOdls9ZOU6vdwmBhCeEnP0EFcfKsxszZ6fjmTJT3ASugYpdGRZJLy1
MEFSF9wVrHch4DHCxATEjd2wFjjkp40HoiRbRR+zyi3A39lknyo8tICnuuzFjQpK
ztlk/KckFgeYfc4dS6ZP79+eWp7RScxTs5vFH60K46Gti52mVRHgD7NMPdEW0h3w
MknhqFXG1Xx20482LxqPTf//OSV7JaGRNXa6B2gOMgHdatw5PIvo6Fiby4FUqS/c
K7xCtQpH2HAz4Wsf7+gdtlGBtEtW7++b/wpM/jdF0H3UrCLeuJptqsNWVtDI+4q0
erG25pJ3jTHcBWMuImk5VMegIljOZRmuVZnHujkIHAvc8iuWolGC8U19Z7PEDoyk
DriaEg1M0r5K6bAL8J/6SZ7fi1v+n+vxz53442+a3Q2NIasDLwv6+/y4HnS3afkJ
Pz1nSkVCGBEqphFxzR79n/j2eN3X6lgam3HfZWOkI+jOV13kjOuKIzzW/BrppD6l
GpZoDYIogjDgkEsDjkJAVnMh9/jLBg9XvIoW5B4m8r64ovmHVNgcyWZTGSQUkTJC
VINu/b1uv+XXjn1HVtxNemN1B0WKSLB8VsU06eJDLaFrH4GUmGUN2xhE8HxSSimx
PBY9BJx/QUkcTNNx2z6xPtvA/MM6yqn+F1EpR58G3wV7DQPwNsfTbY6G3GsMfZb2
7cl1YjkC4+tJ8Yfym8YkHa0qR9wQFGofG47vuElpVqtDRg5s13FloDnvzQRhqNCZ
9na6YBJZZ36WZ9xP4Kf4UQhJrSNk81t5ZLb1hc+x6bLZBN7D3vgR8ymzcDZ2uh5i
6s3Yk6YKUm8vZb6B5h4s/YdIgFxJQ9sOANq2RmqQshanEoKJ2/X4jaCB2sxTaRTZ
SQ+0B1Xk1WalpUrHJOS8LwQKtIVae/lufSzW3zhtFiUHc2JP0JRekMV41h1jhVih
DCjlwSZPknAYQFPQkOWt1Qi4c9l1QKDqwkRNYKMTLshQHAGjxFHlUBRi0yLRAxS9
La23V7XB97LL4JL/YtW3BdL0/K/P+/Fyhf2N3FUJ3j6TlryikncPFGeAi/Ffker1
5ndAxch9ReryoGmC6l/J4iM70e5nigIv0cpA9mXHqq0Z0bbvBHrf3A51isqD0Kxx
IoFvq3v4lWHbItznS2oUbp9oW6nRV+lkYSogzLqA2zSiCV21520HWVcmYsOXXyGv
GlhuSeCmOz/CLytxZiNeAjYbHDllbFWGCfwQKBQkYhrfknnPJqErYEk+xdwt8Vfx
iJoVmkhYaSldYa7vK42uUCjmrdfoVp+j4guYHOMctbJqjNsKrl0H+EaLUpXL+44E
n4WRbICa0U5RNhefQ+8Tv1Ejni1RLa4rxnP3KmC+yXaqQKc7ll20TCV0gU0mp9Ne
jdX69NFGG3fCbs/dZxjDf0YnD8CLqshsjoViEPP/7ZXml+VjGrdMbE1dkkagO8Zx
6/mRIStkD2OvmcHyYSXmLNTjQFacQqMkzZa+2YW8ELCncCGxqwvOCgjKF9dBvibl
P20Em9Q8EvYIoA9Pup2TZT8Ck2sfN6Z9CiDu2Q1kdTSnZ40JcPKGM1Ng6JxrroOq
bWxd+jAHEyhVy9tzhEOljI5BYwk7HWFVIcOZ8ufrGl+iPzZeAvVhv2MLGvoCFKvC
9FZWUpFQqEIrSP0BTz1HwEvKmyDs/DbyM/cwDu9wK7hmYngAQQnq6BOb6vLl/JZU
p7sNk84kug3kU3u2q2jIagZtGA3bvFs9bpQFRV+IZUq0cbOv9zMBaF616VpQ1ZaY
RWP3bjtpqn/ZcOe5sii7VATQ4HTW6YG/CGrpfR8HGBmz7UGsraqQqS84pzfFCt7J
nFb2cyxNklLo4OpjcMjfRvkrW0vfVCoxUt09XkdhcLh4sQbZZbJ2lX+r1qtXjvpU
zG3RuBRXaGEEpRwHa/XhM5LCxl9dAj/DklR00wy2EByEOOa01UWfBNLHTj13piyg
0AyD9vTVwQXyXj48DlNlMe3GDB7SNGG3dCIzWYlbDQSMdpewuIn/fMqPZcEMnDmQ
+RTudWmJMC6eL//YMT/zD+aNDXyBdLnV3bo9Gbtsa7S0QPBdGm09sW87FYAio6yP
NryL0KFRIlCdvXe+U1qOADnniBObiZigqbTQzTMF9aDBmeWIL2ip/+HM/PDSuDQa
1EQmsMP9Lnry3Hff7eUiX5uKVZrYURnvvOLFtlFOqVZtNJowD8ujfLiLqk8ex8bf
2aaUtjb/iO8DcEiLxHgB9Pf7h62PWnhl+fU/pmxYnm4g1meCW1+YnYGSKIgzALEt
L1grq1L45s6B3tqMYeoyWnWGEm0ouAakhcUJZYs1MoHPZxCIYnp73MS/zUOEbNqt
lGbvyZlAlg8VyNcLan8DiYl9YP6JJyX5/PXZFT5YTdVZim8HfXoyZXAmzWQhbJQJ
n2rS737sAW/W33dta/TB4IQQ9IjCa0P/w8baoXyuiZ9Nv15w3l9rBRosf4DbHN+x
B65TnCCExtXuAJy5F0f+WaAPGgI+qhAdaU3+AmG8zm/xbNomY8a6Qc24MiWfswz4
L+OojzIJj48fqM1Bs38Zpywfo4qNM9oDJhdb2/8xtJLVfLys+PznGtoa7CY0PvTw
ZosLFAXoefPCt0y9Y4bT2asm2WZFbaJIv39HAuDTu6TAM+CoQ1EQ3ZOoUBPC+ssm
2lZ5Q8qBjqvn17ItQYHeIrmNnxuEdxuHDTFuKsdSI3Bi1h3EiPvHXglmZFOfK7W3
v+ltsObfyZZ44bw3tKjrkPkrJWYPOtdexcKq6y4q+FaSBDaiJr6Zs7nTzWjRsJzb
XLZHmk2HB/CFSqFWw/pQnogVS5mQ0oVOxEM3x38gL2qL2HutuGEZlLo3/IHQ7kwP
UtTw6e9FlRzLEfi5kmWZFN6/xDrR0F1plyXzIJ5MmtPr6B8q4DCsEtuzm+612cq9
jfb++zebq9eM2YEoTozjjkcNuZ8STMteISnudiy8ur4E0GC1zXjhZz84oFOAltNs
hzkktzX0aDV4LD6W/du19cinT1U6yB+tzE/DOlTVXVQLdPA+vREUYk9vlBvuFMhb
GQ+cdQ0PtZnelZ/zIcl3OPvEKgcEPwfvRHb81UBUla+4HPhpe5Q9og8Rue88ALsw
EvLYZ8mKt6erdsu+dzF+v3rLemn2QIt0yLgX3qRx61QYjex6mQYcvoWBK6KIDg+G
vHqrPzNUgaddJMOtXL2fkYbToqj9PR1dB4Dukz79UElJ+H4LVirXSnOZhfdlTRDF
j5SAksx6QrL2CaMGSOQZWp9+eK9wHZ8R0IGcUaYuNVXSbWEaLwY66OBjuYI3WkvM
9eY2lsFdu6Mq+2gl3R+VQVHVD5N7C472oYmemnGyf0mDaGrLpWIfwBXJmRt52GAO
h/ZVgZsHJgeCOBHL0hKO4wm41Z3WB7+nP3PrM86KDy2DMuGclvL6b3wyIh9gGo+E
sip0PQJqLsyR3VhPeOOmz93cC9PYspOgPnAg0F5ZAyg6Oey1/+EnfZHJooVXrPsC
g6A0F6J69khRxRHYG5vi5vlPzVTHr9+HX7khfoZDRktBui3YGeNBgFzGBMdlF+ry
aD0thRlyl3rvyCTyHJdsF2S06BtLnhvopZEf93e4wPCgyLa42Djtmurf/HI7Tybe
Y6/5/PG7NGnfroxK4qzl5muvdp544wqGssYU2lUD8m8xO4q1PKFluQmSfkiCzZAN
PYuNdGfO07TXzMFfdmaRgacCUx2Nh1Mhy8cimXDAZ5UHOhZbt7CifBm8wdc0meZv
bFP3mNaxyhZW4kCmE0Q1BJ7b9qa+MigW30vgixrJYHkNPkoPcHgMjmi7DAo3tfl6
jswA67YJpQEPsRiHb3BxPKp1g2e94tmps0wD6BU1y8L8CO79/9eRh1MB05KT64Tw
uiLg6KjWZwJF/L6ln7QjF0l4N/2GngV67aXg5taMDOcLYqlrTqOwDRE3Qyv55PDv
L3zHo3MrFvdvY2iwFysicpd4q7qhPlvKISJyNszcuhjmv0iTwDHvzQ/JVUHW68P0
0kVzGAfsUKgeYNF0f/REOfaUSQMeAOQEJIylbdWZmHjvgF8+6dzPrEcdgIaVVGFX
Kt8CO1IKVzbuX8ejiBLKQFCsPK1oYeaEBnw5Vw6+2YZBx1OlF6nSKjqeZ9jY92gD
4e2aElka50B73P11WbvM0vQDr3bT+mezIf+eIZoa6uUWG9oy2YWo/N1dHigeXSxF
cj3NfaDU1hDzq7DMj09IR1Alf1iYl0fxYrZsY7eXA+GBxcEnre1EsdI8GpvyzeNV
DshiYfCc1Exy8bb5+XmeQ/Kdj/+nvT7PPtVrLu5lE2sdS/4RFpZW239EIuo7LKjz
kA9GBp4GqHZXRhZ8stc2A6Fdu5tkYWvcrmsj5pgwEwBgyozpLjyamXznif9/LM4u
eZX8Hx2rgKGHM+l35jYDLrMOsiunXgNOv1CnJXOVYf9qDc6s6AYDwxTHOgNNlFJv
h57XLqT40LIyIBzUmPnSuoB1If4bkl4wtKu2mIDqLN7zfw6heY7uqedcRrZPdgtS
NW++37chU1TDlMKAZY/6obMfNA7Dv7YlvYnGJ+bCE2mC2o+67M2AVRf5PqKDJgti
RlYhv5G/EgpOBV6iO56CefbIEUsH28X9kwl8TLYOraSfPVwOgUQsywpsbsM2yZZX
nXIYmFZW+K/Yg1BCngyaXE2Z4KboTAZXbB7Z5OLUrR0Dhi3KI9H3TrCCNrQgalFM
UZUHcE7W/3pRKMM2IWvpNpVdZGXWUZ5pq8u/ZExX6H/l09TSXBt0sM69bpkosCe2
HrhwDQlq1/efeNhpbhiCGQJldAl/PDCAKhwgmwOYYRzLompAnHqgOP+In4no7Cb0
OvTfO66tKIjgqXj43ZjSVlEX5n97RY3wbBLXFIibHcoGVUfoW+5XqKhEgm+jWXUx
fcHQ0HdU3UvINuJJxIcwhzgnzoHwmJOVq2i1yoKbdPLxfTBOtrHCrTiUjcgF3r8h
Xo7TogDdJ1gqXWzlvkYrSsY11vLAtbatfxUF57CwETlNEYpWTO3ai0Nhxzh/Z2mA
NHXdlspHfFxg1p/etk5aO9S3CYXCdu3WsxiVJFvja1MOcoXVYzQq3VSX/DzfwTKI
pZFtyH+v/2021Md0rC5D52nRVRWBxgS7suapeu8EErj9nsowT/gx3wrlkw0v3SRn
EZMFdcXWijFfppw3yfPZ5y3i3nlv+hSvCUI9JqxH6MVUqziTGEdwjq0dGet/DhQb
quXxOJWCCojvAvbrsVwocRC4RVmNX1tFtaGlj14SnhkgjJ8HyD3OVmLVcYVAAnMT
mGIc7TX6YjY4l1Xjc0eqKNhixQiUS1QyN2rmIT5KWooxcFFaIOsK+I6GwZ2yVPbO
TuQKGdHf+eh/4gvPDqWwS4+GeLJyOJWbwHk4icaSDRl1y6wcHjojREOqwip6nlE8
xEsKoJMc3ac8/Z31zsjrKh7gAd2p0mnPBYHj5po1qnJrbcqf6aTFqQ7Srdb/+hBG
YabcPiRmx1h1PU9MoQz8iHtp8UTvluK7eQ1OTZHjYyznF2x36oPvclZXzVYxaKpE
TO9SJ2GtMfGlX4JvcRYq+5Cq2wJoQaBG5lq4AsXkiXLwwiwuIc6zOElb7esZ2aWC
ft3+AMCCbmsyEKQwdVXF+rOPTtP+/IdzxXF8lLXchsjQkD6knTYJastLLMjqfWFi
6NsrakcXgw1zGIDSti8U39UNzdLLe6rlzchpixDxjwhRnjFGpHGJYsEj6VzXdmsf
CbNj9zPTbXCJMAcl/Y8Ao0W/uJNhVhTtPn6oDWxuajHAf05ZAcmsTQqiQVDucv95
13sAeoSkwsIy/uAjhL1nJIYNMjAJl8bXl0tN5NWkDdurQbqu+sqzLKdU4SWbV4qf
ZiVyGSwf1uAzgdf6NQUJN62d0S1m9XM0JJ6oRWzDLkWgS/a5bKI+VRYNXGCsCOO2
eT+iUp/5AOjXXs8g66M4Xa3cEkiqkU0ohs/E3gdIm8Znnc3Iv1vZI1aOD34qZTDx
TzpFe42+SJlETOOq5UQ7JXgVoxDnQ8MroXFONxR2HuC+Hh5XxhurPBpUfoCsw0eF
YQgMtbHEfWoyn12qzPxa4GFpncgtcpieUWYV6N3gsGBvkS+QOUy7bBUio50JW9uW
cICkXii92ZCiMQNW3auBXBt8N8m5s1ciZcsFq9K0xtjsT68PYM3iHX1YgyQhopN4
ehcjhauLckVc1ImS+7VUq//9rHCh39JGHQaSyozoFyCIZ6dH1pvDoSggY8FxFim2
kxMXtdfwvhCqkCE2MqWxCY4rvAx8mYHAoeYpOTf3WeFsqE8y+oBWm/O/4Zwjnj9m
zbkw/Ah3H/ma4tiCNanqGGByNE4MxZOTLyX9qcpG0RsD9dvV5XW8iCsTTUYH/kpR
17/5VAl0I8tSx9cvn/DREPeCDw47FomMv5pSj72jEjzg6gj/5Pwq3iuJKD2LxhBV
8VbF4LKg+4D+1dYsEgbpYIEqz0dSO4bvN7cWO2uYt7FYMLBp5HK7u3YWEGpfFWIH
qr42xk/2yU2hVhtnIb/6i9JP7ZqZPPqiDbVsD2lH9cd0oxz4PRXZRIReVrVZ8Evq
LBH0lugehAJPRMvbq20Fq+2RJtARMqa8uexqKFax8anfk84FGrzpabX7XgEWzPlF
Z8X+7sXkSEZZ0eJnugsRmH0fPtXqCntH0nOQxVjiNMBFtXNuQ5AFpRMmNvOeXInV
lyf4Wf9mrP1ljlgy+SYP7ymdnMZ0SbP59nF0uT4kIJvC9D1HtemGDrn4b5DpjP6I
GHAeNW/oT1wnTmNXwcysYxTKF/VoyqUtWKXbpQz4nbXF2+WLV7DbUWXO79LAtMol
UdB6CBuy51tiIM/N5JZsfG5wIrZlAK4plTfmJFH+bF7vBDAQf2Xhevc25cGq+axV
rFNlN0hUm60H56bz8euO4kve7CRaxqXcGbzb/ssRenGdgzy5d52TlOpOw6Am5AmQ
EQobS96DYhC8HS6hpsoXo867jPlBbwxnRFNGOEDS/yNW3hZfuv+6Cv+zhbTOSMIq
w/4uaDeoz015RQcjTeZH5VRZEATs2DlcmUDmHKfeh2l0wgtB02e04lgn9K3iv5mA
w7tyhZnzL2wiQxhmqYqUo2632W/MYvaqCeEpghcwz7cCTsRovjIhtgeW1yRdIjrn
vIVwQcXHQcqx5bZykt0LmajtwFGUCbf8oMNAidfBOItB9wl3ZY8Gte0MVMh6Dnq/
89ixMEWInXQlnhY4/jMbfFouHuCzxBSxAmEl21y2kMSUd503YQOJ1ILImXYUQH0p
kMNh3PsZhn4UxXDEOR6ofIs5uo07wFnSARjhAnJC//ELLertwACmLwuY0NmDQgac
Lvohdh2TllwQNosLD4G3hfxpikPG4iPUCTUwPk+wu9fxiZW3YJI8QHOJtMNWwlcw
r5PfMKdI1NsGNSH19qlPgkYmikW+S1ZVWhkS7PeageT66hwsD9IjFzkqlmUSZCBf
FMtuau/zfdJsJVkSXGfgyYf7mclFVLA39zg6jkH1uA6ZEl4HioZi/+d+PAXaT30e
de0xzm1wFooCxZmW+vLJ9ub6si7VFLPoia3m0SPJcq5XdtB/u4nv23ijngbnpVAJ
cwzBqnqyPxD82asqFWUbQjzQ/JdAeZQf9qcFT9MAIhPy6rWWw1Drl/LheSXYmnMd
F8fx5odOh6K6g+9wIxN1WW57U5y/NCMNoY37SJES6YrF2ucmejKhIlZ3PuCe8F7s
IbJS8Nfo/dKxhehV7omlLaippGzBR6UFwLJinCLyKZF4PVMGd7bUWLC+S2VI76WS
wsQnWP+iaWbDUlrqdTJ4i3AmSi6E8UwMsHtfGgdjLGmF+haBkW8xs6iE4HOz1szr
NRjmzlIneR/Ao8HalNnTU5eGF18kGD/6gd6/8i5qlG6LB60TcqkSnYGbBQ482GXF
8LgWH2Tr2VbbctHda9kbnEm3XI2P581CD1Gvt7wi7dcGtnHO7XYGYvZmrwtXnGLA
RWoa3S+F6p83vD67EXD+N3TRjWzXTBzD+XVr4YVG69slyirA3Sl65ykpFz6x2mKU
2kSlVZdJGTsAfmuZA8RkN+ehiijq8f2xuWn5IMt+jdCo2ECctv3tZVSgHAX6AvM9
td1umI/94yIxkPCsQBqY/DWZaVeI7GtW3uTwfJ7si/DnSiKSbVeKCDGn9sYbJA3U
f93qaUrFrdUvy/V+MXJIxhzMutIbXBGDO4PKDbiIK4190GiP6yqyG45ExkBvusUO
4iQisaGS2pEw/wcNc9PYnImybfQWNlCqln9Ru+kY+HgM4xpSUD51uXlkGrXux0yv
r+fGLbaB08ZwFJe80RFhHSjjqTKBvtNFxG5+0lcZvnF1vr3MBgv3mh4bWJx07gKD
kpktFawPm4fQyMHn8ruF52SxUjniHMv+V30Kq6VOMDsd0peeAUmQV1ZXMRcqtcBO
px9BIoofMQzNVIEltXnjQMgSgJfU68MIxxwq2HqGAhlFPd2KbdxeTUiekozK+ON+
0VteHEM7a/FHlaSoFk46RFDQP+LSxK+jviTp+2niz2ip7LgZMUt/CLU6n0mScqsn
izae/UePN7bf8da5pvo04XZSHRbjn4llv84hR/gB5MVk3rGXfXr974AsegJoCjXj
/Evxuwdz2Pqf+n+uRNLWy2lFnVrcGcUNTaCLVCbvXuCe1lLTLnFD5fV19eJocRdk
Bdw/B09Z7V8u+OI+M24EB28Vfps5/x//fkWzU6GDvDqCj22te4LQEdoPv9Fpc5L3
cZC/hgj7Nba6/iIqWUbETEeib/5NNsqW5V3m6iWUBp4WWK8YntXTsFWdJmwlsxGR
QPZIiU+3VMmZw4Q7Yjl0xUn1DfKpqyVEbNfWCy2KmNPQ6ouLG5/8Mze+5cz7uhVe
qW+9x1rPQOAcwSH3a21CgWveRJHo76Sj1TkRTQVCaYRCv2xwa9jZSmb2+XILp3iL
TIimvPcy2DkCmoQliBtEda8qp6EmklnVmTBVbxZjInM5a7e/XSXZK9A8xu+PXbFK
0JqnL+HVTvVqVgkR46WDtLYFEOPGVEOeYa0eG/elRqg365lXEQ1oY6icP9U+ZHU2
IpIX8qoaJJDmFAyth889K0VAUaWl8Y8SZ+Zf6dxlemto1ry8RGpGnPPc3Rd3u5o6
zUdM+D8fCydAzz4SaR0xX83gUhO1QQTmCkL3EUFqvgM23maSrnmPt1igHmmv6jCU
W7usk9FxoDkpqo0cSP09XUlVzeW9tHibQk8xRSe+xuEUrFXRSaxV8lzDWdQumD0t
7CJNxouKlN+mGBxW4YDb9ttxhaaYVs+FQxtWLEdXJHB48QJFKbJ7fZKj9sqXWKNI
HZMDlj0m5pBhn6AcBRLW3ECPf7RbRuRUkEqHWjB1Wj7zu90Viqp2sh7WxaSN4302
jeUluTlOOE6xm5H97sQoq+Lo+J2eRjDlp16Prn8qBzY7a43sDn5htKX0BlmThf+v
dyWrGcrvZ9UKjADN36IyJUDc43pHnnNBWuHKTn655iGkhFtccPdeblUuQgkd+7se
aO3UeXJe5YwUi5C0t/7rkuFrE/UjGyCJ1vMJ4ZQRF7ysQc5e4mkJFuUKbcBFMSDW
XnHd9xKnblSWnxJ6X7S51n9CPyPuqJI/qbo93Z292gVpHdqld4L3FzAJpcNfDwWv
XCxnmdp7aHtkIIxk6LRycEfmlg1POTtOn12T//wJ/TCubVIa21fb1wM49i3eEutT
LagKJMgDeRtGb6H7iNBUVeBAA2dWausG64usHbKh/HaB10Lv4H5zFXC1U4tRuhn/
5XTNV1MQLzUqZtC7TwYXU42G39tLeH0z6NSzc6bAGz/8zXG21kEb51rhNZkyUeM0
QTRiyGzDPqeAh0AePSdtg3d9nUq6yUySqT6OkZyljBg3BB3SdLkOuMkjwV7XY2IZ
rYDcxO8kyRHHho4YNlgeDkkKufgV2ZxyQfZVV2ZbZi5Dsd+OU9ZooKFpI6zj0CFv
Y06Z8f6HerDljcdtnNKhAoSFcJhVuBtW0z/xXUgMlXoEWRRSwo0E4lFwRspxgiT8
d3CPI8e+jx+p+QRF33httxqDNGKA8WE6w10IrPDA6CU0ZZt1+4iMDsOSKJUIbp9N
95bJ540dJKYaRpkxBsYv408PXBi1MyHMKBsuWz5kL6+zxhfHcTKJLH5UK4IYweH+
7pWX1wx0La52f8Hbo86A4leHJgJIdKGLodBZHnoOMisn3MyF3qQVpYYToesEwoOX
nO6fboI6BZJVMstl8fRSnK5rn42kyOqP6QVz/oDZDMX428Qb3KoSaOIU4v7/5S/y
ZjNXE01mjBtltuRfkeVcLzz+J+XSthOwEMoRUvq/KoWZZLLSW2ukKUPU1TgN0+de
FW/BTXZC4ZlEtV7qYF155FleRrUhtO0O3akj604uQGVGnmruwp2y837ZrOlSTqGt
reUnO5sp8pR89if6IRZAENtjZ1iH3pALHAPBxY6EHaPWmnwPvbjWSKq4NtkzO801
XDR+UcVHm/I8eTt9f7bwm0ilYDN7IbhWAGlPo4EMnSQuFwQJl3XxNcoSaa2dmkzF
7m4T+QUCSTDsvYnOZUg5twpCPRwoZ6R3vTpwWOJWwFs3w/4Oq+x9m4WyQunjXNSs
7/ozCDYIhGE5dX9CFtO6BvDa4o05a2v1He5U8a4KT+ypebA3Fru07VWIpraiNrme
zO4P6EgsKEE7Gt7y5/NfAKJyyjPDAPltLrvhAk9+NeWhx8y5tXmAkvyztEQaAdPi
U68Q2j0arRhQPXG0AYk+r8qZy4EXsJfxJNIxw8P5X1So6w6Sx5qXrmZsTY1N4dNM
iOICV/qVOORxpKThgGGXufOJO6+da9gnjJlMBomGzpohsOAWGe8XL2g5D/lGXtoo
ME5fVpGdgqbS7SK6sRbN4/Efg3vLiHcEU3YxHU21BrRUWOOwCwKc1kZCulybn0/6
zPWzJI+qN5FB9VhnAZZfpStyBAwjF82sLA7ChCPuPesGcsJkIl+g5B3rjj/fqY6C
xhgirjHcIlH31pr9ukse97wbdVP8o7HYRHQxJO3cjdq0KRlyr1FJhX/K4sAGQ+IU
qFLcLUzl/uH94mdZnzVFpdAA3sBD10rKoTpsAcgSoFT/glC2EIXTOum7rc9NB2sE
L45MWtXwV7xYacq99VRSheg5qtnruwE8WwelJlubxRTiXEmkNBBDO2/zo8Diy9zR
pe79JTxJXp1N+01HATqCFDwglzwda6XzQqZIb0JNWSMfQDHvGn3nHvIxjkY0pYOF
eDCLXCxQlWwyfaqsrFBb4E464eRmoWPCeijdlsHwS17XDnwxDcoZWDKPonqwdfCj
77flUu52eltchh787Z5XI0r7nKrHJGx2e4LojF8dFu03pcuBf0/MNZXmg/gOLBq4
3nHlp9TMryReAtm1s6FwZDRO09NVEjQfjOAzPULjUnj3BHyO2qxItzY6y7QP9ego
Oxz6w/kG5D252MUmffu/uJPpa7fhalDqBKn1WX0CaUFyp659WVgDxfibABkFMhK+
fi53fAuyjzFK9bXNi+PbTj6HlP6u+vJSVM3s/xAZFU2pXsXAM84DQXzRcuHBL5WD
iRywpjMqdP6Re8YvpUl45unGVYMZx/bpPOybPncvKSCo60mZb+sGRzI9drn2dyjl
zhjLti45jhnYNrGJdwvHzjtodLq/m0nmsmJvdp7b5HUuTqCEWBH3+wgODSJ6Ezdv
oD4m1l9iQMqYHVmmiaQjTuWjCeo/QYqevj84934mo1yWrbHliHMp+VFi9nU7R1Fd
37IzhwM+/4NgimaJFpDkXvCKTIqjTuOi39CUwQMMekwFoeph26oaZH3LBpva/wiO
TCdxSjwj2R3aQDMYKh7mq4XvZZ2tQ7/yTU/MD+1qRZF+06MBvXLdOOLDk2bN1p6b
0Bzg2jQ20069eEyGcUBzhqGZQd6Ip84M4/w/VJJ+9dnQQZAKNOSk4euOckF8l5dn
2I59xc9mYxzcHhfpMd72IHxMfaMeiJVdf4VuQeBuIUt1Pz6s2z3v/K9R1AvrY8GV
DY3/0JNHD73xWhKJ9Pku7divfLMBY0wlqCxMLoCDut9AXarKlQfZtANtUC80L06T
PpqEWehklhpYS4tN//Vqi2SnT83VPJDHToWEqIhII36+acNRfm3hQDXHq6dMvyIV
ijhcno7h3JLs41TA3XokUO3LXKNesYYUQcjFkEqpfHlf1+6d1Uq32RoLVr4DiYRL
7wB0JINUr2EDL8oxY585l13T1etiO/sfK/OzSY6O5P9DFtuDTtD2Tu7mFI6vlKtw
dgcujfZv6FGzt/uDvL8Kso5yG4wTpCum4h+DHIrp1enSTGjcnSDbs0j3debuuodX
UrImLMyKW1NsV3Zvg6FXHycwC1/xHBllZwC4UzLC/8BpeIDCl5+w9LNU6AsIJd4q
7oHemA8M7A2G8dTrTNYK8JCF8lu+AYlA9lhahF5EzInayDq8+o3phh8pICMlhZWm
0eRhn4+hJp+ImVF9j+Ng79KlP1EBl8o0FIMkm0ugfEfB9vQ0QdZZneaFsgTpSVUz
5xfpllICUZ+PzlppfjsrC7bqhHvqAN7WGBSMp4+KfZjtwzqspVuP/1m0ba2Hg1ui
N6CAqj/+BqczWO7qG48xURJSX+rQk3kHHQ2cdt5yu9FnTV5UakwvLllwUpFZYS+Y
Imw6qv7YuEY1pVyNWr7GHhU8/yDZWK9MlsMlrOQTXuixbQhiMgOgpy+kYza3dqhq
HMuI/C+o2R5Am2gfyyABjt1ew07nezJQ7jovMIugbRib7jjfE7sR8O60myW6/oEP
zgdHFoGR9VUcnmafQAlLCP5/Qbz29hlLSAo3Yf5+p+ihE79CxgFuwjF997j8Rrtv
Ca5rT5qswc19pvxwiSAIRhGAmtvr3PFnYvECMljPLNEvkfLuqOQKsZnkXt6F3ezS
GJX5yO9Koy+IkfoAfr1Q55autzpcNdo6BKIBcUo5gfRx1P9qv8E6+hW8H4kcDBLu
OVax1nfGbofzSo7QLQhs52sXGACzsk+jobqzzKLntHf6fxt9GJClgaBWxXEdzAfX
+9zqeYVFdPR/r/nm7ZGWVDDXPddWtS6uWANdBB3TAYl63XYYu04MPNA5VjC/RwdG
lGxkSUQ/e4nqBZNvK9QZb6YncidBOuYYxGM5SnbdlDB6aJYmqpMzd6tkFzkUvN8h
l0GX0kR9MeOWdz4xg1jzeE9BPgGAeUMT+zldzMBE1mw9nq6gDf5n/+wOT8B8NVan
PysX6159M3vkFsKOiqq71mNq2mmx/+mDXNjDTXBJ0zAtB+CATsOuyTRzQHJsSlfF
VGdPka3sgKzaOqg/UgU7Awdxu6VOkltJ+RxTIN2C/tiwSIJ7KKU5YAMOuEKNQePP
5pHJa/pmvOlTnp/tSD1FmwepiowJfejcEKhPcSxo7EEp/FUZa5YPInm2Yqd+uLuZ
nFQnS1Xmg/fAeeDku+BYigfJOB26AZ7jOBZDHHYuddg33buB0VI6MOA6C6xcxGMJ
AvMCfCgDq946cBaupwzjwVjQKcI1hVzisgnlu1rBL3utww2cczNEzRCilfg9AnCh
+67RhuHJretwyCTTmsm5ktDWJvBxgbECrPFZzEHkORhPF4RdZHe91LPbG4J3Vlzt
U2cVdgCMvk11Mbcd1raeWv7Hs9i0gn4cuH2v6zFXFMn5BkmRHfRJz2CWx4y2JCvf
KFZx0qvEJas6fPT8Tp91ey9aeBerdibBRV4IjZUVNoDcpnCbVqL//CJKHqCP9mL5
nYoy56g92yun5hhr3j1YVsRFhLg3s2aP7C3+j8h0y+lMuZdELzgyjtyILBEnh9XS
OmoHiOVtOeHeaBkAIvGDUHRPClEhTF0KBKjjrZR+wAl30aWE1PWgYjIgqNFoZt3T
HofILiFwAbUhZChVBx0nNTQCCHC00WKEwbbzxoM1Odw+RCI9zVIE/fUeghGxcLCt
sFJzARzruMQEl4Lk6M7tuFfbUL3jWSAKE/JvBrbmDv/A6MVYYp2xlQABisO1M4xw
Pv5QM/1YF6At4hunQ+YbujD2d8uvrVU7Kgcw27pQVgm6tlwscL2pO5kmKUdOBG3e
F9PkodXPcdW1hzYD7Fr9Hf2cDmbBiJNTgBKWfWOLtOc7adJM+VfUzfiAezj6JVdE
DfSQP12hNoMa3psusmdUNANoQzjBQaYnCQWcYatGoN8gKSbxgl5HNoHcBDKBYgdJ
xzfTzcK/a9fQBkgYzc2ba9OI4/cwx0K+AIwWejZNku5DLXUXZ6C9f1N4ClhndH9C
f4KRCt/uVwEz5Whhx3EjZ0N0SSM08jmW8LEERDrNaT+sUXL9LvsU+gmItTo9+3Nz
wvT91bTBA3rMDEH777YZUkgGc+fvpxxKp3G06brSs3YP2ILuSaZpqICkraw+3KIJ
JkQtQD8TsGqRX3HJO6uGsTw9KI6nA2d8YrJI7T9JOx6T2J0H7GcomZw/napIEqAj
rWe894XGT8GpfBDeumy93TN1gLsQzVs9h/PwFxpeRBuAtfxCrQnKnyCmLdcM7zhB
sBwH/OrgHls6C+W+RA0pTrDqjiO+YPDrxqJKU5JBaHUzRdNYA8Ts6vgYVqEUwUPL
1nMUv0Hh3cg7eNREl+sQ7ZN0fFDdQOgy2gyueGycQ1AdxS7rk4lPS50a+55+FczG
Oe0OU+lQaojSDdpDDvX6et0NETi+bt6vl6dnyyv/j6MDqwWgJvrk9fCKeZmAegBh
/o4tCZccddU9yiEdVyeAS3mtCaSIdqiQM3Hs4Bz6kTvNqRCK1hFaOq+qpV8xkkBB
mSwHN6zsEYYAw50btjaNxo2lGIAoU0Qs3JC1bwfLWvH5jO6IpPw4LxuuV36p3OOB
6c/wzFuAUXofid0TwCFOPC5+d0KtKtDnnq74A7Cm6tIK+ICH27qzfwDEsQGMoyuo
qmyBOydMST0E/8PYVCl9N+8h1bnhN8lVGNTxUglbseK510ACDDHquuln4QwFA7KY
qOUp5jWwmM5ItbNaR6kN/BbC3sGTpcJQEbLlmP1JXpK+WcmK+CigCc8Zk7IFlqHO
TyoS/y79thFaE9Q/U42roJOvW7XIHoNSJqY56qbMHS1Q0mv97HKNeOoSbwgxNzz3
zsJJv4nvuOSSLP2ioJkTxuYmT1my3jGN35fUtjP8KK+hdvwmdNqliA4CEOAqh1Yc
/FBrlzWXvXTlfnmYb5BdAheFnfV6jBLmTNLXkXuA2JjKhyGBGpPWWyMLFJMJMH0u
FKaDb7lSs74xoiJI0CWWB0YzmfkvJIVarVpPb9Hb/aFnlgcQ0cSlx/SM51oC3k9a
JUv95HQ6OM3B4r7Sj/2ElpV2n7oJtfNlY5SltwCvUd1sDuEBN9D7wIAZ038ikWaK
kPtSi9mPMYRlouClZD54YeeiD8xm7JFX6IKB7ymuErKtOJJBF7oH/fPU35sRucnS
ZXBBxCIbR2TdzqhiBE63YrItxEsgaDxPqUBHG9wgJBUGydWQ1hKSM/1UJtR14H9J
Ox/az++tu7xbYug1UE4Ln38txO+sHvipj9IRutSKORzYo08Vzd6WArQScqRlRywO
8sLm1nzxZm7xkQoh0Tx46+4AAnv2a8EhCQ6potLvTfgysxr/lVuVu49zirwzzvkz
5wbug+LzyWVRyd9an7dClPHIKOevYNzYbCEEcgZxmZd8qpfCbMi7r7L2+zT1CasJ
xXzvQeLIn7/7UeFyGEy+2Er1HVP1gf7GfvWF8FRHyqfQznJf6Pyo+fPpuObA0qqy
E/acHnwB8uEzkmpvCdJWJmKrbCcauS+vc64KHZmQsBaZU5pre88dydo3H08WzKRW
XzCI9wdJe5CfTen6H53FbBjrQuP9vszn5c+DPOBRvpBZgeuapTmjeziCudoS91wh
desExCPLkCXUGWd+/Ngfw4+lXeXTOLI3WivVrl+YfJo0Ozf9G/Y5Q5rYU6vN9QKA
Ei9dhsdaFPAn0mq4s6HPM6CXDE8qftnFHk6GTT6laSjzdne4k7/hrSqMH9WUUQoU
o68sW5p/3bt7Fib2GP7uTpz407OeAXjl0ct84oRSmnu6dsqXNCWYKk0bMIBkEkfa
UIvMeInkrAPo2YGbuD/UyIQjtOibhw7erYKc2pa6uKyKnpucxlZhYd1kmFXVUaV6
QU/3KTPRN4lJQyccHoXJ9Go3D1kKkzUG2TS2vADJE0C0DpGeBPuxrIpX+sTNq7Op
LL1eexTAEwRdLMYMHF/LlYC5nJrsv3GPVhUcCiPi2pcFr0FlJ1BgYc8fnvjloks+
HZ3JRrq8+MYs0zQFDH4rkcE5/B+EoNiwNZDGSH9ucMYfRToPL2I/xgTdpjTwRIU2
FM3w2OpvLc/S2vB2OyMKsCG3j1jK9H4EYJh/WRZS+iJWU1tXX6jHpNJsFsHdrFYH
iOyWLm+stXh2aKOpWPdjB34kk3fevYRxtKse3nrOMJCO15ynPWAkHWo+tzP1mje0
7xpLog40JckxxJW6/aML1U8+c+phDY+r2/vPdUEa89X07TCXungQOIlQMypxRZXN
KR9uzaumCd9Jqf6/NkXAACWIfE+WzPpA4TOuyp917rzUVkLtBO3sN6T6oLS1t6vZ
6O5eHtm65OwxApUvJi8XBwxGU6O4t//3ZxA9K3sfDDUC6HT/4hqd3dcRzVAR9olH
a4SMLUj42A5tAva0vonAly1XpjDgvc4Zcd842mZF9e4v9VmAZcEPaKWARQB+STrK
cBtfof2Bz2arDEhTsmR/vLDdJKR6zsSyVEgzJA9Atwz2r7tk4vmnS1Yelem1uLoB
2hj1D79servTQeTtNSUtpllkFhN2YphCRkYekvqQLYGnczRPyYHcCm9tHGWg2eIl
8h+7mbpSsyWDX6t3SJec1Mf6zTfPKmmGsEbofEgpcTFX5xOpFIRqCRTzN/lxO2n7
uMhkSSUkJhpbprG6U+41VV/3OEgG1n6Yxn8OOObSu42G1jEvgy1wQEN0ak1sS17T
Hf9I0+Lh9H6dEBKMbsOXKZYO6WVbIxpbFXcoEEbF7cJxkQLICMM2KHd+YiILc/EQ
l3srW0MDlWyW7mq549DN1TMnPfkQBTyywPPZR7PG4V4GCd0nfk7wUsgdjLllyPsV
jVua0o6yzKko5NNkAoT/bUs2A4gRkmb+hSQIYtNT+tEzBpiyXCbcNc+FZcaS53GI
6aYFcwDDI3Oeo2lQbFWmDD6phNXOp8XpUWD7Xl79PA1YzfinXABCl00ZmT3DCuF6
jdCvPj61Ow90aQe8aX8J9JH2bAys3wu53N/ZSfCrU6boN0B6ZRbnO+nokbhE9Ba9
AiIgNEirwZjBp+reyYrGRmsiNSY1oJUyjeIYf3PnlfBGrTSjg/9Xf1biO1kQRSco
rd0AqM82tfuqFaYgGpphXMbfj6+T0zW8P6GC4VAw4YfVejpn0QgUiUCdrJUoSP98
VzS8YDPzYvgVN1oufnOp4hwLPxToct3L7GBbt3QYn6TJxQsrtQK7TatLRjBMgAV8
YBXrbSaF+sMgekZRYvtHBIBkyp5iysLz7P9O27xFaoLhpucHHNdTg0VD9s2A7pwL
eO9MTgMpA1KGi0pXTW1tWfJbjOlt3SE9LNy4T9c9VYGYkY8FXjUj7/Zk4CSD61hY
MANel9nGn8t0SPdWPv8GJd5VrdH0OOGx5oWw1gWAj+/uRVSysq/a2hmP1VLr61Vh
ydd1kj7UOFeDnexyrYN7EnkRLxJHTof81rKwxpwPe/qMtlsSYKiQKUwiG3cOf0G/
5qmf5c2ixm6Svr/Cc/h+J4RrVsDwJGUeCvEZQiE/0jLU6cQ1S8b3h42n6nlGsC6+
R7qatFKPaJKa34RiLi1fTzf5q2dLP0O9nOe8tv82+Q+DN13dlQBv13k2ofCXTkGQ
5fyFeJgtXrhV70oaw5Euznd0wD4E2A0b4lb/sXrkIvL03spsAR0UmKjybq0fPcys
gt5YB7yzChWSRx9IekHiFYgfEING2WAjAnilaXtSNZ0vM/mIAgrpGZ0Tw/SBPM3h
rbCiI8rPXmRenVE1LatTeEsp+uuBWbV7RHlsw9v7KsYbWFS2rHRI4QHvmsKGn17L
91QzywdZqIRTxZMnZRciyWrl3wJ0MdRn6Hz6JXp25j5PvZ/cpGr53nYwFS1cvjR0
IacNM/VG65lqeF78dl7UsO3PMbd5njc4+HU8fB7LWsUUMIfUNee80oRhHf9L/i0F
3IdrLNtWEqgtFq/rgaWtClhnKWhuYu5B0p9uQ2YIlPYXoLd2jVRQ8lszaWlyOwtO
k0bWBMx8KU/1vNXGqqc0H0Ysb6njgYMHNJP9vJZE1Ffvt4qbgmvTRM+7+6YTrvtX
fpD+2TJZGQVP41BaaHH6EgIE6ZtwpCnnjH7oIiXXdQ01Y52AEgyvGvw25bcwyUg2
n+a9IYfb3dCjZqbTIWVniuL9oFUclQq1G50yDi3VmjtM6Qmcr77ULbJdp28FI6Za
myLt7zEEnLws0uoISyIRr2sKVaA38V4j/s4VGIqP1wOp7FkUyOm75WOWU8XVLDzb
ppUkVGcz9dMQqYEWGoeEbYX5mk0D+haA1wBv1YWWCjuxG+jGdWCSylju6eQSJz+R
pGFyNK+cbRIxWOe3FoWNuyzYrSemBHdQuQSQLJ8p6gph4OfS2WXzmeCZ0WZCMNcB
PWx/O/2313LhdGX9d8H/PtSete/lItI92ExZnA4KulxMicsb4K5NslHQysGcDSLX
Jz5p5oSRv9qF9IN4I6ogGyC+z3ul/Soot4ZEdjmbp4+khfA1ms8I2nymXGqrdQKa
NE1pQjwyqcjyBifxHYAkstqf4qAnq8gKv18/4lg9cJNpTmEYJ6m+UOAzsL1pnB5O
yQhoyGsY47+dGq+2q9Nt8aKxClJfDDONsBQLn82xfNY2TwugVviCijep7r8BhLN5
ZWFx6uKiG/CX9t3Bq3j8bh50SYnughoA09dUmj7iPHg4D8J75DagrWQFKamTATca
0EcPjZejrBlktG2+WM1gUrCzTdwhhP8zsa2JVZ9zXpsIPvEbl1ic993iS2nAI95W
6d92N+ZmYXIcz66DyzYPPhmkbsKSCSP9T0Gikq4n38Djk/AVsqC3dnDT8mw28MMj
2KzNLqLeAxF7Mr9DH+QY2Ww1jyC24fvT7CmwR0+Q4j6CisuOj757tlFKB2JiTOZs
jxwMt6tyzoPWKWpTHnGwhxHcCZ6aO5B2bOxERl0camn+cZidcQ0TmzBuqaTq6plr
LAsugr5b1f0xJdPqGgaKRLWJj0yBN+DqjnggGJ6rpilrbCxlXuO2FuVqBBJurowG
7k0cU8Z9uoqAaPydPBavt7P2QqqPgtC8Wuoy1L5SwNPPWbGifFolNE4wUM3Fyg5W
UBep6R5SwJ0jm2UnGg2PjVsVtVkcJT3ykU6cr/4YY+dCzwPCWEQWekg5qVlwadlE
vOveIqlfFu/dPiNMaA25HXVwyMezhOYUue2LuvNiIKlKVjc4BsznyyPRfQPE8TU8
G6vZrWJjkXkW7cPdvbzmlGRqiESJbnF6d3gSrwMRyLKxQi50j/8HvkJ8ImDi3qQp
f/CzzM/CsVZPUAsyjep4St6Y7u6xauz8jMQSQlVCyLak4vZFaUCzmiVT4cZGGFQ0
VWsMiHM8Vg12iQoVQlvqG1r7fZeIjJFAhlevV3OuFZ+44RMGtO8L34yFBbB38ioB
mh5HNJrXXOGhZKRyYW6AEXcFehwu0V4Uuda5Tg3ewiKWCrXn1ihcZSYihula+kbH
BN0oJrwtKX5VecXSca+ZX+x+kFjaxysMl3enf1jKU+x4B6QgCZZ4NPMPLLRhjWgb
8lpBSF65skRxtpsvgTIqy6o6YEKaZCyMa+XSCqL/ZZy2SOc8/Ky9V2itwsNKl9kW
34GArcQ+x1E8AX+7aQON5xe4+dqMZL4ybdr1YEFu1fVCZJ07uGU6rbUXkaJSnRj6
Mr+fjZLj7ulDEnYtNUwfXKzVYLWaxAP5BGvGYK2cqh2N+ocfEuaPQR+tP+khxMEj
aK0osph66nbCueQW1BL6+IFEoSLxkDoUSGfjmpfWVMl5Nr6RQkpuHTcv0G1M2F9r
3i7br4r6+KQtfx7l4HUTn4SEEJ3HWYXc82jjnNnamgqk/VAQipITrv2X91S15l/M
dvyeIgzQu7vxuGFOG8IvmiAMfirx65J+CIE4UgCE+bEnncimvxtabbj98mZPdgm0
3LaZiPsI5ocCNLLPIG9Qq3xeVDTJB/8Xf78GhlAVSsZwqk/Ap9cBnSwAX9DvakVa
S32+PZWfflFgTbpMSN+BXqbwBxI2Sau4HqyU3elQC53K3hu/KZCt+zKORKl79xKl
eE/PTwDN4BcySFihPoGEr9XCUYRjJuhHkjQp63cKkvbuay10nRkMta2GOLEwO7J2
FjekSW//uZTdCACrr1GMnPt9pASGmQxkHjf/4ANlrmZU5CN7RO1FxVhMB2Be8yAV
h57ZQQrFPo6vlwz2y9xD+O6fe490RIvQAyoANHHkGczAaPecH9lkqkx7IquFqpmI
s2I92J3wC9nbS5WR5ycTzvRPPQFEr5j+LplHSKz7K1NaPiH6HNJz12QYr9BmCr1E
XMSKWC3Zgjw3r0RYHE65CmNYratsealcXCKNvl+hMZbw0NnekhAq2T5xoACAmPld
UTzE7/W+SdpiSIXvvH0seuf4bAzBtu89eG+ocjHOAH4p5pXXfCTuvdqlvJjgJK1C
b6djZ57wV8SI40Q5H0fnqmyWFv4aWS35qK9jj89veUyMid12g2VtTh4sliTBX2Jh
LP13nc1TQh5adc/GpAtCsCtC4lAiIgHxK7casDz/kmutV85GlqDw7C5uNCDTFLcy
DdlGUsvwcQ1Ne35y1rpCZ4zlx6vAM0Il+njNoax72rsWUgofye2nd/H7kUI+Y4VW
99Ik118zgwfCHO6gSlZmhv3etq3qHnXlT+X7Jo5Ns1FRm0hVjGoDhy05EhJZ5Cga
12lp+Xgt9P7V2BvcNOIzzZKxeC4TpWe+nANerwOX7kmVUqW8i/j3XScu6av3Y0l1
a7sVCgg3KpWUSJlvCFdFJ7RX4fYl7CTXKWqE3SyRSbHuEJUAF0VumSvXqAXxhs6T
tmXW1yfHyE6vgs6jTm4hYCZEVoU3rUgJRkjFRcdHYd/37AGrozr4zbbItExp2fNN
g4oPu57bbHiW5r50lRcicAIrJ0KIT35ESUavTr/YA3jvN6sYUIoQ2nJmHNKRylsD
+3ZUvUWRGDiYVTNRY0IFYsScBqjnygKNddYtK3rtwc9v7XuPa1Xykf1bvth0oJ+E
LLCBfjuEcGoohGr+EpurLSbC751CZ5fDPTl0rDDsz9bdRCNZuH1k2gAyP7+VOVqZ
4kgCRgM/5CwUMLyI5vRh8hx46Qz0csXPQiBBjSsIlNhLAeWyj1E3ofyeFmde37Gt
TYDmnOk563yhNRpt2V9hTrPx0OMardDBRx3+yIew+4mziZ8GeYIT51PhQtI434xR
GNgQupr6vAQspQIYEB9VHCwVOIPf8PvJK+/1iB+pirtU1MolMF+mg3nyiLAzvk42
Ep5mws6mClqVy3h3IAoORFI4R6qfZ0n3lmgBqDtyQeSMT7gLWpgSgZGCgG99KkG8
bE3ytNxH1pUoCHqJq+ouO5SdVVEDM8xu3Oy/0VvE9SPnJUg79e5Z7QIDeUQQDkCd
FymajMrQU1xrvfhjkImSKQHotKbFpZSrUQohIuqUlwPALtvj7QOL2iD2eKZ3ASCt
sPLSW9qHP6ZSAnfVaRm5J35oRrBwEQkKL56VbDCFAc6Ty2To9x7NNeqNEeWfXR59
leFksbu7dJkKDzubPh/ZZtiRwXAL6RnxLJmLsB5XAFVH3C/yuvOdq0rwQDdywF7v
gvVZr2Xb0ow3MU8QNEdgaWdTPp0kBnXD3D38KgPKAK+PwQ6LkYCitifY9JO6owy7
JOiCCAgTimfA+VtcjicazuSm6d+Q+/iE2QiNH/e1W2ANgQEfMl73YYz555BDC2yV
hKGrAheXq9xapneJSnYfLBUsR7eRCYFFyqX4jCxVlvq8IycPL1L6wr325PcS3dlD
T6PfomD+7lvprOokiOYdIZNe2BRg7T/lQldAYD0/bLqMTxi6BARhAS5Di7j3uV4G
j/uOsluK/NA708vrqQKuxTmLY6ICOSS3Be4l7QP7kQ/DZfSlREfCiGtnrraSR83d
3lgWMnwt6BUw+2urQhlM08mV/H4SgzkF37XTU+yg87nAtjFY1bXgS9aLZf6TrAt2
+ff96UigGY/knoPKE4Z3u+w+kO5/Ay2h7iGiPazdfrHlK0hQVNOA2iHCknr5Jv1o
mfADgOq5dvIQRhfMEoYZsYvY/Xn7+WPl4w4Q9tl2m4A6QzTot2MyxS/VnWDiiQVu
i7L5GYgDIGWaB1ejnOch7AL6/PrvIDGy2gIblhKEHQesyID+2xRyFzQ7ynBSv4VM
bCI+dxWnBYfjtYid4kCXgflNZGWvpo5Rxb9s1vrvTC+XRtPqRCw7h5DTaKVUkcaz
iA54PCE5kULlF8Ugh3R/DxvqyzMNytG3sCL41Et9IzbtxjoiQpZnHGuZAqygVoU6
1V+PNhXXzwzZ0n+IrY4fFkdbM+q/O979njUF4HHabT93o68i/7XGvbAr0NPE9mld
YaH8zm9H4hzoGFc4r6AXE6tHaBvg2cDH1pkjC14A6uT4TUQ/tX9l3WrgcfcOF4sE
ddsAUaz/NKLb8/RVRZtWQbeAiqMz0CiAcKmyHX20knNziT8yZYn2FjSQtkJ8JKon
fZPRd/bopNLNqnTjv8Dh0xIWN7rvi5KoVbiyp72ZL+p3g8AMCK01kyEZywOgnSIy
hmcLm1urUuxIsMF+Dd/nHAThsAqqOAGsE1ibUij5PjsE1Ee3xHtzE3cT1f3PeDjw
nezcrDhnEf/pb8IhVcvb2ij3zCY3xPHIScvP0o6YMpiuTs6BVFPqtzwKqKv2LZ1Z
B72/sDdF7Rm4h0NWMQVNozZ7KnAybyyUYQobzu2nImao7QaPKM9JYUTgWVbIyO9u
UJ5c6noxWJLO9gjxiYsuu+0t+aqlDdryKsmzBxfZifV9HdrqdV/x9ZVaMuSXo6uk
98jVVHVN26lRjFSZyZUbuv9RtCFBkdHTFIJmIQDMRDC27ltzuKWCuy6OVElIkna0
vlVWVdFiAAE5WYb3Ui5Y5tR3YPmy9vzLiSvsmfqseumBpyqPABQDxC+unbWrY7p8
vXJjCUvCHbk0nRV8pGjrH3iC84ugeliXzbcblhUoIBER5QlmjEVymR+SnewdxR74
PexGIb6OLHxTaj57YekCKjgbuAhdF4Hwf86d083HWjLBZsrXOGVOkGqO5aGubFiS
0Hn16wLajuU0Qy0NXPPwLF6o0jr8amBWfxdMxnpFOFnIuoQ25rQK21Am3FuMB2hS
x06Glx38wnfCNz0N3Y+xEmQQ/t02EUoKu5sJKXhYydwU3UjU43aHpQAKHnRV7CIX
eOhSJIZ5Bp47dc8hd5v8u6CSzcaMjOXi2E6IXFMegrz3zagMm/VPTvRl/SiEQhbT
N7c4YQbAFdZewrp9N1tmALIx+s0dN2mtJIxXmBq0PPHS16+x+2AGw2z342U8SNJa
y9v5uLEe/Swx7M51Rm7GMbK3RSw1+/mBUESXFL14qu2DEiQjbsCVMSM+EFViU6zt
n56hu6yGwY2G9O4Nl4Vc81yXF4AfehIKujO4q6IPCvbFezQ+hCmxDfNJhs91Nv43
m+TPiATN19EmocpL2bH4D/9dPISLy1VCQkFTgytX8RrTG4LFZEBFFxnvOBi4Rjhi
6wxjRH2mVSmQM0LJKUyVRmFTtykm9IKFyJbnUcJSFOQ57LuLFW+5yfsldJ2137le
foVI+wYxipNfS/975IRViJcLES7d79257pXpNZ580FpmF83mdiz2EmCJZSPWmqiV
wStuSzZIEIpYsSDON53VjF4X2e17LuU6ZUfYQ3OrZvNIflHIgSHNka/ga8tesQkQ
dXpGuTzNT/Qh4dnfnkPWAWA/pkCqzcto/p2Cjmu6lMfBm783RfIeM5YykGfUnVTr
FxKFvukhq0ES4TL73WWiFvyTAug/FOSllhTF2qilOoR6exHfgwUuEqAhqtDo3q+D
lY1LRA5GI/CmwE9MO5uLrNIbnf/rgsOyiF62Zjd7Gv5AHHloaacC29B+GRS+uEDK
zH7vrPupxX6a6mKGyNCPiQp6LNAxRKZehTrogBv6zJOT0xutWwJzNNKVFOAfDOrb
e7zixW/lCxxBbiX6WGBA018GAtzWcsrW09Uj6Z+IixpTA7NQb4d8lG2EIHT8uYeI
n8rXU+a5urta5gyPuuquSKmg5mKGSNO9miEz+2cSRR6MYnOIl5CNo5feNpaXts5b
H9BB96oa4UkXrcn46k7WEA/QKmc4cYS1rhbO1BPpZZisYthEQMSh9XsJue5jZkLF
bROXHABmHF+FsTMy6IUd0r9x7D+ZwgdwKa5zk+KzS4snLMPTkhcBmvg9fU5tDvhi
sZ3T8HhQrlpnMwuUQNWMMDpxfMSufs2jDBWsI0XuzW8UPL6L8AMpotOab6YZ2jtR
NcMLcUpV3FTvYJ8qNOrbEGFc+fkLdHuHh6+c+04qw/W2zdNrO/hmF3tG0FsGSB8K
LDgS0SS1uJHmY3VBob2uK1PxYGXFjkUKsUWrwnneqIWDRECAbnkcd4wGsW8jhjTm
+p8VL3VmtFb/UnCAhVE4VKEXrj2eCOhBpqT+nLAwpHH9MUlcf4Fa1SjNTRJP7J+8
8G9Yb0DNuGWom3R1wMpeRaiN3kqB/8cS0h097WSC9AP//HlJ0iDAHcu1bAI0EnpW
QqCzRLbzu3r06cIDZZCiEfn/ll7ITnaY9t45mb4UJ8wfq+h2ffUph0QdodeRd4Ov
1UqCt/eye9W9D7G5jZVlb30sPlXlhWNxMrDbCZaPJuvVZsXiyrvNXEpa+zvcMrH0
pKX9qttyBOQ56MuodYKyDHKsFhN2ifaMu1ZEf4u5SMT7b6ePTwSIbXWozbQBR+6e
NVqVsVJ+sP+OH9+AqLWEWJ3kRRBwFpxvi/UKXXJhD8JmYzEP46yn9BjV43z34mbH
b02YCrmRhswvmr5/e8mSpN3iKeoXDvRMIWThWSbtE5w+D6sP0pp1rVn3C4UxdeCi
OpNr0g+MfHYTHTTHmjsfF9WA47SMW48LElA06xN1uwpeoxLd2NJJkXMG5EAYI1rK
iKQtRZUFJPqMVHLv2OnphHGDTfLl4hcK5KYlX57HxAhWZ2gmPgeEQO7vdr+x1Dtc
ScsccY5c9IGjUEa1UhD4EPhQbruGctP0LjGRYCPuFmH9zNAV1i272cVVzeNtBMdN
Z4AnLHHboVRcE6z/D50P7gIzqo1cnXXZKxdbnl4rcLEiLx5kXMSH/YCwCDXRNr5o
U+NjWv3b154ikeIlQPsksimupWoO5Uzfn5blXEfdXRnM1T/5Mc5K0j5qEv0M/70s
uD9blCeBR7iyi39AHtWpkrq/dzGKicY+u5YcgTfOaO8CdzoymIa7r8Lwg4VLotUY
1ak9XLtz20w9ZLmiAasy6zuU2w4zVLKFqrOgShNVTp/bz9FHr5fKprppUkmUew/J
hlERrDj4/T8+xyxJSSUbkPe9/NirZvJN/opmfOPjzpcX35mf14/B2g4APxjhg4Il
fEM92K81lbBGGQtyQZHgjfoObmUBUW4w8hukoTPqByY38GTSWZB/T99Dl+h7CQA7
TyPk29p1GD9gHnMq0f3br9fDK0/HrZgjR+BXrCpSNuPwn55S0lLiGAPPCIUm5/bh
HbakDx2+ALo3pF72GtsBEjuFsnGKXjOH+UENhMUciBJP6uqjd6qigDawGypbDScT
zmlAYF7H1UtolSTMJvPU7SbsYkxGj5r+rEJuzsp4JwNdMNhZu4yy+AtVPau09bPg
uppnAC2aGxBYcxw/7/t+Azny17v0e0rSzJ+1BWah3JnyMRaVa95ToiK9UGxdkFbV
5yEk4evs7ahkdXEGrTkra4+Dhm+L5Pqdvh8G5LZV/3iC7HSxUF9sv4t9MzxwYh0N
BppDsEeCmM6b/iDeOjKsEnkN12anKT6QGJqV6p6mjJv+gEYflPB6kBzuZy0ABlv1
CDJJTkGxE05J6k19IMSG8FK2UwzpHrAerfSRdfg4pykMdU5sHrr8EZyrnizF1lrU
`pragma protect end_protected
