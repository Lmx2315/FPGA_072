// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:36:52 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
O8S2Su3LEXrwy8dI6DmJlSbWAnwmDx1BdKGoJ8mC8y2/5UmrsBRj2oOPUdU4Rz0I
Mug2QI5Dl/MjtdgjclZZYKqZmN0Arve0ls2vWTygsR18KWyRJ8Gn865HrV+iXREN
V0VHUJYcnMMPvRkQw25YPBCjiZSbmVqq/VLl9JVecWU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5712)
RMxqGqC8jae3kV0ZfWhaFGl51PPMVIevWuhyBPbe3LdjPK9xfr28qD4dHDtbf1GV
t+MSu81qG00hfpRJM/1nkZplgc5gwDZQZokCxgPj/4C95trRTFC+A0HacvriQea/
cf2Ddr1h0c/Z6MDwTsildN68CiD2LvPZi21s1q5g6ri5qFDIvX3fqKYdnm7QozP/
8bsbyRw+AcvMLv2mg0nW7RprQAPJ+WY5lSTb7YYjEJQmJ/IAijc2jEFh3FKycxBg
pyNQ0zoOjZDOUE0VNr9yZqnaFHEXIgrwnv2K47ERJ5QoGMoQX1vHUXhP5gmrbUMC
OigtWWwsfOBICKa05ia5IfVS4n+jlbsx1p7T3kQuOXmA4Mo5KOTN1XrNTWEqcVXU
7+0qA9l/Gk+MsEEeBS4HPuBt1OCZoqLy0Jd8XVRMP+FtHG0NzGKQywjfNnwOS9JB
UaQHEspkSAK3pvCdLJMj3WB3N3+tqkzohQwbk/xYDrFqfITpuz9OGDUeeAUXcitQ
WZ0CVsgnooCbNluACFugzTm1fJ3NizWZWLvdyBI5JVVQsuWmWiS2NIWRNt88CLcH
CUsFxdKheLH8tI6SX7lnQYuUqAGhE+tj374wip0kY+WVJaDxjkQ4j2gyq7RtRXUb
yaN4e8SnOKqm88/Ax6WYrEKUsVWV013lVI7fWcXNtEQQqJb8/P6FuXniVPnipxc6
Me5pEY4bLZCJyH/uOyvim++mIqhfzcpb2qWLIIpzf5WF5gJGLW3s0KOYHfY2WGCC
FLQ6JKSjQlj9OntYMQzK7KZNz4ssPzC6ZlN2dug5uDa76BeQRR4OW9xjwOLZLkLD
sMeIVZzpXYSASbibI3/R2gL/v5KWe3pFZeGgC1GZQ6dhCuwLR/uH8BsOrMgttxRm
ujx9WVZ2Q+qaPZtbYOGn+CN9ygmbyEfA9AXRoaJcH7Wnk/6nVLh+KgtAyXuiTe4Y
2NEoZdkgFZq89znw+TV0jjeRIoH6y7pL3DcNtxFry/O3K0hoFQClFnFMQDmRksH5
XkyyVsS6yO53b7gfoKRj1gfoxvq4TLy5AVRjTWIAAC85tKRHRbs04r9t4ZmAfLkN
tB2r94PU46CNjjzZc39Vfj6JswCgZStIVuirg9ovTgy6aMqfNliO4G9kQfvEx12K
dyom/B66qS/4HcKhgKDDIAW5eM4YscKdwnwBES0whinwiwgUtXIp7zkFHNui9Wk6
S+aKQ10pEEQ4CcgSZnj00RuSa8prMF/d7kEmtWNq2xl/KRcat0sSGZiBz3e4CYzW
nf03hQL8kJgx0Ex7Br+qdbVYrGwiJ/hlNw/FGyPWRxIdcN2jtMyxOAHmIJ64hIPy
fL/4N1E/8uNQ0RKWCXkogxLQlUnYSdmJg+otMt1dhaCd6KAHp+hVoDxFEUtOIBtT
THWDQCy9ZhbWASVh1SkKHuKCAOyIdM6dM6jv91RWzwdWRkxNxGz4mEgqxtDZ1LOs
S2c4thg2tRV8r7CLs7toKrBpU2GYV3vyrVyY1i0QYNTcdF0foiFgxbJzXCjpmEyO
3Cor8VhgEDmxYgfsn6g7w6GiC1h6fUIzbl8PAFuTq0kmOYDTp32OvFAM4fDKDpGS
WzPe1FVUEEsyxUtGnuwfmNEcQTrlwUP0edinATunSI49eKvtOrzCjVsetetvff1R
7tGD0Ji0avXxEECkV9HXSqE4QqNLnusnnZntN02vu3swtuL1bPXR1gF9j71mtOhm
xHkK6Tqu7jevqw1n5nYPEdMeN0Wlu0DxjFVqONxh+aNzKtpIf3B4JxfWQ/0dNGlO
HKB8vjESkgllEXA36n7Wv8BbTxXg4aNsvbg+xKo+nuuN/q4H3ZpP3g5bK9wzWwPn
j+EZdb0Z3Oglx3CiJ0guo1Ibr5eX5wjC3MxY9A+AyI4dka00fpySkqoXr89iwtDD
IQ43wa2dcjbQ9UmYwte2xCqIQl0b/A8KmiLoRRbtZvzdaRqvxyzkWMoW4GAoCbJj
6PvkHlbPjG1HzFjsRP6JBXtWHk9hqTZzdssbggXOtqEY7/eHTbeXGzm9usWXY0Lz
G4SUUOPi53JderGiz9AQQ560/1cP+H12LeAAHo43fXEjGwms/I3PaMT2uE9IyvBc
Oms8+Q17U9IiJskM3bigurNcDo3w8P6QbmV1CUKNWDATAuqKNICni5afLBLPglz1
r0QLikxCeViSQGujseUJLBXCCa3bl5LvSJgn1yXRjza/65+WpqXv2hvp3BEia372
RQjPqjc3pb2OvespOfyzHIk3fIhPzRExXhzpdlAJPTXpvOXKn168WKBcP5vKJvcY
G1uQejxxYBAOxRCwJjP1JXeq6AYEhPkRMoVtb5fRgZQjjQ6j+b+EtBN/zfjH2mjJ
hUo9qqtJIuxPQ4aHu5F2XPa1LHmXEBbhh86uylgI3tD3MVPf1jb4c2l/J+6ZvBJb
2uxnxeYgJgoa2gkBocagqkUMd+oW2KKp8kMS8iSE51i35X76HyTSPmyhxwSGq5x9
3gAOKFi0ThFswPd4s+fgt/3EqOOkgswOF3mLEcW73EVZ+pcY9Efh+haAH4gcjYsg
2uY2IjSX7qRlgPxXGzkRYv34S0tSc46n9x59hAEibapD6h9LTpeA4C1VN9GxBzfS
i8V2okNDK0fmpvXGjF+Bs1RPBh91itZa8W0Cy/HyZz70LxXo48uQBpagv36R32/e
at6XeE8Kfqz58qzs+r4X/WTNE5OvN9rH6KCp7xWJfq1fAF/I3LehZ3MsNfKa95Xx
5J2cHVZ2x/eL+U6xdDr/RbzpTGogW2soAzyf9caIDFS6GbLU1HxL56AapkG8++x+
Jyk4+AeisDctaW+ScLmYDuA6WJlh6KCs+uHp/StfgIM4ndnEcsr1QXGWa1qYcCTQ
W59jAGpqCx3BQ591YBJRMUHNYMM4KA6In0/3yvJzbm16vsyaZEOCEkRQKxgfZIow
8qd45y72rzvTrxwjxqOdTu63BRoy87TBnTjEk7u2j9TxPk91QNgjPoNPS2DMcqmN
cdHs/OtwpoiKxuzWYWaZ0q/Hmdv1S7iVYZcvruQ7MRd6SpDGHDfD08DMs5C+95kx
4uwJReO1i+srtg1zRJnpVH9VzTfimxPw61+wXYlQRWM9OQgNL2W03CROCl5kIZrG
i4rj50ncDq81tSadhbiw4ONTmQgRUHxDzctr1/UYY1nZv8faeDwshq5BIeLPo5AP
mIQUCUh6ZnBhu8Fp5bEg/H/gmaSoGQTrOysq5ja8hszuTgi6/3CO4rg9DQxhiyge
RRJT1u3KvxEcqghA1r+bFanB3Z+evB1U1qFBSdV5CTul6H6GptsCb037WET5Ijoa
nCrSpstBe3McfgibLf0SwQP9vaoReUU06KMD3dju80EeqTrPX2WgwOXLGmpjkxAE
tMgmCjQ6O9MNF+j9zqVkLcaHvkR15Uam4A+mYbgkvkXHPS/2mnCuZqEmZHgV7PCy
19EH3Eelsy/rg9bgFyJulTxWcWIghhJyHxYmxfZRPwvua7wCB7FFuQVK63ldfoQK
wUIXAC/vsfOgTO16eh9ZWi2HfIK+fp8sYEcZZoO5p3ZzCb4cqrmQ3PY/eKFjcXRE
dHLOBvNUAEjH3UYSID0qSZOfc5tLB2nSWCH82HRsYQNUxXr1l5+RtvkJXDePDKZf
rOdFLgSifxjsTZSblJ1Pn0mqnWbBnw/qkWbsxjcmEkMJw5Vj7jXaqbzy88md5Ix2
ZO66VaypEkSMwFp/AxzGOVRvVqQquyTBobwBMtZU1yvXFQr6Bhmqy3tCN+ZpmhCz
O6CcQtIaZ+QEUgpYzKZhn2CUntvGrjZEEw+PxFXgR1WkPKFSzpFxR3fTW4XLZR4k
oUrvabqDwHsupqSQoRdT3TPqLrVp1BmLRlENAXv3D0juWej8/cO5+qSgTtfprwvo
bCV85gGxfCdfciWkeTuzUBKKd0kg238MkjzNto9MUYwWc2M52X0j39L35e52sxUD
an2tbPGOT9GD4+Ac+/ISvsFG3HoZCjaJcN8eUo7qLMNlunPwijh0Dq7K929rvQSw
ubccswJgAdcIxvXHT+3/l30H3A3mdZPZ2GK/F4oI3SQljCOpuwi8RtDUjwMXt4TJ
sbrMyZt6npTzOy8r6JF/gTHjQAE2a2YKGIJimUBcc9Uibfp60js0ngQvZjh4LX4r
nAJg9jnLjzCWUsmrVAUA615amt75VHv7TvMi/LjbsolzEYrGRi7R8HqBzy6LeSY3
AIZMhciriwwdZvizd3yA7ezPHRtZHM/Mdr9JNoKcWHKa5a16YucxlW++BDCRgOO5
al/W+wjGmnW8Za/8LKsOxZ8bTOIJ3FDnf85O6fKqk462j1dE7phNNpbbSjl+MBSN
8/1X4Drh4lfIWEYsBr/i2JltwPbS+r7IQgm/lScfMf6z7ePV/AqD2zMvsLR5yteD
iLz2etSTE6Ku0JJHlAelLbALD1xyv1kEWkEQmTfPc9G2l+VpUg8abMN1HUYPGn7e
glF2DOH6hF35lCkGAkwJ1xEZRt0WJSIEMMsv+keOvR/I0L0G6tG0zjk4+6xvWb90
jZXo5v4Opx0osKZbMzwAX7eA9+PfEzTPu9zIKmxKwZ97pHzvdgMNDndFWeP1P+ZI
g1GRwTyB8SpL3ZgsHtLP3VNKQgGxZ2fQvuqWldvEm/LTO+eHDCG7TaY91FTyq/rN
JTc6LCTaR0awBO6iPSj1bOTcY6GbS4ZB7pqiuZqwgY4rhbVShb/hVFIFloqd9viC
b6YVa2Nyh1YFNVROCKBAqDlp0rpHmtIFU3mfm4m4wtZegbutDF3E3OIghFmBTj3w
W7+hVGye5Wv5fiGXb1FetIMWq370mdphDDCvjEIwG+4VF4lE44dq6ZUpmde2eBvK
HIxqAGPDxH7IDE24R7oaMq52pQ8Ya5wZEUXxNETRd7MjOTCqpPxOg8jSwB7mUfiW
TKRLyF7f+rWOKT4kLrN1V8VKZSOY/VepjtgDUU+GJ8N+NzoCmgXIedGqAb/fBBip
3S+gQzirBnFmSvYRoIitZAIhrcImSOWYgCZXVhGoi5RnWuvVAAO7gNM1vOLIylNo
RTHs26Nd9WLSzU9yJlUpVgvvBnvdli3SRWDE+KXJYh07YXKuOcysuovYG1BV0gT8
ESkf+OOI8FVcgAFxwSEglsOWWW0Z5xtn4KNCbXXaeadkhGQpAr+R4kg1b4RZapEG
BGYnJdhB2Ch2LEoXiFDXVVkZk/lj0zOj1pKW1VDOPtWvrjHqlpzCftdLjAOAdfLI
SW8qqzM0P0o+aMVFkoG8eNqBBcNnFiQFKGz7uAfuEis5N5ZUdioIjR9PWuUd3Cu8
yubCyCoMyXv2bBQAOXQwALQFPTyQWGyTEXg1armGAu6yWuvOw83ng4g58mgjrOeE
V3soNA7YyuOMcEJoj+3gm9TNU1niwNOvzdA8R//ZTAwEuKAW6WHhU2DbsnzkHrqc
ABuJ2RHqggNMiwBx4WWasO2vJSjCY/e/bGOcrA1cUIhDMpU0eO3B3XrKDcNM2YUo
rkzJfr9awkoaV/ronXZeNdtuJKc/LKuksoGLwgjWglIcUUMHvO6+byVgPcNZ9tEY
A8Dc+RwOgQClGMSP5zXeDkoiOQGSqhWo0wTnBnsbCCZ/QgKRj3ZxCC6fdQx/Cq1d
L6X/1jJ+znSORH/RUxhAF7h0pdpmDMmprWW7wjNIWdC/BM5KhcaAfNgA32XAfuPh
O/hqj8EwN9C0jCBX83RJVOqZI9t/9NYrln5K0S/MbtqIhsVOr819a1vM16sfrRqe
GJ86HGuAFTkZmD6Ar6LFqfUpuCwQPWJ8TYkAenWQt7zg0Xnmc9/9Ejxnr+5VxF/9
AqTdoNg+srkGwf2ZDbsAP5EeizrROlCJoiTLPgaRS4INhgHfsba/4ldYXeF9Nyhr
ToSiyaC8xaA2EqR0dal2qFfGKMjXPSrxdxY4YTXFTCXeB0PjKaF8XKCeq3B1GXS0
cAElPytnVVQnBLDvu4p+VLdwMq/ouNB38/s4PG3nVQkJY3zzz0ieM5yX3hgxFQ34
qA6GLrtXkBm9Xm1bt/cKdpdARPa3QJtdNEurPYcKmZSH6yrg5u21KGFxwfQSKT4X
KS/EiPCxc05q6CqiJ9BOCwZ/qSw1OdSWqAXlW5dydNJ3WsxxNSZKDXAPKemKbhW9
YQCQqqark5H+/5ItAjNHYuzSm/palltgi8CitaUT+Dqi1kn9P1JaIJUhS1/kXAb3
FYnM1FeZuoeAnGtDN3zKQW8zCCCVVBV5l7jqWeD5mNVK0otyB2WrsSKFGd1EmxbN
uNFzTfqVcopmBKjm/zpsl2iT37EefNTi1zCDcW/ipr6txIuYRGNqaM8RKf6YirPW
mZJPqYBefsM8V026rcQ+2Dgch0a4aId66r7Cz5MFaDQoxVj++N/mrkgyknr+u4BN
kI3Zq+M0VIByrFB23yNibX2QBs+ArGlsAWGF17vwEwvbfzhX/Nwk2QskS2nHp6iP
8/0FzYSBYhT1qO2cgF5w3tSLmVgdJAua2p9gutYMOtJBB0kusQpbofQcnIPiCjXH
zipwLNB5wTgrLEri4/upzW+8nrkOIzWGd+ao2LYeZ9u6tDBW7Psz0BQ+2qtkmHd4
4lxuj/vuxQLtGDOU4b656xsCipXAWr7A/P3Vh7XlJFcdR9YdVuzWUf46RxeMHFJc
25zzAJzn7/PdmQs1CU1qJjNWohq5Rtt5pXyWTazteB6Q+Q9gZMo5C5xzxFEzyjF9
VOGVtnVKLd6r/v8A0wiigWxPU4+9E1PKDgFYR6Yo8mHvYLBhIqHXM7rp1XtdHTeM
3ApbwphCuCtiXZMVPKaaTL/eIeGaJnMDp24VmoNBvt6c/1NcW+uX8AGQNzHB+uQ/
M15K69rwtHGp9CD1On/rcYV7dipRf6Lrn77kzqhYhKbdSbN1zUw8lEQiCGIoqJHt
YP+NHefJdDhudjX6hNTmBrgGp2qmpqijWDD4FAW8a03Jr1ObmokDtK73irHUaIPQ
UyFaGUen6slmizyOJZWlhonn+QOXWIz/IVzqSR6KMlKNWgZz8Paxw5cb2tuPLADL
y3nbDMddjC0Zvtf8VdE/pp4NMciObM4rLjhuMfH8lDP3WFUJfm+QYOS6ThujNW1o
cRqB7VGF4UfuxWLnHqQImlooM9WxtNMMl3QWKq6uPUyjKiduRmS0TnG7seIYCSsN
/uMGjgzxQ4I+FSEJr06n5A1R/ln8SFvv/n9ypztwEPT/pSLYZ4a7rSAmLtDAFj0u
mi2+vH0R0NIp2V3YOO4xvK5ncqAu6BqREbdWVMTQbWbrLaHjRSCUp5MWLcpBY7oU
incY4MoL4lyu94h5jOANQQvg3If4dfu8/tRWPqLbdckrjS2OtA+CPMCugh2eGnZS
eFWYhTaB3GTn03Jf7wlSol+Q0Yi/H2/5dCPig+gZRvdse2V6wjwi/EsQOCg+3pAf
Hy7H0eQ08EuF5zNOu+RxEoUEd+kAkcfRYoLv5mkswS0+RjrYEckeLC4q7wF3Phij
D0YxxhNlTs0EP2oLCaIT0zgiMh8JIHve2+0N9nrJJFFrGL4RRr16Ef8rkkrZYc9r
6p7HBtBYYUQntBYOc3Nk5amVXhIQ+aBJqlHckk12MstUtR5fHEsgLsdQ9hHhWlh6
`pragma protect end_protected
