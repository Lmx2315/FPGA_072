// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:32:38 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
O6pddKiPyujonZy1raDKf7lA637hv9HIVNb58oEzpVRWtzUBghFboeo+6Rz8l3aE
lbWxlfFKsWP256NLBcc+BxalIUd8QqCybmdGX6JUmg0lgKGA6K5ASHqBZ9gkRg/v
mVLvTBME0s0Q9K3YHZh6AyXBemXUyDv8jQud5JGitZQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8400)
aoo4YsmaRnKpuCgz2QK8qcfVtCcGHVk14CiEwFURQI2PzUVAuYc0OfXRCEaXVKVJ
gv1PFf0HHY4hpZkcpS+3n0Mlxv8MaW4WKHGzgCgVY5R4KCFd1pyN+86UDemGIHBX
77RVZK8J8smVkoybKEHGBk5qzrUOXakuDl5Cf1IYsdaX8yKxNDfCuI+f8m3D6t6j
7ZWKnRCkp8G20w+i0ZrqW8UMR6xvnZWPF46tMPbaD8xDRX+nS9ckJaE5ld++mzOU
nUKDoLPqZmQqHZfeVv4kZy3fQdzjpu8iRc1/vbYIeuEikCzCdfvYAO6FDT11WnbG
zbJU8zERxc4vDkg+lI5ovsWXj+RPw6608eE5XXCrvD1hdq+s7Tvqa6U47jbDdouj
IRFaUujZW5LUiXOfj05Jk2vTwFIXHOlrvod7QH2vexN2Vo/OV6MVq9moqtBjqHgd
nnOC9EgrsHeHSwZNHQZ9N10wJQb/NW0zVjdJsPd5tn/a1hRHyes9+DwYtI8FZLmB
GUeu4VEwU6d4EourcDCZ5siFQgPD0/LQ4/bzHiKb9Yt9MDxs3cohpxM+DYHFI0fx
zhLogxX6vN4XliIzdMSEJ/MwGrQPnBFBq8RP9NFKwfj5zGtuAwSdj1jSrq6ZGkns
93aeKa3blY901Ty7l3HmJy9cUcRePzm10MCIcTtoDn8SLyXM4q6g1XO/gEjs66DM
/2AK+xHtOKwea8t90oFniZtxVxljT/tSTjKEMLVZONFeFDwM88XIm7vS5B/qTkig
BAWMW2vf5satNsF0YXzA2jrJsKE3siwh812YeyiNNq4Jw01WzFFLQhsi/F8HF7iw
Iu0lFP4n/0CLEHf/DwqSzd+2kn/Y7pOVA0oA5OzYsMtyVZQgTUoHFg9WLx6Ua3if
l8vzj6L1C8ptIyWjyqLN2ltXM4ix/Tw8ehX0OIRNG41dxqU0hL27p+NDyaDe4R5D
/4YlmvoRn9NVaaOOBKadgxFG8yq+Z3Mo4+Gklkk3Wts7jEbZuT4cGdmN3c4IAasW
pt9wCq+S7D57HgNOKCglh9kcvVBjd5Q9809OaZF+clqH9mRTKq95g/AWalVF6yuR
597E/baYjxDBhafVLPXxyl8rQI+ATAKPhIgTGaijO3/7yQgPzEdsCo34cpgIU4Pz
yKAeVs3hC0kNAyOZt73ViB/pDfnvidgPi6FBCRofDhGVmrjH16HEwh7zjgVV16vE
VLASuoQACS2q+2w4Xz4QR1pmfKHxZROvZsh/ysRRnYda3LQ6sEeC/BVjXXInF+Cl
NIomNoN8GEt8gVWZg/GMZoJ2KuMyynfPKOVZVoOOWbw1to0s9ZEBU8ZQtP4zoEqR
bD1IuVNny/6NQ5w05hvu78br6jCaeTxBV6rU0yjPfPRa9CTWvA9he9XwRDujRXDJ
XTY3Qi/+66ZrrEg4t4WKCAug4oQ+34jSgwJODiM2P76J7ezfZMH40+vP89+bOO1u
LFBznanA6/IUvjMkFGPwvvXxuwPEm2w8Jm24JCHH+MaNVfl0v0+bwqFTh5oBnb62
eVoREScURBFmOHkojQ8In394V5vuMFA95DeNk3cj0+qplzO1N77OaAZWW1tg6xAP
pcZS1juCm3ea97tQtRBFEwL7ad9CSOe81d03OFSp/Cl/j6mu510ys+5UgY80QYPz
uiqyVqAlxrHJlkJOm68cEZQE8J6RHCMqH7hJjrlVt7WPUONHW43Gope8C7Mplzky
j+D1GQ9r4iq4XyoaFwxfW/SfgnFPEpcKWlM7U7U3CYdieE3fePtskh13D49Jjq5U
AbWy3zWBGouMVJrDWPs0ClUAInahQprTCwkKQS74Ip+JdoFFYHzeRtRMk+7iJwqm
Q9e40Zjngo1YxXjMSZVwuSEqgdZnu2v5wcuaYP0Atd1Vjk5lT/Tbltln3+gpr6Bx
xkF+b6vply+4DzIqcmvYHZpARLHwbtpvjvGgwyU/9wU5RQzz348hd3pyBlerosEA
qQKbwVI8NDLr+xM20p4oiTBs1dUqpvwb1Y0FCg3CWZ7MPZ12n6C5RgCOW7kTftX8
di4YgT4zcKplfax1R6nx1TQg/+EqcBLXDf5iR8RlRlcy+CrW1WMEgq1BhpHsk1NG
SZu6bOAk8TSqi25Vu6qYxVrQYQVzKOM11GNl31AenYPb87+GDQnSDIwPGJEPkSCD
VfvmdWX+PbyMmC6RKUgJ/KfZyU1utgWFdrurfOtZVJ0H5rN5mPo1dT1cBrW3rq9Q
+1N2Sgl6jlhHkMLhyCULNc2B94Qt0V/Myeg1a76Fm565pKtb1QXUpAZO6Dnt/QOx
2Z2LOOkBuqFbp9FzfH5TCOzoyyoTzdP52FcDC+MM/jbNHKRjZLbGfpA/N7b4UeVH
Ia6O1JIGePyZLyh54Ls4ZySJQEXC+YuDYHIK0Ab2hN240m/0oCHwxmmCmnVjtg3F
6/QOL05EmaIeKuf2qIjH2NwPLjsx46mmI+cpc2OuBNPHhUrf7LgRYXjEcn5SyZUy
PkEVdpmmf8PKK6lDPKGz9xDURxLuP0qGpqo0ETh+8MtfckIO2hU4RMTRRl12JpCl
Jz1Fa+QPcMFET52FcO5EApKVcMePKpOGk+1jreVmv2sLLrL6A6GvBfaWs7QsNQnH
Q8Q7LMJbukeGXpZvaahgh9VfhxhTHmmL4spVF00ov9OmmKB0ehO4jdiaPrquhCC3
UDsnDxfj1/LG67Q+/UiaRCADoPVpEH+WuZ2p/xmmDkbzI4nvK9DeROHb4jTboT3u
5ooC85a6sUWosa1VWKP7K+ZXUTsK2mXUy3aBYbwNTVe86j6RpUn3ToRik1Vr9yC7
M9S6o3cEMYhM/FFJVdvBkv1l8VRGOc/XYiy0PemT9WxH9yLaX4KLhfOGtSdaxVUo
s9CiMC18Il2moCAcOcOj6hJ03wpcmxuVA2D7CK4zriMQAtc+QqG6fnP8xHLxs18Q
MUbQd7I5TXp+djzjKL30lVGbyChj36iX0wOnZSEZw+1ntXtXenoF2SmLGZ/+Ilec
ehqiv2lxoW12MltzUyCx69ZDRhHw65/PcdyBBYijF8o01jJUF3EMVH81bf17+hWH
eoE/X1YjoXx6EibI9sax23YFLEC2R6MDns7nNGsjXqu//ZZh+VD5lak+VDXbPhf6
7WVb+awRrvpyJTuq2fOudFI1jXaXt+XYQQMBXubF3C+w7xs6lDFjYnt89II20drF
X3qr0LDuvbr460L+rJ8xdWLFK2iJISiNBlu6mOFP9n97gN6oFiCW65ntpY0n7kfV
vFQ4j3DeEFqqy6CayeGnryeXB8tWd8ooohpQIWrwoA/QLPmcb+fBfmIgWEvbaIJ2
1yixkADoJBU447Qyi8w4XldU+TE0fKnJtkxXKrYpjLBx+f/hkbe7RHDkr+qIi2hm
aAFcnWjPxM6al1Dnk37bMJu473TicbJu/oGZw0XBP7LmicAJnn67My+jTrYDSqhg
2ERkQk0lLM+BanzKa4yilZjlyo9wDFYS7o7mGlCewbGiMDqNmI07TSGBlB3Qru+e
VNxqflrVTZqxBew42PYea8xkjNF9q6cHhyNbVIeQrlJDQhcTTy8xqsAycfjep5mc
1n8vPqTvN83BzzT5HHzhIN+R1SAz+3H65b4NzQZ31Q8ajzGItYsdMGkV43BGS5Nk
1ik/fZHa3K+YKBGWJ5jGTr+CVuFKgaPKEeE/v/yOIlGp8XRqtoRh8X0pduYxt7lE
Pc4JZm6LOiP1ZwTzAk6B2XFW/1D6XaFGkToEHJ4ClufXup/cO+yJw33b3NV21POb
xns/i8IJ1ML3ooryS0rS0WXzgqajAM3DB82vz2ysHGAJrnVenbAk/WSv9HbhXhCb
SaKX/TJF5hGc8aGJYFhF3iXf6KMza6wpAPTlYWp3whb7VFcNslg0golahBHeIKAB
EoX3Z2gLoe66EFM4i8hzm1oifNA7uZqGAZWQsf908lSFRvEBTxJCTwo3yfrJloSM
twbffK+Ih6YK/iyvexT5G+Z2mdi2TyXXvWs3aoZvEfp+b7QgoC6eKHtfUsqGumcO
4Mrv/GsqLP+9dfBTMXDkPjMYTMK0sWJwpVDKJ23kWjd4e/hFztWFxhPttCpmhzqJ
XqB2mbliEmeDv0E65Td79kZVxuFCGEW/vfs3pblosYFbVyZGEF6TrjH/vs9ru1km
ypla7utH/cf7elg0MXrXoybts17/2SWM+v3V8k2SvwBpihXlSUCU2g2u/Sx2UZEk
idlBYBGkp1DCO3YAQu1YdFfLIwqPuINRuIoLrTx20D2O1eRoUG/9N1rIOBPQuGVC
RZS+S2TwBHgVfmoccMGnqkJJ/qxVv9c+TPD8o/MzWIUvDli/VwhxOgRKaNU3znqC
XJgliFUOK6SC3R7WkgpvUAGTnf8+miai6Tzl9206Q4xYQXZwXKpX5cvztqZ8PCZj
10aUigUInLXAly4FvBAq42on6rCc+P7y/kfXAAf+Prp8bwwiJN7Ngem49synMoRq
ecYdmY2VLJcR58Y/YI1pWoPKFRgkB9HQAo2XnKfLxjrQbxkaKXdMmL/ciRgb71ab
OBJv/qQYC68k9ix8p2oNojRUFT+ROPeph7l4LEqd0y6q7KrpOaICJyntPlgsFumV
cApLusgQnXUcAk35dARdkqXvLdCzbknA5yAhAr6CULV3lsIwdREs6fghVRZDvhfh
hCft3xQMbM8/iI2yX66+dRIgRwOG7Pds6rXeHOJax6J2Ee/39gcPguOVV66t9/Sn
MNfCf3MV6yLpVyc6J70vtBBYoPjYW7SQXBUTbJPleVNj+RRUBpQrm9/bUJGGumzm
1WBaSuywnrJzW+NPAkJbLEbZol8hoKl7P1tIQ7t1Mj6HQI1EBmZRNiP+y5+hN3WX
Jl0aEUKm9aicXXGVs08WfLrznzT1u0LcjG+OxOfMZfpqj/WRrVZrr8sDbU6QAcYS
ZxmWxaK9tiln3QXfNqUrqWc9pIr2654k7mQnpX6w0ScYX6RVporScuYyGalt7ZUK
eiHas2/w/2P4DPdhjc8ZVWCf3ECzp+yZ3pRhE/ZmS/XO1pHPuPr8nkFTSaPlgMRv
UqBWypNKH3Zz+02JDrnTJqLGNfaUDX7g47LL+T/OAkpxsyqXZlEOYfrpP6nQU2sA
8GN2VTMcOZlcL7GZgNCQXqL1CJLdXzuHJjHWMsphQZ1rSiepjkDfXIq9O7xQxlJu
n4K4S1sw9VZW6cUV/hRAaWLoJOcYq1+M66U0py8++neOlWjJaIVPD8uUB4HI2t4k
gIXpzf2kEmg0HCtM0vWahUet/YyXVWEqpJQCR5jgxigEIDY4Dp2w1gwDA6OsSAU+
PSv55z7tXgx+Y/oxfMFCEgee1h8tsg23IC8yhLxmJtsi4umrySZIEHhi+VQNviKJ
KjvM+mlBHJOahPHutKtspfYpV3ZBVrQVjjB1HMByt4yP4FFI2mqTejkGF8l7vx0+
QoESbj8GrD0GaLicF4YnYOzcN4GkJVHNtDgTZQHsw1dPHpbxzmf6fAz/wP9hFS06
n0f5zg0z7hV10P4TGUTxJAMl656hBrzt6ebVq2CpYoqeF8lQNRE3eVufUaZWilBB
3eUQgQbXAxborvBZJ2o6g5AqNQ2oifIDK56f2l+5xeZSMzhnZ0XEm6Dr3OYVzyPK
2dEsCVGklTbW1oJ5Xv5HBz98GRAWATTA6RY2m5Qz7oRmqR2QJ+znkf4+ADwe6tLJ
w4umyd0EZ1QYI2rut60/N28VDeD2WfInWWk/46XRRBSiWatrNVOzXSOhcbvehOnG
DISY7ohN30AB/JwpJdsAMQ55puFvg0V/+8muk9Dw2CrJgnz9hYm2YjfMEd17w8S9
8XJFoQvQgTds5tqzQ7XZqwN/Uaqp0fTnH7s+K+kqCLSJ6JLOTuZo0vozgHx/uV+y
IgEYSf/XKVdnjUgrhX6FwcHxbT/mjRKN9/JNqiGDj6KulKZLuFfUkj7+uS2dZ+M5
Ry0aV3iRP72vMsevtlx1wNB781VLtSDiyKXnTLQi9tpnOIjHIsv3qIUEIPFsbBas
+mMRxUx0Becy4KaO4o8JtyUs92oW9gFyyX65KF9VQJLEfXUg4agVIxWFA2HR4wGF
1BeXuk6OWVFn95EVF+WUou97rIC/F3OzxSPS5iPA4lNAfr3xPcD5NM9BXIL0DsnP
jX0CsgUn/u/LMhRqVBT1IWr5UlsXzKNLVU3q3gYYxCPSdS5RivH41zVUjrn38moC
s60lYXRow/YbSCV233dpNvZiOFg1YHAlLWXHrZa+C8LYauw9s4btedYY4tEW3vG3
rnrZMvMX68D2yu4AjcB7zWxaVEtKvS7sS1vuGOj5GgzlCmQ5eFz7VaTfx7H2MJ3B
W9Ot91AaU/B44nKDyZ3bzfl3egBYfFTvjCnpIW7kSgI7Dde6f1sn0QPFgoApIIZE
eJ1mx2YHrPWjHeUGbe4rq2Jb/Y6oXUK6iT1/1RMDOnL4rfoc+Q9dWZ3GI48sM/Jc
4egFsKLnK5Pp1/eQ1OgI53Ug+1jYN80EHAG2zv9J06BKxElreMzKMkAu3AxUJFpi
TpuGz8ksUusGi16XqUTKLID37Srsgj29RHP3/K0fI+6JiRe06CoIRvDpCU0YXRIg
CurKonqKOVTSQ4MfWQgHkLT1SGf6egfDN9vbrZMFIzF8zroiG6QoishFqgZymckk
WF2mk6u1Et1fHyeKNKf7xeb5GmLZRq2HdlKDcVBkKIjHeoD40V5GOLf1CKCYhorU
Pfgx0ZwsHEj4AEskuJENp6opoKLZbip6Fw2i88AXQwdEapHAaL//AdJFUjF4RBIG
ajsnIwPGUSIA0i2ina3nU+sDZ1aF2Lu6EFU29+xkgt8up6BV3MsAh1xiULI21ZCL
G0ZOBwtUntkklgwjE7owMHkxJ1zlpedDFleaOJknn1dselJks6nU1BigsJjRuQrs
qtWnuenJkzIawg/iwwxPYyUlLLrtcsSTkGht378rv2gTKcnIDPzH7/brsOq/KNlM
Fy3yEaF8f/wGce12LN1Uz7T+jDpIAvCOvN2SLV5KcCxE1usTU2AfSTjGGfyg9wWZ
ta3ozUyCWDfNzNveV6tvJFBx6YsWtX4fEtldkwZKi7tT/xduu7Nvm62KJ5RQsUuL
3l7gFN5xWooJyog90s50uGomHFyuBQDcGfEFBoCwtk34Ptv5yMbiFlsXb3D6Gsxq
h89iQ3ykykBU/2WlbnExsURzCRRox8GZ7SRja9fcEEXJFsBpi+Tqg/3cOZrxnR7j
JXcefvAAKkTJlUyWzNoJLW3e0T4F4h3PmvSNd+EHQw+QzqW6vma+8ht3kl3hOQDh
JaIotw3w0lpnjwsdaZsxbGxVcJzYVmShtWBLQR7QKBNEy3U44CLg3r3L8RLVOmr4
ou8L7HWYljhYVPbd1Y/BF2+bsOCl4JniviCn4e6bKGept9tAzsR/Ig855faXF/n0
a3aqY6sceS3mMYODPl7tMxi+peSihmYtcAs7pXV9DNvc6V7S2tcEqfV2SU7Ei/uM
IErHaytCpaUrnoIpifyTc1zmu9veHONAIhjH9jT2mZ9crXZaPA6AzRNLw9wVbgxL
/SmSjL35ot9Qa447pSrmQopme9bgyNtkq+t0oPNfxGwEuazGLS8jwb1W06/XNQnU
YOIviea+6/EV8rmc438vytZmDEI2Mbu6fzSl8OagqzDGhSqmZxgrJRcKvDx9Ymov
gy29Q1RxB0JnliJqK/g1azuJlyqJ2nf0hNfWpLp2pr3r80HKNcV0yD8JBG3YC3bQ
BSjF5pVGOGpcP3h8+tX6CUA7uIiT+cTh0uRJUlRWEO9KFBtShwOMQgRonjwO5yvS
FF/iHuFhREUudcu/P2ETETqpl3DYlkliWnAGV5E7e3X5oUF9550aobR3btnwTJjj
GgrsrYfcBrF8FZfCOXnC3WtOLiI/ei6ueK5asNEdIvIFJBAkXb9vK7c+7q/lDa/6
W9WvIKoq+aRJscRjFhTiu7HAUBaRM/ZoAoNWYetkMtexwG+EzicRiY+RfKD6RSSa
P7psxgo2lnb2FbHFxezUWKRIy0QgOIquzF5rGFhmCc4as5Tmrx8pv12GappyqnYg
s24YXhW95lkv+yy7Idf0yaWdPGkxZatgfH8+l/7OYCAD7AoSNH0YOLojLvSI11TS
SPzJ/wgdpkx74VinlS7Pb8lS86ZgCWLitLE4kCXvTUF6M46bIgGl6tjEqQb+Gg8Z
nEqc4OToVl1VSCw5tG/vQLVF9lX//hbwG+mKomjA6jwXarFf4Izw0RuM15rzgjgW
lkfWAuQ7EoshlM8qw8yTD1Pj6AVX/8HdyQzE5nE6XwVnVBxP+8mCw1IEfqq6eFYA
TWMckpLJYoCI/8NLyUepKRpsTl7MCs7ZP4eSsQyQUhSxdPEnV17LhgyqwL3umywe
VHqHttOBKGvNLlF9NJOx9cssZnGS3E6joKAurc58DOZoq+JNA3QKJrmamn532F1W
j0hiu49dhClGiFV6kBKpyc7D3Devbh3D/RIC5dw4gR552RszybTMhN1VR1t86Nh4
f2+ZwfVCeJSvi1foyROe03xtUTXimBIVGNA3AgMRQyc8wKqFNCY8rhXSTjSAUqpa
WqvuTmbCee+FxDGONuoqqTAkG6gtlp0Cp+JgrAi7aCVV4Dsx0Dt5MQVqt4PkvVAg
PRgw8Pe/QQWoX1qbgMrDiqW+zu3W7fo5idZaQukllR722IjiKzQSzc5jiC6IrQBG
sexTCNpAfx4gK+Ve482Xa1Lbwt7wVkqBmXQOwpbGMPuKNHIeVfCRkdrTa6vlsCho
jJYeb7AQAtixjPLHvdpz9Cxb9eTinn0ElylPl6pR8AMZBzWZkQn1oabxkv5qX8Ma
5jAOiXzvWpr/SPjF8K9fvyDjvbg5gfFNwg2UHApntFpUhPPvKhlj9ZiwrX5JL/4w
HKugOqQpbXS9+yV8QndXRrawZfx+ZdgnpmRxdATLt06w2hBNJjHuBqdSJH0lbo9f
k/IJ2T755ZSqyHc4yjTRKylGcQSTLCsH+NpCkgMAK1sldxTwC+inK67uglII1WPP
iwrK7FTKtCuK0p7VRD7mzahmAZGjeX/9xbdVo2Mg/2E3j8QCm/9mH5BGYlAUZixD
Zr/U05EVq3ewQHjudC8KgyevF/YRAKXF3yCepcKryjzX0IGRDonKXZzevM5rViNH
/jgwBU8H8Kn2xwrhJa5HTqQvYB5mnDCSS4xjoupIN+5RJUDQDN8o6mGwdWOulrB1
VpT+qxtjxHxc+qAydTrpfr8Rm8ezGsfOsdGf57FJOpZ97R/+uIDiBOjrUuagjFWj
6XfhRT1bsfeXI1iJDAxMV8Owll+2GSWvg9xspexgtP+tCf4vRMyB5zL1TdQRn4UR
1CFloqKgdeisTdfANLnhYmFyShIq36K1KrcW0vkbGDoPgPnALmE9hHTYc3iS+hty
Y7lBznjF6ehj2eonaUI1Bs4w64P7EIeXJCju013gNHzzfA9rMQADOGlGW2jIa3ZI
3FhF4gjEi5t9Xn9QmXRWEgq0Tl09a9XRCRuK1adPGYB8o0Z8la8xHyW1EgKofSf2
FdecXtQ7TyKIyL4hmsZ6/4+perbyBBm7VmJYHwrOotG5+3BHPo4DmTIDjSsdZoLJ
CtSsBsrphF/3bt8aSZGqmeFwlY4NOH7XcrKIT9gFyahDGowDhDK9di1Kgov85JbJ
oytZaCNDnHiuXi2uMlhKLmNgKhRVflxEYjhi4DN19CpOYW53HdXvxTO8l4lszOTg
REflqzyEWfsveaKb0aJE00OBlZ6puAyWP4JagrtsN86Fh1JTT7Vnqq/CRWBqVPp3
k423nm5IVGf5T9j3UQ+edVs6tyxnuV33280XE0RrDHcGN9MOzMNQ0x9GW0o7Zj3x
EaFu3rozMJhlPM4A1XOkCtyRMVuf8NYYSWOTm1uUPWtJs3IT/Lzf3yK8Zr/uw8s7
DgFKewy+cyFZ4vubXfpH40EPTg4kXXAMt9IBlQ5VeM2VWiaFYDxIEeCayBXfSZxp
5A/OGkzqGNd1U+b46J1I7uTQr87lL824+3oJ32TVzlx7VMNKzBc1Jn/Q48nA63sA
b/pQ48YXSB2OaCvjCqssiKpgmMCLMQXixvwT2dIcVd/ATrEiMap/+plPpWj1QXpK
q/2npT0hYUy/GX+rNCECDpVMJKz3PmsEG2JUIuj5hVLNpkmUjTqev76HPDkg2lmE
fENIdMtDJD9KOO6Mu3E54lZmpB/RG7NyVn8lA9hjuG8nf1pbUGHtZQIGPhl5XM6Q
cKYA9e1ajA7Nl6y49LxRjKXCEA69vzFQuglrhXxRDYRxV5P0DK1b+b37TTb7tAo6
E8tSruHdL8RzwFGAWMbCTRe5KEUXUDM6y19GHZ2siPFB60sqqDtGMuR2n/HHxJ8z
F9idk8t0z4SuO7DOhozDmCkhO/krHxta6aave22ucBvKTbGjFWucUq2BGe/GesuD
ASr9e20h+7bcO/YUZjQNk201ehnlqfBLnGhaols12UNX8Q1IpjMS00MZ8M7R07jZ
EKDbRG0bermeh8EUYdr4rPkbszgbSG6kVzqax4ILoy3YDATtDXa+ytLJfJCZzSBt
lUKOYriFbsbyMW586Dmkloh0v/QzAb26NGHfvs0CNfwq7jPZNBFZTBqod/gvG6ow
zWbdlFkjNm8GQdCHTNTkrDMlXsVUzvhzno/qIpa4G2S3QHmFxtU128CRVwIPsK1b
jeL8+704c+TiL9GMbV2ZSJWOyfQWVMrEbS0BJjQy8fGgEAqwd3phrwu1nxDHgC1m
TsmhbPGXVBDbQakK3ptUBjh/70UCERgZgp6olnTkBpbRweZe4Uu36xEXWtf6fuc8
VaEKjQ7/AtEABy3SLKkLt96eWEent8B3CRDjwozF5uiMBPZkFyVEpAbTqgYRmWfK
oQSvb/QbsJEx+qMuK0YLHi5NIJkbfZg8ASJnz+eHOG9C7brh5+/nxxaOa1JnMh/y
uD2/5ExV+E4ksAhTamA07ZFJgX91cmRCBeZ6rQOng/+tsyWJm2oYS+rrH5/kqPPa
sglSZwislJlMHjcqjtHwgr4QfBvI6TcWk18Lz9i4Yo45zHDHZdILqmeQCfk+skgC
+bK3sGNvj2wQgputwAkEVNDCdm2ClsM4HyMmVhRh8SAfgLeRmhdbqii6lKtGqijN
fZHzatLVQ2O7GSotBynX4OeVrwdtCWd5TQhwTNd269Rdcn/C2tScX4vg+CMOk4WM
`pragma protect end_protected
