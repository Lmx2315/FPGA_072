// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:36:50 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
FQffKnCkcjR+oOveGCwAz5rpCv8BZmmXK8FW4WWUjk8ilq6sEYs2jxbiqQjvZqyC
QuJwB5bRjFQ2d4OEXPGkqgDTnI+h7JYQhkGIJfD2wP/1ufrpEk06wHL+wn/M2Hs1
CXczZyUDzya+28G5czvNfzl006wWtYFLmV6UEHLOJ3A=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3264)
ULvvCXEAgM8JloaHmcP4PKlfatY142/L/oJrv5CoJ5/FG5ZyLojmJooaQfr4XM+S
qFiN017wstZzJucTHfEb7Mh33llXUy1k5L260i+AAsSTnbSFYRuAn0Zik1hYNlnr
QPRHr6W+/OGCMZPG2JKvEUg759b1MyeKntTmhjzMbcAr2/4qHxjFKFHJrr4Q8iOx
h0s0mbfL/MVMPVLGZyfnZAr+kvmfALwF+5rXErlQSMOujIzbUJx1l/hIzbdyTbv6
lQQP6Kqv/xhGnDJdGC3IxTlvSRCbjr4CE3hpQhZ6gVuQcztf0QBSv0LoUAEShi1B
eP6KM9G+rEkzkPsLcuFj2HXpR8/jdp8SZN7dLxHKw0Wb4rj5cKNPnqvPscgV/4j5
NYpe7QwIK6EJlqydUaR97/MrljpTq64wCESEE/hVvOTpES3aB7uUqhIxW7Oly8tK
Hrk16JNDdqfrDzLqVVvSRI1452CFwPjKplmrop5mjcP6y6LAGJ4uIaKTwRcLwF7A
R3XMft47dqG3oKvlGGSNLixyH9FcDNH36G3+eej8NvnB04QL+PQ4/SltX6ojjHXW
EKr02mX62glA9dWXUkddye0PEVJoKWnhcT1BQDU2VUQvwD9NB21Gw88YtN2Zmkk6
4VoIzLJ2aB9dkuGBvJjxeE580taQ1v8KB4eQ7JAf0M/T0D17xUVQi6FvGiybcV1F
8C7O+f64STQ5vTf9vKj/zd95mY9n9p2ov8J+RzEdXDIt9SyW6cj+dlQ27jxIYeeY
TmbFBlgsuDlE9Io8xlZlfYsNAisWM4IRlx71tLzJzfh6LnYaN7axa6GK8uJlvDH+
Sf9tQLRv/ujOO8X49UMSMsjOLsZGbPYYm92EVaRQ6RZiUyK4JMBW2cNfCm3XDr7s
iV7HmVaa8Eis58jz030X2Bgp5dx0/c+9zK0wOh33FMXLPjp//8+ZGsfsN88KKX6X
J0qw2iAm1IGaapkkqMrl200NGS7wAG6727vqpiKEm2KtyTxWvbnFz9Immjfjzi0h
Y1fH0Sv+/pfH5lS0QjTfya9ofVxplK1+4fxx2CwIVM+jQ/nJKhW/ISjgYNOksxpm
s9xgRWBRqhkUm7DluUFR4nyeEkhIvZEvwbu3HAC2yTOFhyRDjJpq8pTrUxaWp6WM
SoDw5hLN9BnW+gPVuy7ayAco6xxmeFgtex/H4WPXV0dRLeQGfdumGuZPnHOZHirj
2J+rTYOddtjfITSgh/eLywT0gJH0IB0yUv7puzWLOcrvX9FhoVgl8X1WF70qag0B
BYhZXeh38obJ5G43fTNsWonk50H40N5iQLLjdvRHwnVIiauV15iMQ1zF78hoIp/l
BH9a8A9u6wb66Yjjv7IdwpHoOSqECsvZyZjCslaPcCDNELgZysR/EmDBQyFyK/4Y
IdxVQJs9lPtr/XjcpZtiAs9+rQDMifzZ8Io2TIua7Kvzpd2QqJMHRsOwRhEdjZlP
X6foB9DFqg7/BIrZkvb3P68lo73kaxM7k5ne6G9KjVbsiDQ0X1ul0pP3VB/GHttP
S5JnMhVQq9epNleEm8GevE0lONmmgQn2Rr0WTmCX1bKmoLIfuzERuvhlW7aiCu4T
dN7RuZk6mzyW040UaPDIPqR4IP2Kw4rY9gesmDAnd8ZkqlqcTpRIZ5sUUIPNdFwL
3OHQE7u+o4xVBce6Qr86EntIrV24RpI865Z8I1HdzTY92a8pPY3WOW8YSBKXFLQr
RQhEw+4BqzUazOzQ10aCT+rwNUtvZU7J6foPZc783LZiLO9yuYXmgpSKwo8CNhNV
kHL+Co9ILw3p9t0EDSLq15l27yTl7GCPDdlEtz6KGNfurlnd560RcGBaa7Y57Iav
/jRKKR1gWxHdG+/CFYL1EnJGnQI3CRabi9mCLwKM8kkR0KmNEDeOW8Duchg/a6lZ
dhXuxlJ9CeMSlkVp8fhX5wVjqI8qAuGruJt43AZ0RSMfY0CUiuzj3s21zUe9rEUV
o8E9Q2dwuuKCWLHk1akAHFj8IUWrsV52ItdHcwjJBNTRZw3phHzLr5d88wvlhDVB
1aM1Y9NkFqwk3c7txzv+ci10DRpfmCFu151LRGXgC81csgDM6MeobR7uV0xQhQEu
8YeR4Zhm3f7UhPnrGsv+PF3cnen22txxKKOw3cxwcStvEGFAny4hUDuG2l6hmql4
vQJ6XZR47T6Zz0m3CBt0sN+Taho242kgJJflmPDcOfCnfMbQoyp6kfftUFKUtAn0
UN3hp19c2gJxrX8KZq8C67A3LPYKKPwAKdD2mLaZqHpgGu8EpDNhvD9ytogoORGT
qjSmn4Gj4dwGSy50jdb/c8fswJYCMS3og5sFqn5tbmKUIT63ljkDCGrsgh5IHe5f
dIW4kn9V+aywrrAOeNJi6jaFA0/IdOVWwE46w82S4PI5GtbZeaarLcWZZjXbOhg2
hrBk0/zEyfXLrrDxx9GzFqo1LCUq8BFJM80BdJyXaddnSnjHuASjVe5lGLxw37c6
I3k+rnYC9ZZDDgRG3+RJZ8qkFuV4OW2RwxTWMXnlSpEacAdZgoRudBHPHHJJHFQa
kOQ5QhzEUPMyEqjLYV6cMmAg8e8WA2X4ldEeIpjSbcShg/p/fT83h2B8ZLLvuJ/r
wJo7kifHX9uEtp40fa1buyiDxB4aYuEaxct6hAxGthWJ20Z00LgVjrR+fzmBTVqj
mscdODB2tL6RmH7MZOufWXImVGKUiBG6A6C2dUqmmGzFQqhLgl+23m4UXXcvHWn7
CJuGZoPgrq/by1ZYIRw2198/O/KYqsEcEzhy+YOJ0BNCNRp4/TWfzlWz3tZM1njK
KQVNDI4IMer3AxaIblayund+moGHAE5/LCzUnjn7d55/j0RbXAPQSjl9z/SfEkms
FJp/1Qund5IHylRz84ncuXeCHJMLqSiekghd665cbLCPweWW9UBY/VElEHrLpMmV
hLZrzoTJyvHStnoWmvMPSeUkWRaSha7IN1QBxBcuNOOWHucIfRbC7uEKJeXIsClZ
1b0ihthOezxM7hDxI+JwQ5lQC+lR83mKzAItXVI+1J+vDcY+z4EJ+/kUFc8fldEm
d2IoZASdqMqEEkLYRvB+P96aB7N3JBo6dWB627DBLyYocPy+mmKwO+yBzkJVVrA0
51XmN5xSP4azQuP8do8hHPe1f29T/SgO4/fMN+aElrEPR/xiJ0a56zM5x5MfDx8n
D7bY/ddI/HkctYdCiQdAH9zl/jOFu8xLpPPXFYWtsW4GrFQFUItL+uJGNKN9Oc9P
uTYW8Tug787SCDfB6YHI5iTBlx9EhtByBEXzfPMrc/79H39CYnIn+ZawASkd5sRG
batNvat1P+A0N3n+1ESeVtRIfmoANRo7NKukdtZxZi1zQL0N4ArYGJF6Fdj1M6Jd
Sisn1upxbeaWJd9+dF7FlwxN9T8Dj6CMnnvrpyG+UUM/7xktBiRLs2q0aC4C7fGJ
Rgs+WbzcAGeK1+hNLXfmbOSIAXJwBKDwlJqEwzYzEONfxAlaLWtDqenhYXwPMsnB
2csken5VLfh6olm2qt1KrS09LcCLkG5Lrzqld8o0DKPIv6qySTtdp3S0wjSJrnwn
dh46o1MJHpmfEvjxrqcdWqRbdjlNB6Sao9hVJNuaWLZICLB4iLJDiSId29G/9cwN
1cXmfDgiqBiq5JHDBsG+sDLWHTTJHDpZQAM2SUxokN+3T8cyU/GYcK0bM19PG3yQ
uM5Zge+Z2h6ZxaDfKufQ3MmFdxjw2rCK5n13NT2An6sGUH7JCyrLREQEsLXDYs+n
vruvdFJmy/M74aGwy1/5dO0P+LrvUM02gf6PNSzmKf0EfAShOJYs+WBZ6NyVz1KH
eLQ3Mt9uT2SIFAxXj2NXB5UA7UADxqyfTCCuNskEChWSPh3HuRF7KALfQvfQN9zI
1AVJFdJYnmF0U21SxbRrf2Diyq5OQpg5j+frr0yloB0Hf807I+uKw/VE8dvdYJG6
O3uM4958Ec+2JPgO7LHJcp3wTKR1x6K9liDYAFlvhByjw1fdSg3q50GqWuzgys+T
NHK5QYo79H+dAtXIxvoxO4acT6Q3qasZlaFOGgkzJyA+IjevCfSQXMv/sPovfvZ8
72FuWHoLHpHxTpkDt0YTAOODEZNwsk/ok6fOU3ty4TWfbmiPjLY+3hCCIunaJ+5Z
ei6hfR47gJvhUQPkSGFJj8MEt19sir89A9nhHKVEJObtp/3MqeSUTdn/n1Uuyz0S
y3NagU9+cLxwUSrd6Tplhk0BP6Te+ukzmeHER9khmcGvV/sHMkEq4VIwwI++I961
60tqy55cT0a+WHkZSaCRq4KDP8R+aynB6tnpEcVRbBo2P8SklzWOLbvY5J+V79vw
`pragma protect end_protected
