// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:36:47 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
JnR3lisf83CtZjxUPHPI/imr2U8L7bkEGT5/OsENMOhZT6VZO5Prf4OzzsBJhVhP
TPKObYwA9T0VPUgVeuanc6q14aFxpganjrih29Tho9jstAdTvAa9x8f7RF5DFk6i
VQhD3+sAXgj1FYGpYRnpBlYahRicdAsoV0vAOeDMf2k=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 4416)
/NDUpQ0WFITeCUUhJ/jpL1YxVuc+WvrBuhT3hepuLWgry/m+PHuoCR6kVPgFmxYV
hs8RsqK43pbJ00Y6FXEH1F5gUJQ+5LoBhUZ8tCFGxEtwtAA0krw03DBFaJt0SYxs
A8/++n77UNn2OiDErgjTT327h2CX8JCuYN0K8/49B6xrmnmE9yYoE2tujxWyTHw3
/en0MlAIjb43swTyX0UlsRn33o5IvRcFVJwxxHSiNAx78PPAE3BPR1PoT3OIZsDx
UPfXq7M4Kfmj8QcELnPQz1ILAQ1QpWuY1RQuPbETZY6NjRd7xwDhaYETA44o6h4B
C6w2KTfv63R1MqVxvirAH+8FBdZ/De5WoYYuuPsJg7oTzs4gy5SwyX9HAEnvGlD7
Sa4FBGjP8dwWXAXVqCyhiaj+suMBTwoUTLARP4Og9E2KLVlWuafkuSyjhowH6Uhi
zfoY3Gas3VyfOK6pq44vodpEJkzYOuxtqEOVq/FkTDmlQzIxPiT71S5z1sm9s0Og
oXgi+54mmC+BJDDdfSrE2nqfUaDfqC/nlc5r19SM3Xn2xUHfghkUi0KKdkVrJNyH
urV7juHE93RIAXxGRBINxKkfw6pqC9Yn8UIUv8qGqNqQm947ZqcapgcrA2515SdW
OO2r4q0WF+lswOkkAQJMF2ndvn4FjloGB+2Q0JQJQNMxPmk2zpoT8aqhgDODmdgy
eZg7RgCUOiwLCJZrhs8FoTjhfQ2Jz6erCLWvIpV3fTengVfwsHiPRvgDBHjkyqkl
FcF1Va6OCq3xia3wKAkcYpR8YxLbKK8c4p3Ziw4/xa+Gxul3Vko1X2Xlc7oh5oZB
yYDFpgFC5OFOuohu9YAe1kieh8hHDrV9BrQ9ghaHuWU2DeiXliWL81NId0AUyddl
OFWGT3O7oMbcvRtQx12FweUTeyxbhdVrJNai+29HcEp22SUhOMV80cj0PhoElCZm
U7DZ+8VPp3lMVSWCtpY3hJ9aUS3EY2eexw2FmQJmd8675GnH2Pkacp6rGu2INnrv
hX3wviFbafuxdbDTDib9eHLyBMoq4hAyxlp83vf6Z2yeeqE3jioLAIm/oZvsQd+O
FheaQak1yren+0Ht0oaftBPLWvMM7/ywAuMVqvUCJ9EXxjiwhL3eFG2a+rawVvmQ
0OQ/JSwDfZsKczBDUqSZRouyZvZXJBoURjjVio8+qH3w74TnmVsYVcRyKMqBkaok
31pGf1olxZIZs5SEfXc2pQiLDn26ts6wtyDiASE0MvyzTHGhxjghupQEcT5xIvvr
BqdL+ndIQMhaJOMJt5cPj1F3dlBg/Qe3DB7zj/cjfiuEH5D7ow5n6LMFDX/6UWH9
LGKTgE63o8aUozu5WJlWb9N7UzNv1v/ApRBSBBW2PMiW/gBg+WjccYFvSTKFjFYC
MfOHD5bmiklSieR7Aj3qHYLXr4kJkVjf8KmDbtTgxLCBihR3Y1/3QO8KUjVYh9dH
sJoelKzWTmoNm4iG7scakJbwIG14PeeZiEbv+9f0tmsh7gxFFxkS8TDShh0PlnVz
x+TQMlmIF+qX3XXtns9ebixju5rVAysbhOUWCO6PAywwpGFJAaVEu9bTTsBEk/Sd
gc/XrvBxS5loS03vzvOBTtVk3htA+XZi/GRxBBR3AbY0Nhxcg0JOm8aXtPraSrib
h/lPkrcvCPOT/WU5L1Hba5TkrgdBUTJ7S8F9+12QOg3rpM5wtmUt3H/790hOJB7K
v9qRHdhkKnJRsFYTUF+z42hUnmBeHhMAzivjtqkY6d5OUiulrKn43ISmohkNxeYv
viZ98fggDEFHSWQusQZ2wzQ7jAXyCT3l2VYYyurChCkzQs5ulqJRhFDWmyXaCNaQ
+phywm3NfxEAE/fVRMJRd9pykRokZ8vI0da2bICARg+aQxOiTE0LidxDh0x4P/B8
hHWsyzE/e+xyURtEXh6LiupA61SgSf2vaE5yvSH49RgOjRo7QQwBcBTcmfPJpwbL
XeiywCTe29F5Ny9VMV2JFx4wHct75BzPXn8gmcJf2x9IlMdi/3EJ/2sNXDHrjqQ6
SoV86PX9yNUXrNm/of2Q7wfvBFnr1BBHIm+DOotkBp1eDLNVyNElmNlM3sSvCVR4
m74yohY1mQEzfbpmdRiuKSUP4CZ67WRAtPm76fpsGGPk3zh+9QFgcSYZSdadBRT4
BLNhwPtmh+y2ZjS5BwPCox/RnXj/d6C9QjxEUTUcIF/lVSGOLbEsT5IoSi9GZp4N
W4LVZaQx7opkMDsnGtzR+a7HtyEWaxqMiEJ0h0te6QKIAUACawj4ZKbQwhP25gaw
SSxeBdyE+D6gPQ/E8QUrAXzdc0n2xnXT0pzWF64fxrXRmJfUG9Fk3jMldV5Qmqr1
2Om3xkhcrFdXfs+NQ0hbIzIenScEZU9/+0m0XOWDzCsBDWgZD2hqyzG0YK8KDog2
3pi8XfldDqTQs7+bvPOWAxDm71cylHyRH6qe7A+vKhlcr3T2KNHkVRuwSWDfBgv9
ljajMJ6b+eR4Gnhf2Ln1FP7CRoJ5TOhXnekRLGeEWgtOhnAnCOBXDcLrGpxWxCYy
WV51TJlTM630j5Wg6fFlVTUaWwLKotIk5aBz5OY5UZFQMx9CLxLgJuC1awR0emTq
48i9ltT7ZpqVaZBydk3QNs//u57Slo3RPMtewQhkRdFcbbxgKDVIwmUNkbHr2pmr
73HL/lWI5ctkLdxIupEba9fKTSFej57zI5lwyZqCKZfdgaNEolur0lbzsIzScF/S
w3JkWCnVV4nN859gSJgQiz8oZtbp4y/UCJgqzh3Tv0eyE0xIjriTORC6NFTX5BDA
5HtOr7Ezmpx+ZjQko+x381N7Wu2ZAoHvoIlJSsT2goZr6/kAGnxJKjb4+fGCZvEK
velpWjtSjT9hfiBt6tfqshEpj/UsF23ix3ZskKqdPy+moPT2i03XuPuQwFX0NRB5
1ILdJMH7jNPTBrco9XQ3WlPMRcTpopfS7tJklekj+lcg/3X6G6PYSsfsYwF9ij79
KJQQU4VUWubTMwISboXjbyEu9oq1ARvOgtt2tgM/cuvwWeARkh0aAREXJvPaCISH
pq7KaiFaw/frCwVCdmsvCt4beLHJ0SkQq1tLjiLJtHdrVwbOT7bHJqF35QY8ySYc
JJhL4yIT09ze0mOfheTxJBRhwu1Cuw2wCu7CQxRwrqyUj+Xn0gVNa/5r/SPUN7y+
OXrqXXYnPAftAeSVU0eqSxEKeH+TIo0k+tmUsBpUun3dYtMRhHKH0rLqp2P3K1g/
WbgDcuWWp+f9a3N2MiMIllEXBMHjG+miWcrfAx2iFTa04EE3IArbeRJAtrzyzr6U
aFt+kxsKO6sqsiy6MisSXEsFQDepaPpLTNT+jJXiiIfx69H8uUzH4nWPVhGEVKz9
zqds9mbmvEC7lnbY2FQvPtnNGbFHqHIHSsxDYhpqRd7ZBABzyBCsjTXL2auMRmcJ
EpQRi55FGpy02m7vp3AcFoXkhRT85HAGwzixkfZPCc9Ep+CJ/Wh5vhhuSlk2rDuG
J7xlmStuvfmq867Yg68yXYy2DTsOvMbwTa6dyINz48V7LYKJDZIaRJ2NLeptNgje
aNpq9fGIt3HRJwx5TWGTvP7xXZnOKuJOUMUm0wsTtG4dJc8nklqPH5VNzAb0agOx
xQGufv1xSpuaesQSNiU62daHyluKTq7OFov+89lkY/7egscGaAre0qigz9xCt/Ta
+Qwl+kEqjrxNoRp39reUshZ3XhAUO3uEbkp0qtOHZ9P74+yMHbqbItytIdIy6Cu5
0qlQp71VsSJwUUYBM41b2LMq//yVxiuz6S228znpRDE1p35LpI+bAdTZLzoW/cBD
x674MRsTLfPgsW4429Pj7eXF28UefPGRYqXae6e0NFCWmfcK65MVikI6EDUshIDH
MezZQaXzWKpRdpnhWeIL6x5HQH7v2TtqMCID6vdr9n57ChUzxSgaN+ksn3Yac1U6
IuiAMNNbWWERi6mm5MPtgBGctBN5EvjT27ZXn85Cw9JUd/bSGiA+mDidSmAaZDv0
k3H7IMYU/FjBtzXG3jWt9pt8d5EL/U0ffcHjiHQCA1QHiw0xMOXILQuCcDI/Ahlh
NFT05Fa2wqGmXuAonsjeIOaDMOcB9o0BBW14iFBzizKcojVAH1tB0GCoTB7Zp+Ls
8U5jJ67/3R2FcjyLU5Ss+SVwf3F2U3Hgy0FXp3UthANP1lHBaKcrYjvT/+uLzsWC
ip0Zl0uN+zfl4JVTZLPTJ6RxRR7QiCpKEaTJVwHuujDdNoKkKIZmdNT7kjBe1YC+
K4dwWOt9Y32Y/O6YRBZ+OQj0PoJcH6e1xAgtXEtwsMuAnny7wfRUDITodaxmJHVP
IJEmgtA3rrUZHNG8bJy6PeRNBMHkDW//mfc9twVJLY4TWA3Kx8cckJ3SwOAM8IIC
0GDoDAzEG1WYfDP4mTFtnKij9iXo/YVzyeGWfZRLT/sbP6gtdV6RAj/W8BPM7YGF
zZRZrM0C++rMJaMzVIIFq/ZdDnYXymhcVVBJHuU+pxbLO2RA2d7v0LaYGtWuZfO+
ecfvIw3cERg3w171zpDVsR/d9cmGk62OYxhB3oQTQKF+mRjRZXiXONXTmJA6wVhr
Fcx7oOIZmUdSV1dWXuZ5HrDV3vfT1VaGczcZwJTDHg79TDKXkOVGtxoRZf6c5op5
NzBc6euXODmTdUxtmd6zAMSVx0sso47WzqdAN00PhoV2tjMrY2R5ayx56PbVwqFx
0Npz6y4BnBG9+vc6eDj/LNgxnmsBfmPeo+Jz3sT/py8jHCQgiC0ekFdYPs2LhMWs
HSyI+uxgOKNMfXITGT8WC2adnFB/ZXjay0BxdOVG6NPrG0u4D6rhhF1fQz4lRQEJ
92RTPFG+cQRHxsulTFxfhuZM567MeXD+EWFiD5NalR7eaHq0pWp4OkuPS63rTa8z
JyKWJCz8zOVlrVd8qIpUShDB2tFPWYiKtVu/XfFwWqoUQyn7o6uMMUP/lHRrHrz7
xFbxEVhhdRTxJfEPI9Vuq5Oa1Jn8jSpwwST49fn2urH144WPJrkND0VUKoPaObGx
Fc0GL/vi9wOgksZlUu8pEO2unrbXTuVQqTRh0NRANOWWBF9+y19UUDCK0WpvDh4U
ehKr97vM7R6Yw8aEL0BXGZtfvxgk31GEAWcBTH4DvOXH9Nqe/hKPvT1hyV56/vks
N+cvh6LLpG7QzrOWZsnD6PgheLnEhBrh7ZQ1zreq6pYiz+kz/1OOqostCFWlK8SW
iSSzoes/aRnZKVTxWRYO/ycP/eJXT3VhElcM+4zEKLUreDWYTajF5KyvGJkVrWxs
j0eQrDh7xnTtAAMBSibhm5eto7pRxwbOsGTIo17X5vU+1Usw16wZi0VNfLQ6HSIT
mUcF9J18yTWEdYlBc0VrWnp3PyD3H2am48rBRVYBI9VXxjYz+BFzRO2iTYqtyUl+
/k8vtaaHtvXaWU5xnLGKTc4SC5ew/booJhTBkmsa19c+lMkxS8A2dJwf/T1e9dVI
M7/7q5qzwRZ1wfSHyKqG5VmMkPnlOwPOjudP+5JZqACMgEyCUVMaXggq0mk6SsHk
HxATyOpgz+5k/2Gkxbt8aB4yemDM7F+HhwjApA7U+0epUF38JmrSKRPACa3bg4pY
nPpPjQW9GG9NdGf68U5QJBvUeqkpi5zgS1QpDOrI2fbH9qjiCruTwQOIJxf/tDrM
5FVRzMRW9QjV7fA5++i9TCt5/24g7FknvfnEWwdOv/M/5D4YB7bjrY4G6UK8+WTz
WAp1BfsPOxkluKldtrr3a1m2hkHEvimyJhJUpBs3QNI9zs2xhiAPMrY1NgIswhv4
roHaPvEmpcqCs4LVk1o1cW7sMF0B9myr0eLzH2W4i5OIOn2pigKfxo3JgL/PJmbD
`pragma protect end_protected
