// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:32:38 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ChCLlqyXiiZ+26AegvhaXsY9ux0Lr7yP+X7aETyH1jZGMxNITdmrTnJZmwINqtiT
2gKGPGODLpzp7AvlkEXsFHN2QJ994Dm38TlZev2iYKqE6VU2vD7QorJqMkPj/AqW
bapAgLdvNmhDNH1Jamv5cN2uRENlz5gyA5nazvju8O0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 22080)
wfYs5BiYAh0NCcV9hZmIuY1QcuyBqKSlxtX3Fj0MrWf/sypbgzd+HRsuSjOQsIBU
qcRr06NWfH10WTvT9QfuAvSUhSxBEYpClYeIQywGlozLeBUfU22c1WzsVmQA9L2S
D1P0vwaLNcqgnIBmlw/c0PWPsPoTDfj2jBRcic4MXBihTWjwJF9IMOdr80r4u1Vf
8SfI5TyzXcVm1w/3fivSORHLMrnL36MgCywgJWrGC2Ph/qXQjntsW+zRsYVt1XTT
Iu0aaXe/+AekGbjWoyeJg698rgAo7540JqGmJIxVJF4Y3gMt5frJPW4V/vPzUQp4
vMnCExLY582/uOx0XUsg4/giaLBZVAviiB5DN12C+P2awviHJxPj1zSLO6G0MjTs
f57HaZPP6MO3Vlb/RaduWZsvGrUPIAW5UyML47YCM4Qgs1h/i/faCHvb83embzHD
Vg5YRj4+wSxh1KgmIJJ9KudRot1Z3boeGk6I6AzEga9fmn/RvN5IbrrBhzQ7A1Ky
7HDIPTLLEXC5yMHqjtDeDSc4q/ZYHIePDJd8KdfJsUB9DoeT2l+GpXEBi3zETuC5
mkssIQ4WnW8j3GUL6H122AReb+KexiT4In5kvKqyzbje7rcu5728X3Yja3DUxWqX
hzTx1rHJJEkMmxIbchciKTdv35lvKUet+R7dznlahRomECfE1CqwANM/NdXca9du
12QKYv9tMVAeG8Y793qEusBTZ/+9ZYt56oEC9MYSEsDW9J3j76ElK/EHcGOCivj4
mdNcRbyG1TWHUzVYDzxIAbMB7jMsUfYbodP7alznY/2dz+1Oy9jFkMl2xoRPbsTj
ZxLBsttyqV0VUuiNG1meNUxNE3fYSNSU/mvqxqSyfSp16ZklaJ3Ipm2gzFX482lh
6wB1duuM126z4YD2hz/Gy5jU8UXaoSZeYIgEOIvoIutQeQ4ucY28GmM5V76FyuCT
G1VQ39NKaPA40cBHbpgb2Ve4pOj6+HyqiNDI58L+KccwwDJhN2OD+uAivj2NDkfJ
jBJyDRAeuGOfnWqp8ECnoDKieXCMo31LliCFmTrTtPVXEVWV9mCo9ECq/tkDFcxM
s+1TCWzXbp5eArMrQQwhuR86i5HFQZTk7K9w1fbZ4tLMqUO01Ub3QI92GegDgKeI
kSj94IDdqXnuhTLp9yWGD3ZhJLczPAazqfnD32nruX2POElH0ekq6QHWnLGIla65
tWQarYWypk9MDU4vyMEe7QaOxr/LpovtEm6m3aX318X6aP6Pjw00UAa/dtZPLUin
HT3d2rIWrHeufcpp31UwOWq+JYAFtLu7G7FFiQDQ1andPQa/n5jzupVfp74eB0Ws
++IBSiAQe+FzIo+1ZTlc82nW+nEuPZ8BJ7SOeGahDAYTsip0YcbnyPnrAU+y3fmu
7P/rUhe16xPhJnPjEHvtn1o6hnSl3TA8dByFP4WFX05hu7oeaPDnr4t6Y43dn7gG
h/UgaI/CBSmDDlILd7z4IpfXdxL1C+EpS23U26LiLYK72gD4RwxREtp8GoGQb+kB
Z55lxktTW4OhEu0bGxctl25bSyzJ+RSrYN2qDe8K4Swh8W+ay2BKHKqBxtRnR1Ig
CwkbvZOWXSvLldWv2vxB8JyBUSYtKZQw7QZ1j/8FbjgMzCsU+/WNFfEo1CMJTfvB
GHOW0QvNZA7bsbJgZVmBhK24+pqigGJ30s/vON+0CCgguyHQvG4xop0PXX5xmOpR
BN0E75B+05z/CEujS1b2TZNrtXdi/YyVNdiYGPcSJCxPUsNx09WP1Rc2TAPCKFbS
eurt7G+jMG7hUKV7UQ2DdgGXBvxAnEc4dyRx3IcJcLiTjAqs2efnwzctdmQFWH77
QHgdCMEDcLf7jZl71z1PfrlDdOx8fxjRcGXpc7mRpEWWBfx8vk//imxv7CPlY0VO
vKsedr8u8Mugvk4uHoCqVzly6umnkTFA0eKeg0KlikDa6iGhENYgtIUBmg15/wLW
9/zYjtKllIpU3Vil0q1n88i32bm3XufSB9Ry/tQ5a4fbC8LAbYNxB7YjDXOMe2f8
KA75q2fWTV1ApkyxXGbkfX4N9v2uwdB+uHU+MEWWIMO0y6i/W9gT3ndG/SoIItNX
p43Wk1bgPzvc9MgYk/50aV3eBHy4/bPbmy+4HueNYNaKc++kBaFmAEtU03uhsykG
Ewkfu9gUXzuWIdZV/3XMO/+4CauhsTXRGK+tceX/HP2Qw4tshID+Q0gcH66dnQxm
M2MK0NLHeDRpyexLykIcz+Z+rvfVpo5wV5bA7NgvH2TT0QsW7cRHH2quL/F3RddQ
yQRvUkGUlP2EFvyrl6hnqTUYYttJHH+qiCB+Pfof23pduOso7M4xObkui79R4Zr1
iHc8pUawQ4UbXHDKodXP/f6XD6A3AF/hJYDIqfYghjC7dU7j1vCbsGqKfmzeFl9g
5w2XI31yWPmj0bz6kSJDfYjonb02lfEa7hnbeHkTWfsYsx7XCayj0S1AasrtA+bw
2P0qN9UjuZIJUFz0RWpovkALJsdLQTUnDJGqsbxyfGGPEZuG1aDiWYeGW1ealhSu
vE6+e8Fk2hQnVLzlqbgIlXP2zXO2XfTLjAZYFyp2gEQtxsclCr3pzZlkeKK6Iicw
DQYr1uQBoJu+3vt3yuHUhSocIOEI8dw3WIW1uS+c1FPt5MTDLHR4sKojUn2103Ih
9G3qhNubU0/30SZENmVoe6nBofSLDiLwmQAJiY0DTdRchf7FG+MqBNoHScWUYS9d
yIZjbrmvb8zyoolZPjckeu5RITDBUaCnLDscplvlTnXTaD5kFm1csxgVMAF3NlU8
DY92VQpN3q5hxq/eZx0R3XONI/rBTiIt9ciil03emjSJ8fPyTVKP1JeyIIJkKZGQ
ZeEcT6IEmQyFtUuU2exwJaqSfWX3UuZEPVQ6hCNZgWBzM1fGpwvUdSgrjupcHexv
dWPJmsJdA8KouYcQuE+vuOnJHlwbRjV4RabLzUtpD/P0mU+j/tcJYWC7B2FpTdki
DJFMVBEco9I6HXlCQ17g9pdWlWNsdOu+2u1l+7XOvCh0dKT0IP+F/oYbhcK8AeBj
O5A7Xa8ndVm8+SBw0gAfmiHO14aEcT79TncjkWkJaR+boQDwiozPiz/mCoPQTChQ
gHVkIzwZrnOI/kHlE2OHr0bCeQQkgZSEQwL+rXyIsfDB4C5kM8djlSuXb8dgQZvC
eQn/JWMwWfTs/6LAd1GLOAjhtnvmM3BmJ+TPCa4F2tHBtw1pIGOQHY7uUBfCuXO+
dkR5JKxL1fqGi4KgT7PPD3imSekOZ7PZVlgmtxdTPmPvmj4y35vR5dudAmidef3+
Bc7XLG++5IggyCQrOqXe4OB9Z/wD93Z01nENn5nFfpt4ReAxFTRj6E6uIff9TvzA
ih+khkvrk/s+l3ehHklJk0f9W7HIxp0YC67AiwtNgVmm4dorHKsR/vpf9s3bgpGI
eu3gM/3k0oHJjp8XqkBXLT0zeovMkTPwRLh7qlzSbRv7IxVfhyv1nKyy8HwCbFkt
WyiBa2B9JuF+1UIY59JTv0Kvlf7XQ4XYBhBt8AA2iU30IAb05rEgtwJuuqOkepAs
YDRo5rzQ06AjYGPg5PfAVDgHE49p6KFl+P99sxa1tgRM4diT2in9+d9VBAEXWhP4
lMdsrLCuygWaWPUN2vYqbIQNeglyqGBTmMXBEZBsDcO/f0tfWj5bUVLFBF5l4kXt
5Gl2KoXJpqg//jCtJgQlu1Od0EHyU2U2Arx3CLbLpCtHts6swE0hwqAUe6S8vwH8
VzsEMXVQl7u3nNdC5nH3dturviTUnCWmO2Q6N4nBYE/anu5S+agjsbMK9d6b9PEi
9VzZNfX0DNGNrq3lq0K7LRKl209gFEfuxQO+nyLAwSVpOyv5kHKMxjh2tX8B1RPS
/2ZgOzdIbX6FBRJrkOp+FHkJkTSB81IkNeJu+W9Ua1vNGIwNk06mjbIQKmEt53sA
6Xax/oG87qGcB2dl8eGv6OsPy6khMUl5YmM1ckpdK+iD+t7NnmxVl22Oh2DIpWv/
UzfvCuHcwaVlEBY6IXLDC8KjPdH/Zfg8aa/j9tVmPxuYP+3DL0nDfyDTb90LiPNW
zAO5CClQCMLTowYnsa2j89LpdZPsyklyXJ88Ya+BkayXSBmOygWMs2lVjbwjqhri
dexPsmgluLRVL8H67elb+J0bi7C2gO4/IVQH7v5uM8BGumrYxqqKcd7Oo7x7dsYW
kiXpNqpSJ1+7tYa3jaMurk1M6jMkoovbvblgD8iG78o1PTDqiThTurdcqf+X3sJ+
YvFcBBZLEKGFZB+Jd1OANaJEx8jbRxPxiEXtw2npnXXC3u5hy9pBMQMqaqWr2D3W
cS8pkSSR09Y94eHRx1VDpaP0Cb104Z2cqtnugM00iT6fajCg+CHw40pS04pnGuM7
kdooj5X0Cb1pZjeFC+tgFeQD3A4Azl2v18mIVXfIadnUWCzaTlCVEJnQ7p88LnzB
uyXvkW/AOnrq9RvkWOki3L6W2SVd3Cim8DZZNFY4jigjwUNQ3IT59I8eybhtEUsB
c6aaIReQL53brlF6iFrwhpgfTrbtUrcsISZUeCiiVF96WeCXkyPZcytHCOOAr6uH
M4nvts0ya1KJV5b5yWfyM5rUkO7RQjluvFgXM/RCAsaKdDBm7i1/NnqwnFkvKBNQ
931KR/tmpbZFY+4HHXIt3V6Vz4yNDQ0ptJ87tOEno31qs1n5IhCmt4LIOvuEHML6
SZYPTZ7Oe67PAvuwJUPBvXeK5gOLY+juU2D+9QLqytwqtE6FRog3smth6dbggFRB
nZJQfo16vYN99JpvCnlji1o4lPPRjVktb0CWTR/Wz2E92NpKRqPtj3mF5LPr60+9
Z2IiUxMarQ0UxuAd6jhh8IercDBocgrPUSGHdlF4LSKP8NM3y0+jB4keDuQGiwu2
CFhIlhXm8Clx+smQuRHalcgFwrSi0gtvI3DRXfC8fWrj/tw//IcZwbfGno0o/O6C
p+YCf8p1yPesiK8rd1II1ZufhQG6nQn7hsZUROiFuKDFSMcykN61iGlWBzpfPxA4
1olgoilUAp3aKFn6RBeojArCClq62BoMFMaBK+Mfx9oH647WbUocSnCZf2QEvaSX
ZT2C/8UxCtYYoDzj5ZUwEt1HfcWyOxcoRloL6l1edITNvtwfhIp1Y1lDJU72YKIM
JLIVFdchw2fZjpmn8QQ0FBLhilnnJpkBXH+0HWxxbVrtRNiyzR0xmuheohPbhPaA
n1cA8RGWYmsrFiaNh50bxu3Nhx2Q0tov9c8pgca4SSNe/7ggs/AOYmpf9/GF04em
aNNgCnKKQ9l2rZO7fFYC+X+H3+dvTgOoT+flDxzpTq6klIO+9IJc6xsVOWJkkz7L
QjOWOoYhJKpVDAsil/imD3mL6wTMjQIKA3FEUNP4wVFXztqHxFsped/POzPOgAvO
eZ8bwARSr+NMLvycDmvfPh6ZQJ+b8fj9onKzcS/RCpPV4FX2eyp+dnn9bFmEhdtJ
NJFFeu+kSXAiB9rYjcLzSn3hnm8M83lssxrk8Y8WPOSOiIJRHk38BkORe+gcUQNe
MJRAR/ZKdExht2A1VFQ5hl/B5MZQH90FAokfl3apC7Q8QU+vNi5CYKhlZ8ILB1r8
jAA9gL+dPvGmCOzs0JIChAUdCB++OdRs08M1olyrLoua2widTeoLjiVE7icT2eez
I+gEfXwWBES8iZ4Q3CFpRKAtvX7xmK0DnDcTJwMX/dOZyTIu+L6IV9kocjjTFHZv
nlwcNl3skVJx0Q/XwOKIsQkOZ3b6rc4SVCwhydBk2JqiFDqap4/7Np4ON7ue9FuU
ghn+OXWJmPHWkN+g3UQQ7Qrcc+gvXCrLofS6opSGZBFkmWEmVm4xLkPg1s+XHx9B
EVopitI0V83JEIn56pmlk7oGT2YFUEHHeMHrbDCluu7NNiY++kH7etUvNlseh6hT
4SEN0V6+Lo81GrBkPmFGskHOdINvydrvMOBnkxnQofWiyf6U/BJPujROvCM1+OJE
qP3sNcjH2XelhB/9U2Va8yNgdmRXgSb2YmcYSW7kPwG5PrkvZMNMAhu+nzVDfS+j
ph6k7sXooNFEscMrYZavkuFgvtqLsDajpyqUz9EcKSTR5dIf7HDMDmYbPrapSCLN
CzIkL4eSQcGhO2q/MvjLR27tKSYEy0PU8u16cRQMbOCIAqyX1xlq0qzC1fa7JBcn
moGvcrJtORTo8lskbiZeqx8ybwekFte8nrc2sqgns66vD9e2yF/4E3YZUesLAYyw
We1NfWjv+xq4QXrbBQMuU89YCZ3TtmzwqlRPUr6lYGvbo1wtJlDr6RIqQFPTpFaz
5O9merOeU5fSI9sb9DnoQHlCuOx6uZKkdC3S3TkX5L444YcFRVUC56w4raTT5s9+
FvCv3c61w4SFwXuUeILgZt5ewXSHSrdlx9Igimfmpwde4rEISrbEwRW12YUzokWm
LXUBSiOSVQdIHqQOGapIexKSw8YTaElET2TAfgNcZfAFLGdDBmnFytKEz5aE2+zY
eHNh3oiEMiF6jTFCQCCPC2gOI+KdYvtSMLlbuZvIm5Qzqf4bwJFkPnBACOX9MWPA
rknW05ScXBGvV7UdOpWGrC2lSsL4NVImJK0s7Xl6Kdao/iBF2573qIGLo15eZtn0
H2gFK1qOEpM0wHSJpTfC5l7CuMYngVkxSlNCSCooV9snoFxYiBdT84St0x/Ug09w
GUXvE+hZV1/HRjDFmPg+LajIzO5s2InM/SY8RHmqZm3zKxBv0UCRRl4tmgkgb6B7
xn/rXG66EmLGZ+E8AnUnJ30vCzG3uXAG/JTOmKSk/c7k5CPVY/I5mnReFFpdiAOY
+KHMBcDumhtbo5k5/OzUTsoZPdnofl3I3sFzteGbCNee3xph2WHWw7sBJnGXkdbm
hffzLyc+Snn39JIbqH4mq6uwv24UyvqaDH1SFmh+tXfPBK0WaogS/110oC+cPJ6E
P27XsR/s9aL57AzDkp7amoQw0vm0ucmGEJLSxk18WVCejHofncLEtxr9O9YsNJfd
tWDXM0EGabJwi00yfmqYRlrt5bcU0w7HfOeZjDc14EkLYBSAJpUQmMOd8uHG2xpJ
uqmrYiWtSZSCxlxq45L/xV0JZWNq1mtdP0j5WayFhN107cT+oBllq8xNBP3F/IKC
jjLi9bWHziWigb1Zrje3QxF6zIz92VFRsebXZ2kmpILURo3fCjNv5SHi3kRyBBjo
KW1W82j23rFUNamcHJhWKPi5aOF1U4lXvdIBMmPXT3QAm4lK1Xaf7W3i6oalQFHh
27H15mckxR8HeTD8nfyoxtYDyrmPeyZe7u2bABbUHRQhSAsDTb5+FFlxxRpOQhA4
Guz8xj7r1EL1OQ+5BgTcF/gJnVahHNOSpzu1NrnkhekeG9A6AVHNBuA3T2XXeN9U
XGOrSBc4e002XMn67pg5LxKu/M+raU5UXTFPv+ozL8HS7CISpdxBtJyHNgN0mra9
q8+oTIi3WEc6k7u9htg4D0Fd1sLzj5O9weWvVaijEc7SVwHbq6KHbZiAJWH9t1WL
QHuUpm0Jq2D8tjubJGLBFl8yIGzo6W8hBx8CLQciUCAQVzF1Yt87ng4DAToIGD0V
o1SQbh8ZHbEQ+u02wT7dRKC7w2cTtS/gr6tl/X4T2hu31OSAn7t5j2Us8MlCecw7
rODLFjcYD4ZKID2tw+aGaIojuGD1Fh8Jhxlwu03bc1l/dNh2UIonfmJ3GqaGqzU6
1jDYYMsdrBDAEy37pbt7+ZkYEbyn7ulzFWzmpPUBKyM0tcCFjpoICkLFMdCJAnnM
5mb28uChWl/99X4BNhebYQcFLqnr3zi2f3xZgrwMzdeR7TKxXcTacnD+TlNmk1QB
zIKDuYo/XiqY0BAMs7f3CveLExaL14N8MeyG7HiXNBwhHgcaDtpXlSKKi96EBD3o
mNjxY5fvPqJIk3R6Ayl4wzziG4lchL/Kb24KslYPWa3mkgbCuwc7HpE0qyFykEkE
8EgzUNtIwiVNDiL6YsWkLk+NxVNBZZhx4Z23kYjfMfg4oNKdxv5r8/UmrjXzTsq0
E6AMfhSkWmH/BRQr5ZDBOiUGmquMaNsfBmZuHNGjUE8MD8yltc2TXhuUV31dVhZN
MWWJqyhaxznxWDKjI/4N28JETDqvcbO5UOxWpj3uHISkEK9n5Kw/G9vm8d4JBb4U
ntMOPj2CGZhTt73T4JHyVg7XTiaxz32+fvqmRzBIzp62+iKuMzpPKQyMaSO+PXaK
9VqHCVt5XQEaHb3Jzv1SwmAlKCktc7ga1Fd3KZfHJznWqB1B+tXiWa7vefsz2dK4
Mt5qP7HO4LnDyhDNhPWvAeFnNfdOCLkOV4LhsOL1/7s1d1kxxrlsdJ9Y44YOphLO
J6tWt2hBBbpAjGFLjq+zgS4QS8NfgaRrbxYcIXmpahNPUjbhrN3fPrZlLSmFdYR6
tw0cr+A+sQKeJRQpp3iDkiJm47f2PB/b841a4KzFB8ZX4BZqjNB/dnoZ4Bb8HN5Q
Le/HFcL+n9Fn5RavnxwC+iiPavpOYwvw/INIW/NnXi1pdedwEFEBsboQx4Sdoees
p414IFw6+EbSFi4LLcF/000zPrHJAKjFzSeuvWiRaqxMDD8O9MNZvGR6Yp1G3tWt
98Ks3bofXrFE/+Ev4zSjF8RcI/hCpGR0J1+fKI/MdQKVFqWcqMapBOjj7DRl/JXT
/Vax35PJiuzN+EW+y0kbumKB78nAVe1vk56/UlruGNct7nu927BlTHqBmr1TomFd
piYLuM8uvxSeWPFgS+lTa7vJLars1EXSxWcDq78DL/FlaocUBvddPfHqdPwK4vWN
wWMGvY6lfFHLR2DRjtFB1smFqpXLt5HZky1/U/gkzFEr5vPlQ8xggzeSIlzNmBkb
o7vLbnR2daJTrZhpLWGkYADGEcQunPaN++LlAZfrI4A2erPpSHskJE1w9Cb8my37
6Ifte3z6zWktMt+1pkVwdc2ITD5OKWNtCTJd6Z/nYdmdjPMnJouQw8TcmsFq2jD4
XiWUWQ6Dg7lTs3qU8Ya24wY6rnnV3xbKM5ZGHsEqW9frOe8T9ovA5wqRcTIe9Q24
XJt7BwXILpf1lWFkILtd9xONE9vHSuGsmcqonrr6JtMYUZiMEDwyXCeLsgf2FDAA
mKI1ZrOGHTb4Ibt40oLTkwwhKsrbN1t2OFIXr7K9+lpC4DqGMAzS/OI1e95iLkFE
guFZhIOIpFCGknaR9rU7LodntH3rTfNHdPne7SjipExlMeUy4xIgOgjoNvuwhadT
jIcNIId6b5WRZEtBc/lE2sUEG+oenIXOEvnTt0eGxPlYn5cnU6pLXdQHSOqfu7zI
TfaeaP/QI5WPVbalYeahK2akHPoEtKghxmJUtceug5rICUNfZrKbQKPmHmi7jj54
ayS/o/jX02xetzARlbGkqnlkhpY1syP8c66JjAkya1GagrQqu//oSXWi3EzlmV+v
9ezDYyqJx31yPb+8uQdxsZ1zGIywf3dOMqYKirwRq7Pe5haQNWFfOkKugIJI0Z/O
1tMXRs8l1F3CHM7S4P6M2FAyVvgHb6iEsPdLj2Ubd6MaOFAXj5OSfb5hXZrZOd/C
ldT2rnVAWqazMRIulEYYDbRD10jlFzsiOwHHj5aaO8FdeNuulh51Uv8Z9bY8z43Y
Is50zSIjwRpEldSy2l/ce43E2cjO8x1pcTLrtn/eHdoE4CySd/wl2ZIeBU+al5d5
AIi2OXwKd+ALXFXwDKq0VLGIW6kxalI1EwJksvHbJ6ErT0WP18szrxgTUXGZHAHx
POCUx88wdh+FutLVe3hIncP4z6+ChN0jzG3gWs0id2MpHQugeiz3e+aG9E6Pm7BW
Dzizabmielp1DPuO0JAD1nT85dT2geLhSRtsXNeHhbpaievBzsKOQprc33CHieJI
wc7Djnd6ATmLAzSFnmX9Zjzb5oRk5YZR3UjX9Tcg5/APyBOjuMaV3oJiYOEJI5wy
8X8yPf8Jonlv8d/UUXCqTUbmFZRQW1PYxiHoyq8TTzifJ6poExOfHROsTQ9uTz1I
t9Gb5jvSdnJC5xbXih08WK14FICtfto92WKTMeOEcqKxuEzdNJbj176SUOj29vNi
LoJUOrtIKOJQI7SyGYs5oYyhD9RvZhMLFdw9uWieImo5Q0hP/aAlWnLI5JvKedmH
2ka+JG7U23lxIDKVrYopnx3FVqIWYf10V5hEOvUlV4rlrue5bM7SKB2ZztfZWpLP
lfW11U9pkLJPzBT+y9w80ijdG5fRgUhMSiQ/QHRVNfjYeLOIo3yVUKXw7xZYF1C8
cPueP+ElujqiRk9n1LOt+AqQHcqbvCA26tBa/2qMtlsb2kUD40jG2APQrWGDLERr
VP9wIMIwXwQHUz2nwkWiJEM8LURQtx1I6Q3Yl9olj430AeTEhWc7XItYITLIcOS8
r+HVHBVS1r60TN+XDEwnyv9hMfR4pRh4o2kQTN1aSOZxzb4zdkgRg2F3p39n7ruE
PZWUSzxvoPX0F6tM/O2GXHAMEkbO0e73DpsvVlIhrc0gk3txBTPtBs17NBA10fo9
NL1mq7oSj4RIEjzr0wya0U6fzsBio71++CeS8l+SR4iIl/Lhu/ZqAEZyeMxR6WRM
WM1K3v/y8GeJ6kztrZvnhIP2U0ntV+yJzUVaBeRC2z2V8nfAj1WZqu/7zKS5A0GJ
O+XN13Dmqo5+2c1FO/rtB7PSzZYcyZX3vB4noXOIi2BWvgaIko9jpYESc8pKjawM
HqPB1zRPXeu6vnumuvpNOywNkVIFzXnfvflph97YAh4sJzcO7QWxiXu2EZ9QQhOu
JAXTVi2mwcwSKVV/5Od6fY9h4ckwSXw78ovM7FN6KVpLs+w7OO7LYsfftuhP64P3
HqpPrlwf7YiDYSFyM2gzds46pkGcgrtmppaoWpKfxjLkW78d3CVaDFvK8dVjH3ZG
2XPm/whaY1afg/YmEeekfRH5eoTnSqSeeZHyZPp6yiCttkzpkCEE7FsCC+CZrxxG
bN9LFJDSgUpLbHy5sWh2hnxnKr0SC51R2aI4hupgoCfdIcZr/ylBsHgd5hP4H/Si
1/yvib3S2mujyFjxEaP/nDBUbMBbzqO8RXMzy2XJLmmd9/uG/GapQb8lni+0q/wp
rss/txZ2Lba19C5zXTVV/ZWwDcAuiQ2M6vzgtJR1wkK+8xDZUMKHNnEJsb9wzicL
cl3E5MZ8laCoJxLDEfjf5I2s1w4nbr4qjuWNhgkSaa33Gp3F+/JgSS9HaYjf+xjn
jGKEec0vMlFC67vQ660STUtEEsqAFAfG8Zi4jmM7UYJlDvJ3wRfti4Vwp7UTVJ6+
zlqOit0cNi1clva966esG5aZk+eJhxum86abM1c1/vpQZAh9IXf/6FveNIuzGuUS
b+8dpkEZyrHTvZXlrhwp2R1QHc5gCGxfuv5Z7DBaK4ZBA9CD4Aj7vioQL/IIRWeW
90tInt/G4prdQjwQupmCrYgZb/6qIgsyDocgWR9dJIbRFMsonvsfnkUXq4G7i07j
PNhY2B1dpk532+eNQSXdny6sD/BtNsoZkkYU0Pw3oW1yS8Q3RBxDBTn4SGHLSFlU
KnUQ9S4ES0EfR55Ol578CAECiWxqKEz047dBVoOrKpAi1YxAibh8aFC6rkWI8Oux
Et/Un1yL9DN/t6+yfsI7VMGNCo8CfmM8YQXFk65b8tjesCBha7HES2S9+qEKilnX
CO5qSLlgMalGpwbAR5FzNEzHfUWT5N1++i8KQPW+eMaoLh3wdZr2WvtHXAWyIPHI
pPBINantgUE3Qm9Q3JcJn4aLPIIF19Hxf7wHgU9TGn0+0XeDrIJ8S5iMjUU8AeM3
ozPfjjLlm8Xzv8We0B2G8JywtC0uB0bCRYXY9vyp7z7PB4zFrXtXycQhpNqiFsO4
vT96LQXBc2kSzdr01x03bqhszorW6fGc7RcVQgimwTMvDDWAsNkZi3aGIr6iH5e6
nLP0UI7GzW4KGBjdwnrLL34VBG8sLrFXmJE7g1K4WFOtLYdlKBDaN0AI/z6HqekL
XjFYxQFY01m/5FP1q3t818m9fkm+TspfM+iZSQvYdgfeGde+b3d3ZxS/ml7ekp6E
wrtBc6aOHOiZmbAsyRasHiorBAHwmvfms0aS8NAjazt95LzV1t7GNOQTp2XfrYp6
bNF/aqtsMc+BsBP0HEdeX2L9dl11ROvdZjNygKgOnU9I71DVgfayMFN2aFPRcsKV
mZpHNE2Bi6YvoVnwpGcqVeuiLum7qzc+wuNdhqOrPaC2GCewnEHJS2fdJUyoiwpx
2PlhynA/rnRA3TrbEaaGgnzblvqu4AuOoEA43FGh05rYWhzDdnuoMc/KWu1gqN+S
QbqjR/IC4XcRMzhQYNrI/oQAQvoc4mOqWgs9XVk6gDLdg+a23BHyhal0MXWUQqrE
GBKe7UUjoPiSGrIHcAXwi+pQ7S1xfsOUGkHu6sDOxv4NBMcaGDD73ELYmYjy92SW
99meWur8mXf6DprZ0UZF47WttuBqV5bs9I4PzAs4oFsV+goKfMxfIevPYOuzN6UN
7HMtbb4/82hYcZsd56se3bCImbHQI8Cs/v/sSOo1yVsOFc6NPx3cUjnj9n7HqvCD
WnPSXK4Y1li93ysYFDIYxlxwvg3w64KCIHMkQ6+AqNkTHRmQAkVwmKKPLMeMqAIO
kZ5g284YlEE4gbyWMNwJKXNHqEDws5utqb+FQTogeefUT4EGzkK12XI5abWm5ixl
kloxShZPIbnFC4461tc8OK/81YhtBgPxcDB5o4ATJtIKMgvkyA3D6G+jEVKIyuHj
mAc6wAEqJD+2h05t79aD+TlSxvIJgvcpDiKchYtwb5K81ayUHTvkmcEiKHaKNTIn
kDzvBKeC+7+cJGsaNr0fM3LDV71D+dnxIP97i3TDvxOYmYIXICnOx/dES07HVyvm
5vxUOEkv71N4SAtMHWjIkBcqy84gCypUHLoUiEnhXXEsf8sy2AOaDEkaL0QbP7pI
IttVsearw5vIGAWz0BRHqHuqXCo6UkCe70PRAetoG3jnggrXwz/qlnoAugNa5Osi
X0t7JWlcAvFsNoOPot15hdaDG14dPq9KSBnKMkfx1DXMT1xdwpJgGjo2uFkL5Sxm
WriQBO5FGiGtb77gQ0XLpU0+NaXTSOwcF+rAevSpAR4eezVS5++rWnQfRSWwuXOY
9y5yEIPG1J4I20hujBL5Z1mzdZNxP6ODSLvMhsTrwgmlZrtOydC3VFwBT1gigGGC
gn92BADoRzDq/RLuQXc0LnYPP3M2VcTPJKZu9Pzv7PllEbpzf0Ur8ESxVfwICXhQ
RZQwleC/teT+LPB6tG6kOw6EnOQ1Q9eOwmIKTR8FZWzYEvjRDXcF9KUqEtW/xEUr
fP9vmjDguGt7h3H8Qt/hEYjZ9CpqBnUuXlMAHHzT6d6Uxn16UD+rywl7fJ+2kTSp
bcz67Ep86sXtcBRE/h0u6mz7h/cI18ldy6HksXro85uc4+53RvcLuTJrtGdfES2S
aSarPnoZv6T3O2i/VTLcEwiFoB3+oEE+yb4t0Wa25/kh5P4y5E0rpdeh+fYHWMhs
DYH2hGtyXyVW+T4AnkvgbiK7YeVQeZfKEurPSe/HKLw76HMeE7yNseb8Xbeystgd
rxnc8IRVVGDaCyb6NVVcOt2lGSj1iipLU0ladza6HKn7ajG3KTDn2vt+TtgFd/xq
blQBiUHyPKguP7Fs3L39ThPRPrCeRJD5puD72Wtg1G3OsN+kW/Vw8SgQKxrjlD6O
CCRb3QAQs1je/wyBeRHJs1i8pJY0yD5kVc6aRcywcDsI7ggoaGimSwvAemEhnNdJ
6Sb0cBzhCcRzPB5iPntHNpsU2GpxqagcZS4CWvCmoMOFcbSlo6Af/kwKXDURvi79
3Pa+RZY95eq5p2EQru8Pf94m1BLsxuMiuBy9F4Ifblp7CyzcUtkYd1ZcqfIISx1k
1vCq0YlG/gvj1NkgDtC+yIJ1zxk1E0HbZ+HJvk9i0+VOtkPW0nx+3Y1b8BNjkCGS
nZCtH2dewbdYbKDJFuPJ3Jw5ADAk/JYiAtcqkURDoxAzz5U0TjpNO0pO6EYkSOnO
J+mgANhkEW/Wlxw45CmfefPuynCTRnJUUXSwzZiEN4gd179ufvmB81fDoOQ3Otij
j6evlp/wmn+O22hAm+DXGOatf/Le980MyhDPwqN+bXFwi0OKnoJfS9fvVVgexmXE
+VjOjielo10ZQNrAVqTQTbcAHqE6xdBalTB9iXrajdf4J6FvQhDJCfW3yAjwRGVC
iMJh0+hiONkm5wSKJh8UjEdjyJ7Evn1NFPOAhe3PkBZtS6OKSQhCvnj6xbVT2qHw
KzNoFGq0AeJKghJR7jX+IRVTU+5ajeN+gZI4o2Eitr8Ylxp1UoPCQAEb/l/TmSWd
epnq1LWLo2FDu1W6ATIiGT69Sl79XrfgDNYMqKwQlO7NVouDFzY5jN0w3U0pNWyJ
ntuBAsA8+KQ37MNCOwgiODy61or9viTfweLYKH5t09KedDM0v2IMLnU+CO4V7QN1
Fx0rbx1jJVxArm5PaJTTrtRrG8VqMCbgpQnE601NOGYdo5pi32aOR1qJ7Ug4AK8T
L05BBzD3Bgc8eIzTLUOv4c3ZAFurPBK19+u7moP+yLHRdnhaYM3qmNUERWonpTs3
hkeS7WHQ1pxkLqyGsgiOBdA3PQaKRGfcMn/aE8/XQeky70Ot7VvFJcp2Cq64WzZ6
nD/2TmEBCLZrlF2VXv9duyAzWLnGkki6FwLdqrnGbhtHf1SYAsX6d4UsL2am7S2X
MuxozURQUbc6wyydug3sqfS0LJ5et4BFiF5slRt32ZW3gizu1qlaO3DMtNkx47YJ
UC6EVHGRbmkqV92lxnY7kWUCoU9SA20JUVBC99FVvaS60JXuapusD4cuBcNtqUp2
3ELysJh6AWo1CLqyAe/HAORp6j5MjYHfHsroc02HYcAHI5BdUDWuy2AtXQh+xAgP
AH+Kds2Anwf2yJ4vaTRAi4wbDhgydyjy9E0mAonyvIWqPgE3k9xgCIsCivf48EwO
1vAhknVm+qIx0i4Aq4ZqEcdKJuymKYVzhqasZIdjJaA8FPhKP/Fs65Jjgk+Z7sbp
Wjx0tf6FIjYP/EkyQJ21/rpbzj9axd/9dMaqS2x70hhbqr0ueZuJIfxBNx8Ulm8W
O0LkDYf3Wi3Fqy55TZisw6owP3kyO8J8lbn8DeraOJUcWq/pFHMvfEeOHiOhTK2O
l5LAcwKPU0Mik05NbGNH6yrjOzlqVz+vkble6G1+a81cYP2B7UZWUpPtRZuKTGHb
BDtmK/WTmngUd8GiGDUwxInn3+QpVajOuVJ2RsJUZvIkEw0d+a756lUX8ZcRW0MV
sjlrx1/4WDkhMYTvQlXgz/iSFtAIneK6RBpO1FAsbTAWTGDniyZ5EqMdyrGmkIuL
V7w2Obs+Yj5pQm4/9u18E7sCa7qTaorMeDETUqBcWs0vclBgWI5T5x5P71hkD8H9
9PC1os7kOL7D6JgNZtyEek9p/lVUf+Oiot2QUiIo7rFQjruXWjtuHSlkOV3tNhrJ
lNydLfP0n72ZRjhBCJgsTVdRH8dVlWqxWoqJZPMtt0HuxcY1ByvuLrrudC6k19Zx
Mk557O6I1+vXH6MYN9CxRjo2NkhUFA4VCRWPamyrow5txvTqvu0m+gHVMci/OUVA
LdxHccPDXV/dbpQYUB6fXLkAJ2U93qjBkQ2X2f6137Pqm9SbWngi1mFOWB9sXoFl
67RV2FO9dWHL6y9HGet7vLWV5Sgs8xN/SRpi7+aAtdw25n5SfDb7n1mzEfsmwoAL
IFsomzjIGg0J51FSAw+28BZXZ3TLwmxDkM6HjggkhqhXuQinqF39oxRIVu2gdCiC
4ODiwS0LknT9rq2o0Jr3VEPbDmxurHHz7seR5zzI3Z9jt3ez2RZK6tX8yT/C+I9L
lOrQnzMyyBm6o85NpDSfRO8E45SaNKdnOIa8ys9Qh9QFQg/FmCxYGZX0Db3b6QOm
8gKyOyrcX9l9e6bL4+lNhLZNyewUw9NpwfCtuQTY6AxQE332xKkUlzynWzDFmaZX
8Q7HzCI1CQqImpCZn5YKf27AE9hir2g4nlG04vwvS6Ii09zlE0E5cmy25Ud9dH7o
Z6LY8edImYIojsmxZfU6crq9xEhWvOq3gROzlZHSwizgsObXLxJwZLT0/LE5vDVJ
CNNQQhF4uV2ZPqiF7KWRI9fMNuEO9vcBCcENQChjNLL8mqwxVJYN0Al24Vmx4XL7
uBP0ii1Bjg+ppIgG9+/YSo0LSdASXRjxMo08MpYftfR/33Bz0TWnWRBQdhd5EmHF
7BirC9Gsuq9yeDWWsoW4Q0upEZpSWO9YxkUVbT/SLeUvT7ziZBYSBv7Nl9K/7+Ku
2RAitNp/FtDiq/55klzz0vDLErrja9Mmtx+bxkOfsiU5ZEPE7XYodjJEmILA8Rn3
J3YWLMDdADv18aUxn13+q4oRlp7dCy1XHekqWumTrPj7h/b4d807sLoEm+jRR5Jh
lT63vTEamKTyqWqpSejEetBvqSjBXZe+qry+bz+oVXPkltQlDFiVKQNgsl8Yb/sp
swUlCLa0MvlDVolqtYJGDJOD9VbUlH71W6NixhZbnyKz9oeubW2qkTXod+CW5iDJ
ibxpou3iTXDC0BvaZtE1xkfa+453lYzaBirF2gGlsVOR9cl8DBSF45cr8GFo76u6
ATmFhI+VgWwSJh0pPKcwFJHSP0HHAjdGQAYCXn8DD0KsuH7NbC3zyzut/kp5Udbh
e6MzKpBkwSWyxleOrWuFLN4kLCmS/qDfHrqaYO7DVyDN9dentkpELldbaHFfUN50
aZ+JqnqyjSL+9Xfk/959swduLGKBgFXbBaEbFXths9+TIMr2vw/2Erm5monbJK3o
1THt8vkDeXTTztu2yBbeFOfxGk411CUt2Yu+AwLcxYBeczfk1BzgETUfHAO5GWzT
ayhNAKO4I+DCHQqFr9xvZXCD9rXtgXoY15/G1xlRFphiLPDnsYog1DN1axIG0v1H
NnHajXZkGT9RKOps4BWusbDpfL2F2u98oH3kcaDTF+Sjei6opgcP9rZcd9YIdOBo
w01y2otUW27y/Ncl1umRrFC1TP5HbV0fFzHE00EO9rZSDqPM5LLb5xAHd5X294xh
nekNMeFXbDBLjKzhQuH5uiOyv0CxH3dHx6fabSKg8ex2gEBqz8yVQohXiMouKhXW
pwBkXWCJcnai5kaUT67oWcasZoTBDUDYpNnl3s7Buty7vvL8xlzGPtJgygNC10MA
jpfuk5xWAMWEL598Dt6uUFJ/OMNAWxQCjwDI2kQqd6n71aZ4O3e7ef+j5A6xzJax
TpgelcHcNtv7r7tHOwjgwBRmDq56y0Q/r/heY4HHwuk48g9cyZJ0J3VTAz/vhU5A
gLu2ZIB7fkshyRHixJR7CXROqmqRQ0Kk6P4GeFC/nMFcjyBYRl4xqMtSz0Xkb3AS
vsWlv1twHUOvGw1SLmVaHzLrtZ0CZDFCI+0pxDKZIheOb7HZRHki/dMvURS/pvkA
LwdgsVLajnMom4rRH4oQkVQ5dHRq5Hqz+eSbbqZwnxjpo/t+rkHTplfAcLCV7qpO
nDoo9gkbYq240J5kJcXDTZkd7xWIMmkHYAUXOY+mSEoNz6Gj+XKpQA3adLB6XOu3
2yBmmmyvHt+lCw3msifJ+9bwuiSjciJCsTtNOT99hY+ZvJRrw8pDVbkZTC+iWzmL
06kg+QRTFTaRun5V6OjkjPjUluEYwiLeDe/amU7GoEECrHFMyTHXhWZq/J+NOKS2
gckbQDvhyi9Uy2yDVKGz4Txn4zRMCRRYlFrbNp4TDW3r/c17BAplV9O+DhwpFmfX
/CNpW/dhHMB4+02AyTGHOa9iLkSOm4si6e/kMd9RcHmv+76ut/cbFqpdCMjA7MuI
nOEthfiU1CT4VeBGTZALVE5EJ2eq7Nw7PGceUH+EPu+uhvUYkc2Rzf//M06hVPVM
1W+hrlfsPj2iemzWSeRmDuTBnAM8Q7H4S1tAtRxB8u9mJebP3X7m7+/QTiXVqvNm
Y5ZIGrMugTHAYEMj2dUuWUgAhVtbMt/PzGiTAe7zjHr0O2P2fXMAzo8iktRvVBzQ
bLme1w27itVtRZldttSA6kodi/Q6n7xiBZpmzb7O0brIVoX6WGM6lZg8BymuCDl0
N0wJacmuhdPPMfIk6wrRisQE+6e8NuN5k6oNj3/wAKtW3OybSXM/gvYl92eD8xUM
Z6ZEZVSLb0jbMfTAe351C39edNzUq09vjt2LNqOUSSevnvco36KGVnTmrCgGYMr2
OXD9HhHGhYmAq7M+0MD7L2yzNFh+N8XShulMf+BcixMZHXaYuVCnNtQj0Txplrye
ZG6u9IrbYiVPZvdQ3VEWdBa6xm1vkazRiuxTwz0Czmp2KJMvX4vg2t7mGaYcQkm0
1IH0CkHmdjhDTDGY/bJQrLhXamIQI/cBulMuRu/VcotCzuYNhELDmvMwZEeNuIzl
dhkxHgQyjROYZjLPHiOgP0N44DHFkKvbNrfPvzYEALAeq+AqlF6RAxemRmpSJCVV
JGZHs3PX/5y00sZ+LXkFu8abudf+LEW0LLSOfFQMLincvesvoU3DwUElizLpKXUP
TvFYlMmVvvB+I9IrCHvPbA+fKGWno84Y897DT+d1Um5c4Xof2vd3iIoGabL+v3sv
YLbNaTs7kviIQNJBgz02aL/cFmsqeWSNbGb7fyq0rNMhlb+7CShPrnuomhYjLtlX
65zQYbyS/PN4eXm1qiV6AhgN2lZ1KbBj44ZhCV8w8Ye3b7yaoDpZWR3mzFrbnSVN
SY5PkwSa9uHlq+reMdCGd05r8yjEdrgTILwd9k1IaJk5ghCKyv6ZPPfW2zf20xDa
mpnUuGvqQOVM862Q3+JZFJpNBucCIWIgJ+CKvVd+nHGyTmax1FYxSCaEuAJtIOPC
xoPTYVw+rkr8lrd0RFPijV9NMY6y4Blt+CFREQoKPBn32Gy2fXYEq25Y+ThwuOQ4
/hdOogy6tJSlI2U2MLJFZaqAlmpuaL6ujPbKPZcbCp3CHKkdzGjeklLFXAzkLFI5
BbJ+rsDJB7J+bDSDkfW/JwVbDd1qrrJPK5hed4R+tmbqBNrrde1PxAmLvXeZNscV
n8kySe3iWWazMkFJZTJbs04Mps3vrDkbCPocBdHWGk+2Dv8A2BtsLztDq2dAJjAm
7VYhJ1SP2+b3EHdsDeMxhj+uzamw29Uge3VvtN1yUXKifF5LhDb6ESpTYdN3+NXx
ywkS80yeduioHFdhhTObzQ+EdvLQGop+6FUToMG5X9pKsZ2zPOZjNrPUnqz6DDpV
r5FiIw1GsgWiyLj+SxMRmw5tcd4zzfsvfWSfaYj0W0ciZDD0q4l1GOp1n3fsnrO6
bxDpHD7KCJ+nqALv8lc3eCFvjbhlCgDr2+6q5OKYEinwAgVOsTeuGEfO74/hZSlJ
IGpSg2P/zyh1f64FuVs5MH7CdofwdSpBPc2JVZs/BXdoT+kd+UBZqsmpl6NJ7xaz
PTQJ1VCVoN05+86yZ/L0t14Cb4OlidI0Ul5/S8KxxrjpC1lRlJtVuvGrIZil3+gU
r2PkBKC0w6xmxY2EFqxYofx6dPrl69uhLTKIFWN4kC9ga78ywmifP/cWFV0SI6Eb
JUH8dSGNFoevT6Vi+gAORI9MQxEQFnAt66tyvwkJCux8N0gdomIjdxiHRSxswcgf
NwjMdOratxyPDRrEPQHqaZ9XXVl/yclfvUtz24rgTYy8EE2+n5VuUtlf+u435QIs
nu4L1Rv9XMC+vf2ZP2nuc7T2I/pMASH0RXeTmonBj63Aw+Zy5yBh4IkrzgG4xHOy
r+0J0FsKcaKY/ZrMX08MyqRIFl6y6hn4rgejV/5Tv85hkCttk8cDdnVh0PpUgQTZ
esdVit6B8Km9ZoEyCT6AdZmmXBCvT10w4yj/yjsaaqC8FE1LXhmagSWDIZAVIFu8
Jxc1kC0Y6wzokpFt8Dre476Zx/L7YD8nwTCYh3Ptkd5ry4ip36VMXDDm3YdGHwM0
MISxXtoRnfPHvdoV32G+hQe82BbsC0NlplZUfliNBzDbzI3thnFrz1Cxq13nxu8Z
J9hZWIpytgCW6kqxrgnbP4WlzGYi/VZySgXr5nwDZykFccOB/BrdXuaM1WebmOL3
2+xsOoXoM9xI1I5n7B4L306Fr0xFQaRNV6+g9rB59xN9D7tFqWGHLSOziopT5ZS3
g7/m8WqguUwiG28hjPFIkZg33Wit+z/StHCT5E92tMjoOuf1aKwophtpEgqMTNLx
4RjSgY6K9pblbKd7tlmTuFNE9PKrvk4ULy8W0Z4AimKOKNEGuKl1N0erCn80lDOX
d8S2PHbLEEkYckpGxQv7patNwT5NEQROWEYBPuXrab63hMonw3EDagkdF3qPXIKO
8g59tFUN4PZiZKxg2coTKZfOD0adA/b6b5YILoSbwmkTmZmdilA18VaIpGzVZsK9
P9hE7F8Vzj2RSFAEgtgod/4E5GWkENka9/dpwEid88dScRRNUbMjyxIHYyyYSTdw
y2voTf1SOUaQK8LgyvZAEln4CFiQF/YuWx8OC8RAUf3SO2mXTeKVSFstMNcWDUDv
oIEWhQi4d2dculyeD+91EQdYq2kjqXZ6n6ma/i2mAhB/wU79tlfoh5BAJPGgsSCY
Jap+G16EZmWV/8jKXShSUIZpx5EjX8oqs4wYnyalBuSyjhJ6byaN8OlowlEVw2vq
8Sgkg3l2Lvz3Tgd4plNAilGZyze2TvfEHp88Jy2zIrlYkjPtspkqgbOv+zqeEgSV
I3ss1w/8nDyx2On4a4emxnl5QXjgq0aSOiovjc4VOqVtpaYUKRhGqseIHFD5bdJ1
n6nBw0dmPCe3YdKfVwU3oD2obONyWd85vNqMKE6HN1KByresHp4hxiDD1GcAvj0U
aWF2pmXQAtQHtGDUydqLGqga1rv71Gn31Joc/rB47bddGE0jUG2ysOcrsBirX42m
V0DbTZRjpu3g2NP3GySW9fzuY5cw0D3gKgVM+7K8CMzTyG8eE9SbCd8O5Bcs/KOr
Vvi6kxeprv1eCT6/Wqw1L119EguhN9rMd/tlf7BRxPBGFojsIfTZcVWpFqfiQ3TE
Yre1eIKWl6kDhdCKqIn6qM1libhrOfOlP5i/ZOzeA49YNrOrXaxNWzaRDxD8Qn6C
KOGB2iEdc/51L0gtWvU9ttxo7AdHnqLqH0W0zoNqfFQhKSqI8htzPUeLyNcS9Neg
RodE2hg+tziqjYu79O1PsejFxMwq8kRJLdVzn91+mLt+nUAFj0vfDVfDcKmvft5+
Iusa51JEFhsEMcPmXhMtuwMSn4mJK9RWKu4GUfpNnTwyAoFAkWFmrWsLQAzx1A4Y
6MEkQ7YXadBolzvu0JE7bqofMQ6twDdbDHMSUlVZ42NV57rhAWwZzbQjtXm5uz3j
GAU7Gtonxr0JTmEezDlNmu6X5pk62XSKhx2Stml33MpJo9GoZhIRN0m6C80U58Bc
JFYmsGn8Pw1GYT14edBrAMWtN4KZ4ih0IB7IbCF4WN1nTDwnXB4Ls8AXh3xLpOqg
yaA40a9gmYBASUbK9HTf1cGR6BvLfxdwfUkxRBURR31nHT/IfSKFbM+BdHqT5X+O
21OwdYH2UeFD7WhMobmM3w0XA7DEvCkXqsADaybQOEVUl1+6wIRyKAiPE/vaSzs4
+LfIUvn6KNYSMCn6drSB5vDRwfpGQPSvIrgBOyBDgSL4pNCV9UEPEsBVrsv68nWb
vss4eTo3Y3BHOhdZkBG9ZvoybWOcsRykzLphULzH0J1VD4uEW2xh5ktPlFMJR6AR
lcHqXZdiCJ6DvjTEDf+0GXDgsqsMLGy9K/B9p5YCVUf/cW334DNTJZjDPeneo+An
rfj7AxVya17mnfPUzxu+mvv1Rm5S6dEEMhfsPQwaxBOYhotgXMdqboR80Ziraauc
otezosmUNROdYFbdW0uJVTUqvnQhHMT9yNdT2hE5XCq6Gwu1nd/CRQdUlUniWriG
mVGHjbIvT///kkPDBAoHUGcO922O4XDdpdH+DnVwGrgKBLrC88NKBwvuBtqJab14
TEbUhSKpynHVmEv1+0346VfkyvmG1PtO2MMs0P14Zph5PricBHkSvO+d7XaALn/d
11G3cHDsPteyPgJJjEBVVO2BQqNWIGBUV9QCer70r3LfAkGDPcyvsM3bpfFfqLxt
dZL6Jtw4upkPfYpUyATOJB/kuvbaIez4W89vpnMIYst3PwRV2vCgrG9QQRuUeFBk
nWM6+Eo4PFNaY2CxJR4y4wLBjwTZfcILIHCIdiQTxFX/wZpBHbqci5TT5W906M4a
iQwU7TrGvVwe5MSCOmVIwbYu5YylGdHtodk47KJD/GXH3G2lNmS/eFdvzgJppwED
dPWkeNYI0eyu4/llfF1gt3Dy7QdA0Ugtg17OBZJ1A8Y2vpl1UqVGK573mWcS5dHU
zutDeSRg2gIQZdLaN7Bi6tUFbLBPnWKQCg9sg7pnXVj1EPijArxn3ve6u6eeZPQ2
wDFPkeMS2xv0DwTzUVQW/702Qauks5hVCWjxr0jChcyRSCbb5UF7swQ1lpICHPVl
nud6SLjNXwsZCpaEMxWsTeaHDFtEJ+goNHZ4K2ToQboi104klsc8zhCIxFeyIvfc
Y4gqAwezVDEEprvHAbfjCrps+nHIJOCon93P0+jPxdeitCBdCUz7jbTuDoM3laXP
8GxOpMoyAdL5UfwLXqWI3qSeJetO7cFR8qsmnRUAzPKgxXkizsoDAUWUiZGy5hHZ
fNSDej3DST70MqhR0okO7mEt8zqmG3vVtnk6s8pIsD74rAwzq29NmvRjcT9ovJyF
xJTBfolZonQ4z+MKMH/0luI1Y3WaO/eqZGTzblqxM8LBln/L5JCi7baj2eA6399C
limQlKEnVK+BLh1cxAiQc6SYdFfeeetdad6X8a8Q01hKZ4PlYOD9T4S904cykZIt
2+y/dyx6XT4CtJT9MZIqcCjocdN7bvS9KnI6Fjejv2TJYEAcvhyhD0Fq79WfIYK0
yBNK92Wxmd8/2yXYwj/mJaGyNg40LL4dTGslnELkYu9UoSN3dVqtJOQHc+vz2LkV
ecolcKMXnWoQpuz0iT0Xt88pzRkHKxmx2Z+IC2a08sZTkWWRut3AmYvrnOR9FK+T
dw9fstO7Epov6EuvSyJO4WIjUcbis/DamZCLPOpfMJNTTxmGZhjnVij2955w9gCh
nJPyIa0dVY1cJ+jSJNXbHGtK5t03AmKzm+JoKcCFVfvdKR6e8CDR2h42O1a8561J
v1LUndrT4asVpBKViUFCZQc8agJJW4ViA0zAmP7Mp2q2f7Kz3QLAsGV7G9dMNA6Z
UKXW5X7XMhZxIWhnLdjDNgrfcBVB0ib330zAAMEJuHdM4iefXsgiVFWhGU5PVptu
p0eRcO+JyEQ64diITJkWrgdfT/3JNANrccyRWeF69veV/CY7EoHi58B+WuQHUP7b
Q2WlvJqVh+1fuJsRr/8OaIcGTu6i2NLt1D4wkOm401cxbSmjZ51n6JOO1ZWzVbkG
tE6LJT/U6MjWpWk6kFtMCcX/swq/x0mO0GfM94ZdnDRs8ep57jW6SSN3ib7tBLtV
KqxrYwHez8fDzPXtuKbv6LI8wp1jZNbdmB49oDCyg1DqqOQwAMk2RIag5ePGZpn3
aKqFv9ChqUtTRg7nQGCuhunJ2TTl5ZMTWZSvT2lBNekogitosVWTAsK/ndlJ9Jvj
k0Y9J7F5oTaRCraRvONqWzJZbv/66NnK4QH4oYaiRCQ3Map1jH7td1neN3DI4zUc
17wk7IyjiX0ecXII7MBBvGHrz7SMFrMYvADML+kGt2XEVk+MFw1mWloqCAmwvSeF
0zBoNfHjW0+CXqMlhq24fX0n+LE+p2zHtN11eKv+ORQ9jsxQgMPlK4TJUUop50BC
wyWs91XOYxwUnUNy4OikileENCYCrnWfr1BwHOcQmIejeD9dAVgK+2FLVHwpcPXl
gkWUePTNQp/0ygMtkCgRkrUxe4fxkON4VZY/Cio0lHHbIksgbX9uL28ADTZwhzPR
FPrCNC7/0LDvXjd5JKhaEQ2x08aCSvAwtn9SPONSvMCfEw1mt29EkBnblGoDsU03
2CHp6XluAOP21TN6AFsWUNPl+981hkYz51AJBHORytJ/Ugn9RNITxMH2pAaXpqMh
w+4vj6fW+RsymLx2bja3fkEribcrxzvoPIYHmHR204WW3rSidj/kFkJmb2OTP348
yqTiTJXMR0EuzYm/+NfYWtsJtJEJ50egKKB7iwv4yXaTh1qJiJr12i+WMi2ljZvV
4k2UtsqEEgq/1JjuzjWKd9ULn7KS3MYIMHNy4/SAGLOA5J61VijUan9omg59qMjD
XfZ9+Hb2/r9G8KVj3v43Iv0G3SqQgpwG8xX4c0C3WkKHl7bMrJyJKxVqZLedMBQt
eRYOcGJM5rqJMFdCR4m8tXpTZ6sGEY6rPeqEdTT4g7Ei5cmSzHM4xXnHOixk3H0g
dWOb6vIDE8eWO3u5oTTZpTtIQG09coiGjfzr26RmD1bQ++289OOiqK1v1MrCAoml
nCdxqw2gXw0eoizMKE4mzOYGOiCdjBIohwiLsNBEchdgct93+ESZjqWqitNoPzQB
jRbIfJNEjk+690TA4x1w59tUIdmtNS5snZzFBxgMF81e+VCV9VpCqt+vkoDS+N2n
k60IMviwp3w8BNWxQkBMfnBOUQosytFZWuBBctf4zrFsZ/bku7sRoqQ3neZGPuC8
CIrvxLMCkgWFmpce9nL1NSiAw7BStNDomNn648DsidXsEkic42ZhiQa530ozwINh
99dO+9ATGgLVYtWUJ1qi8pdV1512Wcm2yWq2GOyS+wKg7tvBdI1uJUpC6MXeIBnH
zG/pcf/Jh2VZCe/gRpK3V69WvVU9ITc/St7vORKN9gLHGEthVpnNZ0Nw20bcgV1D
Z9XoparuABuWZW/GLM+iEYNAq0PFcSnBlerDqYsiD6lV7Rth3oBwhay8/WUIc2RD
BEkWxZmiTGsjT6gdBOEIqaQSsAWJn+uPyl64U3PdlCzrWqx8Zf+aGD3mL4hI7elH
7xCiImZAmvnJH/1q5Pw3z8dZtYNXptLlp0vvO0X0x21CEmwSR3aOSr8Q2L+byTzZ
aEw7Cyf2kNw6PrWl86CYN0fe+Ad4lQcGLraDZpYyUrh6iSEo5kPrx+RDbrBDBg8B
8yisgPPAtSBqSZb/P+DMwCH3jsFVBXx5eZ7AbVsGzWVOYHsqalBNE6EPjmNrrt4G
IJ5XM9mgxYPdyflF0v9IjB9RK1OR9Qs1Cr/pB+1TRax4HJXC4foaW2YmmuB/7AcT
y6ikPQ2mtVCB14UG2opwJpzOsAr0aGDf2DJRWkcCVytKt4485slWjuCLp/AAOQZz
+Djaznwr5dflI03nOlF9sQo+I7BDFY39sXHEvwBd+LkD7GYQbAHnEBi+xLpsx609
cCIjH/OTekLAAAyTJhPWMlGGnnw80X4oKRPK0/6MVjv0j0ZE3jZhUev0G+sWoHdE
TqfALa7vAcYJ6C1IHf7kA0kj8LLWfevWOvAtjH0yTzQfQQpatZ3kfMYs+oyn1sSP
M7M/MKKFmW5goj/8jFg3TsPQLe9Q/UoYojs7e5WfPqBjkv4GN3JV4duAGp2vkMUr
8uxCc2+56A8v6kRYHepyDtcHbu9kN6Si/GUHLMoWR6Jmc4f7gaHaPgYZM0uAL/vQ
liPts+AHrbuVZRlq9r9+U9jfcx7Ac0sT1mLg2+N3FMEWv8TfiWfuT8KAbMMSRHeL
MdZi3xvxISgub18L86Irn8598WWjWqCukE1v0R8VPn8U2IdNmN7VH2MSoftgIAHk
pWnEBffpHyfObYKMTXOQG9p9LlIFIkqqpJrXSg3UhM3Xorq0VL/YogYmZ9ExMhPw
9jSZfCv28tL2uEewV0Upd7zYrDfKSFv2Vqm5j4iqwKjPAJl0AFA2Nde5mpQQnB3Y
AIL9MF6JTR4ah6JQ913COhDCec3cWlCnIw1PmsZ5jjXPao8Jfrz3BnKax0ojDp8T
Rx7o6tkRIIeQwYAmQtEVDQcoauG1IPTiwA/kd0KYDT/NTn+eN4lVaQ0LCweBKruR
T4ihsIZSqhCF3bwP4NGd2Bwx9AB6LSWWY1vzAxwb3QeO45BwbW4pzXS8L2Sa4oKL
0h1GGiubpA8O6sJNgYVrdMBrr9aXdpdkpQeKBa3sK3rjVMAjm8fGkMV4D+ywxIwN
uHpfla8er1v/85N4MhZAjdGqQNxO1E4YRLeP41ivaFNsDkLEG9BtJ+HAKC+Rqkng
bJvbm9hoJxcYlXrnJ+0NiauvjyPIpI+THyo5ELReasss92owOmI7/RyGK7dtSa4V
dXOQbcIXSv0uVokBdzzmF5iyJ77raJlDRUHwBBy6bPfgEeSXsTYfpZKw0iQitGdj
vtkBPCa3EVNu1BocDIT3BR/vXS1BJp/9+a7AZxk3hCJirGhteC/aQKFbkYRQ3jwk
xdjbS2J6t+xs2xMqHUeeo8bTkand5OPpWrRJSi9N8zc6mk6i9Jp8/9OyLLPS9yTO
3CbcbLOLGBNQ/+Z4olqqvJOprZpeMytzJ4eMDOpWd92Xpor+DhW1CXHCIA7OTvf+
M1HlNMy5tHXSs5dRLmg2SnllhKz5GhOCNPocFsnhWJAE1ryqUCOEoVI73yHfDemw
qZLehwL0/JGNi9ktVyvUljyt88NxpHkyHKchD+/U+WovTBV79nzNRncBt2ThK658
gvRDeH8Pr7ldzHyUVX4K3P9YyD5f5bcSMmVsESLm+y7l7+p/lGJav4RT0PuCqECP
/Nb7QEb3Jd1eCxjaW+U+Yxy/hhf5f7HKueT1ltUoCOvi+boZLRDgNBJB5bbJ1ZW2
uVqMobLoIOBigLLIIOZ1Sr2EleyIK5XB0q7wnTt7KWWHmMWvsiC81JZMr+ZplLbx
7fCmdX0vboRp2VUDd8gnXN6rd5NOoA6Y3fcIpWCRSCh+pRnHHkaoCBPD+KRDYwPa
DQpD2nIaUBVVDh2iQsMZ8qPSqpCm0XGOspw3mFjYnMkmiIV5yFIGqkFZgDr7cBgI
kjQuPc40BPOKl5gzYsqF7/eHNjHjt2jIPhWEqvajbOkzy9Bdrs1uzsFKtNAehiq+
yEQL13RsqU0cTTOitTMHk+VPwdr8FKl6WfnBcSK2odP5SVX1YPltU35jOBt+0v3p
KmzEs+bkI6kRMpGxPUAVIQcKXBI99VDdVDM5Ugta93/6lVdhjly1TB0slqa40/J/
hiQi6GOH9qlNrVzpJwNhHNT8EDMra7PzFmFSJhRxO7qLhNaS+5XDiGDs69UgWSa7
agA1nrOBk76OmcijCOvHW26VQYAnDYmla7J45yfw3V4InF0NkLxnDpk9Icz7bpxc
hVGwJ0PmofelSGRvqJlcKg2RtUPzCN/GFCby+cSarTrzKHoihffoYvnN/5AdR4tQ
p5So8SnAnozh5xrfgEYvUnLpsaMThfzoGZ3gI/afUZ3VAJOeGXEF18oTWUvLvwrA
lD9EaIgpIWCEtD/zIfIjQ61LHnNIO6jLeWo17H3QzyVqxGUpu3Rb6UcE9WFxXLyJ
l+VwmBoRfHlRMLsP9WZI+pMxYz9/XYftHhxeWC5hio4fpLBDRYg9l9mlvlaylxtf
QlZHhFXu9F0UA07GO+ISzt718+kSFBl8bIXVwmu8dd4BMH0rWJ9R4FEg3eU6gw/8
i8c/cacn4X/b/Ms+W8EKcs1uY4adxhRVQmAowKDEIBp7Uxbg2oBUFaQ273jxkqv8
a6catPeFmupJVHYUOvY7IXDaB3IRWwT/cKCrK+TZsc4BWLeMWBwE2hfgQ07ilSsD
cKEzmb4jn8wP6JaAPqdsvbWk69wa+oNDFWl3gvHMewJoasw8FGihCQE7zMAhy4ec
A5q6r9OsJNbfdcF0016ijtJq4oTQfNnbHl2XSzVFrtE3/r4e+VI6i/g4VlAowBZd
p7VrjN0QxCoUtdwqWJhQb6GliNsPNTLNkNAhGKQKGRZlRmm3QRX2hGIRZnhVrR1a
m4NDmFquj8VdqECuk4muZvy9VyzZmJ4P+SEmvLfj1hAzAM2zZJm6ipBWm94HcFsf
WVrktqGSYV1sa6NiJBrHM8hLX4uBBiYjaLoSsrh0DDzRxI7wyhIuO2gjKaiUYA39
uxD8GkvD4ylBwiytnxVq+Un8zgL51ESUUnn/mMC7h/fSOlJh2gJdrSyDRXePCswX
sZSbcNJ7mxInOZ1ch09tqL57fMQt++djP9D0dWZdFaFNvDyV54WRf6ReiTgLfqdX
KEFuooMygUxZT6BCAKvfi9Klx6K+lOqsmck8WT6+6uresQT+It+kraCL4Msc6YtB
w3bxdSThewIOd5/AcaWLoKvMydnyCxAwVajH7hXJetm1i+PoWpJ8+JwEB+0fQpIb
DLZtboYzAs0fgT2nOPHQPHREgsp4fEWg2EK6ejXeFKnwTe3rzngOrdTEXeo3Gjri
g/ISsoAfXKmorxKNcuBq/Pz9R0VhluFrZodzgSIDuh7Ig3UJ3k6PlMDoekJ4HoxH
qXCeWtAArV1ulgnoCc8K+PUJyRgiqNeOLMsASF0a6jqPGW7QEC5or9XkziYrCWqe
5p8hJtQpjuaQZzJRADiFv1FoEL9tco60tVfHdm3c/fmF0cCW9Ca3yLZ+URg/rbG5
zq1sTOWV+y7pIbmFogNEWC52WvxvOR83YF9g/Nd3hLLwwilINGZlCVUJkAKkU1fl
hvDJfQQOjNw4LBM17thO9DVHAFK9YLKgXweTUbBbVmUeSGKMMooVtrcafOc09edl
7fR3AOnruZnk+Wv0w9QP7bJVUFPhOklgZc/GB2Zx15FUr72IW1ToWDXlxtD3IvEX
LxIoR+CKFqG2MOlgoL/fgRAxQgxUfBjWsaaFhxsxA6FUuVCRBc3ZLrxZS8ZRniFs
0n06EKenSbsfGTZl8kNHyWUIhJK91Gc0vvAz7nMkjasUpV4tNRhtN9KsB73C8g25
rlzTGrsObwj4ulQ0JlGTrFwNpc8REiF0wEHcpMV13IrnbtbEjJqAOjgahh6oDKoA
L3iC8Uf6dSkWOqrqZhy3QqAYesdGrM9BFL8vpDazgXivxq2UBtXqJBIrIKchN6rj
qcKzx7xgWXlFa01uFXh0FatJCvcwyiYZT4U2nhdadVteV5fOlo8UtPTYmJsf8eir
DbZ4dTP+AhiIWaL3w1dbeY11TlzRtQAsnkhB8vG1o/Qn1fzJgSl2mCXTwJ7kjCzp
43AXd9CuDKkHgKAc8LIvPh1o9+Ub7ApsrDyXmQEON++DULA3KowpiPqc9uXFOwvQ
5BlYvBymng4HARG1oDB+evrMCaKrdrlJiO0WPTSyvomTRakxHVE5QpBNgZHKQa0q
CuRQhcHosTDKoUGfFyd/5xNP54SaOUMRgwJvC9iV4uVoRP/4UcqhUN4SVN3z0LLw
`pragma protect end_protected
