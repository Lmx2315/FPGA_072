// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:32:40 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Vyo2EIYamsUfBeiiwTFbDAUTpfD+kW0hi2gD8j4CtwTCdk2bXsP8dXM40PBIK43p
CAFDNcqppUvmH/rcZ8VAH0WTTxNg/W2MCSS1XdcDx+ViWiqjAHVkt0kBbklmf0H2
7z19EllkDZ8ajZHQpRpReikWiQcN54piZrBSVpamzz4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3040)
lOfn4yFqwA2E+/dHdh9sYEMkvhap4L6W3wnRkWfy2vM2SGyZFLGe0JnbL0hiXRXE
47yWk/1hVDwcYYGnmDgbnwT7d9IJC9NDXKKiUobYWo/rC16/bZaqny5eXqwGmnqa
HJo7lS/OTqV6NtgycgU3YoYGASBTN7EueYsNU19qGjusOKbygOTyUw+VtfX+SYfS
wYAUp6FlhTHPexDvE4Tqr+sNG1zo9PmJ7G8GJn9xmt1yNL6dOFI8NFiJPQnR/nOs
UvZ20sy75xbf3x0X6qZewcqzeGKyn97r5rTvQhfV8Mb7OEk918kRxRD4CF67ACqU
1Wy2nsZzjqZowogJgxFoAanb9oxmfjSQoJyH8bP6oUrb+34u+t1q8bHVA7VMRkqE
iGhBPYGbxUsUX0FNyA90F3Ertao/X84CIQOKhPWNvsOWX8vwa5e6caPMSrgeUlfN
4yYiOCSDdmvlBPKseH5Xqj1Ti6fgQGIAgExZJ0hK7YbHRkjKTCLIQlgvK/jRSA61
C+r0EYcxKmc9uljlKlfwpocepGAL+II9PExm+tHfDg2qxmSM3d9yibV0WDWP+6SF
0RykX4zdQykjbiE9mDNV+OPeDQzYtynd1zXKJRWMBlkvKfFjr/pCRNj5my2iLid/
rDb3E0cUa/uxXCiiRixUJMuaqxpJ6I+LKyV0MbcR3Idg1pJ/I5R2VS5lL+Xbw63Q
GdCu6Vaax968K4jEVZW64xJ6cPeUSfoimHZal8iIZxq8O/BB6wFKOt0RYtMmaRvJ
XZiFRUprYiAVmPOWIlOptJNg1TPxHUlUixyYeJVtb6hLUpTCyLAyankoZ53lDo5j
McK67TQuGkNYVaNxG9lZaxPREBlvp72CfKNsrupha91YtYidzV8ZwHU4UbMYOBiR
+Ue6+LRH3IZGgn3qVOCO+F+xapU5wHQgYFo9OpbJt8rd9swED4cQIgXCFDE10H3k
SDqEcAksFKXv8k52AhWCuyGzzHw2apKa7ap++9FgKYk0ZDnNZ3zn4CJj+NETAJhs
j6FQgShQGyUM+jgXvpoCkZ9MNnOkWSCfjkwXIf0WqBUmSkqaNzm5fFf3StsJPsCW
b1O2ZGvk3C+YTMHTIFpwu/V3zE/ieztXoozIoUuCTrbdS7NbXLyEECLeHXiunBik
zxh5dcpuaHEnBmzrNYsouGW+K9Aka7i3fuDRXDfX5iMMSBKIIsf5UQx0XHMW4lAd
hBbzt4F/aQbUXWh+MNObspRESgN74k/XvGvPhxpB/+DvxmOtyTmb5FoygX/2XoMu
UbmEGYePGMZ8R/yjtL3Env7fQluP6DVFPiDCwQybQ0d5hLwl1iyFFYlon6OORgrt
tDKenpNT0YsYu0PmChub+O7d39GNu4fLW/MlN3YhSBQrYPeopOo69rDKQ62WuJ9f
FBeZKSEpqUMmpY3Ldvp3S76nNT+qD6CDFlaUhMXVnYeXqILtkIyRK/dkalZuCexD
rBtdu5Rkt8TjzVc9uVocbuCm9dMaUymLN+LTVmUBRxo18dU/rRneQ991mBrvb4Y4
xONBjHptpMQOWVqvbKuJwon+TNNFley+NYy17b4l4YRu1IpuYIiQ+B3rghHJf/L1
yq46vUIWX2yXj1rP4MhGxZlhUNbFFB/Ah+mO7eSwfDCRxwA/EVV51XyxzE8Pbkjw
xcZERgTvbRR2F9pw+QDdy8cIbMTww+LawDdC4Qo6PvhyayBHvZqoiGwJgtDkE+7n
j2TS5CI0WM5TkQ+uo5YhZYa8IkSDsR3q0jV81tuiFR2ZwyMPzSVTfOo5zhRmIbyC
mXL5K40NLmx/LzibPeKsLo7SS85+no/JiEjX/Pqyqv36wPNgyMuw1aKu0CR10NzA
gsWGVIny4CAA2xDHwEU9Lnyl+qeonkji+N+b8+YAmj+Q+wx8tTiVdeLohMTkwMF9
ypVe3TeQTwFgEH6fY6r2Fy/bTkj6ki+I4scFta7DsFwk0TlfbVmK47AHEIvArHbd
voRzv6xzZIbWMV99R42EDgCGuUzCiiobsSs/IVzOahLogBrxhkHf8VLM1W2/Hq2q
XgcLVgUfLogPb/dGLwY6w7pChroYawN7h2eVzipg1Wn52mtw2khesVk+/5hrtah6
2EzEG60YAeujmbrK2tN+Sro/njgxr/sA9UE4v09goaOzm0B6j+5GyDHhTyDA1rT2
0uP3ceH4W/zd8NtD2nH4ku2TCFAf2Oc4JWaMjGPaOP0dHEphmat4oq25O2Vsh3xn
TSOaNJL9mocbI+WyAxF9TjPhic/9F0bK0d6UjzUOziAiSGcSnO6at2pxzDIa9bZX
yPPACnGGwdEx+SpuLMhXWzS0flNmWX/q66dTJU9pc9K3J+kHws+qdFpuuOHE2jPx
Kt4l5/Q/tfNPyzUPiL8fvwhwUSo0yJogXxvMP/zqGi6M7XSUb6u1e7iSt7K7uHmM
qaLKEo6fxj8WSUtbn4K66KRYOkdkXqkSZ9kRGW7dPmXrjW0xpz/wdxUNPL7BjHDO
YZZUHWrdaLt0F5OMXzd1ez3OYJwFa7qMLeH7q1raqYTxJF7rOdPb8xu0i/I9Gl1B
8MO5fndKL9hnNm4y821hblD3HVa9mflEwvuGWsbm3T18miTuxyqeA1hGgjDf2TSz
gKhJQvCc/gKIYsXM3lz92hmm38Y7AY7is8j9nTajihxp4vxurhhZZmwhp1tzpjB8
koemFC3KYLDHGi1Fbqi6cCnjNVLlfRxFLabJsXERjnSzhrDm45VVQ/l1S87/pJ8E
FA3twNluraQ1ViAGjde3FT36/nuwptssieLV4PDsu1DH2hqDUhG8Xfab8depmEnh
ZUSCDheMjkvwQ/ivhMZssDDbR0u+AHm8knPhDa2A/Ot0bYDd5G9L7uquDQxtgsrF
seWCUg7iBApi4g9QNfZyPMAuB6XJoMBNVQ6CkEzFadbCDRY7R8fUWbCpkKrDSHF7
UE5jbx3XNfS0oKxGBFyb2yFaOfmWAoo7P44iy17FopnDt4BVtrlgFgWnot86F4J6
XIdZYPfj/X77AO3aMGtZRpi6Ms1q/B0QU2e7bgRuWaXtGs4p8yc9yeZO2XxKRIzP
THvzitLk+tgqQQW5+hsZdRBuefAQKcf0UmcehAxDfj0paMNTuLkXsnxnmPsMvy62
5Eo1rzVPsjba/1kfyZ/+v0SKV3/Mb3eYTtZeT3QavXJhov0+pWQ+gdYhaaUZQFQY
7nRhj7/BN84OVAHeqWNdH1j/VtW6Ab2ru3CaDi+BLtx8cl/s10CwAjfHzZZYWmfs
odO/mGAwbeOvPS12UO8OSMmpXwaTLpBTWMxuWSO7N6R2rgkeBrI9bJdbxQ64r0ng
TPAD41QcPcH+IzZJw492lrM0hauNYn97h39VAArpBZHnlp22IpTOYfS341tKxTbt
0k8X3UbCyPRhlLfSv7V9ZC1eduOVP1uKsqLduyPMF3xDE59dE31WQ/nVXJ6BIsP+
JE46Zk+nB+WXSLpsvsrizwZ6ybRmdj5WAza6yy7a66d3dZOwP4tF7XTYd884XX/z
MZhrGx9T+pUjj+XJc/iSSzpbk3IzMOZoZebdAYHudRgQxMihw92ae75G7Yfur6Nj
jPwHzBseu+a2+pD4Ot6eOCK23ITpCrVlZ9hH+uSrWtGHO+wb4iQTnku6xmGv6gEk
kc/vlpz6fGcBUbdWjbjeg16bCncr1xHBc/XNrimLqPISq2Hfep/CbkQmXaKcgpPu
zgO7sD+GIWh/un7x689/sf0OjdYbaedZXXYwbabQkq7l6+nZGt3jC5z/VxWgGMBM
zedQRBIsn3BcO9ZQlpMSGymnW0bPUhX45O3gB0KjwrcXz2pwCHlWjxlqgAykzkyY
xcbN8rWusXVIji7/3+TtgJoEvyXxZB+Hsp5Ry6kLa74VM4nElghcqQ4caiAn2pa1
v9z5MxUahHn8ozZofMc0cs5/rjtJ6h7BS2mcJaosbBCmBUZRGxEJJZ//qegdj0tu
XGmfThBpdFsxv3PvutMgv9FrS8MRbA1p3m2awQXjzsmI+59wKsBChmhXTBvS1kIF
Hyt5Srk7z5SbNtKLX64rng==
`pragma protect end_protected
