-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
l4FqE1m/QmsO8hmIPooTeqp4hFL4Qbi1G6SCP/6RXZvl617QQQkwJXNsEw0lnHGyI0LAOOUk9cyO
B62H+T1/3mTItjZvUhwgUtT2bwiA4s3JyTOYCfa7WTJP6eSmeNfDKq4cl5uC0MCRB91xg41uLLNU
WbbuRvjDaNisF0d1pnYyRFlRco9SyVxFGAZfkDtceM4RbhgbRTYO+sV04NIPkC54vHcK7rFptInA
8z59VukJWKcN5vKgEb/8qvIkk4wX1LZ8s+No6M49+foIAp29WiIR9tv3+HHzx4nqZWuIdJKrEfL+
HmW0cMf1YRSTXaiOAtYrdkhhXK0HJga/6TR3sg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 7696)
`protect data_block
v/hpW43DifoEc0XsqFGEZmAzL6qnWVdLnETZdc8ifR8E2hZK6f7YtxjjTA1snrX7bzA1yi76RmQy
eRTjK9qM+B+VJ3Ox+uhK+YOgmhQvAMZT5m5QbscF9M2Cl/Ap1+Rh032FEowOBPPCnY9hjXzheDgJ
GHBEucMWLjBC53/YnPfyBy2gsVCKUXk62gCIHuPA2rUyTdWihSRKhUOLOPpOSRzzpzT4lifV+ren
VU9p0EYJIrFy9NML7yuLZSw34EDS4e9d+bJ6PQ60W2A91kwNKpPpWleNyNN2vVI7rqCm5II7Nre2
wycKOOZr60/v024QSgzoc5SpkeR7s75iF9DkwUf/rMErekT4/SnxpDbHK7sRG1Ej3FCCVfhArb1s
PxeVZQB/wjYcmTxEF+AfsRe4+IVfjbcsAoiLojB4+DE6zNTsioDIRn2USC5YuJy3xlJv9/rcKJ0m
a3aS9A4F2XAydMdDsz5bnINosrfN371HXY4z0YSOA9v8N7OZDV/n5hhTDh3UWWFgg0SjJFQh/wJh
sN5xH+We53HEYM1DiTrO0VIKOveb6tCYmQRPYSQh+qIrqxmZ2FtegDOlGNt6uKEcyXAZ87nlgCC9
EROEljoiMDZP4pKvsMA77QnbIEefU8hoJHR6D6yL7IFuC0y0HlEQ1fJaB8e4pPwIalB8seY9e+BT
26EE/jFLXFzi7TT7ioai6Z6rr0JG23J0hYeSKArtC8RTp+TeIb/0cAjuuQWAsyfrJyjVweSxS5EE
qcVhjwZS+/tEOmFDCKCZmXwThg0CIpfv6pFH9WM1Je+9Y8vDrnctr3nEXVti66K11Y893yN9+nF5
cIubDKcy+FqDGmyhQlorfYMLWWaKVnWs5g652AXxKX2FK420dBvlFFBQyJM9n4v09EyrTWEpqcpc
9tbmtecxcloRDYB9EpyMOacx+APKWtLCTLYMa523lc7ZOWRO6SqIXbndtCE5UNfWxOXaECVidsnv
sTxjhnuYTRm/ci4PkBAtIGrO9kxvV3IFi+I1xYyRTzsgneSttkIqmymLEmaCdQ8eRjX4/ddEbpfO
7gojMI57eAY7G2nS1+Szwk7qIlbzRrHXYY6K6GFv6Z0pNWPdQ2NgRyr0xLBBQidYdcig8mtRNw/g
kYlS5834lgbtNnUhXvRwGTaO7acDFoL27v7tn5x6CS8t6mxGsxT1xTm6iKPg9eAMipYMlRhekUjv
jdwsmYg3KBYnMsJ2M47vd9ERmfpbL/l2obO0Qh0T/a36EWkPZMVqG8WUqWg5jwiLT17G5FVFc0bV
fAjVd6tAr9sYpsvd+/x+G95p/fN+rgX2jqRqB6PzVMPCQh3PJZSS5S31DuAhAawqYanc7vgzxrRw
4g5REe9081M/5NX/GS0BJo9kv3J8kESyStti5hnItF+NOTUmv6+Us9qlCClpeRXCpEpYAiVmMEDN
GcjRiKLmnKkTWpcNK6od7wi2lo8l2i+8fH3tUPjeSCVNbXvTobS15bsjsXsydtJD/Sda5gXEy1T5
5ALZM9zcWweibTtXBWlzbVFQUj5Pp46qdOxxj3hvxY99VvZov4gtCfvOyfH3p5SBWCm2fqpTqgd0
GmyLhosPPcCB0h0gfNAssQsLd4zaC0AzM0rluPaiiOSWf1uUYMcXbib01fHWXGXPhE6/G4bwxwaP
GOpUNJzSqH08TsQOA011xoGfhM33JjH0awQK+qutvYemL+6pbeFXptzyoZCrZJ7KqMUtvtC3qOzG
+ycVypSxWeoyH2gcM78LUT/iEV+8RN3r3f8GalZXLaRyKZpdTZArx/B4BLbfJKFjgB7+4Q71LEAv
uyr+L/bC3ZtYBGC1ulkmu7T59OHTnN1D8qnc3EjhgbhJtSUOrQ4d7f9J6JA/GmDLWeV3FiEUWDv9
0aXrQeeo4gAM9E8/0h4QzqMGE6vXdx3uYhCbOdWyUaXsj/h+qqyCSQOjGUAS2k8KS7NPoEtEH9E3
h4AhKrvogm/r7AhajmI+JL7hYggQnZuaMrD1r9vkgkdzPAaigEEqhAuheMfpG5N8YyYeCBB7b19Z
zU+Axp8KdYklTwlHStD5py9e1gvGGDuJ62eB6zjK0F/YuRkLX0+WKFIiUO7AelLEUxvbUdDoNyv4
vfQRO4t63GNk0EfD0QCEbrfR5D+ic2ze49RDgwiczAkpPZ19LtHuOunOZT/qX1AnswLcjL82aUik
J0I+PCpFxutIGlwMAC3+tUT86g0V7YrOR4Ye8RA5Cl93/V6+I5CEzdofriqfI8+wgKDct4FIP1O1
rjSPCdaxUOfu+aI50pKUMN4FCkTv5oJpz2anJrDzt30qaCInNA1VDvmGASfc/i93u9AfgsoAsniA
FEr18fT9rGu6ObzoRcC0rdwXqeON0NlxMil7ejDu4jqRmLY8FRRBdJORmlHzMEYxQo8PtYYvr5vu
eST8OTLN9+DRoyDfRpnm9DQn+DQEbOwMemhCeyy619gfOQWOTatgCoHOv+tJNphp+aZOiLDq4W9L
StuqRKIQ0xk92BITp9YgcRL2zAtOQW04id2egUUbMASzWsYGpI8wswsWtDwknl3LD6+ff/1ZAT5h
TCnqhkXa+a/NyjIe4WEgB5P5rOPhvoaZ0eqzLaY2kK4JZn8zZPWBN7FgVa0R1PgwD6xyytBEiRY5
D3fLPqQi8NOZIfR+/HJqXLNUUf7LEEQPDd2Ot8fbOR1lqRUljs1qI5LrqvVMRiUqlmXnkv2uDtIr
SDesUflBo1qCiiETs3q6f5hbX3XnZ+v6GCQsiTRayqJLIRulpnc9vBLgSq/lP8uY9MWLPSW61ABM
N2VQUVeL5m1W6BELcuetYelkugKYcOkXqxrAXni2MjvLmL+LdKTSVpVvOLKcayTLuD+ctbrmP4tg
x5jM15wgbEbau+AQf4nCmpZpt/PjnHfHxplh07qH+Oeud1olypOl9QCmyt0tGJ2ggAOJ087S0+cy
Langc3puMyxVe8Yd5tkaNKoKfNqHFgka9Tt+1nH052YSt83y85LOHo3KeLDnR+t8d9ppzY1PXj9D
WhGm9eLRm6nylKR1NNYcuS3RSBC21AtdaNzr/U5xC7PveLo64DaCBNE1jRjum82gwvbr0lQbji6c
hg1bvaP8XB8YNVvigtZ+lmYk6pj000a5tVghlwH2ja1sdjuwbeuyFp7wXX/uGDxNd48aNr/wWAdK
tJhWNP0lyA/GIB/wRs9DMf+9OFHT+Gk5+B5dLfgS7HSod56LjSGf9Uq5K0/nzQDPkeHjk550aPCM
oWyvaFyrW9c9T1lk6xo9AheKhVzXnD1O2n9+pfNBTKCEYoW76/aCDHNEjAzCnE0Jdlapt0UyGka/
h5jzfDaBQsWV4jsDLms3W7zut64aBDnIZ8ifJUa41PGX4KAprjNj1rcCKzi4puBiGksqAaHTXCCP
No2R7aI9AXIF1xDMqs2ZR8rW45d9M4oBwz3Pbn+SXdUchue6dQhZ403v9pxb7CKTbemmhwy7UULk
2cLhuoj5NhY4RJsGxu9bygcxyEJLKZ1I+0n2xmwODZnDI378dFHm/M8fekiJZ3ZU0oajuL4AG3Zx
yonzbCJHyKCk1thhS0Bf6gJxhpqaZ5e7sbi4DsDRmy6S0Kfvu/p3OeHRsDDpyOUBUILtCOZvE3lx
LtVDQ5pxhwyhr6VnKr3QblKE8FvYLprVJYhrb/XgViXBnGE3vk2bT6aABJpVY7gjCAVFrWNo4kFE
rzLUBmWASYYxEznENqRR53LwGbOCckXLGfWZ1XIUrBMGpd8KI7W20va/9xHOobdQYSIW/1EYq1dA
aOlEiGccJCfrg5YNvTz2fCW4L76g5mLjnqOBPBZAAYroiNM75/WShH4S1qQCXwyMkRrvmaA2ojRi
JyFcsiW+hd3iVUnhbvIf+/cyC2WOjau+KpaVz1Cy3uz0eJsYLQuzTEN/qkijhCZTj/qR+b6DFJ9j
/fsmYF0YZhSpxWZ+vG6O1y8zn1Cu5PX65T9kft1fxvCqFlt6t32ivLUVxRwEuJGWwdmyuGw6A9MX
/oB/d3FHwUPCqwKVBQ59/xvYeAAq3heJMmGVfDZ1g593Y70mBUoBFihECwLsMt45uG7Zhni+t8up
uOcGM1MaVIsd5b8qpzI1Y82Kl4PwF7wkLX90+CnTLLAjVDlBGBWLeGdNXYVNl8S8MKIt2vu5/3mq
GJATjn6UY4IhKqozQ7mMXyhDPNUblHGwOtsKrOlI8Kz+uNy2LYekqx6nQWm/Fx9KOf0cB1gxv/VB
Q2ylRuE+od0JMoHo6xeZAz0Ksgc8PeGpX0f8VSZehH/3iIUuOM4UpwEMhCX7HPAyQywLklmSImtX
OLdCbEDrDkjq1zktAn2FrO3KS856YygWk7pcalNfdYT1K7MLx7Rfrm/Lf4hZ8qHRKn8CJVX/umU7
jeF3nS3irCdWxzdteL9O99Nno18RRFmIiSnjt0MNVJThqdkyzghNhPXW9frjnGIRdO4yKD29OHhr
iA6uEl9BPv/k3XoYo3VLcUuoexXdzFD+ecUHqkjknVsOP/+qtFO7lfozeX2cOb1+w4bnd7srWxvu
zM/QL2BU89aHg3j+hTVy74ZIqgb8PkT32OpnYeNBbaEiYhfhaXfgeYFwFJX+u5Km9rL3wirbwWIi
qXV34nIg4BUxbpPVRP8/KrXB22ttKjaCg/ZPF47qd9IM7xPfepdkZSq2DmY5dWHgHavzeEwHOiI/
Jmqj5r4Wjh7wuGot8Rs+wIo/JgBI2jqxCXOoXl16HVnSSz5WbxxmF1Zcn6B8giqg/xjb4XJGIF5b
wX//UxrQo1DnbWZ5mBUN3vfyJYIwYxiuawhHPqBFjAqmAg7GjR5NUhpPa9ug/az4UJwW2dJvXJB1
uScL+16EKQPtkTbd4QjcKfV7UKI5O6+3LXCJoTNY7q+glkwGkESVKyi/vWTPiaebbCPbrjSwxmxP
QlboUyz0rAGzGx4JeX3/u1l6McOwS8qMYGxme/DVZvF9Cc+PxFDF423bJl5A6i67e+/7op72m81x
e/vkSKHht2/1WY7dDzU2qlozUalNJn9rriDrxjvsTH8XQnx6YaNNIrSbn936nmUaLwJTr546vwYy
Te4JWRxuv5hM5APM3IqCJu9yOCb4d25OTtPK89pgMwTz2xOhVBXwT/nj0luESHu8ihUxmczf5Rs4
GHD7FE1jfi4Xejt6K8/oVXLVd46fW7jgVpUTn8Fjz4PCuD6AAQzVptqmCv+E5lL3McRmB4oW5Rkp
bfUe1gbxsYb1o6nwKvQd1UknwA4dPDSzWafcxXO18f1lhYMyC74Ix7xaFFc4YUftG5PDHASN+LX+
wHdg2x+Z/JnltiJGI1QaOom1n3aFhNU/qmz4DC4WkBEqhqQsJa3h2FyqNbZYt9Un47Uyi90y0IzE
3qO6xH8fALqZP57Eq9AygpflKpMppbnk8WqKvDbCvfFOv28gKL6NN67I2Z1wCuha2m+8bGyozONb
9yXHexmBycPqXb7rKvGw1CVAA0XaNqetwTB+LIf8p90bvRSPgG1uhUlAAUMvSOJY8jxM+46blX5T
7/5vtsAndnwA0zkpfqYw3DwF862a5F1iXyL1zuaO8mNQ4mlSCdGG0TgpN03DTLFomJGOxUD0Atrs
qjCld9/n2eK6Bfr94iJ6ebx16a9Ec+OvjLlXuGaj6LgwnBVd5l/JUyVBm95rX+6+4/kg4eiKh1Ng
bjZDpEiOQ3lZKBM1aIPDJB+NyAUyFWsXM0OjwNGR014E13alr+ViiK1+O4r/rmA0iqH9DvjC9G88
bcUG1P/TnDG7AjBzj9MlWMCQ6iquhbxxhk3poqRtZZtas8ya7UgA6e0PjB6eLMmtii/+4xBTZpkX
rOpsBZpOiP1XGHphu3TdvoSNtZYEP+t8o4o8bV93BrGDYGGFcVE86SFMSl40DMe7Axdrdz2Q+Z6B
cCE5wUK7vweHhJtEQqL4HUJHGnTzvbexC2iT+sXaSNHrjgqCT4DReRZu7pb9FJsrEPj1SwXNuL6H
SAf3R6vVQMH7ZgZdZmTfeRc8/NDMUIWtF6pZzey8j0EvBNs/oFrjyyfGCbj/TDBRFXy8ItQTCa5j
v8P8lwDgbMJ5Jakp4ryzTYqJWFK0rD52gXrAgZCnR/7LRbxS9Rn0ucoyJltieXfFoadgz0aA9DV5
HOtn/Bmng1MyH1ylYUJqFN2pJbnBCI7/X0fzJ0bfgNYwcG+ANw2iUy7pdTgvpApjjObRGU1pE99y
6nOyp2tmomUhYJthIhTOwMdVYJf/Kf896c0S2mRmi2Dy0XOZ5+/35bjqOibLXnsa8EJSoEUE+Vf3
LQkizIv028gZkmv7ci9hWnq/jLDOjE1mTM3GwqSYmPr6LODPTi37NJWRqdjr5t5640AiFx4FCUm1
cXHja1+O34UilT5lhobkEf+RXePYbdfu6D28iigzS+VE92SdjXh//6dG+8mSyI1OIEiiWYerZhZz
tjCJdht7KcmG9FVHezsSanKr3l+o6sM2Zk2wako6fbpcKX7UbwPqJQ+DEVV6DeYryIUmDf+fwL66
15fx0gR2whJDzA4TlOTGrX7nkw6PPz9tUDPcPkcL7aShefdwLiptE1O0stCmRuW5vTrpGT3fZ78s
t7OM33t/BWX+7Xp+FhLvMj3Oh0WaVyCrUKPby+9yAQ4d6pgyqSkGJvrQ30z/QFIDJ/GM6Eq2JfIl
sx5eP8sqzDQOTNCUMJPFdkYql07GVsVQvWBGWjfffbGmvc4GMk6kVqxcdDyNu2K5kfMEA6LVXOWn
wy+XACP6sGo2aOIeSU1hGdCqBB4h8p1NcQsD3/gbk2z8A1ZZl3LRjFuG37YTyyG6+yVFCMQz88Dh
6GRHKYUfUBR6vwjMa5uSrrOrwhUTtkG4Z1xCnYANDNYZUkR87oY331z88A0QuKK1V2/BWfz32HjW
ssADmmTL0UzFgZ7WWUdIbceQw95PmqEIwowh9OtF4uw+ZMdpRE1Gmtn/WaHZ0Z+iAbsVS8Eitu/M
OI1/oTf2PJsI+mX4j/zGfDMmLSp9TEBscttVIU/aHgXX9S3mYn421wTVjJksapf5173gc9BsG6Il
XKnVVCKX+zsP5OS40Ab3HbdhbFdbw0NLZIEvty8KYIjrZDTrOFSa1q8zSAzC/By95VkJBE1RFNlJ
tZS/D9xt9r8TIRkLzvdB2MZirPLnSRRaNsunyMfuOlJQkZPXrfqS1dY17j0CCqgnVoJ3TWCf3UOu
+9QI5rlN/hzlf/SPLcPl5BQBIAz/hO11gDUmVRfO6v7uyV5eJSrJf3yz8sh5Dji0+4us4o6Xrvgx
kMUZr9uv/H6U2OMYsbA/Bnxcs/on26Up7yKrTBshQV7IJGFf9pE0V/VXO+CXzYo7VeQIeh6thG/h
5Niei+sI8xDzX0++RnC0+Beui3+OVZBTUe2tzXVL5UKOzOB35H7tJb8P71K5eiLTXDlhEsCdohil
8ahcUxvZQRYLn6aIY7CHi5pjiOnsssFIuWRZ9YnfKBpdCNPSo+BNTzrqNMDz1oYWfghEZ6+l1Bf7
Jn+iWJskw5R1r4/d4qZdEPOGEHfDoRC8LhOKZVR6Ydb5K3g0oYnlWz9GxbEJdJW+l6fpCUnV8kc9
SWCp6WrJjmgx3oxO2qceR+5TEp2z3Kp/B5vyMFYIu5xa6TT9MdWV7pELTMU7PwxQwiimBHvgICg3
evm8fWqrBcLgBKGZmAnYEbTWIClNwVrH597AixWW5jDn4L99l8xQ4CJwUtHN+ojV9qbNms95EGOi
mBr4MSQMQNnQ20BJNnwPN2rU5rzBZkMDy3qlwq2eONOfEQeKznarwJYQXNo2QBNZlrs3Drhv2J+h
E6D+d9079/b/oA5TCgzuQg8KuN/1BCkCo/HNVqP2WjT18IWtQrTPmHX0WzMdF2cBhcsvu+8+RUmN
/8FiromhqRPJgws0YT6oeyrapB3AL3opeFiUhu6xXwQ6bFOWf1rPtfnaJ8hqQDi67CYvwNMDM2Qs
pgCFf8+uKC/KlbK9C39g3HE3JIZbmtq6I+4NWgHlMM2ZQZn2XWUpkr4Z/KVL4K0QZx+b0sIYWILU
io681u02L+a84A9yi6hz3Q6y+p+NqcYws3Qbp89l5Hu/EBkHpec6z+mTzJvRuC6q4onJMiXiDV6p
/ozou4odgY1Tj7VMvrbvih28WoPX0MV7PC1xiCC6Ita7f9s4NIn9eOtc0PdnDtV8hW/zyL6lCoKn
GeNCAphADcxMnAaJ0lm2EBRtD1Qubn/MWcSKORyQoPPkB8Fgx0uBm/sUaZAn271+YJrlTSgWDHTM
bIZfCY46gFx+YfNK184WTuI1McnnebZ8f6toBiEfAT/GhG3bwCmiVB1+bClbwHEuv6q3j2DM0+57
kECczqZHbomlJJWitzioRptgV8wQM9C/tcSpQY62UEUQ2SInI1c/roVLzrLa89pCBWKByHNBd8iA
TvLMIJgFhG1UGCUJFH82yjBWn4Z7LcX6KC+wjU3H/VE0yf7M8rmtMrbcafojuwiPCh5CzUB7RU36
yeKtzx4U3AA68VMxJKBziwEe/41YETAHYvVA8dr28mz1MS5iVlUbH1pTvbihcDzEHj/JpEOryOiv
qV1n2ulUm/7xOnpLj4UufDxqFhuCM0dLN1w2FbFCjh/Yc9UpADMqyeCj1FaEzq8/aE7wVGYKhj6Y
LffK8rkhND+TsVpZCoQ6n+AXSZ487+wwvyAMcBnuOiNvQA3pLB6/XL8WGuAz7fexImX72Yf3iGbT
fvM/OJsjcPrt3lcA1FfjmSNYX983fgLCT6lnrz3uuQyQQpnD4ru6O3PBvjkupIYZJHe8kCRCtiBB
rrc9cGfvjRupg2KTx2YF9zrUKrUoObWI3h3flmFdlqAkNBFQTJfbQyndNrdvLyh7xhz9xsiWwkgN
bktpMFFR7JUFV4gOC0hYoiiyb1k8rqpqF2QoyLgiprb1pT7LsC8x+PBVVDHdZf39ahe5LgG4tTcT
s+k19SIXk84/ndgnyuxt7OHlUbr9ZIlhaxFtKk5NyFXWOHKIiDaDlI3zfk1A0A0rU+Ppf9rXP2yU
dmfE4o3cjrNXPq3WLP1jjYWAYzCl6vx+m86XF1aOrkxScd/8NfeEziFmnECYqdcWrFoKHJRnD0Zz
vCO88ow+T7lobOkLtrKYG9e1wDe013Q1WA7ywU0O1Wg/GYanNwFCiViUpZqtPZfT6wx7+RzCArUn
jd2oEO3i4yEJ93OpAbIaVsz+LqQVPb3auuOi9rimnYATO20yzDNjntlgEFvA44n2oXY3QFvZ0z0l
XaxI9Rn+MRPKuq5tZ4AjAcoMPg+G2QEg1PXU6rdx/fm86OjgWe23mvaPAQARDaZuuXRVOk+7dXtg
17l4jW5DRBozkEUSf72pamowQ7bST//YJ/DD8LOwVVI8vS7MUn7RBFwvSKvXG77Dq/3ghYPSObjo
rk6B9gQm5hHwrfpOogKJyQK2rPGwqbXbPABTmqIsjVEe1v+Z895fsgrzsbsMAF6vMlZW6j59tmGu
XSl9Q6aTjESLA+S7wjxUDt24Kb7BlKdn6P+Vp4FDqLb9BdP/gebtjzZ+AwjZA2h1jso1j6IRFGxs
/szRlT/Z4cPJxeZpjnnMxWD9JED8mXWbOzosQRiapTeHslU6+y3/g+4q4rMK8j7o7hq3F2IX7QRB
p4bYTOpKmzMGEV++s+8UeAL+6cMk+Ky6KlWDuorPdllyz45ku0yOXrE5SMHzdoES91VRron1snOp
DOgxOcjTNooU4QuK1qnU+m9KQjVY93w/Kqrv/kik41xVaCAtQ72ZdY5l+ly/mBoNMqIm3C0v6L9n
wz3szPlXvuaWRBy0XaXqW1j3kAGVvSi4BbxF7e4ZaxYUB6x9PULBa2TyZeCtde1A/OEtwIKhqx6Q
9/f2NEJ3Zxev5tgjR0XEAXiby5Ba+cYtTMgJEEAuaj0+3m82UFZbYNvBEPqQW4hGLhgSIov4/Kf2
R52PcjZi7ovCY8wab7QbqvaxAtxYgWbMmJOUpRM254f1NaAM3ok+oTSgaPhWqiQksISwki26kmMg
w78gJYi15Ylr7Tgq/WPnwCvxCsNgIwM33Dhv2JjBstbiHsiF6lRq6RaAo4WN9OkBPLEDMGp+WcY5
8NEhdKA2aznwgBArNcndqGhaO++++1IrrsqrkYArtgPQk9nBCKfOUDIWtz21givoNUqIm63wY4vK
kIVyoKfecX39hKWCqQIHO4SEsbvSwUIFf+ceDIuBHX13xp/g7pJVZz5ZKuOlVpgRCAsSi/GIZHnY
4g==
`protect end_protected
