// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:37:05 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
TmWDTDGyw1ZYdzyiSdv5T3xPmFPVy2sO3bEg4lI0T+Ab5dRT/osJNtmaAxePG/nC
uN4U4fuKKhcmqP3pr2zj8GW6b+scaMShDLz+uOtkMWE0Hr80KSrKtIIP03Pev0NL
pSauaMesHm6WOG17kRihEzIFeaidxoTYT+HEWrD216U=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 22912)
k73ksaEOWm8+qMqRxKGURYx6mesbUT2Mw/i9leperl7uXkaxnpGr1cfT7AUUMP3q
hfgkLOmw9oUh7AuRBD0zZsqfhbwDHV7tJ3m4aDB0dZXn6PJQ/2/bBnDhvQrTZI5p
JGAHJYbzNcq7Ybf5It9IvBNxMlQ0QfAogGynabTr7hFi/r/xRM3iX5Y/2m3Lq2U0
jXUt96ov5LLXbtsaffqHUqpFouJuvAPRSsDHWA5CoOfsX2K1ewpGb7uRCjP6HzV1
XWVSybl0z9nSK9UUF9rAhn6AmMZlAwUHXW8SSYA/8VYCadKLaXXYdWfm7t6xazUs
ALRoOqtrToe6Mpo8jD15NB9yJibNvaGQeFymroxvy6dpjDA/6O1xSW8SPRVqgqcN
SQkafaAf897WT2aTpsh3KieglqUZpztipGH+dn3BuLR/bBda3EIF8znxyT4MIiVr
TXaQogPcG69w09fapuPLp3grLB0qA5x0Pdkxtrt0UqumxSmZryiSLvq2smbkrQi9
ZDiaf7erLU+FGptGWBGuoAbxEL1F2x64WIX4kq+mpN9VbZ4ddpoL+VVM9TFMAX/R
cuol9Z90GDZF9jxrz0tunXNwhETamAhW1moHb+9duga6YehrlhzaKXL5V6HVQGFH
meKFTSIce9iGHpuI24B3zEJBHvDUrrMGqMj64YbmmssudQiy74AWZIm28VvSuMwg
VjyDTPgaU7bUM+UDIeMX4Wfku8Ecf50tRdbDcWSK/DIuvBBeEbYY8vKap2y6Fo85
d+h5dhpvk02lSoaDse3tpqMzpQWV8HfzoczRWLrdYwM3H7A8Be0hccey8rtxcQn1
E2jO1XSrn/tbqvUY7Yq6FyAH4R6nZKfgDnVKmbzkE1ZC0W0eWr5zotrYG24k9RNr
pT7LSECM28pXTe48u9PbCk2Yi1HGOZflD2XZ2xCLDEToVTmBQFpyWpQFUkKL4o04
cudMosv7SQDF8o1MPVAP48pwb7FQzFtGtvJHYwKQtK1lRUAD/zbZAV58JIqnOmXj
CMoSqq+1RxCYS+AyQHEGjHdH/OqwnLwN7ubyVn2cS8JUw21n7RrOMkXVC0JgpxBI
uieg7jKYJ4PQTT87ZMAxvrxO4cHNp+4UOi/7jKZMDkD6QarKhur3u21PO6X0nFA0
lpoicwT+GhVYBKTDIGIhgQb8S5tSdyFxLkpCHFsTcrgeIPwv1WD/kYpNfWhyXNHj
SAXeDLfauTFrRS5IU/k3z7CoOz0T2leE/I0QkmjkbYfPQi8JVW4Qtf21hIlBznJH
3kHnuJsAPX7uuFkNXqHxnfPEsxR+ymJIQ/wNQYiZzv2BJlQDzvALWmM4N4MLhCNC
cUBFIfYmA2WWfCwOyXiRIdHSjgizTnv1AiSANunMS3xmCmzF9mA2Vv7rGydxgpnY
cnERK9bz88xsgVxpnWJhi/JSUcqHfAuckvPspO1ousCdtI0B5QnGSKWyLSMJLv/R
kBubC+7O0xc6Fc+zKaHgnMbfrBz2m+p5/TyJ5nMPnD2bjEKnZzrZD0HRBf4eCO3Q
YrdOqwkK6mNai6eBMRYkUS+DZq1aeaykw+af4jqgrnhp9ozcodl06MHHc7/LVbUB
aunCavVS4h1mAwfgcnZaO7HjHTin9Qd+DIWAAqWgp06o1xNHzlrqPDnfaO6iKfTR
mQn1hWB5neEsZTNm7/j48HSdKEvUneOsLKQqC7kN1yOUP2OA0bLuuVxba9CdncP+
DwoyxG0Sj7qOxq3PfsmbEoJMiCxujJHNE3m9ie08ze0YchoZ7W5vew5+Ie79iv+3
I+WPVsw7edETmHp6XqI01FLBjh270DX96WxvMSTj7PWDzdqpePJ5f9n8zduSHlL5
sKnOI1T8jcOeSbixloFQmys8dGo5NHz22fJ7EmNXVy78W7vWysCT7IE2pye1lT6z
jyXgbA8aV24hUnUEgi9ollX0+fmYIB/0hrLdUWc1ur7K0fvynKBzPh8W65tA+k4e
/P5rfavKTUTOejxoOu94TYhGpK2avGj9d6porVjW3u5GgXBRbCzW/GMFapWoBXOb
jTkBzdP8DSYceKdrk+D4hsfVj8dzmkESqAVPPMbTgnDdYCGN4baVQmryqG/Uvn3d
zMejO6qOvqWbBntfoeCyAs3Do2Xf6JgOCbU3PRzm7RnWA33ooxhfCH6qYtXIvLMy
T6aagrivoo8WpH2cpGbx8QfU5LQ42aCM9gwfzSjAymVPnL//J5xhoeEOlaJ+5VW9
fdD3wz7ERTnM6oKR00Yb4OxbIoXtqDc1vMqhfA0Qy6L9cqyQhVv8wFJVSTCZeq2N
bYsl2gUHZ2odQ/CEMfYXL/v5JnCnMjRxDoTmYHPfKLYsY0f7j+MHrIhgkV41t7BX
duKHucNjskXVfk4BfdcW0DSga+urtXR/5D5a0m35VCKIO7TArHwihZCbtMJyBudV
e/jCT7NADg2Uv6Qco/Tm8CaldgOnRynGE580ew3VyTNArl28mjQxCZ62g8jHiBEq
rUWrdc08towSEVEjdDFtHBPnm7X9yoEffxAEmIqleT+k6JlKqOPBwu7cB5rgdNsK
M6w6tyskxolagu5MP6LMGrkIqD5XgNl971MD2yAGWKJRDICSkTXi43kyUyh9qLk9
5eO/FQ5HuI0DQufi9ZIQUB578utnjOaVAWbXILQFWd1v+PMS+LOorE5nHLCWAjiO
esr0fY3LOxLkwCqHHJIzyssC/aQxjaZ8kNHVBCPxlUL07STe0Z89otvvWY4LCIRo
vkMn3ZI78Hcrjk6J54OPnjC61oHwYXzCCq2AEOj/4rmCnSrMqqBWtGVHBG+MwZ5d
VnDmjkhTStsNl7e9Uq10ZFtVncpQ3z/Muij9XAjnr3oTlegXGKb26eRPKhzkktqC
paClWxh+Fam4c4gZGNZylPAMKXIgCNGy2azXVdDrj+PUsVEReUHfgRWceovozXw/
LNcuVmZ/PRu54NrpBrn9MK6umISVaT8eoX+oi9Hckipj22C3/kB1VTlEkGEzKZUz
y78HCUF1KemDghsGr4x5RrtXxZXUSAw4dr0EjdBpQM8H7ksk9rEJpV84QJIIzTPm
LYco3/HlthXUlXZqCSpaSWqS/ZdIqO22yPq5pqbTr5CATqEHup6LKYNLEA/fODbP
YZ3dxFwpIPp+dCm4x30MxSCfOHs9XgkQd7T/iWo5B3fUI3Zgc7bz9tQ/TaHGhbEm
UreOHNI33DC5fOMxc2m0n459ujsF5XjG+a8U/9mnWRB9Yqh23kvi6qnbwli7tk/g
aAvu0WznwHrUX91pgt8CNLRnvjvt4WtSmR5ZbIlfuIZA8IjcOKDbiuzPZ0Jl/ogP
Sx70f41d9a9EYLQhlWFI9PAxs0EEybNyXb2CUdVWkDPGDmyUYckoSC/t50BF04CE
nv19rTP88sOKqqh2fJs6M3Q3rVLia7Dq1WOe/Oywmxu6Ypy7xM+F1VbspRK+wxxU
gO48a/dh+LpJdbM5NbU4Dx3e+be75HVc+t1a1NRVvIsOhLwAwKpQzqhOE/8rqIt5
Aqe0QoNBOg9MLEcKV9PQtH1bb8I6SAf3TKLWts1qvV2MiuISQNxeUR+3uXzWyBgu
OUs4da4QPpApHYoedbeEh0ISc4uclnmbY4tw9BvkDn+cXcvippH1znsXeDn8Iqme
L2kBIL6f0M3vsskoXLSlP6kNaJZe9beld2O0QsIY68IhpoiD4CVJ8m5niUek5OPG
Pv0J6zPc8hZiRW4TYozfCRSohb6bZ7N0NxJYrf/mFl8oGxjxPLkz0IHS1htT5J0+
X93XLWBSwlw+s3xItgVfTPj+cQRwJlWlCPJQmcjYR45xS1yYJKE8S7oHezP3peyf
GVa6k+tWCA4lBsHCkotDrhUOoQOrJLy6L8GsM8LtvFCm8a3p/+T+VYONWTDT/vb5
h2sTI5RAXh89l4kRN+vgEjEm8kfdr+YNw3+uIGF8WPZ7ncnivc3C4rfFel6Hk5Bw
hLsoRaVHU1T9Ppphmg2HEXjpg94H90E14Cttbubr0OjzjqPau9jzd05dogBIZvW/
9yI9sEajb0Lf/bYJwig8kQJ//EQqJPfrNSCtfgl9Ic1Rnlr4moHD/N750jNO1us7
ngakiwgaJkSxwuMaNwm/Ht+M9nQUdWbFWbKphueQycZ1PBg1NfTwjoopMcBQvDjc
q8Jm9Hh6yHBAHS2HVhRUiTPy4JzWmNjKHI9A0yS83TTRC1OO4WZVj9Klvf7wyIlB
ObWlt4YY5NucW0vPg/39UT0M51IF/WP8rTMRALpUwwZ3yRQT3yUsZnilVy7cgUss
BiKcLSmCEolQGKXWsWR+HdDvC7vFWTPmhGeH7KI6RVj5slHORT8K6WeFDrgoydNs
C+VYMBwSXGpl4rhwyH0nyOujJFzRJ31AOblN6QNsgHY6iu7hO61tHZicjIOi/NvP
quNf1ydIsFQ213kAgxrJHmWXmQuWESTaa58bI52+E6y5IwT5R9T2G+bZ4HlBouEP
oSonXl5hvGsfbyiYzwFMYZPhW2Z2Iq+HtXC+3D5FmNY7RYcy+k9kpxIUQRo72jMR
Vt9RJjnegZkAqyb/2Dd3wa/aSuQ7H6PzzJzOxlK6zJcuYDxgXuFmWqqWvi9htcwQ
/3mWTXrzZt2ETA3S16MkajNN7mITI8RsCeSEd+t7ky0HsC9jQwC8yI+CZsYKzRPd
0/b85hiayWwnN6o3mC07TGnbnW4YKjAEwQWILueELAt0hW/6pgafxHqQblhwo1CU
fdOQ9uzycQkQTzZQJ5+buW+hEm5RZaDghp70nwvrZKVhwNunT/FtPcIql9W4quw1
n3fobJNQiKL6yoV8Ya3NyOcq3XeN9dbNuCpDv3vRx3/xBIoaHLHjH4IojL2JFKna
c2zUVitZDUYm6UD7UV3mzaI3egr/VtXrQ9gMuUQM9h1+IYO2e9bp9LUd1c80Pd2F
ZtcakUhdFdbv7Y5XVdh5e3g7ch3tuMBf7cKJXod3G9EOhOPBVUEiz4Y+SdvAW4mb
wYTVRa6lL+J4b038xbGgEXOEUYGxwkkZ9mr/xeVm55U24Es1eUkbKTd/kves5V/G
Fn9vj9C3K0pLWlSbRw4BdT1OP4+WQmzCvxhSpQhMMK+57RoU47brs0Fz1mdgldke
Jj97Foczfnhiv5Km8TITRltjN5nIougmN25ClQgxaX1m7TKcJ1RHAR8fo3Z95xjI
V8yd1plSHiAJKfTLYSvHqLjNo4VCZkpJ4SB22ItbuHhy2vn7eG0KgADH4C3T+qZm
f313AVlfyVXpm/+rFaNyP4gxd2M7b+w2LMOJ2H/axq2sYdHyAJu2cprtVf1MAVCH
AJ7XDeWS+S6/4Xv1wd6tCf21Sk5G20b0zWKySf6dFc0w019UmU0N24wmIQq15oyy
hXsAes6ZrYJtWLgVC6FE4HNKgHJk5jld/s7JthBuj5a7seJG6cYgC5ab4LGTNGGW
SuG24LdlAXuLCAijaQnr+X0OFPYWu/kBeHW3MzEnZ3NiyXiKAaJWpROZ/DZxPYvj
JB89Oe9yleR76yo/J46/UZJqZdefh3hvCmSYtAfp4xBIrhmoGu3MmYXwLR5/LXEV
reukIt8LwVFSrkXzxuMokn/4Fx/yPXcWWlouVQxVMR1sk8UJEBMwxQkh+GTJPQ8Z
xARtFBoTvbwrs+5JvxpO8NQErexy5bFd1Wp1ngGC+4+fgNV8MgYstzE3M2TgMZao
P5Db3BG1fxX6+dZxdggSj8I62AIkA084YuV23Le68BFkFp5hVKjg2RWFI7fT4wdi
vyO8GfdXxkXdyWMqkT9x3EbOgb2aRAbd+kgaHfGXOsSSC82TfairOl6qrtVeL7uj
iBS+AKTMAAA9xsxp1QJY961hsKVW7EKsSCw8yvAKDKKkfHCHoJox+wVRXPGZAWGL
ON1BTAs5e7G3YAW1ZTz9kIC3qWLvtYiHXE1ruPoH63s6h9aK+Ydw0DPo5qILncsM
u9jFF+5lmObcC4vDuSF+W09SyDBl2Mt0EGrn2uq22hQjC9VItUx51jwGGk3UDHN1
miBaGKLcGQ67sU7PvMWT5nGFNR3TJihbSMESsmZnfs+ZTXOxAnzNl0jaq9npClCA
nE255kGpKfZLVcU6/dyRO8wJg1D8s5AJ93MXyjQjOozpaM6QIi5Y6frEX4mVTOLX
aoQt8ZmLfeKcO0MHE02sPfwnjkTf+VLhQPcLE5V4siCmf48tN7rXqXnsyipx4uEY
uae77Tl/LZk1bBzY4aT8hKEUj0aM0i+wnHVLdKo2U9iLRPyuS7OJXhJKqfhCRzX1
xYSWOe62zfKoMMX+9ZZr3zjFlVOg/qBwHwaDPAASzgXvMawNJmWGzPjZDHn94LVo
xL4Fi7FOkZhQqzGIONzNfxuJKsyRBqAtpeihxc9RqnxI/N9La/yHurQq7oTHd2yN
ZBduZ18aiCbaLQriFgCBiS+11weVCGIiWE3qPvtDRsy2UCzzlSjMsT8KZ8y/4FNX
YWHhlA0ixu0BJj+yl7C18s64LzaBOjtOdEX5lypQD42ON6Fokle27jirM5uJQX/L
gOZDb7ZO3b1UEarebEuK8d80aYo4yHkilpaQZpyelere7cgPfmQCx6N8WF3KX0ju
e0q1/yBQtNFeUrFoyKuJExoGZu2gzHwfBQ6yNzh0k+xP3LQB/1yOeDIIM0S1NKCB
he6yQkCc1Ff0uYct6fDekwGsah1oBXTtdmVl/lBbQM6vYMMAdXex89xTV/0Wj6Kc
ymITtHaWPMzU4YR4QTkZxpfqcKlkRWh/GYmGJ8ShHZrYYhD5zBIb1Pu8DyjGJtWC
WYm/gohP0yIZ7LozJvD0Pqg7Y5BxUJaR3AwlK8m0L5V0LHHn6YZ31AcQRltMKczt
MtqX7K5THt6YP2Ee/6MlBnP4Z5GURQpvrvN1Y4BVtB1fwoOaWAVsStz8fNzcy2Wk
rRZa4dbETURXxlMzToYr3bGQkonl8sb7/kIPFQPpT2fg/jVuh4G3Zue2JoD/DQJ/
thGTz34K4ZN1liK89p9I4tfUe8XnW3sR/meB9VKYQB9xjQWMNx0v0H7Ak5QMY0j3
I20ARrHfJNNN3+6FUdeQZaZshhz1kcVs3MT6qn5Yzvmc6YgbprP5HHNTiXVE1Eb4
8A3mGn6aWogbBI5uXkqp9nhkV+wPN0h60aLgaS+eICtHe51Ivs9hNPbiDTmWbcVa
5126APAhpB8i7B0qAXt5ZuTbi1SREIgeyBB7zfb9NEyRwAccQ+/g9G1SPn0OxDFr
4H0iHuHu3cCyMUmwSBtnkP8iD/vnpnMlFalsKYD7Mp7lGlPXxsVPcGncbgiHGIy6
euNW2oy3HJZc3JHmsDTOlXN0SBHnAXPEnV8AYsxMmC/WDRYR2XuMCbH6cl21IbsV
VJ2zCDWTTqXeJP1WR5H2lSX4AQZ1tcTpEB4IBaubdoKBhVTP3uVbN2oLVd1lDDwV
N2MRltx/eiiXhjaxsGYbtYKrPjkRcfTZZMG6SUKdP9f9UacZcX39V1qqF1VN40Y0
Jwt3SB5MKXeFLcyI2mZTgVu3XwkHZ1FcjgddiB+E7Q0kiQB4SL70ogjyULzFyKVN
RzQtmmzjn2+TPsCjhPdJDN9TrCarBS6lUF2bTtNSk22U4Hx64RfMzgGEV1A6R1o/
YJHmu6s9QaCcOcEIh33e3lLy02HyfQtZn25T08DGfsj2BdG6pVXkw9N5iAaN/4Cf
qqwDKY1IaLK2HhQQzCFSxv/apWaPoNeZf2uSZTtqj1GgJMHfimIOFeRyfQ5s2QXu
hODLOxw3sG8ukWyFzGmtmMUFdW2v5rlwPqYjPBDgNGjEAeq/SO+5yo991qRbuwjW
AZwfDkgnFzA0ZtDXwCuSLv71SSNSX7LTjCPneiNf1FBPozDRW9UGL2wCcLcGix3K
JZlzSPQTpuJ/X1bkTXNvNG/IUJsUGDLrxG25/W3NTOc0pYeGyzeN4y2N+vPNNVF5
0PADJLvbKxcirfr14NFSUsYwr6VEaOE4e0DWYT+qfySnBMs9NYoCJqZS8GFHVUyV
PuzIb/al6t8P1E5OdmoxyLTuah723b9IjaK4zFj+lSzd8uE5y+e5FLy0fGEc5IXs
46tZabWWcEDR4OqR5CDSDQ1SQ21Uqm02xr6zuqqI7krNaEEZ3v4NzzrJR4I0QHEU
NxMUQw9fFUYmMOXDEvKsNhj9CeXBQepu+jdXJgAJlfNp03D9QvQOviJuJm7DDhhH
Y0tF1+EDZfxzQHjVFlDAYKgdZUBKa3M1v3cuky+jc0aeN6IsNoLbkkfzfofIpxC+
3LnDZRUInX+2LlRjD9ZkeGA8nJLmk2OzubohG2y4SqXCZQ0pDS9hFIQ9ZzmV7Jih
OfH72w+e0temqFgz0MtzDhK0LSHgJ099zi4GmGkONfVn6/Xp9BL2DllJKMa+Q/Z7
cdiM0atC/gZ7MCd2krWL8nI8lRP++XrwmGbEju/uHJhHybzsdo2JIXI1vPjuMfDl
y2UqTjgn9IMnDbiZr4DeK1Y6uhzLB9NyRJhU7Fyv4K09LNRDBIN0w3sISUHvizl7
uTBCc7STMYA+tcWyv6BAa92EjPLrLh0j20vE3plb3edIeXNmHJWEEToowq2J8AUx
UK5X99bkjjtCriEczvsYkrJSElQPJlZDEovWnw7W2XfhnC3UtUO6CKZ+1fl/UntL
qfS7alychPS2E/rIrVRWtTdYbYqGtKMzMEudt2lzhzprPF2sw0xXxNGg/605ki3V
80jQQIhOp/+6b0PQegaD+Hh35KljS/LicX5XSV2xRnZTh4AbqBy8Rmb5fO+DtqTQ
ZCbCghq2+T91IZvXnKCmtq0ky8rx/HtsmDTH+Iov/n9P18KByifmlyQwP6NwDB1J
euw0zkv9KPw1EZI3/BPKivdYqQpoIYM0+dCB0w6WeN4YELK5H/TFTEblLHYm9XEb
AOpDkf9cz6kjDNVK/DLlUj9f1vUjxihflVM8/GAOoNPB4DFzbaCsWmoeqCJcHQDu
Lt6I6jm6TvSGMuvHMqteLSTa3ZfVu7LkPFAnvIXiWdaKFeDjmlkaEFlp4wWso+NT
wD19vKkLQHOK60/cHGckDeQgIAdF6SfkNRwSmFmwJosmmv/euikEPFrUbc/teF7p
O8ccu7tRTiu7LtdpINeOQYdgyPJHLCoOKl+LJoYZvWf21mVaABUGX0D1oMpRpndf
U2yrk1bH8Zs9tOcDCOIENLQ7HDpkv2O3C51ndAxuWCdQBWWEFHTNhZQVPCaF6RcB
stSJUbfOXLNrs+LZ6BWFACxgEMOZqHrB9HXkPn2txf7NtyOMj1a0RZ4KKbC8gt2w
RU7ELouqqsshLepuEFFaHNwi0PKYdEE3zSY92pcppkkBVZZVFtkX0Ji/3tjJlKOl
SH05HDI3brCjDlzjkW2n0M1NZc2q3YhfWa7vi7mB8+7W6vLBbPg3a2KSXk0XxJfh
S9RVlWEz4inEIbe9yRHCzLJ67Z49KB7Q+eYNiJvxHZVh2lQdKdHm8H1mHtFYyS+P
gT5lDl29ca/wGL4aYZryfm0Qg1UnJ3Qq1+1eLl9B1tShK8fSnGtRG3P3UPsnPtAd
7g4NghTeGGPhZgVzaZRO/TER6tItID0w3NmjP4/TYGVUhUHnm88tg0LYSAjP/wbl
rVo+mXZB8nvULvDFlYtooxhZ1lvu90Tj8dbpQP5Pm6zC+90u1IMMj+0JnTnH4EQS
mK4kEdS3/pe/6nUDKkR+r0m5C3LIftzNypeFaVa2IBW6KMbD0znkIACr7Nh13SOK
SbXyQS+KRv01sloHg/1zSiVeql/3JedwQd5Rl1WTQGMq0Z4DSqq5A+Nq4UDqsKk5
/QvvGgE8QpqJU5cEh3YYsYENl5cNdKnE14xdEdE845Yx61Lh6SEB4KJHnpwkgN2C
PDhNlBlPx6ZrD/ywgJp2z6POeOgtwMc8hHlJh0CiZJfrl1MFwIymJjl/gn/sQlrQ
6iWHeTDRefn0+nEv1NyGW2Asc/OGLrD8iySKsgjDSG1BlsOxNBLbyJT5c13Vy65U
CFCtldBLYVGF7oFKmw889ZDPsGdOTKVgrZntrVmxDvLSLYzXwQWFgjZJ36apVa3I
CCJOetSOjpiEQ1U8RolZJXVIYHNM1p9L3e5Qs/0jsLRym78eUWpP5CG2ZWPDgA+L
11TDr7Kmu4zVNXiPOkfTx2FSaetXCXj8QLmwXokR63pf8XjowqfutdercquZTOBf
n8LGX26K3sMwDNtHleS3ZBsFL5fKkzlpYG5D9IqXRUbyYNrBR6ORi9qxaTOIvV9d
2RYaA03FDoRH/TKD+sD0yozIWYsXl6Qgg0YNsJfZG3vHvjWyyWxNMVg0t07GCflD
jt5eSFCAPgGHFz7zI4vbuk6Y6bSsWmfbC1ios9YT/ttEM1CriSVPR/o+lX5j/Q3W
w+vQITCk8tUjhzCQQ4b5grsIw+SlbJbHNa+c/DDydmHcH3ShnOM1aLCHeGSRW/eH
IVfhVIg4gBJMA83L5/TchR5TzkT9U/GEyDcrDJsS8xr+w6esA3oXINxmkDMl6Mmk
PwMCZgJIFfIEtFv6gadPIwwC0imy8ukLojkgdd3ZuFmY4Sr+Whe9Hgm7Tioiuok9
UHoSvfE8byqXFyA9oNCTyP+7hOABaR1GPxfZH9wycfeRtIZasN3OG52QgW4oZEhA
zSnZcw5EvHBBp7gxdWhLUdgrjrXTOfKdOg1KOqAvACYcCZsxfGloZ90Y3x9B/cuX
QMs5Q8EXZ/J1CQ/uXbM/ty/6DVwFVNPmfcHcc/vJ5NdWoPeVuYF/kCEFO+xOxyw4
COT8rkUdmsRNP4XH7GV9pxx4P2Ha1yE8psN7rpLX+a8Jq7uQ3Tv7D3FPECJCebpQ
Lb4C5jeSgRDRTb5RUfiPPZQbMdYsm6lhX54W3uBMf/DApkkDKiNIway7yOuFcEZH
/VwAiT4bfuqu3TI4ClzMLbNmPv/x3sdFBrb/0ttr9VZQfOjFf/2syPZwrn0UyOYA
qRfDAYh6+TrxInS/fRidzjKyr0E9rzK4CvVtZZnBi9howIqpbnlGIDyaBVouIxH0
sVq5P3o7JElMcT8P6O6utivz85Bs0/SIJ6wpeC4yVwLf28Dn0kb5nsP9U0IXQtIw
oSHx1jGtkA/uYh3Khwd8VpagKOG9Z6eFYNbW0zhZGzc6My0cbXfbnrx1Lx0RYy4g
NSoR2VZlQgvFWnE4pn/hrMgrDDKj3pApR/UqGeFBxW8Gbq3Hl174BegtC7Z4m6bP
NqWAKMRGhm6IE9kq/3LCK8gGeJbwe/DTn4lRVTLG8HTNsTxmvHOKdZhvJygLpsn/
SoEXwYoDvO6Ynn5ubMHTAhYNvx0Vh0DkKKyFwjhFXY+8hW0ZLR4Axvb9jgyFHfc+
lMbqYO+CYJfCDHTZUgC4RuI8UBJ0/NMOR72gKB9F7Ifmh5W/pp6nOTOgxNz0ce2r
MS+6IItG0FXuP8GHSzkMuhRBgwW+OJ2Wp4NVEaKjezF9jWQtKxsHX7xQjWKkwcGo
7HmRieIqhZqhNDsUrBvSCoJf0ZIuVEKBfZiXSQwnPvJm59zhbdVb8XFqFz9Vuycx
1TWEzcQgHQarCTx4fA3Zv1YRPlmwqpFG0ug9NB4lzlYLziqayaa6L4MQyElQEmfK
2lwUW8S43jzcYNCFhHK4e5OY2THCAYONzM7GTxLD68xiCLdd8xdNSvC61U8kWxIi
f2Kwbir//6EdaJOus/QjNQwUqOTxS1Ltk7PuXFhb1ATpj/giFrSUTR/lusi4NOyD
a+GN4GOMf1HYOlrKFfxkqTY9rueADsCdn9jKOLC9RLX3PeOouBqW+M3YKBcMj5Uj
TRgfhOikgDDpOwrn2KluTKiA2P5uHVU2xsRVR+7oRBrbOLoZL6rLL2zmV00+rODV
/dqs6ubhujnowZRMK1ZFjTyPn6c/UmqgJEzKi+IkDbuCCaKFD97Wh6jD1ADOK+iz
t3ZJAz6DDHAwysRfizN7+jdOdGhZGe3xMCOl32yvIaGzQZbLx062we+tNNa0bWHt
dwYEe4uQhwz4miU/ZbAw+i1tO+oHbkNwfS1ilCGQzi45+fsoJOjFxS2btD/dEFE6
P+p7mRrmyNVXSmTppNcq8w2XoMhP9t3JHVd+5EsP6zaFx0zk5V4vp+7g93IUpgpu
gFR+iPw2Hc8JEFOA2+J4/tKLOcayT3mTdCg0S9QMb0ye3jmeyaDbW+1Bk6IeCRpF
A5GkZWWhsi0aPUJ/0XeMIh3T2MAILLxJ22Ml8beU+1lRLCStLC1Ua/VRRiPr1bG7
T1IMBsksaEn3ZG0G5qrp5TSoZ+L8FzMIk9aSLOFjcUE5vNJcn5spvqi/TjMcedjn
hUYAGosWeY1LmahMy8kaZJY/niaDGgTXgf2O/eAPVTYI2uf7fYXVNzxzqQIE4owO
HH1jHofkDHL5ugVxkoVBcP+MJJYhH1U9QPS4YzoHwiSFG/r/C8gboIxKrPIw6xi5
U2Q2VIbdqYebbPt1ECODeoN0fXUM4g1z5q+cOJPqCQ2k4cZkTLKhgnEF2+nE+NGs
+mRclTNYsWQaZPkyKIJN2+XqYi3oxg1SLuBHBaNeImTqUlu+R+C/+VqqmV8yvBX2
j75JW3EfYzEl/5w5L+DMvMTGp7RTlYYZAqp+ujJwc0TDjh7ReCbhYzGUaUZFiD8o
x9cfwBOWjxkS+saE1IlvaBC4bI/jG5DQV1ruQ0vj3DbdRUOcwi5g/X6eyF/xwSP8
D66J84I7OmmTgpdA7VZWX0ok2Ogpv8uIack6Hiv0iuqU68Uw9ZYtQRGIwDGFEurN
KiGFuziG0QxUK998clUP0S3UYfcH064I2rUyaRwHnlTBkV16jKjXVep4OcYmfd3M
4OvsUW3PaI5XCKAw+TDc4wPB6w8BcUmYa4mEZ9kYc/G3OBUSW2LYr62oA6WVPKaS
5RdDmXTMp7YH8mV9BY50GMCYJMts2hUS1xNc49N2/gxejmKUySVtyitDT9x65OhS
YDIyoLtM9tny1UZ/vN8nqx2vxKtHs9jkjS082OT7LSaojVnd8+0+p3mcDKWhodKM
mLQjYsjEUP+iSsh41INgDSV8+itXK+ReZ2AYXm0xYAzIui8sRYE7EdNLqIvFz8aR
KH/mgm3V+BbHd6HBwABGgfpQQ5qhQHzMQqOhaL2JndocjbA51Q2pGqq1yB8Q9/WI
PXuWguM5ZLpbd9DPvELPEocXSNXThV00cTXtVidfDvOVjJxhdDZvOuvtYY8gnDp2
0yd17x6l6UeAaDXGYkRsxcuXJASP8HJlvRwKZvWcZWk58/SO4cry3B4raBalFBdr
c94yX2LkGHLPhf2tG5ZGIS0mncNAnNcHqrOmKYEA5kuaxnDJHusw4lEyy+2aW1jk
L3ucADPgOP6aUf/wU/Ls7M3F9pGMc9yESOgCb+VUE2cmxjFJtwfUPTni9IqLXYAA
FY7JGI0PGAwY4x3geF2IK6Ot211SI8rkxRiaNWQC3M8eo1ZQs0XZJWGtbh+9EUky
qO28yTeCACPtSWTCXz7x9ytZfwghOJGFj1XQn5KyWAiSBdJfgulLQWDz7hy/acae
vrjY1b/dSvN4z6khoVF71thI98FE0QgPiwjibwM4QhP4b7bRU37eXyR/MWzk6Q40
Oj0akfyXDjDRgmsWA72CYwTjaBNgglJDNPA5DekqsRGqcrMsVnUQckZv7TSJ7I2w
tiGIn+vtV6RLL1vkCnOre8d68v/a88CJwji2SDl3siWPgC4xBeC3qy0ZotrrDdma
d2ZeSV4lrcFXzJAQQq+G3reaQb64HvkberSPtJwoVoaO/0qUpgwswvN3fLsQ7B35
6vahmbDqi2FprRFHIR0WRr7K+MSGiqe2mhGqY0cjDJxGBS71moyXQrjZpoSF84Um
bG0ije5EW6ZDdvgKdcr0XhYtayP+XDIG7sBDIDwSqcdFBsJQ0FWPWJJGSPTxb+YQ
86kUP4nVunC63Bp8Xdsj3QEZMLZXS95P/f+9U1OR86jzUA4AuUud69DCZckRUO3U
U9OhnRcUcHYyHmwHXsbZthxR3SF0hthwgdwOP/EW/v8oiB/Gred5KstQ5cicskkT
QcpOUzX5DTWs7Z47k3t/sWSV6X/jbH1e1nlVRF79NlnIU1wLQd0h+GZX8KcyHrRK
HajntcXEfs6yi3eqqlh+SMi9LteYYuJWVneR7QEh0TVg3tYnERiJ8OuJZ2pNXfMG
mpMxt0reojAIx98ZftQYxnJo7XoKFG0QsKoJJ25ZWeisCIUrRw3Wtar/BlCWraDR
ToY09NtpVrMnK/SqGW6bcrv5iZqgorBRZ2GJMnkJ19C7QH4rozIaxTbSPgC6qHJp
1SGc4RgzvokiadLAlL35E/ZnTklAwiLbl1vzTLjoOLZ9W9pZnbNiggu/Z9lU44CR
IJjx08Wn+2c+Tl+0nnZtw64BS0Us7UMcCfDz8SX5Fmljy7kLW5xGe+WEE8jP3phE
jH/3WwYUdHrTfdRrCXm8p1b9yGFY0i5ybYkl126OvwhyJbX3dCbBRrAzmxkj4SZS
Oc7YLO+6mgnSS4vIxTBXmqFGul7LJKV1btsQ0j9R3RiIFRJ73iw+v6o6aJOa0pJ3
i6OwSYt63MYoqBtvSs5bdXDPAA00gNoiO842/DI5b164tfcl/zrItD4ihR3PiCwq
AygAQ7K0Sf6DSot2MqxgJf5eSVoODtuHz05CMoMsjytxqnW8LwcVlWritsUCsaqT
hxJ9zsz9pGFKAg/ijRWKpvUPRnY1xGqPbsd5Alq01gpHCSjX3Z9yx//14TJxCb86
iMxu1nLMfXqsbv/E92aHxI01EFkT2iIlHXPe65ldXRxGtgZQZF/C+yPwS+yyW8Bo
dd0Fb/P+9Rzyd3i0IoGkfQIdSdzw3ouKA0QwbZT8TU7cZ4DGGbWt1wPfDX6a+NzN
CISzB7Ykdsrr71rAzrjL3z80DZJIahgilk0eG1KPVSDQxdFcRUVOS9XiT/kw8Z15
hWT+kLd9VtbwC2hCU6qRJxVS/snGXFM4e9+OePUr5MtQRBRcwCBzvDQ4N0EPNQlQ
UjY3Z7ZsVL/n7ES0p67rr61dOuC84ni+d2rCC31oy6mGBAk22h+fbk4iocU4af8a
u2PcShOR6OWbIvOnPBrziy1rNKg4wOFIkmeGTbZXmMgOCyAX8OkzfLJ6We6kBL9a
LZMOauUcW9aQrMsqX2S/WcUMFy25H+xlPX5S3Sc+VwS54v5i3+LSIocLZ1KVwoE3
h3cYHBggG5oDlNgHvVs0o+n4mg2ZZoAFBKmVP2BeGbkpH78wTaElC74FJHGpIc56
hmfgGaQf4Iw0XsUBKVyNZKpqto8Relxy6gkpnqsl6MCafSjBj5gniDBNSezq/iaW
HG7ovg7or4TU92TKnf2cZiaKuzR9CfE3qJzpsKoH4b3l+4L5qdtjevz774T0lQZb
Z20J+ZxnzKv7kgBaxmhR8zapxvnqWqJSIVwTEPVYYUfRt0PriPPgvxsqOj9MaEX6
bYTFIxnLjCoWTv3C+KjRh6QK6ioQipJuOQaBjgjxU2Ti7RVWXBO39Y0anmcz42pn
LSsWyqtMqy/FZvL8qyoqzdz6vt1mBTbgtMkDRyCE90uIqOYJq4egCP7aSLXw0FxS
ps6nBIv08ehknfWjutYMEJ1DqD/Mn+zW+SvrK+E8QhjSBBJkIlkyE7w13u6mpmEJ
Vcp4+ENVCrWYtzkbFvYIQzhBWbPU0onoUQAdzDkm06jbp/EfJ3LB6G4ThA/zg33I
CFGmpszMxDVYRTuexbbarhfF+j1DYBfN5WTvea2QdqYq6t9bWRVTR3XbV2hHV6sd
GyMuihBqgJFc19nGOx0XIvPOIkDKOunLI7aF+QW0wzLO2XScABpy1ARJAluWxRYx
gZozMGOlVCC2I2TkOfhYRor7d+1j5SyEEoHmKlLG7mMD9V84M1hM7JpP01abMiQk
ndrbbs1JzA/KQ/2FMKT49GxVj6W0jEGP15wL8gMqfAarl2ockB6ArfDgRDPVeuIw
9iELqscjarD0FhpKTxM0QSQusdrIskkzE/zCJ0r1HVmqp56YZeLjOgplgBw7z8fk
7zMVjBnEcZLyD1Umn3+WzpBkoCuw2v6ui45/FefGqmL1PjWmWknJZzZ4IG6AEYN3
5i7J8O4aEQpQQvQ95+nyUELhVlotCarBqO9cmC0D+gvVswsgezTiqPPKxoMZ+gL7
89RmLRzoWATg+bzKwfD8dFT+zHNxazbyaBEwZWITnDellofzp5SFM0bzaLnwoXKB
oj7PlbnKpJL8BLjSjgIDojnoej69V6MgGIWf9OPAn2ph2YTKtoMQXk4sLMSpNKH3
UCXLLOFfWEsimax9/G5B6IVNuuZGCr9kS6WLheKaZnbzAInSA4CTTTxDHG3Mwle5
9LuLgwSUx2lULR7Gyz2MGCiObZfgJ6f9531e0ZqMGJbxgBCTa+sWh5ZTtNnof1i2
Mm2Z4uW3M4UqhouPQ0pghWVXQQPmHyYkXcF/Gt+RrgpfWEQhs9LSz62THFHdRnE/
8pUNmiteEpk1qn/ke/1Glpggn56g7a50kzzJq6+f2iYIFyb4lwgUdvW1VMTP39CG
rfAwYPWIQT+Pa5Lu1KhIH/FbqNulVH4GoE8JmCcbp4cRI33fAu0DymsigEGg2JGE
bVyW2Bw+0R1lJFtRgqN3lwdzUMzBJ4taudvUY1JBmokWz3glNwGPfVTWC4dkE+Kk
PBT118pUp4+dViFkuNqWFxTvW9T3qabDFwSuvFGq6FAEBxTdi4Im2sXzDeC4KGKY
2PFwbJvaC6R8xK2lQa5FI5rgWTF290pqNj1lND/H8HWCioKE6s4yCCXzT3MPVqj1
bWWdtEW6Qd7Snhd6OJpwg7nXisLGMv0yKbdbfV4HxiADs617GKhV7XhXvWfYPNbC
+uqaatnguIRmXZ/hUoBmsMWNfaOUz08prHQCH5W7D3f7DZHN0SRBIMuXKVsjlwmF
9aamvKh5F6R6CQi7Z7ZIULkh/SmWpON5b/k0SDlAq/Ykm+uCjY2brUbIr3SJxvz6
ljhuuXQslPoVKQ5l2kAUFHc2dRq2EAHYM9zOazHZ19KDCWXoZTEZmvUOltARqTwO
q9+PBRP+qtgIrlGcPNzHrAATkZJe+o0xIW0oyYl2voCvVWnMUD4+Ps1qi6LwCrEW
giKl2b8ZZcFf7vJ9+Y6SYsw+SW9FcLD7seNACG+lFmebDetzFkPDYhNgFcOKzOss
VaimcxpEjw7CCqa8RtAPMksKWWjlIGqKkB/QswPO+/l4sSkwZj1KNrNT75wfca2S
CiOFXe721bXBbj6WI3Mn7fPkA+tPqbzWB7NVeQN66Gun73eFko5YIRyZER7QlETR
kyTuZbBSnaHP0wmDv/vS39fpGkOae/teflAMB5+SM2Ftb4Y3Zd7YryNJlIT0jfmN
k2ZU1EO7Bgyi74/kMn7nhM0iruWyidoOziseR4XGQswHgHkCXcN57FPN3OJM/6Jz
1gzgbXISKRlEh+iA6X4PCk2jcRHF1vALTBlxVrsJy4Ono309nlVEUzMLeP738NIS
gZIe/FH74uzHx0Vr3d4A+zBZcigGp3nPhzRmcgpvciw74QEtVQFFhXHQ5/Rsb+ew
4Y4rQlZFjAiqG+tP5gw4v7etvGMgpakSYlIbRmDwLJrlE+TpRzbUV8cMxMBf3a0q
S2LrF9MaxmHpKO4KcMP2rWEhoZF7/FzfQyQXckzTHRxNhi/eKtKjTdXRDazIWEEb
12CfgHmdg/WhH0hzOnpt8xYasUspoaVhTWP8IKi6b53p/Sd1L4oDkbX8lUl2Owa1
pYqf5COU/po1NSGUP164UZ+4YoomAcmJuFEVtY+1syF3XLTY0Jw6UQlcIHosrVbP
bP3GBFdZmbjVU520l5zkhoHsIaT0LJa31ZzeQrMT3+6W7pe93qynkMCTs7jwFrtv
LOlJbBg9hevT6GGY2QgEAYUDMSwzf5xPBfbXjWlvjg/8+e/UCyR5N7W0xumvJkiq
wNy51Mk8FUxgB3kAWzf8NPw05lZ+zwZsye+pO599keFl/iuUoAN9OqfUZjNro7f6
rzI00sYLdkEgNRtXjWetXpMg+cH3qqpkqp21HOXuC43OdMitpUpVMh44QrGBPJBk
OVyPRMaRHIyS+HMfz45TlvBP6J13ST2jag/3Mq+QTLYux+w0cy3QeBeKfP+ZlwAz
66RCT0mcfgkzyfz9jG4W5Iy/0g8grtBHx7GCpJCVi5Bpqt1izXc9YG5EGUKyKNu+
QVauLocxFfKV+y6+TcQSiQpMWqkq38lx2jhqtjODybeL+ihzqNUnQXROnx1iKuSS
kJJEtcxAjLkY4hgtC3N3xsw47h/Bs5yr2n8NjxoyRG0VvDf7iRmLCki1PGyR/B8p
BvsVz0rDRt6cBvG5m68l5UOtxaP6+LEu4+C6OF1/H4JdOKWg8iPWsi6xdtikoaJN
5JxjHEVWHajrM4L3uX0uUU9AQOsRXAYMW2uEKvJ1f0gNbQEe+g1faf15o5U2BTtO
ebN0RxT+ZaxJtK55VACgSQtQ1LjQ1emO3eJ22s1y1IcOmrLza9l/osVB8qMN5x6z
li2ZzvZ68LxkTbZhsqhiZkt8aOPmOM70YLj5g1M7YY906apW+jlsk1tUInFFD1Ty
sFKC6rdcJk9ZS0WorWZQQkI/PEnnV0KlTGE9L9A2+IjJ98ZE10tLirPWAPz9jXkb
jYuf5ULfiQr9jCynDd12AIO30SYsA1O37selFU50AvGBmHHy4JByYl+4+fewlfDH
l3FSDx/v6eLhVLjtDc8OGnySI9p5rpMhDKUjUS8shgC+JNNgTdC+oXJsTRCFSTRK
XndSyTptx6w+e16Vuk2kRn4rHEqy5GbOQRTPS15K/8AS4sg+dmxmjupE2VzkspyB
ovZgFzAAySd6DsoPfqFXxjHCE4yAo+ALl7rYtpn/bI0Qe4bXz/tyQKRGRcOnHW6D
B6SdvLTcgx9vCsJQCP7Tbgvl8zVFfqDm4FIcUihmI9KytfsBH3Kb8b0v57o0Cf3Z
dXuSUrWrknA6yDfAQ9ok0SPrIdQttsq+6WaOFMbaqxj3e6wR8D9d1f6D6cCEr3oV
y8bdADQ76eHRv6bPuMTi0a6Olw1RQYvdYZzZWtXww2YGh6miGzKAUgxCGwJtp3Ad
LKzLBXEAPBxaLIqVMRu/u6AlMeGbiyxpWtWpx7JqIoDfN7p0WWsF7uLYtfOwWR62
TExIhQLeuJRBfa7SozK1w/D+iH8jU/J3TGhTK2uiYD7N+eXDkS5QCqzYHM+yWZ+U
2qo2Y7ZFWZrzO74K0jTX+50YRh+SiBvMsVixL249ONkQpKeM8mG6kdx83/DGp1+8
dijnm8v3WY/e+oNYzpqc2QPOeq0kZ0RDgPxfdtW0QtKAYIYOKgELKmK1eC3hSD/w
zu3mbU2URpOuXUOaod+oqRdpdXMRH9gTmNv76MBV1+vQYhp5CrjxfWq3suuViMee
auyVrhqBgAVujOILX6hwEPm5By27e9TGAuM1o/oVcVZMuhNj4nkVFMjpjHJ5VeFb
xHRZYBgoR94eFtl/owUp0+dNpFQpYA/8Mflc2KAhNYi4vwW/35iUXk6KNH+t8ZcT
uekqSatoOfhHhyT47V2yLgvftQsNXjxNmV3Dnm8Xcv7fOXm/rCkEUEVOLGVjpVuj
nUmslxs/DG7t/dXLG3bsSph/O+MlQJS4zEq9+yU6J9g5WdwmchdeJ387juD0beW3
N19iLUwWqxrXMmqUTyD6VG76y/BsOdI4saGxraN7lEFM3yC9QcQTxCJvmw5DbnDs
N8isfbisUSOeyaYkrf23ui13OSGsfA4n+1D3FiwJBdlBsMgC5+UPMxijfSdRxiVn
2ectXQp7asRJJ6XHcffIqMdZNOkfbh1BHJDTeij+sAO780m4JCs0IpoSwrAwzYAR
fffHuzZ460JIP1xLv95rLNCqS4lCnqcOEQTY7f4yXQTUsEnMiExhS2wtZe7f+qA6
cPMi8jtrI/OM3obdhJSZ7HpegjuQzRCEFVUo7teVqFMP/JekvNiDMoO+gdNQDtWw
k7bfhK4ilgA56DzEn+q8AT8npgvvYxlPvHXuwikZK1Wyqjh5/FrWTTnfsfWhunXj
CYYcpfU0lCXORyJOOclpGz2rI8DcKYrZIPPp/BDftg8hVsAyoxamimZ1vomn/v14
PQDYsPwKjywI0ZAFub8AxyqiXQs5w7qiSiKPir9lEG20keTBYS/ClG349Q8UtbIU
UUJISMMusqwQlft+9uv0YisPg2fX7mYdWUtRzRFoJV3w97CwLPzLHaHtfgD/MO8U
6ZTem/+ItVH3YN3a+7iE3PaA838N9qidX8/EZdRLNycim2oR7ABoZJb7E1gblshs
l+dKhfzen0XcYRG41q38MIdqnAVVpI6QU/Db8TC63wQPQ2RfTUNf50BFaVwrLwWp
WdEV3uqxDlbUIzEp3Don2p2HLxlkBRZZrmxb53jzRmO/oPzg+D0yfT/jI6eY5ScJ
9BHVs/wmU6siFh458iU9Ze+4PonYsVaeIeJhwaNq8X5a8dHE2LQZZsxqVzb2ZSo2
GsLr9R8P1ek9q6YkfybE0A68R6tgpS2ZF3uLqcDVN3S8lMW91pLKuUrVsFP64WIR
Vg1M21YT6wAQHE38MWl/jo3CD/Ao0dGS2U5VsVJirMzFKc7+rEp1ZNrfrUefM168
9vrMOZorOcNSW69/lO7LcgQAasWVTTEVZepLYxxPlFEYNzEDC8cMTKw/kw76Jcil
z9su7ZqRS1b2C0RqP8on/44urtsb8i0/eXBLivkQjXaHWO2TqUs2Q4oaBAU7pyy2
WXBu7swx0RjWCtHGJkNbNhCswixzFWA9EMbf40U7OGrIAXD6Bi+QjQmAX7wJP+7g
PRden02IfLizQ51H7gmc78HKc0Hd/4rU8jt6nFjvQZOn2SkSKETNQyXyRaUlkZYS
QMXvFie0gtTnWWmFmxv+zOZ423OOrR62xXMiRrU7ieJJpxlm3Ub0Jd8tZm2W/XAb
9MxS2dmvJY/hB7y6etnSPN2MDdlNaq0N0rqlwuI5BAVYtXVZTzV2ndP+aLf9eHpz
gdggSsAPcDaLAynBhG5UWMzmFjhvGOMGmLjVtl21wXBO0vj9kUxekiahdrGZBtk7
AF77imiRJ+oTcVsxn0/WpYbQq+5HD5ozoitjJpJF8Lnp95MgDvB5fDfvUlcfeHpG
zkCpUjSArvLIs3PGfsybmfAPvZLWrMgWwnMiMeXvnxK4it8pypfGTPzkjOFrbT6b
PqNmkmPMjCRsZIoGySJ0AJ4s40y7r31ft2kKEWPLg6gu00xKTaykGOn8K8DB9TiR
HAPdFEECSxka1IzalHQ2P++vTyhKkbj9+TrB1d6Y1/FyLgau8CNKzurgTVrVzK/6
M8DXyYqBNOwx6KNcCYYaxO9NsGzHihxjMwlx0bW6C8267Ocagq74JuwMxsifvni6
C2HSeXJbha6DbwqAdtIT6Ne/g9gxEKWArJzML+qTY3caIfAD977kuUYwhdzfphpi
+twcZIbv6v9teQ1CBkGnPmXZWx7h28X/sMpduytSj7msabKNBrewF/LfV0Si5vqY
rOxG2Px5+/4ReneLCyR6EdDQymwwwoJOWrcLvoxQsb2TzvOwQQts1Gi0YDY/0DBi
GZuGv19WEwa/VK3nOE2u8yCmuc1rk+zJ4Zy85DBPRQ/8NKv4aC8POQQS7y4dRpHR
UOGfvVxYXf2SOcPTVhqp0sUotYVRWtUhWlf79HRQNyBNeLKo5EjzpoaIyO2zmuWz
o3BwSbck2KhSll33vPCXcGgFOauxlVsI0vGwM5MJ+iiVLqGVQCILET6DDwF4j0Wl
xI1xfuzns9gm1rJVv7l91fYDa9PrEpcgbXaczatDxfDp71d/NurIxWn1ute9tJa1
aayEII6+EVvt9PDiZNonq6MCvvW3jwjJhPWdYpK083IBJmsd9bWVyYqjO1CH7eMA
35T1hq46brLACzbd40Jin1VrfIg3E2/QC5QzACYv0IVLlsICXq19L0ft1MN92EvR
/PoTjPFln+9wWIrKsH8snv2TNmZD3klzaK+uxagcua6ia+Sq4Oi80GDb+122Tacm
3wZ9td4RNdVtORzov7e5LClfIsVDlP6IAzSDGDI3AiCs4VkvnAXOn4Y9jEVbfcNN
0G+SRfYoxl78en4+sKv739TWg/6W+ooteJQ2h4VAr31pj+x8MJWeUxrg+0h3was4
d6Vjh4fyi8FXNsgQvD4kmuxusOMgLY2P+D2WYKH4MH/qcXRy1JXmtnQADBgAgdYA
WfG1OU7cfxVir3nVom5CvovUvqZgSTtus4/Jb+MclFzCNslJLGpEEQa+kwk2NhxF
fRW0TZBBebgM0WrHZl0zyyvmS12xK9fKoDlTJiYx3KHLSyiyjprPncnOMf7zsqvx
z0HhVmQr8FKUozLbpKA753Dy8OsDwSFSNh6ib4YgUTIGeocz49SAPKNF0bha6DZD
AUEdkQ7UfmMPfJQ3TPAg+vWtDgIi9jzb0UB8LgA3l//bhtEXknX6GO6EBjx3iCR9
ubE7D8YpArh+J8EfGcu//vbaZ5iUHP/wAoFyGOtadt3Z7XPvxNoTAx67yOQqsVsM
rB9afMs705Aopw+2VplPb5h3znqJ2EKjFcmnLPwR8nyZWekt3etWo5gU/8l6JwM2
/fWdqEu0DgqptdWgdkTj2HooLYa8MFVeyFoau5W8qpS00KwPnDQbeOlNmaV/rM0S
+3pxQST+cm78XpFQozdzanfGTkMHej8WEMuIJXN/jMm4defu6Soixv86f3BCUim+
d6zctQuL8RQoZIwaH/qqTtwwafCBuM0UwwZ0nCio4eiq6PZv+ADV1BAc4Nx2Rv7B
Uu7+Qvy5MskrcllbzVhSM57LWJI4qGBoZKI8naE8ctPBwpHOiP2jhcWN4lvoUklY
YRLGVBZ/wT/W9AzuC0vUpyi+jhwvLBtLMK2RUW0ovKS+0uVgqxvFjR2MTPMHDxDn
E6l2JBw2bE5jWW1CUruNf3kUt82Cz/MPcueKG+wt2Y/SczVizKZY4CfQPMZJhLRF
QHGcBW1muFNWh1UPYu55daPzu71b+jiUP3vDHC35N6Y2beGt25X3OGCGwdTk4K42
cQzN5E9n3OaUFhDJCkiDcYCtS2wAaGWNcjBiBHogkLna0JQrW7P+flkkZSlDDrC5
bLhg9Vm6fXusLcJApq95qGb0Xd3mXCaa+AL8ecfXDwqz84TokMSjkSm8toIt8j3K
YCxJDxY6oxPpOXGY0jbsvsi908U3nZJEqbcZaC2qviioEDU7x6AOc4U7J2nKTL/6
cukKuiEAGNYBar2vLZofFPSHWvOgDQiiZC2fEMXBzVr1FuqyzwflsKOyRDOc7EFH
EFoOVfm8Q6nlEwtZ7DgEZsf/XNm7OTuiWFXL+zXDA/inWTmqZEOz0bCIZum/NCst
wOowommmxTNzbupc5jh1+CMFyyvxR1W5UU4jaZI73MgvuPbBWIdLI+7nnnXYXORD
P78T6Xi1fdlmaBQYLYR86WiwJ8mPmOLFkxymQdlrPF0gXsQRCv7zWk31p3pP8dG6
ss/88+4jHWTFy51WRVpYTN0KW/+n68D9ztB2X+yJgEe6GrESh02EdBhVD0njrcu4
iNVYjt6/QcF/Fxx/TFnKTcGmq4DlKahpsCM4ipynNs5ggPvj+wRfi4d/AlttMiw/
4CFWEFCv84ySu1wfltlLn7POOLQV1+QxIx5TQ1v70KLJQlPMvYqXeMmmJERqcd9u
Rv/woWaN7QkzyzHYAUClZ6SXCaapyAWXPrFnH1jIOA9xXgyZsLlCw1PskIgXFy+H
1ZZVyMUYHZ3QJgsogMkVwXkZEw8oe5iGmgFR+51lnqWrufgP7ygGnK4FMdPzlCEq
mlmAJ8oWDMVAtTeM9dUgujUx7i/2FM61PjDOz6JDalgP0k9vA9EQvwBZjXjcoqdH
jsW7hgUDTu9LA7GEGf3uJkYsBzZbY8a97wp8uFxAlfTZIkGyUjFn/CGnxxHOXVEb
Temd+lMpd1MmmgTOLgUw8Wy/rDaDXmPA7TVhNnMtDek768HeFfI6cVb8bx9nbpzN
o0q8iNpKSZExv3CWNxPxObnM0O5K62MsWyKhMybcCLNYTNTFIhhzsVcE4uvOPU7T
hkJQTg5/b1Ng6OV2RPoolipmGTsx2yp5kPNT+2Of2Dzwa1Kd0Mv+LL79dsY5Ff6p
6iZJ9t0HCqiSkuzfeMW0tCAr5JXnyA8NUlxgvnel2PYJY3MXahh2JSs2H0Oxslw7
1bFrHN6HyTUzgI+GenE3hyN6KRHZOQ4Xr5fjzm5BgjfeiJux0DFJmFDUpjGTSKSG
vPKI1oCi9vQL3nXqZDmJ6Wg8LIi85Il6i69EuMaYLpH1Q+otQgoBTS2wCsD/Gniv
jp/RCuauUeRh5LaxmI9vE/aBE+9E9MIusD2FNiMoUD5TSeW8dRVvsmia72eL4CmI
pIROIe9I/be+4LLh+itT+IT8rPxUXf0MOwNQhEynthU2UfgXF2zPRXOi2W7Esvf4
WxnXJXeBHZBhqboWdKa/5DagBdYAeSg9deZYeeTkrIu2WkBaOzGLa2/d1kc7MNjF
YzRgf9OQOyGXvajYxouSFxp7YGxT12cOeuoSu4fbvbBo6T/+KAa/pj4HUsHndxK/
f2difbgnvPuI3mJcQ8Dz2XJzcO0pg2W4wcd6I/uMGVMofnv0UKdrYV5MJzi/KNFs
iayqjAsNp/HOzbdO5RmS+r1JtB4cChxODw8BYM4VeQX23tpHyT5iXTGGF8yIIr58
xRX6TYSfAU7aExXKnfU4gXeWWlyf5QtJiavkI6cxM4hLHsmj7XyMIEQE+IMmJNsQ
FXk/pp2VOcyOOev0j5CRR4jsyRGeoGtTnGehrhLFvsVQaEiVSEbM0Uij6YLh2PoU
Pdhm4xCxtugLRK+QTjStYxpWqZiyUb5pjbx3b9gOFdxM8IlSYkiLUD1/e6x8n5By
egmjx2NArkujxRdG5g9FMhIUgK6xcZWqD0j8sawNVbVZmky78VKct7JrkvgdTqHx
vmLF6rfSRX5zRnJuYo4HR3zuAyF/t5flWTTtEHWNHmJaQW5PMiNiXvzbFyDJpYSl
8jEfXGy6h6aG8OLsV1H+HbBhXaSsLbGCtbFNB5IfmmuYOffNbRiXUUAbVTdlDSRS
kuTPmUpXIcD0aTsB0Hrjv5mtsJ7P7vnZfrqt3Y+4hS8lIA9uLZq6nzyOm5JiDuwm
VXiW1a+5g4rTHKqvTwwlC/4yXKMc2KvMQAdi78uxOMS1hb9uF4/k4pf1TCBdasZT
i/zlWMxqOKb9wwl4ASbPknD7ToqNl3k4rtO1VimZXhr6clN5KmYKtzI42vCXPka9
8r63XshhH+Plb5/rtMgUjwJCOSebQGk6J5tGjivDIB6Twwneo3bUhcSBmV2Zzl3R
r+GyulkcEBnIQFOnBmNxWdtN1MHYWodPJyAKHJ0pMWbrec9n3g6b8naA+iCDHoFf
R5mWkNvUtNKqNooI6pWhDo5XPeMRulMPfaIok22sxPbOSogn3hDQixy4x5wzoh+P
hPEkDZ99BlLiBljEZE9YzZrAupZt93/epjNCqgaosa25ir2q5GrxSsBR7PqNuCAR
1y3DzevdVsjKYpRejnJtxjELJv6K11F/2KRJITVLq2u9SiKILxycmDP0bWCnylan
wyi0KwmVR6ejAjiGDpxSHpwX9zVb/fYlgjRUVjM3TwM+tJfKPvNCa46t9wcc920D
uDtp2+MK1nl3veg10keOCHg/K2k0MgwhyefPZGJScrLt2lVPyhsQIp0lZs0u07w+
zwOXAJSaPl4oHvtqSfSHQxFlLnAZo9zHWOMsx7OPoPPD1ZJ5s7vIU9jnFbmsw1pK
JqhiO1JqWnyquPGVQ5UySd7wCXPbX73lN5mHmBDts4Zwk8XHexY43w9dA5QKnbfT
jdbOyEgmrcnp70F/QDFn93brKBp9K4JV4mX9TPCzFH1LiegYExcA0uGOfFgD5goH
xkpA1gBTCqlXOpCJZ3CQNfVRE8WvIjUeva5qfBqsfANvueBWuf5rg7IV86RXNJSk
KhU0NCvO9gF/F9VILJ7SR0149Xe0rAX+O5QZ9sOQEoQRu1HIIMnH63L6buGjACIa
ESOsGrPl0InbE4Ib+FnIe3nGQvgJ1Qn43p5IsEFzpmtCLoXZv71hLk2lzgMA+lln
qY0hyoz7SqsifiIarSVdxt82FjOx7MK1vW+7HXwemJ0sdMddninKsum0b397ET2f
gxR7H+0KRzNurlYEipRvCVrglap3breQjNgAmSLpshYb8ipEbo15ch+bb33uVE/3
1bAKZWwZup0ZoyNhPzPpAtn1QWNM9w+LO42puALsVoatYKpTmaRGPyVG9kdPeVoZ
VjfllV8wFVXW7XsEkOIo3tocXM1wZPieV+Rep+Ynqw3r65qF785Mu7NNsBuEPt9A
w2eNp8FEanCJxvXUmpuZxVFx6VhKBxvwXT7MrIGVYOhE/fPyNQUdY2gUL8x25Fwa
rZ9Aa/zlxszOLDDwbQNB2O8Pgcdb6WjrmLnauMzGj5cqtgigTt6SIFBH+TeNixjw
Wel9TcC65PQylreOhiltaGHPyAIUXFVHcIHy+1kg+E0upP8zlXZOqtFxga9VS8oW
GBk7KywnnYA5V34wosusv3vLsgtLf0RfrGyj6mZmWDrHVg2rZ2P6Y1admPAzWg9J
ibks/qA0np9cPP5pde2oVS6Hw86DYMUA0eBW5uRiQ5f9js8o5vOxDZKAad9Md2A6
r1ncBwcOLOsMtq5XAVgg70ay+BMMvboEqYV+sRsVMofTiaEgUrokhOoNowpihrOj
VaAIfQ9Li19B3mPLL+DrKrYu2/FWSAkZI/x73spHL9ssNUMumGt2fuZi4V77ei89
NrFUc4UqbgeCiLWAQnDLdlh1BMG3FAbwB7/Xf/TAWAgfmEzGGlWvdroU9R1UnQRr
u71unAbgwsRFbjM+Es4gSWV44qPFqlFPzHFcvLJRLb8YtrnMf2fRU/vyMaww1Mdg
bV7r4A3Wjf11iOe4syTQIhGNIjAipqTf6EjxHWq8QrBvb0/4OMJ5mQ/KWY12413Y
m5DuzDm61/UxRgNwjsCSkhbWNp87Tx5IPV0X0Q4adkZ7IxYHWm9nY3cxInCkf2o5
0gaLM4zopmli9V32XgfsBco0Dol6TjvHl3G8taj54D7LQxPylYGLCpXB6rXRgbFQ
Z/JcYSixKe0qI75E+2Yo/s682AFWea2hOADyRVaqQpmLeLSm1H4UtVKIgyl+AZ82
vgoc6nITBVZ+wpNvt3u3cN99p3Aoy7WZpoTi1YLE7onNhOnLfi+g25A/mtUrJ2UI
yiJBpNarnirgXpxFBrO0ZitUip3gsj9AdvA4p96KnW7y7yknHOOeci1CW8Nz05Bo
uBZ8g2o/HlcjkptoLHl16+dwB9Vg8CtI+KEbvL6OZflnitO1V4Cd6FeYBP77USVP
saeaNYzKU/zUmRCkI9CEK71uutrx18p+DEje7xzVi6cHr6NNFJtQj7lBhQ4GqiJo
bA0wNQW4R7VPed4eg+G589ZkNHJpHPxKC+4ZX9EVtm8LIqdq7cDRU05TJe5GbvK+
IRhuBTR6Nvp3u0ybPHjiu2MLJGFsaJHvRbBgOMpEIMXvOXMFhYrsrlabQ+wmZ5Oj
0aICmvO+t4XqwDvmfLtuQTq7cvwmUcUJsN2ctIhlAWzXFMEibI7pXFEQ0hSn+yA8
xX3YHPJZoCWyIN1C8Q3zKmBCrDqqrKSpsKqBv8ufw9spGzROEKxzKHaV3V5YoFqb
zRzG2vGJ48R8IluqNI5V2SEW2LXZRkxem76zmKO9oBFekQ2DvGh/gjs/ggdoBbj0
L9lnfz9DUavqL6hCD90xaiJBgD5B07ZrRia5DBrIdB9l9RsZ08HinGpqfy3FmOYg
Y2eSR8NDvn39ubf9iCmEVh4B9lbmeb2r3CU3YOJpupXlbj7mzLjrRmSKbBPu4rvG
rhzdA3hhRqeixvfN+pdXjQlbqgtoi8SnY7gmo7CADQwPBryNQT7GyJxrX3S0as2l
NzTFBua3G/GtjeqtTSq4B89XF7ppkOMr/WywyzO4iIfV+kc+OK2EvfbeaTVoB2Hc
Uy3DukGFR++HsvGuVuFbnFup3ScMqRBZfoSNipopKVt0OLa3rCCM1rl06j3duTkm
k5yQIImxgDROA9e12j7ch2KPE2KOWVc0XfgNZzZ7GIER4GSg7wFwsEfcfflj8uAp
4vx/E70z7t4EMcWzfFWHkFvkYAICjADzRLY1aH9lVmKqJzT5EdsU0aVIkPld9no/
OSMJskb7SuAA238B2pzRR1BRCwcQWY5qjoKg200PcJxw65xWjpeb0j44tvYkhxSs
USFUP9RKOBGjuigfMfkw2GqlTgIAlf6kD6GpjbQ0ZufS+zwevbqbh5wsykUIIfeh
m+lRRodrUasw1If17RIQN9iWa09dSz8fzHT0sZmOJ1jxscwotbNH9DZw2SJ4xByH
C6MsDuyNnoMzMfsy+sQH1M7OfwplldDxAsRo0imsyq+PQ8PK68N+gjuLdw9xkivC
yT8W7gMDQvhgrN7AwE+jWtZWlf0fr9XT5yJzVhNkQ5anXt0r5N/9rAD9PHMV8Ne5
uo+oib1k6T2UKZedDKAbjUKhfCRYlXLxpQWG9NacydBVIfwSzLn/x6wFQWqkHvou
IBRuIOnQgqGuSP2syYNkalBC87wHQ0PQXzMdc2njsyTUf4s5hs/d5a44/Q3Jyfga
02eyHKRoVfleNybTENoll0erQWtrr2ImXy+RNd0S61xBVpRzKi8sbsraZJpe4auw
HnvbyaFcBFBvuHFMeDS4nUcnpEb8cTwcn6MEnN3P/jiyN3EAHB5ZrDuq5bD1dBiB
f7A5XZMkCdJ7rcW9Y2Ag5HQEXuAVrU+iOrJuhfVST+owzflnPK0DBO/5hnk4RV8e
BlAFr5mId/PaQ4FvnM27SSkKEYyYGR893LY+mJxfpjjU/4b7LSqdCrEfj0jj3K9h
z+JwbFJYQKkHjpfdXIyNUj03NdcvahMSsvXpxqCrQOmzmVOPhvldEN0EvF6twzI4
9HT4NwIhEXjUe/uGo5+5SfC1yldufKQqQAXEBxqcYw9DAhx5iKbdBO0gDaG3Q/Ae
HOMAQ2PbHVuvSzQp+3cS27G4WYlmHWnVgEJen1COTkQh5l+tgz7HpROSaJ0T7C3N
yxVQqR7BpQ/h6lyF4iYnHk38F9m8QvmKv5Q9s14pj8Efl82U9vxcE09uvHR5eGv4
wcxDYaKWrBnYIfP7BvvDoCZBTqgY7WCxBrC2xQuXjjq8cYVemoF+VGxQJG4TJgUz
POVOq77ykMKv++mU0T7yX2thbYtI8biDLqKACErZnRS8qqQ3GYj/9qrVq+jllvlM
dZV9MWrnMOyV6AwADcv5btLb2uR8zGINOPzXX0YhudsHMHVIU9Qgj3GjfBj941yj
cIqhdq3TeHOePFzJAkARuUVRlduSEUWmYmUuDVAVeeSRoKZsYOk+HHdfaQ6OSSBk
1iwTqFGjpOk/vQ+DilB1DGsL8ETrPuggExWAU/lMdZ8bqycgpUnebvmobwj6pp51
hkZgPWh/8bLNLlrmgknsRy+sjSi9DOUgJTQ+ddkLsp0g5n8L3DPf1Pf47MDTybmb
L8csCL9gtyA78+TsAzC8vJ19y9TtzghtIF32KvhK7OFoyrYUlaJcxnKe3vfIjzg+
Kr/vcrsGl0fcga1VaOJD2P2ffN55di9pWKQADPghMJtiYpgGH4P6JTtLEm0RP0Nt
TF2AFvF9qxsasSmaq54hSOzlxsRvCFTrQv9MyM3Ecmuh4PQ7U+g620+IQf0O5h6F
aUIoEzD55MspNuVKlLn3b2We2JpnBCKB0aHqTWN+OhWamG4n43p2Fj3W2ivRP6HR
N7q7+bcnYnEmHJJpFFOCEL0mau5dM+Q++xIgZL9qiv5Ro3LuHuaT7OGhSz3OSTr0
p0p0o/UCbZnkWLq+4BnkeoZFMnesEqCHOHJxsmKRxqBcxJ4Zo5qbQ2hNOYdoszPC
+9Y0dU4FlUlBlfrEwmJvzB1x4ED3IT9+jJZlghnCSWvY5uDfmdrsZcpLDTKRjEtN
HJPTuSx3S0LhLxxK5O/VYLQ1NSmBl0FLRuM87fy+KVqbC2tIvIoBHRRoV7BmV/XU
0qbkIxbdol1dvhCJW0RHRQVUnwM1/fVqVOOaZhIMVmRJ/xpaO8PUhWdarwPxZGjT
SE4VoQwICyMN3i9aLM9ia6ngAf3SFlDsrnPfAmFM+hzVqcM3KG/IuaNiWNZQf15p
6r/nWAl/KZPPCUwImIUYi4p0W9+9kS25sPoYqloTIgLRCOkhbn2wt2M/3gYUtZ1n
tweZ7KbkNskLwnDdFPDrqk9tt+PQZzKN7GjByFkR5aE5uKCRQmdePvFhFs5pIrTF
Tqxv+nGq/5ZrMEAVXNCgWfbKqY0OzlY2rT3XssrdXQctHmsYJE8srv59nmHGZbU3
5B3iQGuPszDdIJBTFVl5QYZOTn1/nEudUovNbnkC3SxpBOtz4lxvQe7toWghi4BS
16spRY01OqiSwV8ppQ3tbPL+mj6SHws3cC3skEqUXol33uAhd/erecTe6NOYCR62
G3U+7BykW08/exVcaetSdQ==
`pragma protect end_protected
