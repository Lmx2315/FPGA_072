// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.0std
// ALTERA_TIMESTAMP:Wed Apr 26 13:33:37 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
P9PhKt8LFvM+S8yl4AhupqecKPW65xJNnj8J8nTHm4ACoq/7MNGrNgdJ7/5sB0lH
uVqviQZy2l8Ff9SAeHcIcue3+avE9vgWIY3VSAvQZ1ZwFsq7zWEoAIVBdmruHXG5
NQc4aCSfnzTh7lyrMKLYHWplcFoya2MRdVG7UP8S6OA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 22080)
lufHipShO0p6M1KmZ5+d+Eu8157sZY5tFJEdfgHMESQYUoyto3nEFuaCstgr0Upx
+uhKvEQbeZBKeg1Ts/xPcH4uT9qAi6yR0xPMlGeO3q7Su3DFV4M91ZWJAvzjBWn0
b7PrrW3bcrapacbk75kxeei4RtlIx5z+T8Vkyf/3r+pjb85B6NK1O4Gta1xDh7Be
wbb2WZS5Ven+bAyZs9SHCjWGbcr4gA5nV0eh5nSeHvp++PHsi6PR6J0aVyGUF67u
ykcbMuqRvc69wG8Hq/zM0FOXgGP15hTbBWCjgdX5db7hfWn4PhlmTWJ/v1SNG7Hs
O+Wnvr8gLnYNPr9nlIwKXHbDZX75uz2K3iDAYHm4rwf2U4ue3e2P9mlnF4tYagxR
vFNXzfk91exVgiJBkXK5j3duoSp+Qf+E2+4IlCrTeGQcxmqJV4OePO4KYEu5iH++
hgrMrieBfR/Fp+8mY0Q5esJIF1cSkrZr6/1OZJzGYLbvy5XVFFmHrv5QilhSZ0rn
JoGa8xxBepHl7eN78wwAHhUzjCu3eriA2B4Tsa+BcECrraxgG2CD1ALlIdqBiNhV
EFngZDkhKvCgsGrKYLJZNcqBcCsfbzj2uO2QDz9tL69KVwS/0EYhGySsCcjmnPND
Mzn6R0ngEwzVft1iepLYVPeOIPQgRfFexj3eSjsi1M4cEKxPNnRKwc0Uew5ouPcA
amDtx3jj9QsYYjYl0u/ET7WARf8WniT6uphV+cnVrUEKXjg+KXuCH0YjCui8ia1H
y6Ug5z1AObb9xento6IZ0sL+T1/ViZXJWm4dlwpT2C9AVtiEi8vpEV5QvQa9s50c
T+H1ON5j7bG0htcGXF1swLdbeWr4Fm4BW+jzW52/F8c0+p7VFSfY4Lg93QT2KccC
wUPYKKdWWjiJjwHuy+RoMRI/wm8yVmwQFL1hCfq0AHq4y39/ZCvBEsLfCcvzB9de
S3RZ4cwWCPNehDu3kmdD5qvOO4g3wvgiIp0iiS0wU17RSx4HtJVh2RgGzQpPfsrU
DzojjT39NNqwiKtglilfOXSrCFavqQYMC8fzUfUSVg9Srd8OrR+Gg+osJUl3fqkt
HL8tApRji48Qz7mSIpDlMCGNhihA9rNbcfIylo5QLmb5RoTU8NvPM+s/2L42slpR
JTwgIT9X2aQlvoakkH6k2FHz62Z3klnCfKotD6VUvcZ22jKuhEYKzrDDbSn1xDl+
INo4W1dNVTiFKFhXOKmiaTYd0YLi2TKbiJbzbTj9Y7syzcr5nw5XO1C0AxzmRK6m
YFstPbRnjfkDni20t47RjuDUBmGfpC/OCJd57PdeGc0hpt2ATx5j0bB+vj9mPR9r
mccqlBW+nuCG85mLzmqglioSpuuLEfmugFbVK/fsStWEoydKA/dcuY3oXKrTHyHn
LaMfhVk3oQ6Euo/MXd3YMvyISsCJ+KrljxY5eOFEyCZEG0Lf1gUc2Px/gKbucYeH
c55tLo496wgDzG+2Ws5f3i6rrzszGIlWRFVySRQROr4xPd26u1CHgF+ucwZpJRmd
6CrTYORZnDwijCnrFQIyzMBV43bxTacskJ7BJl/AmESEBKJ4SS+Qf2sMIyLvQZar
o0OqjPFtNtKHLrmmNMLUB6HhRLeEoLYDKMPMrg0zjZ9hfZyq4xCnd1E1qaae4syS
SsdY1ZTsGeXFp+hYCWwxQjRiReWKWycL+IzC5BfxQN4yZIhKdLd/lmt+7z8A4UiZ
69z98gW04RiCocS1emJO9XJDlXXinaaePb2xETyjQjRn94xneXA6pCf87A9MNCG0
OHLdPdq47fS3mfag7GMXKQ38L1LCC0i3DZnvD/XS3EbV+wHZgeR9+jNgh/1edgSO
jpaRKmDjR5pnWgoRpydSgxcIi2lHhe85JOQux4tR2+xj0ZrwHWtL+WSLXdXfKWVU
BTZwX73W0FwBNEbHSPnayE3TfEtPUPORolyROYVfuhvDk/7Kmgxd0dxxZDXUbSpJ
RPpofoioRnOtAB9qYmfLyAbwAa6rOLWKoiOqnYa8xLw3rbWOQnnh0vvRZI6hLtmn
yLF/yuyYgYL8ID9pOoKkbZ1E2KJ97peIvSNoskvZKTp88jwITlC+2nFdJKhrNhYX
Pf9EohgeXjuhgS+ewjVrq7oeJPpNxsYWb71/aqXrjuZE0BXdv1IG2z8emJ/rRC3J
BJZJFNTR2lsWRtwD7pKXunqRDT7ScnZkG7VF27SVduDR5K5sA/ifGpCtFSkaBxCm
3LgSnIEqblYoptVWNS85jX3Xs/oQVDFahjd5uNpygDLLZQVYxp8SFrrqIvBqENPq
h7t03+PPbO+B/4+CBbSL5KwsqsFa5BYyxyPjhjVc/v3zh48aisjF4lnCx5UsDMmZ
uwXrP4IdjSw16gh8c18aL3RYpYnuDDJIWmMh8kOhcO21+Abc/QWIad6H4N+WCpK2
vxFnJY4/yyrkqEMj0NXWX8cro0hDMAGga4XeWwG9Cv8ZKrcZ+XvUomYpI4I9ki8k
EYCk7W51/KF/AJdcoWgG0yiWQ5lOMdp/w6HrgQ+olI+Y4VbXFpAnZB1cC5IpictB
r2ZHGTicFF1ljDMM1S/1EMRV+6Ly3O2Btzo5h6fkeyLgdWChHQRIIVxbIOKoP/ds
SZMIfAv5dHD7gK1gN8P+oHJIk7U5MFUxaF+jvvnWIEX6f8Rw9WH3cPgIAWdNVo6Q
sYPQIpfnB7+q9xjaZCTdGbwl9mLl1v77Dd36UxjQKbRaJa33huLcpwwHtZjsOJQI
iI+gzBLr5dH1bu0Z1djCQfYgdWmpiknkiFSAUzNjggTvR07bxvhP+P0HrqtmvMiV
4zw7+lZxS2Z/VhP53S0VpRlSsGsSzrhlof1inuqzr9TGDhH1dXMNuHAuX4pshBRU
9dOYuRmCDbQxRtYLqaiaGPmVCcOpXokZULkY76WlWucZ21wjgBMu4cDJpnztjPbP
/6GCKxxWovr+hYnPK7aOrLvWyi30q6+Lo/tLaYDmx2GqCxjsgUc8diUK5FXBAf7i
WJ2EVTR7ccqqOjMPFWBLFOlR/hrNWzKTg6BtU6UDxJK59rxT+hzCT4b5iHphKDl5
Fo12iB+T6dJMTuPcTfGNmHQBg3UB2h3xBwy2oKZ+GgZMfTWUDGo2/osZQ533aCxe
1CJ6j+1ZdZ/loy9+9W2SBUmQDetY+Xa//A3YQI9tmSh3iJRedUzf7EQgBKk8ryxr
qbRdO5f+jPJkdHku3KlBXBMabFqMdM9d+BKArKZbJ2Iaxl8WjP9RfH1tsvnRDnjw
iu19yv3PrXzNDCZqmpzQyoWXV2JL4ZUNIfk3Mr5SLAj23C1NSk2/74tY4uHbRwF7
eIgvfq2p5D+cVZ3gCmfIvq0LWtXUMXIDinLczBdV2VoXNupEzdpYO8BJBQtOmObE
Y6d6otKuPpOUNffhvXw3rldbtgyYygTp5C9jQl4WKlox5s+TCqZPkllb/k13jNGp
MdVq0Yxck9V0JLlEinx/fWvWuyKyc1PZiMTodpX+q/ZnvIGS6FOMjCf9YHfaRBJP
EYgGd5na0w9JalDDaYxrb868il0yzdnidmdPJMOq+0AEuHOrAaP+EkVo8V9Fjdax
3fdTFVN9MSBVcnZfV2WytOEjQoIzOE/GL2Vk4aOZRrIJsHJUZ3Q7i4yfF1lPMXnt
3N6keXY/5cLLv90ACWCETu0+uSdfwhzeHeJOKIhMsIR0F7WNx5q/JETCu6EkuUBX
YgzPgA6FubtVYI/9owRpxHa5b2ER5ltcQoRGOdIIxT1Af7/Zq7c4QuiGiRA/Ez02
JpPEO3naRbHUttNzcUIuMsFdMpUBOWhMIwQ1qkjKKwA4Ac61ndgr2UmW24eBi3y3
AMO1NR6gCd1PmHoBnPtTCBFq0DShwwsTnVL63JZcRrgv5ebye3w8AD40zwHZ1EnU
q3md0cTVv734Fv4Z73sK6nA3u+D8BknJOW4MatAbFa9GrH8+8mMoMvgRJOoR2ygI
VVjZiQEvuo8we3OP85rDoGBdfP3XhFRCIZNl4wYv0u3QJrdF535KzCZXTu2yqfJp
X4nIvkADBeEPB1ITqfZlqKDjBAnEAzNZwUYGm+I2FzItQui21fr3zG3x10fDwBVW
KvRnEhPzZfOe7wSV/X9J+zgfBXkm6LjiNE6WvFNxRwJKDdXG58LJrLYZwOVIVYV4
ELlUb3hWB+PpxmKv/+zMeKl3IxhpI8Y3CVeDLgPfz+c40mPXBFUJLBOQyMhfS5+r
OCmemzhF/LxFZrp9B1BzP6EIBrR1yl09UAUIX3/ca3pp9W9mWKiUQjkit28l+OUh
EP30WmxsmBEmMoskzUNCVBrbNSERzO+YFjDdKXvNXrHYm8CBgNXKqBEoJybKrXXp
Smo73NsuF7FGmoNpQ70Ltf9jLikAW97fRVwrfv1SOjCi9Wnd2idE9wB8GvoT7euZ
EAjK5HHa+BnVEt5H/qUIOmAPJeslKVEXCPksuW6kOOB3mnOzSw12M3xGk6mAUUpX
HiYPdVCDze1NLp65xC3tgOaXqNdaLTjBpXsjS+0ULLsouEQSt6R3GrSL8DSf0gkK
7jwL59aMvZLgyrGr6ozwpTjomPupsAtmGrJE3d6uc6Eu0PpmLIt053OYRkUtrATr
1t7lgKhN0958sIPjtD+0vAur3yInWsa3FcJptt0tqbHFjvZ/xV58nukb+of9f1Dv
MUe8fxKIJGetLTR4qH7Yq3GikmpPnrDjIgzhe5usQNOGWYXCPOmn2AsSpOUbuYub
osj3UHr31XQBmppqqJpATRdE9CcT8uAvxg39r5kNm3oOypBor7g6EX7tCCgCSKBQ
N/0s28mU9B99MopLhyuBDo/ZT+zVHDEvS+jcecuielIAaS5LtbH6RhSkJ3KRPMDx
bYX3i1xF1aEDap9iLr9i/cPTGXwjN3e2SjPfQ/wM1d5Ix/KVjeUfS9XfwCz+Mbd3
0qey2GYzPGWiVtt5LGVum4Z+bDvKWIXsxhY1y430BJ6tscsXeaoUwH4npBbobvN3
WT7HhJ1u0GIo8Yh+acD9XvGUZ/0EDepCQLIPXu4XH4vr6yX870XFONefapp6fb4p
vzDSS6DYphEWhEXIPHxIUdZrUs5L3TW0J8Mu05Y+xrjiZ5bPluBR9GVXrVOQtSSv
5QURyVV5yxfCX2qMGqypHLN+eRhr8QlocVvoqNCMrIPJkX0K3Wd1ntxf/V+FKPSb
zEAKubyeKoghziJIQqYrEiphdl9SPjuavehcjXtWQoZR5l2FaL/pOs6wQ8tNvU78
ZOwe56++CGlcHp30ANs5U6GJpPhzRoWydKS51hDN2x0LF0rZdH6bMQoP+WvJNKXX
Hk+3R6sTSx15wNfjYaHhuKhXHEjpRp6QHmkm8sCdh3/U9x2xEM4pV22RSrSJtjG1
+2YhSHZTj9RvNhtX+kvOVgyqNsxxj3XTdBC8uoYngwl7clD/F8paI/WCe52aGpkV
aKmveEEkzoBkzKeVWmEHdABimGgOtkrd/IDUcoNaFNk9kIWR7GUNpG3rQMARKM8t
AstYF2vatzPBMKhr+5rbFXKubcHQM9yHZrm8TmdYKi6T69U4lU28hfhWV4V1sfFi
/K1GtMMp3P3xib0ltb1tQfRSI3UfHVKaEDnnNXZsL9n7RK0vh1kcxBrP1zq9mE+1
Mhuxa5MQZJZcJcfmDHR0p4BLmyXY2RYmrg3SV04tUn1H7ATX2CTfFaymneRDXlQ2
Z/N9gIssc6t5BSv8u8irt/ibK2cdXWkjFUqucTKO7wuuqSeSrY7VpAhNyzoD4e0V
UHtPtsdsyzx9sqmsXcGdg9h/Uoaj6KuZBkn3nmDhdM/s9zILL9uFLOrBCTg4NZPJ
xwAUHzgHGMCWi9iiy3bxnkirt9OgwjjZej2OzYXvg/B2qIeLX3K/EaDH4ie0hrCS
L5v0u1DvBl1m5LS8yE6KjQdINiMzUuIaQRKeDw21LS82ozLAyM7eF4CPyGCU/Obl
YDTnHaTi3yAWMrAPDcJHcxa2bleVgrMvn4KOWFDFfDGLQu4kPyL0rwMxoGoaRzJ/
TF9nHqGdaQfaDgBlkB4Ow8/FrPIBuUUydiuU2T+oC+CMFdCFqf1aDxJEJJnrf3pi
qddLnVUL1R63Vq/lRxlE6hQmKUPP7Uzj04JWiaLvstldt9HRG++yVAZQJ55FUW/W
xzjK1pf2iN9RS2LRnP00ZX71iMYQAsaEo0Crb8JHlIw+/+FwsvAS3WTFvarc93N7
UvRHC4UgdnwZtYrwjkNrfhfjdJmto+Kcefjv+6CNC1uRoOkbRln5PXuZ/IHF9wPG
0Pq36oGHYIhi7v/U4gTARbShCKWqeCggpJJOccAl8dU8B6y6+HBLbczCCSCJtnth
a6sQQKVPxxnl3vYouZSUayJWj+6INXKv9gmIjbjoLF+4ryhS96xajIJLU55oQwIA
Qw3q9M/uDrjkS1BDg/gWMQb0EKPBoNeqGXbyoQl/wY8PDMua5dfLXOvhZPg4FVse
5CskY1qJEQiLSF8wvtaQ83YXLOGvwYdmMHFSTjsC8Shs0h8aKEnNkBpo161tj/30
IOfqvt0pLIRCWYZJO+UL6Bkv8rpPzYcMPnp1rfJwMKWpCkqjjbeOHbwCIV4+PQUw
L0oHS9X1uGxzSg9Mx7mlo1oJL/AYuWeacqGG5W+M+FxGasvOiNWkWxnWTXKturbP
35k/ZpRXFWnvNgiGXIMoiwYNFFa6wbRHaRr0lofD9gFo1XLpKFXmsv0+lXeT9/Qu
J1INqZtCUNjsZWRicxKxuKsYKoYugCdwEA46H1F9Vls1ChUjgTarNhpvB6A6fseJ
5HvcrTKe9o1FXUSN6Q3khKQnjdnHmJgjPDBB9JaNOTRC4yBKNYWG+3e89miSmIQs
0cW63kEK5fa90bygUur6bFYHlxWLabEuduycjdKf045/Qqmoeb++cLa4/jbLisBI
1xVhmaEK9IAtBuS6FSFppoAKp2ogq7XIygHSKds6Md0yK3kYQ3CZrzXojQK1hH6Y
K6Q5GRtuxlYUXZNrJsFT0v3loyYpsc/oWxLd2MSfoY9uewJ31q6wb0QktitM5pI0
Pl9p8VwK57ns1WAmc6TyOY1BMqx+8CfYMQOhZt391j1FW+lm1NZasVrUSeHPORWV
IcunbMWlN1l36SOO2Uj3l9Xkz6QzN+j2nZ8kMzh9cLKnUrhoqKeOuOSvVr1kHJhS
cz7txKQoUZk4am3b4oyp1rjFIXQvC20MByEb9tMqoqeIl1UaG5jWQKdo9iOPwHy2
jjVtHXuubmoDN/XlRGCgnuAdUVdP1Tz0s2JYBvAp++9YUTzjX3qK8pnsGGP4eV3Q
nAr8FG/CGM4W/0laU20rDgLbJvnXo3xxKhq6gnd1gw1/22WQbqNrRNBB28RKNbM+
hWHvQ6huINatbn3TCe4USG1UOBT6uMkCEbYN3KT0JlAHOSgMIlXdgKf9ENMeIC6U
csQwPQMCH4VPlSptWGcYTJv/KyLo92JFTT/IshDADAxHOqcJS6FSvw2dqY5qJX+G
w1Sh+6lsDmP0DmTGOzFyWB926ZrcUpeN0YzkInDxRJ0I5pcGG4vQNcx7n0hS44Rb
xKrS0GHk3y9xaLbL24EvKpZgz3JVt3IuJR57fUZtRN2t3H5hbHH0vtgOptSeBiPX
zGkNJawi3N7xiWDRRucWlIImOX721qFaPpG+1kLV7XjvvYmaQdVmdWk0hdW2gviR
r9TBbNQMtsBT6MvHvMJsRFf7AKFQ2+op3n1tDVe881qsGxdoHWddog9+fqEbob6N
iiTRykzFGNNuwsFQ8/8sL7PqOCQHuu/BtflxNh6KHCrHSPWabznfi7WSh/p7sox1
1WCbGnTpxWf+1SZjJkdoxP1qvxCQqYjaeDrlTYJlJD+m8G/ig1HFPublymfHcuXH
gxn5gMRGqh8zeb1JSZRlfpaKUeQVgSXr7F0wUn82f4JzeJW0UqXCxbBOXvnAw8Ak
y9y2df7FzfA7H/ZRJQABV0I3aKEIVnazu8SWkXO+4Jogz5ML5KlcRQe9WbDelXFk
1UWgeMBEGg38R+aIkFL5M0a4X3pT4UbPwxfac2vogvNfJKm3vPdxn9rMFIVGgzdT
Ldp+UqEMUFE389ps7+M2CTa2Pl1Ktvl2V4cHpAw4wWfmVqfkUfV1670QUYz2wGE/
Rc8eBBwbbOjEEA4YlqdoxhFfadRVqmzEWXDx+1bDbgtWCIbKiKbfhmJNhdiwHGc/
lP7YCHV7OzzRZS0Ks/RTDdtSyFn+6fpagjH2/7lm+ag9p7WLCGHYuMOvTUSoy63w
I5EV1puXDS3oL8gqxGEwJa8/TGwKF3XwdsZ3nd1JnyeMnMAI/hI82RVqHsSjzIY7
ZQ997LsYIB/FN9YmnIGr6qHiD0rbjJSgeQohu2Va5o4XvvKNLCr8mBhRv8gnthbW
ciHb1Ai6s6qmjN1ZlXpjBuyNReePc5DpZ17QFx5WuoR3Gb6VPxeIaL+b4F+lDgo9
77rASm3JdZ7rqUKshReOgvX9h7ofTeOThcZM/CdUtYYYdyceNL4JlFMCiHFagCPA
VfLO+6gijY1qw9TnKo1CFNYJ9mT1GBqrjY2LxZUqAuf4DrthXhN85NNdw6yHE15e
+kroXrg7R6LO6MDQnDTURFwyXT6AYea/NxB+EAl22adMfG1V4SJsrbqwG3AU0Qlz
rHM7Se9SxxUcyjVwe8XkB1CIkkrqMe1RmdPSUDHSKLCxMySrPCO7HPnzaMqlNT9m
NKU6bUV+lXNdJmke9dQyKXyMbMbRyJbZpuqYzeZXp5onwQU57EvHlksiRujF3aIl
4lBd1CaCPwGEgdpSdsZOXLD9Y8fPSQOy+NRotN4e6z91co8FGGAxHYSp6LdTyEkX
G/FWDP2kd8bifF12oKFAENWfKJY/kHCewL0Z1DJDPDy8EBmAwsA1FrYKJhpeAGVB
He1qOCCzj+z6q5ASkGSu+MTlG9eKjFx0dl2/BVCwJBIiWBN/dxBOasdxKQ96IXS8
zZj+2aM4Vh1R/Rv5au/vp9QYoVOdpUq88Kj7xMyWrgC9Eix35N+jBbX5Ch9tG+Ol
fXazi3KIw6m914of86xSn5J/gPGu0KmGsgemETQnSZS6heaoR25OWXpDZsXN80YD
VaxTZ0BK6/IkIetWAbWGa4hqXMYocjo6XKipJzw5BA+nxAgC/A53mC/YDLa6noAT
Pd1q8bPqQnd9oVdLsBNEKSP5WGfFCUSRckwJ+X0xeNprTfuHbN+kysxL5tIyjxj8
vAHUQfftg7wvKzHZNwuWzRmpDuaiS7LkaPDsBRt/3hV3fmQlxBz+BJa7Kvi5SYiP
6qOANqvwYpQY4ykxhGY/rB6d5kZ4lmSWKe2jNxntUzQI5C69ZVCOz0AEq2m8Wmui
/iPI0mAwuG95h8RyL2sNfoRwtepaIpgObkcg1RhQ/rXAD6kDEzs3HITWE9CqebkS
dXtFSg36iOoTWI3NKotleVBKUOd+P/8ldbVbH0dg3zSAVgDPy+LFp7b0HUaT0V4e
tzOe4Wvf5O1Ju/s3MGpJM9GYrXcoIQMZdDEOSnFRmbnyXdmi56qkaywb0r2VYvc7
/zB13BPwetMaZNj/F6c8BvoObh8737EHIK25YWxtGGvx586vlnLairCDIcZk7dwm
zgEhctdjx42jXqhxzrZYyYjhqqGGOMkcFdmB2fFurRvCDQuvqIb+QvSF3VnjffrV
i+yBwWD0AisvttsajT2PTEQj7N22gfasMIFuwwOyYVrLgdlQuMlAxlXGM3ZWPa78
8ckCoAf1pJaeYNG+kjFeaETAlnGSMz6gR+oOaGlKyqEKOH6GMTXM34ca/h3E33Zk
e5qf547hb7iW6y/CUKsuUDfh9YMhpli4qY4zAPCh63AUmt/DdZLvw4XznZORYLPZ
xWmgUoXHNB7Dotwl4RN7h8p6fRcA2Y14trLcGC6/tB4FV0zGkForxu9QNmCJRt2r
VaZLzPdZ6jE6G/OvGhh0ZNQcxqK9ymhdbFyFN3tSi6Vyw+WEdAuT/3NMr+mtRVQV
XDaPMK3YHwbnqkNf6F43zii92JCufrkcOiKznfgo1HcWYIqu1omzOLN8YXEledbj
vS63kKOcrtCI5tfLoislcG+kZJnp1lCAvNr9DyAIHLNAS8OYcSEeak8yGuw+5SLC
WnephBlzxi8NNWN+IZvGbbVgF71A7iWqj3AgYeKfdRB4BKzmBcmoU/dbRlDO/mo7
MX0YEFMXuK/ymkvHIRzWlXAuQYgbt1Fr9e1gQQQTzdONYD04NN3qNlyMKuPhpnGY
MT/iqxrzAUOta/M7GcSHG7jeLrY42tUrQxg0ZGUZnJGcqY27V1ePsP2zJoZVJ6s8
6WCrInp5yb6A6yYfMndaIwRvl8OZBOex0cgEeXosvGnTfI1xihnLas+ASMOXiLgH
WAryH8tlQb8QaBKIFEbOvp2UPiUycwDnsy5XLMk0laIKFdg/NNwn1JQYSHpZGUIY
lQ1z9KjREwvlzk4xOkHJIsS6DwkXj0i0j7N5onHmvziWa4k8WAcbAWVCRTpjHTyI
1KXxQcdn37Mx+puGJkoESH8U+sExyt9P3LRUU5IxU70nB8P8zS5hLnk2DfVDgHUv
EcGGVaOkucWgccGagpeSPgpFYRGiaxUGckBeuGsxSz3TwBGMbYkUapO7NMjp58k7
vNtWvDfEGUZxA2FUbNnABBni/noChcaAxc60lWTwLvOAUdvAXOlZJZC5GAeot3CU
LIFVYo7wVC8o6MGZx7FOZiuDmlK18e8U5n6KmT8V3jqk331XHSDA+N9mJoqrS27s
Kf/jptMXXr2dMBZunb0kYTJ2ZPoOhgqVggIbBI3An9U3CLU+5Id+ODv9n3+vLyl8
z3w6ipoYn1KaH+tMXQsZ08hFew59QPDvWISlQ5Omy4Nc33kiEaUvMtcaWj7HuuDN
75Y/90mFqrrLEmX9kbNP1jyKxa616xv9Bnw/SyAZbPglAmxf6KandvhDsxGHVHYR
ibCOoD4rE/rFIPUfwEt5c2mXc0+Y9eV45AegP7/whRBtcu3vXh5kUPeJZyYm+hiC
puFIo+Mcth5j1DoY7/53abaW4ZUeuCt8CwVYq6OSYT3ofYdMqNp6thRuxfAnj1+t
QErHSgs0XCFUBNQxjq/X5EctVZIc7xpE916Th7vQ1q2fq4+s2OGyylRYeowgLAsE
1mndFyDw6q9tOwW6c0+lmBSotLL7XBEg6e6+kfx4Ste7kbfg17FVdeIFxbr3743T
NcoGarixWyeDEHg6c8QafmJ8qMq6LBgR71woV9o4VILO7i5JUBCt1v4OmLG2e96V
983cnOJfAvAVN2soSoGnYEhhGpOWNDlauxIckqB9ry9P9AA1Rghqm6NmZJGmuLkz
YUQaqMAb0mpd7xgQJ9qzEc8Kstdw25cLtqput8fdPRfsaBuOJNcKPrb3WMr63Cy2
xFqk6fZn1jLGrUTA7L1xilVlXZT7D1LEhSLs21piPhLVuVG/CmwHkA9J/ntTUWIu
K/iUTK01DtkbuKJmAb9m/nDlBHdvDcDL3nfYjKrUnmJsWFlLMe2OL8Nni2JITcdh
BfNQyzVgQqtv8IIekzPGpVFltF3kpt5UQ06Js4KkRDrk/4yqOqjH0F5s2mmv+ErL
PjAs9TykRBTSBW2jiYCzJgCRKTmwgSJplP7bq5+jFYDiqYMiu9TQIUik8cMvBFj6
lDQ/qxzXxEmuvTgaOHVTiAU3IvEZ2z+UjsyJSr6nCzGtfr4uvLBY73+Q2NB8En4s
iI3KwQH/6uwUMv29k5AL1PLke4HBhDqVhbI/3nOdwZOX09cPOHEHKv+KHo3Ux4SS
HViUZASPvd7tQqMr84IqYrPFbTQdFPkGzEqhlXSu26NtcAa6iRnsUzQXvNv7O2G4
7Kq6/ppsDLP5AkFEKmW4bOyK4kYWgfQW0HZg30f4PtuFO0PPOZMNVE/8gqB5PDFb
ttHfucjXMX7iF9Z+OFOpwMkSywGXKMKXEPFxDHMyi7bJ1qbsFEl4tZsvZP59PHSk
36bamVlBqC0e/1HXhhffjLXIcP3z9hqQl8lUKLQjykJOpG9CRfpqb6yF7JYc67ZJ
emd8S9haMwWVSIOeus9nYN5MgxboR5I2luaA1dbS0KYxU0ryuyo5BpF8jOhPTuNb
YsIlqN2NgowdrT3kv2W2gtLP2U8MnDCC5JdxaobdZHG93h/+w0Ql9YoOX1bT/lU5
WLGBjDTDWb/ey8uN6IYuDv7g3mPVJZin7PObbjpZRDSYYBopnd0m2m9QBvAgL2ek
4koJuOs5RtuUDMoPT99SD+YlAEnvCC8qBQd9gdW38902i9/t1wRuWR6mhJdCrSY9
Z2hJ9CcSn8FvA8iqQLz/DNtAGHxnZYhcX9ESBYXmupEv9kpSi2eRjuT1bGghDzWC
P2f50AD7XvDrM/Jo73tTaxCOR1lQx4LZFJSjC5kJWMZgSsIRUSoZJHt8J6s7IGUK
W3hsIFWd5DJcMgEoe5SKikgmQZQ/k09+G1hztTZM0k5OyGgfsYvfRlNHyLxKO+yS
tqMz68tymUsAZNMDWcaERJ6oglpB6rAI09FBXO9NgzvaqtI+MZfiPn1jn4GwRq8d
gjASnEHLOnXWn3ark5+sdsSTXwKPhjB+FwHImINhuySyTQp0Y3aHC17J1TiXgL5U
DYiWIcKAo8Oe2WsMnkKx5CkMQukGIdcfc7e8AOo5DZT4YH974M1K7ajy/w2OnR7j
FW06z7CGuZqkDrkSZFWfle3w9mWDY28uNl9Cgu3WoPZp98+uz/nyaaxq44EXwjcK
rfx3PI8ONsNyI+fS4N6MDqcCdKNOqZDckaWnYtqB5qm9GPyTUoo9esIUGvssqj1s
mJJW1ROSBGThAMF5qavnVk6tZClja789b8WiDM9tP/MbCAw4Z8042tCys+F6IlhR
BuSXgrjBBOsF3YFHZ7NJcBkzysGHN/ADZ2HD+SVew6XxlQXreEFAjA22buisZftG
Qjr+g9u0vovBoq7bSdVEc1vkSbKX6I65wS7cZRyUfQhK0Jo+WpW5KiU6FlNejEus
vZIlinVJV/fOEwp/bsJsAP59kDDJRVy+Z+iBkilEyq9nv6Y60E/BJl11wIxT6mvj
I0DZPFoTf9EM2ipYiuCYbq5RSd4h9ho74UfTWmisClj59xwQps0VGZZHhh3KeXgj
GaocGajo+fLqiFh+noPTwl1ejz7xn5OHwJVTYf+tjJjQijgSU8gtmIx4PtQigzSr
iszdPnigxx6i17t00XBYPsJQjyfSV1DT8RL6uaxmRoxUta2DfHmyHMG54dWUKlIq
Oa69L4isi5LO/N6yVVyvAtzjdjGX5Nlchawo2ar0/8GQitnIrb6PpnzCAmkfauZG
VvSM1DZNlFX+YBQ4cFDk+xEVJ/MqUlxTbMVZLR7LPCiFBNJ6/AcT+EApCVMlBsZ1
0UJKGPsIqMfSdPo+iPHpUan+Fir0frICkDCErsMlA+wgoWLMuaGpV5qXpgPQ8F/w
2Rp2LFBWkH91VW2rdxe3vTD9NtWx1CNME599ljKsrwV+zEpIAdpPNqeowMyic6KZ
FO/ZkY4pi6rK2gKejPQYq0/xuRyagN/LNR2AM95PDcIOWqJZENfOCFW1uOF+vyxm
m+icbkTeU83h0GW4kFD0eTlNYWj8BROceR+R1vuQE9xGVta3nvxHIM5T6x5JpxiD
+M/Ph1Y9+hSp7qPfw8LGB/8aRD6xgtDjqeeeoGXfgswdaZtmR4iy5MIdF0r22gT8
zs71nPLzLVML1R3i2YLNsSMjR0vYjSMOVOzOI7NHemt5Jtx0l3S1OlsSr81Ph3/I
K9iqUqJQN3NyBltvhifBFf5Z/ydW+aQfOT2M2i6HKtbmg7otrz2OSHfskxbFl8MG
AZs/C11kpowHZK/WQvTEYCzeHGn4bgSuuXVyFdKoJsRMaS2ZSJ/auNuGbMPLqh1J
2XI+RxzS/oUrYSWUnCZdyiSll9Hil2e5HHFpexZezlza+Bt7aYku/5ogsHD12I2a
Uub2aeIevs9O5iiOnwKnhJMYkIsI6GCmSm2cgfPZZNVrS9CWKuxKVgtgLtOSKtZl
vsLr3jlsRiU4FGI0hMRR7/FGy79+ZH/71o8E8YB4G9pFJYp4ZmRTUKvrmmrnZzJi
66oaAv8471pZ3qW7q3V2BRsmn26DBFmIlvcpgCI+FlYQH/g0+GvL1LISslf0AMpq
eHqE/3SP2l31H5S7Qovju4tcKbkfFhU+mHYl8pR9XXfFz09oiI7+cpwL2lWrm4Gl
XPK86yEjCPPEbp1s+7QwGIqPpibFAo3Ywtk8uNdpedMDOd8A/XMpECMxxHF3wJVL
gkJm7aNAEGplUUffVdwBELeg65GDUXYRuNhN/5yPk4lrrnBgeOcDRMTbPPxz7Zsj
l+aRJjxc9DNwaHzgEIQlQ9aJvopkESSQzRmX/8ohZ0i807gzMam+CUpS5VjuSBy5
ds1l/8tTxtD8DREuh8lnxtHhU/lenuvaen3JIVb3hdjn0Yt2ap1ayvmpKYxe6MQo
sfWWrPvVaJFLnQyEoTcSPIT6YGZ6XzuNVmX2Jp8w69TtSHUGed2p7pZgdAh1/gXb
zbq59euclrO9G7cYtDa4ycR3qZoqWxcFxcSUSU4042OfEXvYsJKNhSFnUwtUQavs
Phbkl2UpHmr4ra7kEnMtEqemyOx57ifqu19EAMir4ZkgKhigXD8/r1kA6u3OLw+8
f2ZIxrX3+rA16KwF+fq/ZCaTMP/02Wl7gco1oK6MRs8qyjxCdeZgg/otGjYXi67Y
CzgnnShM3XHkuP2Rma/GRVEUH5rIVK6YxIfo0CtqDphgV1b9PRABV1qktxmAV0WW
UE73ueVUfkfyQ9Bz7Q7jTiHhRdPPiRaxNywLjHbnlhGuC9b5IBXyTayy4ARQpNyP
cXhONqBREKG9/LDUUtC1Go/HlXC5fB9Gw/e9/EMq+UKfTL5VszVFjbmaij14GE03
mqNFIx+CbYzMHZq2sNI/FHej0gq1TOE/egFzlwc9q5nFRcDtgFOAj300o5zHRmHJ
P9ChcG1wOxke4r915WFuXKxZANckIpydLmYZHfThI5afwwxgRjmR0WK5RRtvtcvb
j7qfSvRGM91L92cKDxPQ9VRDft72gOJs+bEB9ap9wvKxMVhmCQfchpxsnCfmuJm+
ZaZcxOWih0iixBpO0LNoiH/FVIxpEEcNEu09TdsV0y+JpzanBTNmS2TDLRigjOxu
QXRRKcXdhvcrVq4NRLR2UZiqIeXtpi0Zw9SIqOGxWYUbSbDGTUJCZRP9tpDeZsIz
2EN0KaPn+A8//AIgvHLXyxNw7nhDU85PKxtOs1gVM22L6hK7QwQ4SpnZVzPP8uYS
E8B4CEAdb62RvYfuNrkWqmEdor1AkcubqdO3nJ3gyv0+sdsJWAtiHfF89swbCXgi
BEv3XaUaMErf0H4lr9bM2++L5bE9XOoTfJWZu73IiuMfS0bIcUAigPIFqsoVuOW7
bf8gLj4uqS+3ETDA4fuB4Rf7mdIi6j2v13FgiPD2gDHHc9+zwEB6ammgPS9cQSwn
R3wBE2+PNntUyRHvH9J6RgaujqCOz1rub2SOpk2eK4tPzLrOTR44VBKimL1u+n2Y
oxwZXxx0h5BhTV0pxlAg/17RJyhEB7zJ3v7otyNeSuNk0cS41BRksxWG/y+hbRXQ
AJ5BNWnbQzOz/vDwe7+0aSZDQoygWdcR4gLPfxbFopbd2rCBe4rOvWh61m2bPZJa
YC+ReoZAYtAiMAc0CpW6IEaK7tZXeZ+9z1G/uL3cSHLHlETS5l5Cw6XPNgnkEgiE
Sz7FXbZ1Bh6ed7frVdNy+If2RQJMgW8kFUQbNBNrf5hxhX50A2gYCDqt+oDffCyK
N0TVJ1IfZirxuYI10jQzvTrwmVALfyoxyNnlZc0Pg1B1LE7Pwh/kA4SharYMxhmV
BeKLUWxoglXYQdhrLsZ25UZXhDE5RfbueQGRu3eHUvwdrF4mk0yNviOPwIc2CA05
nCq+NEbQlVR2VP6QbaJH/ad2y281h1bIiAUt55NR+Sv816KxOgHl1NGPz7xWmSL+
p9/xqo0bEnx0nrP+bF7eyhNRyQilXZJ15FmIlWvYvILqyk67ALWUfGMYbRsSOolM
1uf1JmIbX4+r9yyWWeWhxdoqFm27hpHc7CFck2kgK28G36gDjrwwSePb2JTiCuJp
rSI5pwRnRuUKf34+ZNB6YrG7vd6HhxeruK4NK8kPYWL1f8cEHC7cUh/ECzhwhWU4
beN4UY9w0Dt9mE18udi1bdmf36eLjJO58eOXOHDdXz/bqyoVQG4FU9nOYTkP++AN
VHg+7EePoKkIdRxC31BIVWDpbECQCcP1kkqBmRG16RL8dVNtMuuIZ+ufRv+X7WNz
rO+VxK67NvjHQDb/VlFPTzh8Vx+yo2C1XhxFR5V9oxFtSO9uL22v6Mab6yP8E40v
Ql++zAm23nQsMkn/Z5pQntplTypKh0sFTCGOCdZsUjjxjuM953n9ML00a9jX6rOC
a0UZk8nuWM+WmR9/SuzVMJtY+WY8tHJG04XG5FIBUfVjd3HMF8RHr0fJynn/9jA5
zWld+ceJmXgi1gppyESHpMazso5eonK7mvsk+aev8LB6RxUie/JBGcJnp/cng0Ib
I0nKWsE5wdMrZw+dzJ6druFOt2KMejhYXmqijc/y/5Qrs89euptXwT4WZG4eVaN2
STo/pRseuWPmNxzXNQYtUAFJpypTOtSVQbLvcwFQgeQXqVwJJxxjs2UcuYu3IOWQ
1eoaqpDJX2KFOQKw+5JX4bEZNW8bjSPpYv5bdZ/yaiFJ30jMID6MFfMV/SQNTJDw
9cCVU72XYULLmMRuri/jCKhlBDoa8nPXLPI8xvFrHI1QKEgav+2vy6WNFMhuRehY
lNSoeSURafAGyilnrKdu/cSzlBih94iVsqtibD8PgpFY2k6iDyaHro+KV47rckrW
q+qwce6fPdoF1PtLG7Av6jcluhOr8HAcZcs4nk/vAolw7m9v1RSXbQg1HIAak1Fb
8WB0RFe1xFsur+5DRhQvgG0aqvPt/7dswdMmNuwEMgHIjPsS9HVhIfwtWKcmKkue
IrfoF+ZiXvAE823Jngv1suGCF7OHagroe/v2lwo2Lbq2iodEM405gp3VUhRdVMKH
c8FMdL4SpABUa/KrvX6yr7xoq/PZDa78SZlIiV/pBEcSIJRVVt6bJ2xZK6zFX8aL
Y0P4Jyjq/j7NwUULsDnioJRiv2IALdQy9CgMPvPtNFzJZhJ1X12ezqrzS7i3dV2P
HpQ5DnUii/zJd7SvuYRcljNdbJ1bJQTIHuVuOSSLGz5tO8bZHEWgbWq8stdrb8iv
DOx1YeeWKM+JIWwpO0J1yMzBu9pZzQllDjlEWIdT9UdYaOjWtp0zBHn2RT5Dv8aC
FG6q7M50tC9MdSEHrdS6oAELMqjSL8fjPUaYZ3rfv+FT7Tzj5F3mkLcG3SipJ3YW
2/J39WKMLF7MqXIviDARXjXiLYoHI4rF4acZh7m8IbUiDONOomAAtH6vNZLVnlTh
qT2amiZp79B3OwFXm8445QTI93M3JybAaphUNGR4YQe3pIoIbEMRvu6t+UMcNW16
0cVMU6TVt4kw0Y89leedfFwtD7FhWcKoonXp8PjyJ106+MVF17Cqk0SPFVAkfmQd
AcThU3TxWCOqj5gfty51e+cHPG0alXPrZJd2S3KHNFe2DR5fgU51OWwx9HKxRt//
B5FrmdezLLYLjhwqoHrGByZ9M3fEOLFYVqp+6EXcB2OQvKCdo3LKGl9pCnrULbQS
EEgy5xGWZ9cuVLAFjbk/kUirP6i3nGAZGZ6RV3yAWXoYrKoB/v5LzeZ1wwmjPA9N
tFBrJ+Uvi17SURtzIZ1Gnbylp7Jn0+29/nGn0p3X+yzHOZ4P9tVgXnAHnuAFEJLM
3tKH6mXlxdS08Vc/d2ef4G6KKHN7qtTasY6rISI05k/8Uty0xm13cUE3aupCbJ5K
PqkdY28Af6JytfI+wtfxHmDvsT+3lSMSY8ZSyFziFe7ZN0w1b9VVXNEfZf9MFg9t
ynLYRPFM4ZweHYEnxYbonHTFS59FhjHxzRlKumv0UhbiBQOQJgCDTEA0zxGP9WO6
6HgBHFbpGKn1zlb0JC5/CAdKZV4TXgCxAccZBSKP6Vp2EE6AKSFJBUn2IfS96b7r
rY1tq8wosx4n2o9oC+4IxLbVF1jpUF1Zw/4GUwuEZloPNNDOQwSlpp8DCl985He3
RHo9641YZDAv9XkU/T2iwSgdi1dZ1RqGMisJltka9OCauv5+GJy4hDw8tWsAgs6Z
ZYnWeA0jynkLkE5tQPWamNbHorfV0B2K0RppZRtB64OJMR7jxm6fY2bEs4FQRjhU
JihvGylvycVYNCjcZpcck9JKEMWTGv4aF3tScED+pTI1Vs7V3eUVOJPEbkTM6ALY
9wa95wrfpZO5r9FF0lWlJG3cCS6nTFAdzIWXfIYhuADQT9kFXCJuIrWQrkaCJhKy
/7po7ns+6v7ufCI8N5ATH6TVwg3kCSQSx75ROrsKzSCdiePAlDuEcqUvWEXNvBPG
fPA5WTaIB0oRWVm6xbsw6bsClDkKUWBh77goIZvXSqLTbEv9/uHRpMv87PogXDwY
IjgFUBebVkQWnO7hBPbWi7PzdQl0was4lWJQofbtgYaZSZyzM3bOtUTXHH7JUCsG
pgTOusPnAklgb6RecUuWiArRa5iWdeLM4fI2UQFOw3ZxDfcTE6qZJr16FrtfAe0w
rpJMsVuw+Q9Bvymo3AxfzLYmMjbGeVPslmUbAY/4jUoxYE2+dsjLShHHDPszY+5q
2oWhkeWWMbOzebZafH0RtouA+gp2k3+p18Pa/DIDjvaOqWp+rvdapIWaPAlzFuRT
4vfcLihBFQKOD6/HTYRWphfzeJAMACj/5PVyGbf+6k1ewNa1O7Hsh8vhJH3qKCcZ
KADdvC35MN/UBg9/o/OjSRakL3cMx1A4SGDXennTwzgxH/gGC/juKGrR0Y3MV37d
vtdHo0YQaXqpn2HoSI+DhnqFevBoUi+Z8o9K8tbnmwsK+p3d4eBysilGmYBKdLDf
2xxgxH3/P8GS9V8qnysd01o7J1jhXNZfqay3JMBpNQYbs+wPsNT7fwFeG3Ue0kOx
37GEgzxVy6JcbaTzmrhzLJxOienc7FdMyrgbO56OnPDFoQsTSn4coTnvlbchF62s
BFXp3X2cXhxoBWWMhztzy4yH6nF/eZO4QtFONsBRMjpdWLZhPdKPrWZIb+4iUaYP
BfDNZHfEotNQGQMhLuSRHJhFvZf6QRvjYmMT84XhqgtEB/BDXMwesyjYD+Ss2I+7
eII844KiMGJ7/mj3bawyKGkNVp2aR5y/1wrj6hOiJeGoPHzlqoninr8+h9nrzsRo
T4Z4JcUYHtAwcwFE5VOYrH/PcRWdPdN92SRBqnJ3v6jt3uWX+NgZU0m4qNCVARPx
mMqqVBfn84QLTHBbKPVf6l9g0o6f6uGKzyVj0KUjZWSVLgCIB7NCmSIgnXMoDdHV
EB/BsQcSCEYcHA/NypMusfql/qM6s4Wxn0+g0CsL7Y2y+27ewWf3bBvni1H0f009
VE0m+DE5bKdTz+RHMqkghihgOybmeF1tdJi10Kzu0F24Rdg3UkCtRTa+tBYE9QJ5
fUPRse1jwnlmFNJrWPkrp/h1gHAis9mElj5XbqzrW/FgKN3Yz95siyAale0HP0qZ
9BezuVxgV09LT6r67xwVzX6CvuCwRXG0eLoN1jKOUgLQu0ki9y2/ehbcEskqOwc0
EnwhZms1NnPCsH/6j3KeyRcddv9MjukNgFfPKFxZue6/rnSbOw/b4OJq5ndlyrad
WvxL/80GYyzwcTAGicyU+o3ViUHhxHysZ8DXAndWa/l6CdiHClkQCvHuJ6TOMZXF
bdhQrrV8J8RoIlf3R2hpaRsDlnnD5zh4GPl2t+ux5wasb8l92TBVluF56AP3rW7J
1O5hOI2oGngzR5bCIOBwOJ6R0xeZ57CHP08MOxz22kYQ9UYwn5k32mRMkSb3W3Wh
PLKNpjm4Qx/uo7OYDebpYgsy2snblwv1iik4WWtIRNaBVrXjTHN7YRuGCtMQvXMn
RMO2ETnsXQL5WEhf0ZF/wkuHXpUQULk89IOdR/wHR5btK1plwAbdooP547fjIHOR
MQqr+HLNkwcr19pXHLSY9sTXsW+xOpD4QBF+ciGX7LBPeOANzUOJCrAxO4KIMMcd
ReTPpqx7TePdkry9GRsXIxnsY9K1dGwapj1OJXHW4P2n+FIPCIpV5Ph2LgUczuN4
I6J+prXKaEJd6fszeNSnwEXWLyWNiYbsxKsZt/7sJcGVPRy0FDroj+EXyu74L3ld
OjelcXrWY5R1E1TDRnKWiE0HmFYd1bmC8abNEBtfUsxNa+sWaeHzsLbVSSsoxxDW
cxDNmNU3n6AcFJXlQr79o8cD18j/1COaUIWWQx45bQR3OJVLnd0oQGi0z3dBin2x
KGxkff7n9FaqfMe9wYvygkJYyz6+Dwr64+vdMFwf1CMgEJxtmLMuzFVc5ToK2k6O
UPviZXc1S0gpcmfgoGoq8saSQ/EZE6FQtptrlEPt67iltwLHx0GhyWewzxHjVYfm
2s32FjNgQFpIMx9wf5amyUI25KrgtYupBJTXLM/NCREui/K/JGa4kmf3WOP1njPt
hYVP8yON/5XhBQiSGCCEUNO09tz/lPt9CyImjIrEDdjSq/f23Sox9Dz8zbEsr+IU
h1Sjpl1gU2YmnU6zxurzsKtgiRhInGlosgS8w1nDSTGWmN3yJmqXYlmiM9eATPwG
greJTOw11vMQvwR5VlMF4zDqkKuyo+i6hlx+qIrPZAZ4t3DSgwDd3QsRt9LIzes+
GGXjQqAjZHHh3jx+DdoZrLm5vxaIIg8itg6+noEBAuIPMP7dWW7irPDrZVEN0WCe
FkX7IV3baAZqSVceg3P1y/QgizoERnNXAQynS5x6s6BM/seC2WB0qeAXOQ5av95L
5EuMwDfXk4JObYJ2jLOIe+tFof8v1a2+Rt0fBGGCZsxjNIkYSU/FJG6ZAynApSPd
U3HvZhrb0i39RNXqq6GfyY2cincaS0JmOhcMAlxIUkhfkL7heDaDSDlW2jnKuYgD
sys0vS8Q6wXk2tJjEqZKKwibVGAjJybXw8b9jT/Bp39N80beT3UtD6ebky2JIusU
fqFwclZfXvoT1en3ehohJ0z5s7rVKeXKPmi/vAfYvJF5nihiGHveH7YErTC8geVl
NxoD17oC6jUjmSWgvq+7ZKEphD4hgyzuN55bENG8QXi3ck43a6NYxKkHRUTjfRGX
E4UgVnmhetyIeikLQXsGT+P7kxVAoAtQhfbUaCJ9hY0r59qv7jCWadIzTriOSxrr
Yghmpl3TbO97/NU5QPzIoOAZbGMjkPgizdXQo3KRf5ln2720y0nS5QZLUtQ99bKP
x+WHE62G2EP20rld/WhTgxfKDYCpMXQReFNvgJQYvx7vIvdSf7IGCD3SkKnrpVxn
odknmOHRbf+s0xY/o4I4arXkAnvBiI4/TKTIHsue2/j3Fhj9WevVavdFWo0UrB4R
Os+cOWwoVPdV2JrRKqEUZGlLSefP/0AGy/AHEvjOnkWXKucdpZJVkLwf6bVI95wb
PLhRmsv9Jx0NqIgwe3DWY75CxYjtzcOYOhtZnQqofPFdajUjN+52cy+81viCfIh0
Tfpd82I6SS+UXHJnMs7XLQOwlCMR/zgh4nzlPQdNh9zYZYCSmjId8+bVVplzaBfZ
/qQ6ODeBjbXhS66MPUWHLvy53pAkvZP7mruzSC/W7+n+4DbdyxZmZBNBsQZPx7aj
0awh+xnkNWjsiZeMCfgaRobbVq4n57bkC2yvOmsJoYN+MJkP4CXNsmQesdqr2cjG
1++kfkagNveomekRpx2b+nOo9wEFICxD54CHKqyaBy6LiektB3larIk7DLrpCM5T
ijp4foZRus/1pcf5ghc0ddDEMWB5vm1R6Ty73fVNg61BxwCQ/PAjqFr6Z/sG5Zff
opxNfkx4Qt2LlYrnLnVK/a7iOW6MDbA+tD51z6ABv7bwKqc8j6ok2nfYsnXXAuWG
wGGWz6Wwmsx8OaE7IjuHwSBO+7GgTSMiH7BU2dCfgxhG0H0pcs0Uk2kHE/yVuHjt
COKh81IIL//T9CJ6s9Qv7BH7E+elWKNPLZhvvME+SJYkV4RRf/nmqZTK0o5R4ZXr
68fh3GDoU1JXAkHr7YEmfKiRQRasVgcJ6W/XbNzsoL9ki7dJau0xwFjvza06GlJv
dn3z4+fmmoOV/uM5NRYsOf0wXYcTfXNPHb+MWFU3+yGR+yyFPDBfNnWHTGHQa2eF
vY36R22dlhFtNUOpH85IiIPQ49zfPe1SQJcL1KN2h8ezLUzALAp1Ajh3yRd5zSRt
QSISUfT4MHsPnAJRKzNssCdAPWbReFHxpXv6E/bHy2YZG3JF+xHK4yF60cx5Pprt
jttcys/EZOZD2xHtlWAviIVO+mhtHEzNRUNkIOXe0orOcthg3SVisvdQT+mQ6jUN
I2emj1zR9F70sjGQcRWkVoKYE1XE/RbFntJ7yiK0jWZQOZf8UHJH0MTzhP0EZr80
RUZfycjc5Qem4MuOm4hMuNrb6IYiQA86g5ZHnyhhyO63ry+0vBXYqtnOLFoUEanZ
1oMzMVyevIJch3Bz3PLW3VvOVFBk38gr7E2tDS4Cl0b9WeZ9JDAKtvr6lIBM01N1
/BzUJdiaTdujOz8ziSfan+0r0GA0ux7wmmPx3cFWzpRIBDmpB1TwRxSmKOpJ/jEO
yu1eqUAXOXbl1R62xWyMmO53QVFNmZKGqbcP1SRYvVDtD8V2iTUSlCCExC8D5eCn
7bo5nLN5ivRWUDlRWcNaWD0mfuO/G3bbpSV0qm0rztCAdMkLnG2s07NsV89NxriP
wvOdURp+wYRvdzabYz+mFmetPhnJN7TuNbsiVce8U6kS8Ic8EpJXqRB+gk2YtbcB
1U+jOwF3esn8STHzPDvl+J+r+iDiZqCS9Jt6P/61q8Tn+bKgm3Ax6ALLPfjUu2aD
3IAe/+MBSgvfomaqpaI1CAm7arJi6ARHU71bxxL1un3bMZGbsVh5LSwn0uv7YUd6
x45DoAnWIgcdTF/tFvcUv3ZmuCEcB0RzNJnTmYN/Ug/5dXPLu2FPryV3DGjNUvTe
Vt0yJCZ2JoyyD8WJF40wRGVkbcvuyzA4iI2eKdcemKVZJ3KMlLM/6HwasCrRAtEU
CSgzBrWgG7skdsGCFjSIxGcrj5SVLGnmXkxOpjDRsb8eT6pxJNjgg6xne8P8EL7+
evyTNJY2bLvEWj7ogKTY9LoAKciq80NyXJs2nmFinGCePCPArZlVyY7znHo9GL8h
3eGpigVhyZRp+jSPv8aDY/LwBnbizTbNoN6sE6Fp3IzEBEPqCo+wFoPB1ol8Eny7
X7fSVEE/Zn/Y5icd1Iz6SPxuvIn6b0SEk97peQxX1RLW8/0y8FMC5T+CY7jlP5qO
ErS6fisx8ei78e3HgEtBN0murPn/W9PkXhQ2PLkELsghHE1H4cJ0KyJg0jDXyl82
gxS9LEW4qageqNKRH9YzQFNUbViTpw7jBn65HGWxu7S0ykC6Hsa4xZEFn0XjdV/2
S7jdlMKuZOeJCnJK6m2BD6mbAj5CkgO3uY6sewPHUmnp1gr2n3M91EhIocv10eaJ
O0+jcrt0o5EQjitlK3VSP0Sn8KFCjVLwdGjDGnErkf8LQYtjH/Wc5FGde1/56ZUA
hvbsj1KId+HWtbQE6JsuV6wpHNuGtdLNaIqi3ogmSgTrPVkwy/4x8NP3m5KHGBxR
CGrqY8o6RTgt6v0ok2ot5VtxcZsrkrcKeir5gnkTHRopAOWnVJq9l/AZibMrvjn0
czL9SUULiE7durZfLyYbIXfg7VSSNid7B2m1ngSwdsXsgwcpYPHkz05SQbOm4LKu
WJD3BwJd8dW51CC5svl9YKoDhBV/D1TW7iOUshfhrMrgzq/d5jQbtq20ANCy+v1i
0FjJp9mvOFJldRRh01ggE0pf2+bAJaqeD90H0K7s30MXHmIMuM5NhuxqHPXcSxXa
Il0T/+mIVglX/4hdNWdbDHyIy3duFQRguR32g/D27cXMhb9RStl9+lDZp18PGP5o
7fEwlhQZe6Inw2HgaFfV8XlPD4o/9+sg0Ncpi3sSey5SK104hN3RyqqzlBMGDr2/
uzLG3ZA+2k2oU/1yIeihvrLzgYQFxi2q9K6NNQN+0WfCvQ7YPh0ZSVv74MGLwNHJ
2ImPytIMlTUt/E+QmwDdVVRkWt0FxNbVAA11tXMT64GFnZAsHeDCS51vU0QwjxOy
KNWrS+5z2uDOep+S0xt8AZ6Nl0kfQhXTTKwJZpkXlpvmeBi0VO6bNclr92mt+bZQ
zBeVu9ppYWGQcpk8uAmUi9/CNQoVLivoqVyZ1Y4ECcsoxq0LCFiw23xn5ZQjLsfb
T/Hk6rJ+r5mfUp4/rYXw2lfzXNSTe8CHgiHZ6eVreLC7OuT5DFnIC7wvTCljOL7K
FPRkZjt9qdy9qsajKk/kDn/H8HU9m8dgyni+lJ0r/FWCw1tPRxsZbwqrVEDcYHuH
9vj2kLTvLC20fxkVCTTblblcxzjK4/2i2IKuDel3jYBvor82/dRaCySamaVK5ofZ
zudDfFWtvPsOBkL4OfIE1tedeYBBnQUSwb/eKZWxs3h88GSJWl74Ea5JVj52Xrn/
6K0fakxX2A0iL8BYJGmeP10GAQHZynf6I9vG3QopB9wx2jAXsOcy1TY81KmBcmlc
/ygUm0YSlM04WdmoazpZ3KZ1BVq4RvrbCum4MBunWpvle6xj49WHRuwcCRy13bDM
4A52pwcSUskqurA3Ut4EtYGkOEcfCDNDPCCpwrod+rHK9tud5JEiNB0yBEqklFG5
cQqGAr+bF4NdeX+0GCk8SP4ef3I/xYKrlaxlUwATmh434GoUvwWH9MEI11n35neC
5DxpRc23r4ShusEHQJ3VkU3eS6Z7m0HWfDqhQ6oixC4j5Fa98BoCTIGIvCWAcc3g
PvQxRMkZAJnxzpGu54qF29ZcFLVJF89TKZWWrb79lw7WznCw+xca9YQsZI+o6GLb
6rd3JUBN7QACNPoV2Jpay9qC323fJxEuGMdjzdwco4V4B0iwijoNqxQ7+ZnffY0Q
GIIU5c5xJ+0LUORMe1Dhs7U33YcZzG1wUozdABwZEimaxTMSqjI4oRSna5mPj0cR
pYRwL/IXVQ6upqrRvvoMAHPbUysIoX5MxLRpg4j1WChbM1Tra9wl8EByUscC1v1k
6vMUknhj7T380ihWu5NlvNRzpWot3Q/t/ggA5UGgT9+fqRnqmqiBBFR7knEr5sM6
gQRIxbIvkLJYs85v24XPPE03+HK2yqMGVg4NiMqF0c5mBq8CnyihjUVqQY0BcWCt
RQYhDCDxzrCevYWI2qhYPoXEGDbXV3C8sHqgqDO9syEDUVzzYhjp7FntoNF9PN33
12yGbJMrCfNqnItXLKlridgru5zTOpUhvYGmv1htrBy1Ydvlk2Rk38VNcUEujAai
lrbwbwZZHPnYV+dv2LSVDCJhKxheHfqlg6k4FNQUJuP0KJVeo3rBEh7CEHcC0+ZS
QWwodBtYal3A3NH15b6iPmX0qA5EUMFTGJA46Wccwfgn4W+3EuY9lUfNBTu90iZe
DUlVKz2JMaAPWOJi5O+1y93BeReRaoVepRn/rv3p7JDh6V4i72ppR3a6+RAs86Ih
Nna5IUfSUj95JeoUDQk1I4ohQukvYOXFgezIAroW9tRy1aQzQrn3TtTsYhEb1h0h
HLoANmGPldHhxiZvHA+uH1kdK60lwHn65MoCAiRIsBRIAtkyoD2h1I3ixzarQ2Pv
GDr21/teH+DEqJ9IJB3QbbL1NsdWTKLZ8gzcc3cowdG88yKE+kIzATeRzJxq12J8
4rXiJc82hzMO/lnPtW8dWcIlvGPfJtEeCbz8Yc7guny4dqL6kWlY00pAjmKvjhN/
eqHlsfpxtA4+hpSqX8FkI7vporq2zbzeoZ/x7hhMvaeZG62nh9YcgczJ9fwJD2D2
ojx+l9jhTq8ZVImfG5WGbqkhzgovQeA4zRJ4W0T+FJNSz2QNyv429AsTjXHqICig
C3+W6056C3q9dGpHK0dMD2CscMwC55EnSZrA0NLYBsnlYGciHbRvWe45OREGSAHN
C6brt7GY0ukBUt3OhI1rZGG2bR16W/rqpiND316wtiHfD5+5+/DuaA0HOFJ0QlJs
n/R934f0aCrMbbvgmH1v67jJkggPnb4BNrQ4QD3/i9INtrexmeH4rmxA/jb5Lg4F
cx46TsT17/+osRu901vc9sU8hbT7rW8BREJnPCBvCqzjnjnQ7Sn98TgX5Y6o1cEB
GA/lx7DDwSHkBfuLfUKOxCZH5DOGH1Ftz0pAe52kIlHcyld1C6/Ots0BBNCqDFkc
b0l9xP6svffWKFQRaptz2a56hYLLoCIMfehXV756y5fh8sB4wTnE5ECXZFExKJpL
RivcD7o/GzELtdOcR2L0/mWmAKK91Xwb96i95Uzn4QgUocqiGhoXJxa5BnMD+5S1
Idsd2q9hJzmcXLw0DP8xtb7aF8DFfx78NcwJ8olmcSeJb9F0mbhbFRb89Rcq1QeL
UMOYJ2qrOlQGuYPJkZ+k8DOQTa+C1pSklo7qXULJTJGujwpVXj88wiswLE4IhGwu
pJoDZAaCb5vRs3/9Y4u1LSuKgoEXJ2wMl5187535IuE8MLLrkS2h+2YbcWjRrxcL
jvCvCilZ8YiT+jLOSAihKKLy+MkHtbCTEYR3SMhyNNUftPcY3KRMUQN2ipDwVfKs
Q3xXAxPSn0455LjStd/4FrjG7DqOw6UDP+oJ5PvludJ1512gcB5cf6kVsuAD2enx
EMvKpoJQ/lxj9fLgkQf86iJfj0t27nWgzcsTcdHTQ6cMNAhzb8gc5ArPTtTIzZs7
ogik8pjD1rP4ug4pcCs8Eih8LjrHxIT4URfujlsxDVrgQ52LAR/uQbVWvQu7tRuP
m1cd5A/nMX47hux5GuzbOhL1SjPCg1wb0kiuTU04ZAV0momNoqricP772+OWdrhF
diBGti5712gJPKKVpLbq7JQbMmyFXPnUNt8nMBM4O1VUOZbo1NcFZk6x2Xv7r3bE
Z9bNR7qlwUdeC4/Spvl1IBq8HgwTzKyVXXZPU0gzyc35d4oGdtIa2omtNmkGlwZy
xO0RuaZVfhrryMAUqN6efuABYpmQSgBo1PiSs9x/nIKbV30CIrJiCAu76XlMDoTA
1HGW1/4VbTXlyU+oc+6RNWY1WZ8DFB0sIb7UsB6RB8tJ7d106IkgP9pcxEx1WElv
L9z7uo5OnoQCA/N7Wkmu/RsLxmwnemqKeACYNVluW/AaJTBGS+PleBp81dUAELZA
YAruL6hXHQ+E2XWcv8CXqzmjkbX5YZ5bwn/hevup+Uc0SjetlYa62tMzbN4GTH1H
/mzkZyOWPld2LNdPxCfIIRczxh/VdjrZsSx3JS1oAdYpOWgkWdounWmLLOdC66Nq
IA3blHQ1LbzByUu+XO3ryssGHTuvsi6z+sFXxcv8memhzjHVX3QEXkKmVa0DcIYY
Y6cmwxByW3AvNv9rlSDRA/Fz0wigrGpfaUYhCrIKXeAviplzYbMk3bWmIdqHkqJu
WFtNAsw70zlI0z+OOZ4NOlpFUCULpaRkWWKW0JUda0IRXmKPIo/9iNGtLrQwmT32
VgFviGjlRYNRtYdOTfz8aJaHWqw/sqVvt+/bGQlOfjY308e9u7XwIksPRrB2Psv+
AmHXx0l6eDIcWYuAYvw8Ex0ovRFe06yGz2Mc7hB6ZpN8RrynA6a1UHP92a7hHLQL
d6Qhe8OT/tTu9buCZJBif3UYksPcxw5/VkkLTkEBUQ89oGBeW+CRG0GOhJm426VE
8m7WLHplsUnwCIZjlMDofF/1HhhHnCW6F6H/TT8T4PybN8pd8tG1kJVxUNyzi3TM
F13aZTFSK29ZuYKQu5NdGzSGyctXnSDM09dS7bYraCD1U7YaqkYKJtq9DG3PkMc6
WzLZnBEGQNAG/K6oTe4eatSe1IlG7waI1SqcsP5IHHT2eCP9ET9foNDwrcyQjek+
etW96SCzQTevchzJuwYnLw40QzoznozTT/NIfI5wOdXceNaWb4colFiIOYPO5Epr
sPOkaeDhlkZU0iWTw9eIAaHs9khxHgmBfdTqo3lWypxEoBFcMKzGkYNqSTkKnR9R
QeY2MPnUQ4K301qKaLaT2Lkg79U+5NWMW/CmdQSWnwnVHdGh7joLPsuSQq5+/Kln
8tOd915nAlLDWMeram4zTGl2ZfrxOcFDHENfSSmTo20bJ8+OLzx99zoiwGO0mAoL
MLFmeW5Wcxw770ASwQfo2s2j3/dg/ZKxlHqSstWnRwm6cI/5gk2aq591xPrqdP5z
8nVD3+QkY8jNZDRk2kkKEXuSAsAPT1crMy0IxRJU9yyooB6eBAx5Ggu0mezLAJBa
N/L/QsqG9gRSIXrbVvloey+wctn7AGVoW0TAKszwYu9JCtPAFkty0cLAaD71wdbv
xKXV8DLbwTaEShl3TV/wgrW0nqOmcI2Ih3E4uS6+PHuQ2tKyAQdrc7IOjTzM9Qga
iQjIacV5Vj0djYyJ7k67MLHyLMPzy8+kxHKada0En6TGqa1NIY363rqnJZ7/bXGE
Ud2YoDz+B4V3uM3swIpG1UhWCQDBS1TKI8Zi9GfynG6KLqtS3rY4N+I3M63YlFtI
rUvuOPirAPs4WwrVm8beNXN84yah+sDkhWRwvJKJZADYZr2FsSWMAyZQUTRyCx9f
2kefv47WlMu2TSSMzfW7Q7BQ670NFbbguc02KOBDtqC1ROVvK8YampUR6RBrfqb9
Y3+9XYYLQM6nvSv3bONS/HHTNpFngg8Joful/sb9NXp9iBjbiyaV6xKe+ZSXfR+A
AR0+ZElRHUglhaDYzl+JmALj9hw8gKb/lI1zRPgW/hsDwWI/CnPkAjS/SX1PgpL0
JGiNhFUIzfaiIhcRJLdxrjinDFqm0SC5K7+No2IgI+jLHqg69vOMF6AjRFaAh/QE
wv2PRQ24L9z1T3AwWdGakesRfeESObqbLH04rCq74Gj8831erl6XQzcnrkE1Icgz
RutIAe/yNgSpsmBoXoAmjUbImNdc9se5VukR8L2GKvWfr2288Y7YFAdnOs8ACltQ
rOx/kDNYG8RXc/WQuBZ8FHWrq3OQ2iAT70iOkjN/9tt+ciOTy+iFsF+w9ZDojHL3
aR46k/gRuPNWhLXnhG58x/db3Bd+JpuPDs4F24/rgNJbI+L+Dr4nUHoYhIySuMcn
/oqmGN5QyVmzQ4bHlWsFkg5lYBrXqjI+fgkb10CidaZMIjXpG1ANQ4h1aFB3yTHt
ZEA3PdbO5zfslRNfihFzKmKGSXDRwDd6OJcIoM/FOOJ26N7PbkYeIKao4wFYVsPQ
sDaA5Z6elC4oPgd3s0sG9qQhwP3j78C23NHm5UxiJOK8jWiqUwnIkqnHxFk2w9ao
`pragma protect end_protected
