// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.0std
// ALTERA_TIMESTAMP:Wed Apr 26 13:36:51 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
MZX6t7TyJEF0MiIC9rNsbOgsgJqlDE2AFaBgWVAsDe2JwmI2VV6yqY6877/L0bUb
DHyG3jI0M998vINLjFJVXlIbbcFV7hO+fa+oWIqGHy1LO/Q3IuH7bbqK4vUU4vGv
fevwMtPnv/Mq+nbSzKnyjgsAu5F8AJ2/A9Rr+T8m/nw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 49328)
AickYvD/aRUQl2Pp0gqGZhxEdjLlY6kLeXr37eg8mRCxunuVk1NHoPwj42DQugfK
Ab9YiT30xr6Azw5aFWbWr4rp3oUBYuMp1o8PEkOpvK1jvr8IOI/NUu93K6rbbeCn
hQqrT81Q3c1FcFCU3U+J+VX2HLSLvJVKqc3tu29FOcnapejli8xLeKbya5Sr0fMY
iPmrRcu24c45s36IHViNYBoVRyCoKUdyI8Hs9y8S6HVFwdQgGLcldYJdJ1Lc+loD
WQJL8yofcnQKcRX/U5GE2XOejGdOjIgZC+UJnd57H3RUJXt+7quSglYD3BybeFWU
JCBUTRXL5NIW4JspxuEXTWTwTld3PI+wWVK9p9vU+6NbvOXHeNfVeYNl786WW+9p
gxm1eIqkgrCt8sHDtVP8eX+HZl8kD5etzRoBe0xqzckBgY9wIIYLsVLJrEwf+/g1
k+IPBB+masJ004Y+yXeFkeLA3pvWuzsfgqeThmy47794iJY7B8WXe1VM1oIjICMO
47O68ya66+kCkdrdvnuag5+w1VvMlen9N7nu/XPGksdsQtwcGSOgj8lPGwBbxrNz
cFdmqiV49i6IwL9gJ5QP4ZrLrAU9kER+EkSKQTJgLXBdrAMvHVFL8vtkKAlElC8L
iVlPrfBGVd/ZVH8v/yxhgN0e6b4aiZfAedjGTvibrKsNbunzdGWwRztpISdI8TA1
3R8ZqzA/GXdytCV/BYL8QeBPHswHHJcgCY7y+iM85Qycg9roet7uoG5SMZwhnTZ4
QduLL76m0ZdxVbn4eDzTKfdEMFDLBoa760r0BgN8h1jqafVYB6P18eXUT5yR8Ls5
UYiC+iQr2wQFmSB4RRIp26hXIKAKV23+TMuMXWk20rBLVeDYX6zxoM6P/w2NqfkI
1I5Jt2PgxFR1wLwX+B5Bx3JAX0FU9auWsTcFBpBnp4TBamcCwpIxynkciThNFkyn
8OvmrRhgaSdXgrP2TjPmE/SNxJ+dynhQ7n5olNfgX4J6MDpuRM/lJ7c7omJ7HX0v
CSWKWpJ+6aVrUY2N7rRpGg8R00p9UsqKMhfbbef/26ghFbCadkBDRbXArAqIvJAM
9ekALmBUEg2+cliHX3d70m23PDOVXvkLX/mCX97oDwXrecNbOtebxW+NSWduau3T
dSkdfaFrnojB980IHWQu6kRABahU26hAnhd3R6pB2cZTHdcNbnJiAdj0khi34v3R
lnSwQ9dnbN/GSBzpj7Kij00xKlf5dKNOSdJM9qruF20G1R3YjGyWg+TMtTK/1g94
oAh04r7FT2+mcCdPu3OtDLsan2HPKGGVlljz7iiCdfwnIQDihIvITFHv0JZPcjic
NXcu+gkOgKGf75rn5nt34km5i6LBIuGzWCB3BYZ+ddvvZGMJNve3F4EzQUGV5UeF
8CbAyaYgyCn+FO/ISSH37L0KzrHXLz9XdfaRMCGO8o6iI4cday8VeEPfs/XvPwJJ
vRjMLJ2urW6dJ0WuELqOQnViOvY+QWDn64XpU2+YT/dTgtDX8RmMrsaJ4beGXUH+
6dQarfE39Idz6UnOpwU/6JIOrcDh1FonahMw38ltTlG+ynZXy20PdLENjIt0ADCw
IpZ+q+LzoXlEDkLJedDHXSdY5+ncRdy9HftpDjAPHak3xVr59hMx5mnUTNI4ibJ1
YfssZd00/0Lq+NG1w8dh3QP3XR3ib3F4LHNW5vy0Yt9pLnbd9+461UFJsIj8BN5F
caFP4P9wyzcqw1HupYhk07EfI0BQRzUhb9xEwpW/+S5LP91rqebJV5WfRHBtuK5v
7Ooe9ghLlsG6iYIGyERhO5iBJ+klvdmXqH5oSYEXu7UKbuzeiDGxTGKkN1yQ2Mef
YbTB7vugZDZK2VknqERRR6JUF6+ucfmUL0+gJPRAb6d+zvXomC90SxpOZAiEArFD
EEJ6O9vl2CfVIPQfsJvNBG6QxSIiGrlkx/b7UfbVoElJ5wBVrpaqfckcE3pwf+Ip
ok0Tj51+zud1yJ9T1JFKczp932oDv8EUvoype8Nlx2HF+meKxkEIbTpAxIWPm/hO
hL32jugGkYSoWFH3GhcnspsEiwxlU59mYDWi9wde0BtDvGmyv6in+7piXuRMzqDx
Tbg0dx8KikHW7Un8kw+AE8ahYm/bfdX9bmEm6zjUMbswfSxRlLAs0EAyI2Yl23Bn
XEsMLEqXOiyX23Q1XUJHl8haIGkhmbGkpA6zRf10k/UrY42ry8W2eNHBtq73dIBh
/3A48ZcNzB8AHgJ2aKP6xvy698aVaf3JmTd3Jlvb2nnCQOr96IjJ/d1bNAkX6nzi
8Ru+Yjo67df24f2Bm9F8//85C7tV/oqRKsu4L+XU+TMQ8nLtpQdgCPixHxJE1sf6
9U8hEspGc17iuIx5nxi6u4FOn1e5wMfDt+FI8sRRA8SXI+dXKmP/fWZf/SZwwPj4
HwOAk++59GkRFyNoqKNZAoyqUlt2XmMi8jwyuZZ+zTy2dQelFr7vehvk/AgmNnoq
h0X7/l7ke2u8bUO0AAY99ATf34cLrlpTtx09UYaiZz7VSqUmMBDKa8gvCfwPnHE7
wP3qLCY9wSxAnDiw+0IKkxYH9CV0YUFiNXdCqZFUf1rImCcOBTI3EVyFMeEXSPv4
rWPYnkeJLQqTxKO3R4IR07NQdClnGsBipGmiLjvszIdTLg5Y/JL3up9t/KNDvpYd
Jq7yHN8cVVEpA/S4tnKRiM5z9Ra6kRw5ZxHHSnCfxkrEIsqIgGRLW5Z7G/B3Ppqe
FnBlxNRYAIoq+Aa15IqaJ+88abzj9YvSln4Xpa1Fc6ibPjvN2FpvxuinfIdTNUVn
f6OadqFxxRuboziMvAM4jTYawxb8j0b2XgyBDN+SeC2AzCTwihtPVpJ8AnqfqrjV
v2mB2N1dDhbJinSH0AXOxXZr1FVKDHvvUNkG+stPIAfCNL8pR7iFIS6GGsOH49WV
E/a/aqZ74rkzZkIK+ezPkQ/38QRh9aVIuWzWjcfmZCG4FwWyH1EiOumKu/iw8SbF
TktVdkbKWp5BV9Adb689UiXAgeAKe3H8DI+CYnaBfC4Qq997tQX41aXLr3X1VgWE
k6V2MBT+pEOjPlFsT1bmxE6SO/8NiEMzWS4Pc1Z/tqj0eHgrO5Gj/KGly7RjCj5W
QkotdjlfcqJh+kZCsYS4XFdHTPmyI20EUnyBGEkf4yRn/vTrpm/7bhplLnNd1+8r
qu6HW/LzDsFaVnby1JAsH1x3i3zYIKKrDVdwtCW053TgEd1WnvKoxQnATH9cRUA+
D+20l/z77ii4Zzg44icpUrpudFq85n4ykRSabw6kNeWOM70eE91bV+QgmoWBzcj5
VssSZ0Cl0fpExIcmAQ2LX+rbAajGprhqMfBO7xn+3ox2RW43XRvEJFU4nmr4mjKF
W1F92um8y4KTISJ8auj9xjd3HOgP8UBGJId1Y9SGQN+SJEITyxNJHTAXP/BEVM3Y
LtY6OpxDU10CxP7NFwIpPW+VX8i3UENOyfqEVqGlToqZ8iSDy8pAWVk2G/GJaXOm
knsHBtNcwA8IX9zXgY3nxdOGFjiLMmuBXXf+5aVe3q62gyZ9thEhAd9oo4ODrMaO
6EbqBjZORI5baLM7vZNyPh0yxXgoQKf3Z83pxefCon/Ra1dzJV8eEbLeTQPETpqQ
/rsVlisGbqFm0/LlZZjCGA73MYn6/nUoXiKKuqu/7UgfoQgrRwdcyCIcbIc7gBOA
n7I7M9VkTdK9pyLcIwcH3jLK9yVJuO2dZ01HnE87eQc5syob19EMPRhkBW2StHIN
4i7QlBV+G2rIegyfaeA49FptuFW2mTjzZ/PdgJt/v49I3FPHZoYnQpjy9cLSsKl5
pnlME+sgqVDNrVuxGfAIdJka6vmt7JPl/WrK/oj1nFmFl1Hyxt42iL7uc4woBJBD
UsapqjebD+cZDaABUuVBnGGGkpZ8OGmfF1j28ai70fYbaiEEF3tw6L/iO2hQASA2
nutbAR145+zTo2S2gqz3n328AYg9rJv6YlEgJj8pJe/ZhopD0PlSNx/10UASVV3V
FVi/EsUzOmMA+VufiA+LPJLsvn7sOh7P9skja48AIqDumCVURYSHcbH00+NCpain
mDqMnWPKD54Z1d1l6ZiSczT+c6fpdhSH4aaC9wumJrTtabp/th7A4cpjzNPi60wL
KefgaIvyEewLfJ9n/1U6qzIrV1eEzrHE86pDoHyrJpNkwnyOy+RHiBfViKss85m5
2agT3vzn8jGnxVPWx8kjfLDjQvRV6lH2an2ES8vqHc89WkAafAnGAT/FYHPymqqe
ubdd+h4Qd3LueSXfSShFXRASjoqWCyGqLUQPc1wRDoSMaliEsxRaOSTb5VubE+k9
yFDaUWZT1GjJ2E1t44tXVHFUQQrXs3Lrz5mtFwQViGWfkpp8RfYF/w/AIvN8eVUj
dmEagDwtYgLAQts3yIvvRoNJxOW+bewdTk9ImK69mIMkWu406FiO8n3YT13tsZRW
+fJ7ixsvXVrv2yMafsoC76G0VHkjWD81ITA3LdEzsQZdmx6ntXqb/74+LMRCJky2
g5Nk8Vpi8Es7CXYZ76D3jY4THLUSyHerqCyvQ3n1Yo5DdhdIrJaZbxPISap7iUbP
LqBxKMEW6eAvXy1wZVMm8jpkay+Qqn2iW3GypcPepPeCUxYKDpP7v0Fp6ozeQ8uS
ejHW8RkqigDs/OHn6vWiDHl6qaPy8filWeML+r8O2yHtxyFooXS4b9LXkYPJUDWs
eevntT0SYcQ4Mg052D7lkxXT69RjFvv9XUnsfF0Jt1DFk96/mUR0i97C5HTmXB60
rOAUBV7wR8F2W45rfk0rHs57WDIDO2N97SNDmsuPp44EDsnXlOD+gEDpXW7hoBbt
jspXc1j8PkoW5tdLm8HRXIv8OieafZQPDj7jk2N53nDzoIp0fIHcSaYUjr/y2L2L
ap2B5oP4VTX3nj6XPfsTbGMXsXchacrEWv6RBz3eReGmTkB+nQzPjLkuElFu3eTf
Jtma9OFoTuM88tNfH+xSOoClgIpUwYe0v/HIk+M8CX1QmJwKydVwoIUktbHfOGiK
mDXGQWcQ9S8YhRiCHxcXdxcc6Qskvj5pgH7/bMMagaiu28E0FL9i7nxHRNn+Pzit
b+sF4MK45Kpw+uK3/KkTSCPSkW7JZjMhYeHxt67wYORACP9xovutn99zsizQrBkW
P9gP8RJzgVySB5E9/yS0+4QxGBa2cicW4boSAFUvjGd1U7GT53uUCcG8UMpva1/M
LVpglG+Fe5iZi1WHgv5O/y2Dq84EIUnlWdzCzjGIHxlCRAzZiO1QQ6/AtISBluP6
qZsm+pQ+sH58/8nO4LGYXfNJqEpnYN57/LCMQC0GLNJM9ncFwzSoA5449cHKW1Ob
neQT1k0ocJd7QZCETmN0OMHBTJ01Ql0PgktbdaH5ZEtyqP+0QRxXpNsPhiiOAVhL
E78rciYWF6zTF/EukEBXsU5EYdAso3WOxIWU6MFoLChc2n5fvRdXxffpLPF0uuxo
oTkGpB1dXRMFFOdCNMx4h+Vdv1Il8rup3Lu9MPAmGewIoL1EnS+A8XFHD5F6ragW
M4ftrrlqSDkpvFrtkUxySqdWJVKeQlqzRa7Bg2nhJ1uBpYqTfMGlmwziSgS/zlff
tbDZVUI/Nx3THtmuU7F5b6UYblglkA1R7qh4Z/DoFfHz6hn26mJZictGXTBOK9As
tZcjEqgsin16ya8yQuqDi7m3Uy+59gCuvgWu3kC1ziD0rX8nicd3+l+6a4fVr+7I
/e/nNDD3ouH5n26FOsi8fToRH0Q9CbaNNbh8TApfpFUgtJXXERtyuy9N5Tzib2Qj
HArPY7QnnC9z1wteLuYS58ZvAabeDgdaz1EjYT9KxC3vEi+gmIUw568nSjVeVjS/
OQbXP94ezP9Zyut6onZ685WM/YyROkzHzO3jdVXqWY7nv1lrG1WsiZQMnrhq0s9+
KpY7O4f7YAcLH/pxw1LAzyEXVeyhHpJgH7eUiSFcCizW7epo8WrTbCQSD7N4UPQz
6DwcwhwddEsojfiIx3MjCEUWYm6Tml1TQWVFIiHeIgrh5BmukwLwmkEt3JESRrUD
Oq3nxPjpLCOc6hS3oNSAO8HZtVmgtQBBvYkEM/YK6XvV2cW8CiDQdHYSuEZIdEmq
u89KyKAk2ByXzgpEmt454iQJcdOr9EzQz/al2DJ1xcdiXwE9EWuv8nP4p4UZFt4b
4cPLc4LX2LIKkBzQHSKO7idQr9MFEa15jhabkqwEUInwan9aFS/u3ZZUkW1rimMx
uXSQULFJ9VB3u1ciP5XJj2d7RNP56+46bb0leN0rd1V2tmk+/Fl91BJsp6ddoXXd
zKNDRzrxQ62cDM8y32Un3ETROnmXr5j7I2uvQqwDHeHwUBfLp562x7nHVcWfEcwz
z4E4Zjm+tGIjCi5K3kKMReVi+6cE4n5kqTfUje46w6ilnXqD8+2uzrtupU7nkEoY
Lu9L55hrvrNRNBcv85S5Mwu83k4StolzV+YFZALChL1cYIh1gf61CqknydBa4k2k
d5Bh/YK5Z8Qyz+ON6Tog+GxAcwyqfq2yYpF5J/jDh7QLqriAtFQ9+MYSyKOee3vL
g3Mbth5aGly1c6TgFdcJeMzvmD8Hn5eASmcluYPOnSj3X7nCvJ3T7o2nH0igzu1J
fDW1a0sRs4+eEFH1b+phc18VRuHoJWH4xhnriDKtAgPNktIK76YUvVHf8OZF5nYt
0vTvzIxw/XiYXn1YhaoWZjrfKrHZxF2v2Hx9P9Dy2GsYuzP3TN6oaCliEM7rvF3J
eS1D9Xt2wIG90/dxFPbdrRGgvM7x7+jOuvyd+Gijly5IZCZW5/VglSmqHZTTyzbH
9icrHCCM6RcTfKs9sZGz1RQGBeUMmCMJB9dMakceHcqxVxQ1nNS1PK5FDzAD2Ljb
H9RsixzDtH0NErxSY4vp+Dcwkywk0XL2/yI55UA040woaIq9iqeGwIopkC0HMzYl
YUAEKSBbWymGX3Y/zO12hAa/kwDB2XLbXNewtIm8lGjM0bVSqdoP4bwRye3X0Kyd
0H4DfFY+H5w7SqcVrD1QRGn9qgsk9G+0CGQ7e+cBKI7yKDqRHWKCYrYRHA8XkaqS
0zIntoO0FRyPk7kQDn6LW7YpSi2Uj/uKw36zSh1vwvG/bC9uUZ9OOrEdOn/5Lv98
MM/QExghPJLmlU0ZbAEv6wzFdYAq2Mtu1EEKb8fNNOGWGUS4/1YTUzHxH+iNPVGv
ZNwU8fArRWwcJ+YkqGrL6jd1A8HqwJhqHknagjT1xgQiqXYv9xWbu8T2C8aQoulf
RUaL+ezuHzc7kc/URRyz/C5wYzLrEfyAMOSc1jAxrwGQ8XE0nK0b5W+7tiUMr//H
E2hPWfIPJGjj+/XGV7CKI5lKbqq98f5FAiHGMs81JMo96iqKYTjFSWT8FX0jVyie
3dXkWA8QYnovpiqmpXwg2IY2Cs1QMK72vAmxy90R1vcNLFRJQLf+r72X2lDmnBg7
QWtwMWndIVnBBQxrvymLdyoMOrjeaVxaoiax0o9aMJrk/s1dWGtgPyRKCECRgx+x
TfKO5N9bAB5ivT2TSrP45gF2mrGdFWpfmjnWE7Ezj+w1kIWc9M8va6pZtf/c7882
2DpdJujJTOWaDUypQ/B3icJsXdi++CMPdk0c1aVlR7pvWHPxrGg85Hw9AeqYosgm
YCNifL9hPUbCbSkjYo9iGJ5TJC83zHShHbhH+a884f6/SQ0Y8iVDyjrd7v/a9B0a
O9MPoHyXzQMjyfE1CTSZrSZIflQaneQgGH1a0crtaMbhPXiLOkNLX5ohrJ9wH5Xp
yMW70AqLNlEdfNXit3hBG8AdWTfUoNCxmLUconqxtJcAzq4m8zbskOsczMrP3aCT
Qjo09EW3DoQQMyCjjzJSLYfwCabrzmyuen7yBx8uVQifmdwHBV3b70rbiQHwsbGl
7mavU+UkEt++oy09DNDHNk6x3+X7GcViJKdWxRUzXI3mr1NsOLuBXCw55ZM/3Xgy
Ffj8EIVjAQU3jCkaNiL2onk1GAyFnz7AZzWSA9+Zxald5Ua6yX+cwaTmtzsXGtaf
9tWe1R/7kj28mXb7Nq4sLRFyJq1E+r5rjgxG7CPfwZnCThMfOJWVhfSd+XRIj+Ae
gRVuWJdXggKuEowrjUxqmHTxwC/jbGKQPD7VSyacYdbdKPsD6Zqhls6ryq5yhWrA
fJImxYjDLhU5Z9N74t6Dxlst3w11+0xhkosIDhjU8QDb+wUyJqMr/808owmmqnI9
IO2xU/hFkDCtQQ+r3cuDtcq3rrEmBTTZ2jCEPaF7+qRdm+q0yAfxEdi/yl5299jP
dLs3GuaMRo/0BY0Ft3/cq1EyHedixiKXb9RbIpzlFwNpNTFEKU9WokVJAnf7SxTX
+yCcPqaZuNRB3rnifwOLTqj0gc4Vc90kkK1aF8Bb3JG7vjK68lqVT2THzWyqjE4q
+PhPBDAOS8PGeXq4HGT63jrFNeMiYRsUttNaymugHaicA+iVoRJljWvPJgJ/yjil
Yk/t4ZnDkUWquxG5n7W54R5b0FnWr22WU7aHyJc5fme1QwJLWrGFHGjW+3ClVUYM
qXecbW2sp/7dfCgjTZa7s+3fmJt7igxmh5uvJxjpwyHMNLbYSBnc3cR2zvBROx+w
4bGMgnaLgAE0KDbUO9G0mObjloVgpdRRLDtMOjTrPO+Ej0/LxibwJjtO3TqIeQS+
nppvkRnA4FelFYu/ymvdSmQHQYK0wfPI/5VFuK1ebLn4q3vGAFzSBKd3TA5r08FR
OmTxP+A8zAV8tedl2FqPg1jNdS1A/E6kfrUROqIL4XCZgAz/Zm+cO8awuCtuzEpz
sHo01xwHqxFZNc7VI5/IG5cnZR3txyI1flfxmXaVOwwKPMpJ3nTfizHEDIwEZ0Js
5vxkJNkzBbOlCmfFBHCOFqj5B6FhgTcoVwVQXl7V7140SJu5/Pt0kvoIq9PDskzP
ogC1VwwAAPYoygo/dUUWAooIv/czj64qPgHcVysZv5NJINcOk3GzbhHGJyBN+V/f
mD8TBh2zOJX3IeL2bZzxkYbNZNeg4o9GAPkgP5lGTEVYNkaNL92JaAnZTMb0mlcm
xBQKncwrJUUSDHAmSbV/QTZZMn/D9McvNBeENe/XvkudqGeKnhvpUf8avmhNrovX
a1ruM6+i2dscS8uK2AVSd0m7gX8uTprFikmlGYUp2Axmq3nzZMHXoU+qHmSCbOas
cJUWicZ2GMrD160fyo/Ei7IsczAHdaDjJgKE76mWzMGbonlatJgNCGAbZMP915eH
xiVukvee0UfJTFiTe67PTg4x02Zv1kx+Zy9N0j7XTwGAM6Stg7l/8dRF3RiplUc6
MbAECZupuvN5GQF649i23dYKNTGJoIU/qAv177+DJrssZTaMJbFGu87DMd7nptYf
6fXSg+I1r71DNZwDkT9AOoRMWRu6OeDsAl2rY477miRWGR6Masnusp0jieJXiDAb
d8bOCyvg4PPt+BXcScEZyIrZ7D1DjRI2J9U1A1/L0sKiXN6AsGAbBjPDXK+cCVKm
YFmvZZUeTUgoQm9rDZDETgoGowaJd29EIkTgv96JK1eZs3lDNBavTSi6FXV3qiM/
/ryvqqfqOyUGHithy26dAsMymm8vt7/za6HzNMequj8hBjmcT/wxikF/mpZv35qu
6UmWDhgigfW1/OlVeq6qM1+lXG79q3tKUBLQRJN2Ixuc0LdBH4t6P02+rCZyUumt
ASJ59g1OKxKLlKGJdbhf1Dx0KJM0s2VCIAsYUzTXWdj9I/eUer9PkEZIc4eZQzup
lqirWAJ70VeDAjnHimhR9uP2JPvtG6gniORJbFsgdEJJ2gBQUA+5pixzZ5aWBrnF
bdykGKFa8EwrSYq3aVbetJkoAD0YOoDQoKYbJ5QPdn2RFExjwRQm4H5T/H249jYI
U176yTQkpRrMqsrVR9HMQtAjaXPmGHw4ys/9uI4/AZUY6yxXccqqWngC6UUhw2tt
Ck6ETeKnpK2xgXdtAUUEf66acuM22vFmCJx6PJ07TKb+GLE4XAaQCRfjnYsCh9iE
47btnw5K1dwsQ+BmSEcu/MB8s1bfivzI7wnL6nay3gI/5VLvwYDUlRFgmIe5aGED
FsuiMt3Zq5B+h4GslPoFK6mWUatDOVbQVzB3G8/hvbZgdKSmhcSSibO2QsMXfcJS
QlCJQisXapAQxwaU9vlRs6ULUPIzJzApxDfXhhVlsnQ0FH64402z+tO5XHgz/6GU
nVI6l+GIPvgJdM+i+JTY1BY9ZJzyxjzZF+V+3IgVOAU3EYtOZvcp7bAikmQbAcde
YzgMk5Cylbnh7BMhekUvrmcaHj35g7Xx8Mj++dESHJbGU4QZys1c7MJ0LxXA5pi4
IIq0FD1+GOeWiX3hsUoXbXxbB2wQLvKC5UrP6o43xLPrqEE3sWI5z/Ww1u9bYP84
0DDizwNcsGR51mtMoeWHkQiS94nVGcpry0kO5jH5P3PABge63+ZrP0JpisH13SN5
POAN73s7XxbfKeLHOyUzRRJtVtI4NZsIDecjkUtc7kBTpW+EBUIClZyDtLcUs+GJ
fHnL/bxk4Twqdgt89xGR/Oec9vBz18oWLXDraxbgxk/49Di2oWcBcg3crG7Xj7xC
SXbp49nOhgc62G+UJA6FELUZjkdlZQt2ndK1C585CVQ/YI+6UgOPhnemeg6gSMeh
ENUd6QApSkS7vKL/kTEEnligzTWYTqDp+hYC/+AVRZzx4hqAiMWefs+9CbGcLNzc
mlWKuKA3dP0r8QUvRXXwqqq+Wl5/9jFhX8ljT3jmAr9pvrdfm12dj5BW6V/UCzWy
u64Fj1T9VbDT8ZhGAVONSK3VsA6RMAitFo4nlyh2/dFaYpux8VjqAERmGax7nPHU
dXtbiVZHQl+ZWvyJWJnj2pLEEi5YB1HEIcUpbjr35+vVb+0IB3tSeyB5XQ0mmpO0
izqT1uxhCELfOKoL/CM6kP5VN2aoeTBPs2lcvyBERywwLQPi1fCHnO7kywjVOM2g
IFaTdLOr+WUznEbXHrr4Gw7HJOlAymcFi4XH/qHI6cqgVj3h5qlq/ZeOeeZ3bYc/
qZ5n2i/H1OfjIqKI+EU0qajMPd/ls88RIyeKSP//hpDBizW12woBNA6gziCxQewn
nEFK2/FWLDPCr6X7ag79sdmdd10gHua+bHyH3iJNWeXR5ohxU/D+nkubWIAwY2mB
5e9p49UwDhVoHA9OunlDcj79hmxQFHiKoTWDnA8k/Nv0YXdZogXnqPw6CeN8iyKU
bszm1ZY0CVwIp44+RcxJ8Zu6WSbYsNxXTKYxLO6BreFJFGHUxf6/i3iyCFtYrfD3
zSzG6QNmYGFHj14rv6oMcwg8s8nJBeW0YCpX0JPcyptoRZib+GNdIwtKRaD9Uxxd
3Nkwo2N7lovRcVsbhut6uwrapdRp3j2dj+0Abrzt6HJ5/nkwGjO6WoQTEbhebYn5
+mMKshGr168QSccW6ZywDcSPbrJpPfCTLxVdEJtd48el7C3uomd8/VDBVRFwaCtn
eIbnrisbvAAChgj+zZVNxzQ9fh8ovFLAru+jhucskKR3wiADDs6tdflNVjnMKti3
5Tdx+eRcyax+dWxvHhSijLZal1CNRsITXB4rKqSfNTxKpeOxFrmvQFcY8QE58a9b
m9J6l5ENxNsqJL1pYFZtxiGWnS+GVUmlthKC71Vm2fV6hgq+R3FwBMBZGyGznPYv
TWeVhXDvt5BXX+gzvjw1oksfGiyGt70aBY78UpDeAWxjS425x7MPWruaMRxXnhNV
szFZNGpnUh69k09GW53W5jtzzToizUJ7dF4lAQwMpyGJWO/trLNchJer4T+wp0Mz
mx1kPk8Zy1yg0Yq+E43y/XObkgJq3IIM51t5O53kutmZn1mMP7KibanCZ9NNQKQb
RUEKDrWNLP0heJ4cY4Xb8xvn0wIue6FNrAVqlSD51tJmJZTqXv07ir4q6QLS+agS
plmU1NQSgUeJYOa1BaroH4ZatAX/5ulGFtoTqbI/New+HSNWeyI4u0afals48M3C
yiDVTgSItr0KgwxwTFX8RlmMErmcQt1zOt5tAbEhnAH+ZCggJDM2OhvZCaz6E0TG
PwQlQOYjSchIRQcedATB5SJCTmJn1B1Dhfln6YtGXE+c8Mp/zQIPlgeHYTHuR8rD
jza9C3/H5rF/Zb/8a8x+7piCzcr9CdOaelgBHGF1HhmNQNbLNM0yDTdJiLA0d9S7
XVa0pXNgKjhzT5T5+kFYMD4/02aApRx5qhb7zuxu55VjZpnSLuR9rPwHWt6qrcD5
UGhRJogTqQwpQhuDu5mdKHWJALXHB+w35Kz2D0b2lOgLSXOMR5u18TysQeVi9DaE
C6Qz1M4IJ4RRzs+DSrVzSfsbyEE3Cgri8ucFf0Lz09bLDp2MxzjiQx8sbjA4lYbq
jVAIBs4rJ0YiaQ1U4xyDkwVLrvOfpVSmig8TMS0DpJN15ZjTq8skTRQCZvbL5SAo
13APsrVqOw6o3YuY+c38jSyPTIWE979sIpm/6WuJDpb34xiQ4JIe6DkpnIuoo0dz
41xXBkVyT2Yl6Kn9MO1RAxggvMYbnhEQIN/halPd1hQB4w+T2Aji5xj+EpNU7+zQ
00s93x9aPRviAn++7CJrY+mIQVnnGEaz1n0uhdSbSrkWOwssjk4LlcYf2relOLjb
60Eb/rqAMSGhJXO1oiqwY91a8LKi17eArMkiZdXofAFSbuntAM5CBrLBZLFSrZFv
ZmtbinLzqN26/gFHARE2ATuux6TE6EiljxaXoh2VNGY8UWp7/VBtaVlmZ6squnkP
BivEpMbUX3QhfLlhc6+C/43V/O3doAXGng3zZbDH8tlL+HWI0RpoCYURbMwDhoRC
4M3C5O7Tz9O9NR51V1iHOdrqjwepO//NiKRbeILXoP63IreJ8nfbGFgscnXERjfH
0JFPKX/CMgAgnjdDH2v5bOpfxNFkNgZsCn6o9VKT5cOObUj4pVc4yHcUjsGzohL3
5LDN5HE4PImvGQdi52H79IR/X3+MRAKVzri3FDjj4UquzN4Aykvszz/6LWxkcI6n
jBYled+l6h2GE8Au5Ffy6zcnsCjq4m/lyBB/vUqN87tAfFrG950Lb89Lky/C7/ES
HhHzYM56gM59r/PkxpHO3gKmRXAUbfeAkYUB5jrCCctdV9tU5zSH2AFp2McBRGKl
JmkUf6nSBja8DthAgkXtrV00FAhDH6AWpvEUNrzdoUP+jGGq/t0kEMeHUF0xa4s6
qlMO0WumNLG17yVIovVwpPZaPuyI6goPwW9o9v6fXOvjFv42X4ZdO6Z8Yq7g+tz6
OZ+rpTTXBxVn7LSFoFWJGywaaiYIhGcVqkGssa9JTtPS4cCaQvApExV1GPNLEVQN
Ti0kn+RUTH0NrVC3zrmCqdkPxs+cudJeKEuhNa3+NulCNW1NJSAPeRgvOuJ1MdgM
wUkPd4Jg8xQuSKcMj5hnzzi/rywffVmUNTcw3mI2lSoI4L/QnwRkSFXhlYffaMiH
B+Y0HcL54s1B7VmBXcxaqpoKND6mFM4Ye5icHXJ497wOKpqDn8N50ICtJ5f3xgjd
ZIZmqIWZxy88iV+1EQDy4hxKgDn9nE16UtbdVYw7VIuHISFjWS20vQz7xsY8bU5D
bfL+pZKoncbyjbQnCcKHy2yM+SJxkQuGrRJuWp2ipeuoxKn8n+1CnAoJxSjlFcY2
6Z+Ik9L0gIgkesUYoA5XBn+Pmg+TPUjihO1xKgzIjcDapNvYAKUYIkCXo8ycZ8c8
b/+YEnAVP4nEuDNRWnbHJ19n63fiCrNEDFI3c5OGtcfRbEfLUO4CCJAQ2vmssFRp
/ym3L+ye0ETph37zmS4/h+/8QIYSo4BDQkFGsG6DEqZ8bsnIrJmVXkFBEUUUHcoT
9vCJPLmvjIjI0/wO9YMMuzp34pEidTllN5n2oKJTLcprmJvSlTv2UD4zskpeka1J
E2D0eQS2XF7ow+F0kCPmc0ENIUR7DKyak8/B0r0806Eca2SrlymhroLCsmNd/dsg
43HWxk5m/wTh8wEiup8wvQeO+TSt45UBSOEtbRLeA2bqtyQzKJlpcu/y1jcKECCw
RzKODMi5wBl2TmeIMoJbOozkAdUTdnq4i/PQlLtWOO0x1FxdnKDsYGqfQ+UVSe/0
q7SGoxcHTXWQ7Fjfe6o0ajHcWXmyyLmImoBrCsoOAihV4pW//p0+VicrkIy5gxde
hSxuyLHncpmQLiJRm43Zsf8JwycKzJRyiehb2b4RDXU1X1rfTKKkIPA1UmgChuY4
Z1mD45dIiz/zrwS9YXK1+nzmFnb6qWBUr4DDUB4lAuJ+IPoNrzBki2GlEZil+wG0
oEBI55LNjfcV9YzJHdFgLmxn7W0mbizPzN1Y0vKfDKSjrDebH16B07ztxOBn6Nmz
0SD8fKezTxK7R2Ie3FwLGwMrgFhXn6zh4aqXfbwUXT7Rvw6v7yLHcspg/ZC9GFm8
itquVGn220N/5X9ONuIHAL/3RSe5vs01kw5v5w4ACsgQkzCWFdfTcKO9TkgJBGmE
601Wm2oyC5jOfahjHze+pbeUqxU5FasJg48+Dit1nqU9BO2VipErphIH0mL7hU5N
jx+X919rmS83tiCuXhaA0Eq2GevyZz/Uj8qqO9JCIe7UKyvRe9AdQxPHmAwzNOGR
6HtGk6sWYDrz30BEOoGuxruR/OIgWxbr24EvWfcqRSdlM/71U5TtNrRtf7aIjqcK
hM7X9T9GIbar/oMtYjnft63zRd2vO5bD4kA2vLc9nP+BGQVrSL+6V6X8pVLAyNKg
xx/IsMkGW1++PvxUlWV5FyGVnzxf1lHRDkuHsqJf6tWkTgMw13QzhX5Qjif8IHGZ
+g2NsyomWyGGcPHaBPD6WnR0gRWCfaCPUt8NCJ1veCI/jLTlxIMET+Lfdc9iGUzA
xEC8ukx0qU2DcoQu+cHskG/YWj8XqqSG41S+yXChHJ00lFcs9/MsBO1MUvVWAL+s
H9OKhMVg2vlz0kDWgNalymQV+t29836/fevNWm5156tZyu0h95nWepfKkXGKikW0
J7aWcSrKGdzfcH7KhQZ+Yp6i5e/J+vtQ/ikmgWzqvSIXnqfJ1UaODpuMy9xG9KW7
xfZfg6baab+dnvGdKcLgLCKy5SoDyBILSRvu7QRmh2Div41MrZeqnmOuMP+xWsoW
4gz9sTrVB7/v9/ltqSLDaNNNT6sp8z7UpbM9+26AUD4Vn8MxXkrz+pNO5qh7+X9x
szBohy0cpU74xliXRE3PUGcLdn3AfJ7S66+ajzg6MEjSx87JU+o+A9EkjSTkDo/T
7R5aavm+9WEaWxICqtAQyOiUoRpWrd+74OCpQlrGZ4YsYd0BemFaXjyeYkCPTJtY
j3LXpab6SaMUTrwOTw99spI66RM12HciOWeGCnl3LmmngKjJiNaCbI0krrAWvGRd
fNJiiTMoBtYVjleCf7BU2Th9A3hlsBYK+rSeCuc3pKGY9xGeOCBZNOfumfHyYtp4
xL1sCi/qzYxvDZbdOXjPD2iABJXQGLm6HFTAuRTOFExTDEik2T0j1MRuOAtxZL1u
4YPRGgJ9ZL+BWwDQOtAHMd9Ps92eATr0Rb7hjrtQlU77Hnxzen+M4xYBjG3vpoSI
2z/JRoXhPAoBsgh5rhiBo88cCAmi1L5nWTkcj0jWtWVF5drj4aK+pTkDWQPUIV0k
gHCMU/F9sgSBJwkw8FZshITybNTwAfSl1r2kjDVBmFNeb3IAH5/ARetrCpjGSfjI
2BFc3dskL/0Jx2eSkcSmdqXhGV8GJAJ/klP1GlXR0V+pGRbLwOWN8Byu+VFoA/2a
H8jOp6FTgPiy1S4qVswuVETe6cb7YIeuxVGMNbpWaR56R1M1zwqv2sPp7uOgHaYj
gZcSW4SerDx+67asePUC5bKXUjHD7aMphJzvYKeCmAqo84qIpk6P8ymaEXeUrp0I
ySpZryElEv2W0P1CDY+y7CCsWhFyQD3x3gZIcQiUIQn+SRZMUutID5ysZnuhN2B0
PHy/O5XFJaUPQ02u3GdC/Zwv64mztn/f5LJG6MsjkwhybMJ7GVufgxN7EkiyggGn
s19WD6fUp75mto3C5fwqZ7lAlaNa5osvmX4TUmXbCHGDmcgNRMszKkAS6Xh5Y65e
ciZCX3P4sQN2N22DJEx5/N5s1V0p/H+Zi3W8jp0AtaobtVcAkEUj9UPYiUzqLfJD
h6ZgWOI2o6wTf0viHgFteZC/xMM5ynO1NmqEuF9JDKNdoHC3X5fLIZWXoKnkxeqq
IVAN1gs0f5ZwN+hqFaXMbkWtCPsTSpOnd7w5sBgv3NKDftw2Tl4+zlzFi4VMZRYA
qaxPUZ9n7H6CzYXfD20UpPiZH0Q3Bz+Lno4rBLAZwXY7FqQ6BvzAK6FP/4VcjYuh
33azO0ekdyCYnrFewTWKt5Hv1KeP1TuAyxGZD0e0E2gvYxq9XGRVSy22CYF1nuLG
AehhzctGIqhlOBeBHklquT73c+jCRY8+zemXWbxlDLQKfVG7GnZCKeFfxWe4Uqph
y/Sx4lhh6NlPKDjmgShh685FUlz0dT9EmNhJLs25irfIkWGXV5oPO6Mt0agIMY9o
pTvGojAcaBat5tDgkKN+17eL/ZXGzJJIFe7mYs4ajBe+BpZX1mmcvzyl4a4OJgYR
GX4s3pzs5T2HsgVJJM7SMu7rtX/lwhONqjT+ZaZtKEbP/P6QHevxR5KO80TJZlTU
KuVnrlDn3eJbVnw/W+nGD+3nqP4Q05H+a4Vr+tEdnVae16CQmCHooaF9R/+XmYaR
c2qecsG85RhI9Hs7JfTtLzAea5qLVRrLyVG6SQ+2z0/dN7QLitjyXQ1i5vDm8UmQ
F0+P/cxLSpUsWpjIzfSbms3zH1ypsBMjqomjoj0sQnwS5/BAJYw3GTNdjCVpnT6b
m/9GexhcnpMjCxK3FMZq/HnjLFgMBEtObyCCglkw+xeh74E+aMRnWgSB1kfJVKqN
JiNz+BPfdPMG55QqL1xMGFAZUUzcpugbJR/gNGAttm8Fo8pMfAjk8Nv3pgzjIkcx
I+l5G1va6ax9gqtrcRgcoZZvkHQeaYfFQV21t9zO/pGZ4F8Kujz76nrd27fsZ+cy
Y+iZzC+T1Vz++SqhqqnZjFQC7GFYy9cqAxn/5IAk7imOK2qc31x3QBIdzq4nrgWw
BbzPRs6Ceae8IMUG7QZJqsA9XF4gY8vGPv4A3ahqHpX+/QKA/hKgbzkhf0CLNemh
n8TGOQsWD71dFBtg7Y2LM0twNQSKrJ9hLc3/LKyXKbtNFmwcaVgYTv/+JmbQwYCX
eqbyKI0auARYBW8AGmPj/3cFjc6Vg4kyi5Q4k9EJt8vLpL6DSlisKFnlezb+eQlO
6YLcdywkUMsq0zsfcGjt1lEPCB0/NUWIl9DuiBSaEaDYOGP5Iey1Iiu++Bn9dqf8
GQ4lL6zSYKu67l+RSqAfpYgPXfjXa4GSwwN9McPnwZ+qBdFKNLNiD0Paq7cbQ18r
0zve2WPfG1vMrJjg3dK3z0gHXZUBO4cnp3I1i/bgUYJMC+DtLHmj9PJwwKPg/CSa
99sJ6wcCg2VTN1pvXJulxwNuocAbfD3QeI7h8OtxM0Slt89R8+SgIHFJW5Qo419/
Oz//xNeHuMkkZg/0aosURuRqqspyJte0CGAfwq2ZDlUdMZ6y1vNovC3+/+tLsQEe
f8Y4Awqhw3d5SCMUXko5cLa1HoV/dSpkrqykoTFnqXeB3q9S+Xc22mkcyq54mvH7
zR6xIqGEMSBnTI5PIiLGz0XHGUg95cZto7Mf9a5u3vCqhg3P9op2+14OnPCq23KN
MAb81icJlFYMQEXAsJYYm4ytwyG4ChEW2vF4C7gPZL5vub2fMr9+rzWcgLYWlZIq
2Br+fDOjb96mxg6H975jl7HCx7Xc63evXdLtUW4C0Y5ilYJNHckjXZajOkMIBshm
oXUYTD+/uW5Y9JrmMiIW330B9bcE3OzeloXJLCFL1x+qky5zKAGYrVeWLuXLKUPI
1hbzlI5OCMcmTFw7fZ1hwQvjmuSoiGN+NvzkgVaV0Rr248ZI/UhQvhuTbbVY6yBu
xsxGS1x5U2XTEIdheYLCq99Oj5sj3BEjxXgnbz7lwdLdU+7PecptRMKCmROZ/tWi
Jh6xWFjlAEvan/w9CFvlTDBVkBu4Xb/4iJfnXEITPdXWATJ2SfBOY436fINzz27Q
8UnPZhYGREyIVM2TgCwnfQQe7r3tGAyJIO/qCise5/Dx+IPyvOzQkQskTp01guTE
njr1UMno81xdt80tNMjw5MxCv9S6o1aVel3sluFz0Mit/E1n83cNXSKU/7TcNqvb
ZYPh1KFUKlJE87SIGD5lNVrxvfH3eVRMd5XqEQNwyCj6QiQmTKJP3nFOUurkqUqn
CMOAWmKcicq1UBr9jQ07f9bX+nuYXyG/zYH1y4vvPdCFr/kP7ZkSGO157R2BXxWo
EpDytbOQrqshRHwXJ+FzHaJ9b/d1oHrTlpfFBTBieZ4b2HyrP04g+GxeKLBSynSh
Lfl78SxDc1ysuf0LXZIL+V3Ji+2CAB/EoRq2AvR+Frc+N431wuOk6gj/Ts67rKeI
p1O2X7IxFq2jVHDpEDCQfY1xKPuLYSXUEWVphC+kQYGwpQfRqNGF68lG7p5Y0kgB
bWe74kfLPOVZmolSpHa8YMOVWGyVnsnjUn6tg1PkM32lNqimjqbIUQfKCaUdk15b
idpUki0xLoybPUVTI5D2JIHwD2djyKGm4PIdfgAAiJSYya2uptfUxxbtqkt8Yi2w
UpdbO+eClTF8IgWacn7v4ifNi/J+EyTP8jgxJwLDmfkzOIGtDBNZybcHpS5acX2H
p90mYm2EpXc2H5vV6OAkzhvuMYQnlOl+LJioUciXKOIu7XVem4hfomj0yh/GymLz
MKxPvk9tsj6NKm1P7wyfw82NZcvKswYtAvO9VvPzoyqCYeOyxqt0hqTIyK+QfLEZ
O1Qv2pw9QA3zLfg2E7WdGK3p2DJ0Cf4Xqg599pPer80xZ+8Pi6kYVl3zCOYcOuSv
a76pLPl+iAoOeJOTipXLkWqoy60efcM4UAMSHm3TN8oUtLKsN1pRspD7Gl/Wz3v+
jVAF852R0sPnd9QVoZVBGr+d/aBEMZMDOE1mW7mF6YYEdpAfhtru0QnuzFcqX7DJ
XjiJjU6LvOaD9XQmu6pVG0B3w7aiiqwz20Mg0yeicAo0L3VoBIPSrinEcZ8ni9aO
UM8Peqp2z8AH0XVe63UUq9J/UX2fR+x1RgodfgUPThCUihkui/B63cmWQijtqGKj
T1SBwUP43MHYaNqe7vUEVbNoVL/6l+nbB1XfzDEAab+MCX10AB0hZy/ch/CxlIGb
TpYHOt+7P90RfUYkK8ZvzCMSGC8p2J/8RWLsMIjNDDZC85wKDsIQup4dlSRt1dfp
dkRpEibb4XjDWw7EuVaWwxR8NsnSRxbZ0acLUf5lMvjrdnw6fBdzXe/Q+oKDXAwJ
u5J3WU6ENsfWfg0wRToG/6Tr1bK6Y7QoPhEulOIzGBqN39XHe+QF8Sxu6sVvxf2q
JHEwTRTT1nmx8Rftsx7t9z0WoNOj0faPfNZVV9U7zmTb2jAPbCVH9GJH6vjr/iTr
l3ok9s6oTJg/F8iFYcIdix/HYtH3WtnXECSqjju3v0FPLdPRVMCnevfMtmFrJO/g
pdpVWKYJImTkzXDkMhivLyAvLcBj4+GA7ifPSJvxtJn1DpHaBgEmPgnHtXT/wORQ
c4JC5nF8oBK3ez1o6bR9p9TomyxTrpgmGzuun1WlHSNxNAUMsjAeHxEQGM8hN2td
hTP+TCHrS6hcNDVWrBY3TLEAKFDtO3PGdKsv9uDcMO5SGki6TUKV8OmRcQmXnUee
MRKevmLLvKZeG173WZf30RAPCmdA4kjb06ZHi7se02PeZtOks6Q6ls9YiAQ6oiZw
dJIPBXy5j0YxAE6xX4pUOpWCwd7XygGrusSZBW6ZOfMA2Qdp8JYiIyA8mkj43k7e
OO7/z4TBmtSychIexmSy8fhXcYCNRvL8wb+u56lCND5RjXrZ/u92kEtk+3wS8cYb
dl6nYxvYyAV2CAB6wnwPTVXgXnkSSaGkSzqQOiY7wAW8S/7DCAS4r5QU43F20k7J
JdtXjRB2FxHBUZfbh1R6QKWNl5b414ThD7Dc3qzjNoIV5vn2V0OLCmtx8aDkFRak
yZHLXPlr55QPgRxQaOuBmh577oS5ibIjX3jjZUdMlw9B+2avzJn1Qffatb7Q3K9J
V2BYVaeeTTMWn2r1+TrwyBCeGJLe/ONzNFJJCyxuIJTP6wRWs26703QB8ahJMHMQ
bBE7C2iAzecOfYLxf1JlatS0xb64rMsQ/BghRrwlLybF2ijN7zDaTqNsW2ZyVPtY
x+tE2QElEwvjTVV5wM/Z/iSphPoxJE3ii11CTNebCs3wBzegxsSN+rey07IBrbZj
hZF6NuhGLL42EewcOCbEP8n5xrWpMYxNNHJTlU257hgQ8WZl+2EOb+mtoj5bdRjb
SQ30dVIiMfFaxsndUhIAVcb64fzQnwjF0WUGo7dOJ69W3f+F5IGpF0wNMQudgn2P
07SD/JQcPsgY427f83ygQI/k8osgTbwS8qFAxloLalmH4hviV5QsOzwZFEGtLQw+
5WkbG6hrF7theCeTOqwt89Z8HM76ae9czhTUsOtr4QTE1iVbyNpsRp/Y27mYv7xV
Fbtasj7s+0x/2yEox5UVqk6djb+qb48RCmO5AvrKxnwERcXk/sAICAO14FhXGrUd
8gz0oKN3V01e0z/dtrZ5ak8CQJonElw6t/GJkIHAyh0XpUMJoNcXfTDRBWPCN3+t
/I6jX0DFWNId3ArOJYo60QxZTQHDP660mAZbjeUUdrvdmbq+7Itmwl/TGtWMZozk
Du/tsq6tn/Y27WXFKG64qpMxPSVoKvxPXATROD4Lnncx+3OUPn1HGKdbBXCUUHiu
bwCvmIMxcYVzRaacz2dBT/D9GLzz46enIqv9PXhp19Md6BhBXCeyB+OJviE0F3PM
mnLhKWoZyBSVFDcOQL4PnP4kaWwaSqZRSB5mOwGMQWqqE62ZVdqIvXqnXhaYe3Br
bHSem97eYh4z+QmSTIt5K19anNHJqb8t9ECNX/3Xmo/VKnnSyZjJSsLUTkEB92S7
27AGxJTcUztKSPycGrS071hyQe+xlq8lbs4wGcw5GJ2eg1FZdBa1MbWM1UO3DMPI
gmo6c+BEPbmNgbtPRfgjS2Js5aleJFSPrsa+Ew5iVselKR7HRRVePrBkuURJfP3C
45FqcPFeGrTVgj/BcVv2XRGrLiU7hY5a05zmn7BtL5JDwAS+Hir/f9j3vHF+FqXu
/yMpyZiRKUIvOKYH+on4R3JGIyezuGtJ/JIWjokBe1ekK+0kFIJkBh5aOHWG1xuv
Zhf6mVBuj1x7RjtXPXL89u2P3G57cRmgveS0kIedDdaeoMVN1ufm/sqkzTgZSwPY
MBYcB0znCVPhvPPRj1OXOOsccrABKIStaqEHGOL17rybcJnQ1G4qEYoQ6R+DJ+aB
jBTfHTsZbkCBQIn+ZYbYnsgDnOwvw5bmXvHx8tbMRgRSDyLyr3Z5yr1nP/KB8k2f
Jl5tLXM7wDK+4fNm0DemcP2ab8/Je5W3rdMSDnzHpFuqbdtYeqGouoGgljHjtail
6VrGMfccmsU8QkoH/Br4vLMyrjcE8Pg9JHAoQ+Fg2WHEmoPinwk0fnd2YlzjS6Ef
1DFhdvnk7PLndQ3wz76akKhAMsjloit8RcedkzxVWHnRMRQqmaq6IPdUssQOyGHw
Zgi02QZ7EjmJkVVIAAJbX2PNhdBd8yGYVt4qRsVZoMThsf7LNEkdW17lCwfSbgRw
6lZ7P1ZFCIhcC+pl0vSix6slSOltZbwvxqQjoagaZClr/IeL90c1HwZ4kCBDciAK
U2WywdmWNBOEQC++QxE/FaE9IRjQrpcTL9yOLVqfsq09/IRS54a1vDh4akYSPsGr
RV2XCeTcw0dkmQGyw2y6x9xlwoNmRHqZpcZWoBfRxlV1991GdI272T2j0rNBtThA
kDfskOyntU6p6kyYN62Cjy0JmsDkkAcvHbuORtwWACqUTrYRDWm9tsDoMp45g53e
uW/NJFhTfFtPQweqdbesCqGKoRkdroXmGPAVksuQRuCMQUZcyX7kotuSDg6pxc+c
M3nVzNYbUxxKml7nNTQbIIzexTrHvB8Zy5SYGZagt0jy2ISQzEERqptkZZNvjhXE
zIlv6/X4VM9cQJ6wvvTbcTI6GM/CbO28670KwViqSJYeVTQDk17otOwO4X03a2ah
fFaPbNJvwU+vz36mPr0nTON0nbd1FHEukbPKJwQtLNJU9J7bFVH6aOX9hvhK1cDY
RBRgHk/RdVLzsqpT5gCZfwbu4rM5+ONusel9BZa7Fy0+Pm49xwCMssRX+Pv86zHd
iEZxPbDRfjmnH6x0a6VkhgrT9foXhNk5Z+oxudbVkOqnPx6YfpsAMHZoQo5vZnlX
J8uhqYwXAMEmlLkAeBtPal3hMNNoesk5uDsCniU7ZHXs+oziCVZc7g4XgcSJE/26
PFAybRGSpaG4llRp5rApovtyzn2+MJdphV3D2Ga81XKKbAbuPHGOU0qJvW8f7wHF
V3hpeVO9jxIXM8s3hd96mAIG2Yy6OB3GqY2gaoR3rvgNfE380gv1KqToYWGOQOnm
Hr+oobD7+syGVkKiwT2KkIE4pPlExglIWeNF2O9+AjIFGHqkvkn4k/HID24Zz0Nh
OI09J7u97ioNrltRgCgwcdSM/DCm/jpIsrnnwyxBnh3P684pQvIur5OaFZOfJ0tf
jRdZc5vRImdvKIeL1g5QzW6pGV12MFJwdQFj6HhLiMFs93EQ/5ZSJwC55yEBOjp4
KHHeGMTOqc+B29rd8hegjdal49rcA01iudmpcuuiMmxYCDObRAzrXaaeyG/JEOPg
Sxg3mceXOdeqOmLzuArUsQUnoaS8baEr5SR1qb8OhFuegfg6hmfAwsOKeH2x95gK
YGXTyocuhwv23u8rtyIQzAEdVKyYXe3firPkK6iWaZJdCzJkPE+a1RlefpUDwesJ
iAH8PgSagclAPc4wbhntdNxVkfcFufvOkZCbKhLE1V2HF2NlV/xYIr1ouDQglDuh
COJZVCwWCprc1XPUba/SNedE8HLYw1Fr9F20zHGh85pPa6JH70PrNYG80ImMu4bn
kY/OiYcx9ypfSQsXQG8J+mseW9g9Yqs1UqbniwZxyDRYhXp125Iai6RTKZp0ZBzJ
36M2ACzc0HvOEPBmRSGgqbygjFroCga7s5Sg8+X+DtG1egLxUHKLTm+LshMf0VlG
au1O77kbJCJl1oJ18hCQqOHfZ79ZRvKE8m9NnKsBJ1K31ulDJpeE5rnBhG0lpo/I
FbLCLoe7jRpBapIZid6S44R3vdlbbMALEDeMYJXjvSrmwcLMRDzXhoyQn701p50L
IOoWmk4/0azzKQF8mahoe6jK+4LLna2UcNGE+S6wFYg/S6ceq2NzIQhKTSIWot6l
CReLuw9L3JOhuHNKaBD3Gkc69F7yIoNR4UF1A/RuPJjtpB4VROKNRn2g42lTeYPc
BWnR4z0vLLtWzHsIdzQWjKRMK+0aS1UpqGYn6pZHrCXE//N72Yd/hlIY6cQoHviN
G8EcUm4tQV3fAtZD6wr/7SGNPE/88OfSu1w/T0Jklz7dEjf0vC3kXONE7stoDaiP
QHN/dkaNcGq4kIunnCL6NizSvbqsnt9EtEC6IGNgzNNZ9uKHS7nPt5r1ZBz44Cp1
KjrBp7knD9OTg2m6uTobLWgOUPOfyMRO0DVU+3RXsAp9SE8FLws3bl3+DuvA2MuA
0zU4zpvP58fgFIims6sCv7X0cwMYwRO7MHtcG4imeGYlZ5ntlj+9wrKz3qpuFtRo
QwisefxkwJqdsInqE+V1qTgqiOJWKXP1MrfMGzS5LGqkSZEkCnpYPwejh36DL4WB
w0i51Cd+4G+CB92yBvj91qLrz7IZFH2VGLxSSPTMAXUinjiiIIVFXzCoLyL8YRBE
OTyQOQJ7TYACbn+UDk97JypqfAkIltj3ZtEZnSt5SWbSUqueOHaK3Mb+2159FQTj
iqPmt4tIaJgTQdHbCPjv2sHW/B3puV2ZbALYmk3HTaQpoN2VzsJ+GANBzq70BCzP
G3Y7Xv1xei+BbuE8bR83Q+QgJSYenFMGdaXu8Ap91N0Ays7iAUPq62sQNJCZbE28
43y+k1rCK52kjKy3Ovl81pEcDL+qwYLEwnbF0fxdcfkgPjKNzUsDEx1cA5YOGuT+
5C1IY1GvmPxFLrHozGqL8VOAwyax7ljC9n1sHWumghw4CSb7BgtDZedT3oDkyCmN
BZzwqknGubxUAsMrFj80h82YrIX3CFXLxjgUE0/cpcZ4DAWB7x0kmPfLJt3poLUa
BX3jcKq4MEbes4Wkfk2dKEBUj7RmUYE5XOKi8m5q/jFIdGPrJGcag84Je4mD0qQe
aMEpHjQUDFdHySQlDMwr/0Tb+7V5w5wtv1vyapxkrSth2Zl1aWAfG37tepoAciiv
1ux6evrMM+5/fQcOeaOvd1QO2xvEdUDaxuh8Y7Rr14KhYK1CDaW6TSAGUp1gTkWN
/d+duo2C9oFszUNLwSIO0fz7GsyVWl7iz0m6/L4JmrWTgpJZcY2EP2N7cJ3AVzkK
5SOfX3clc6cwfvcuvos0KEQPREJqN1zwbtvPwrCZUBVzGizTWEkDk9hkJqZly9Nc
sxY8z97/4/fvBYCjMcW62A/H95I2c453+HuCEKcepQUqV7WhABCGidfTplcSUUaH
aVMzozvGzimpmCLmENszYQlelaONJBBNg1Ch8e7laI7Oe9pscmtT7I/N0trhpWNX
gScaDCBfGSWh6jjdxVgfV/eTPk/pzA/LZJsjhsNGmPThHYn7FDQDDFWI1jDp7He0
fTbrX2FxNnlwYLyiW9cZPRmqyl8qkiesoodmE/w9+0jVIA+b0BkenG8k5TvhB3Z0
vRd7z0kTL7zpbogKybnMfaSey4hxmsK3dgCNFF0LPqjNrh8OPj8QjilvmS80Q1nM
28uJTVyMoO2qPPvW3mW+5S5EcD8tl6bnJPmicGC1HtDWOR1Ojj1b/c428MlQg//V
z3fwzpi1wa+Tqtt31zGUTLUfPXLZmIT3oSmdljXtEP25Ihp8WhNxKiGOHLS+3L2E
W6dTOtuwGe6U5o/RCnLbQlE7MNGoe8oRQ02AU3ZXyn0ZB5gZEB5hGeXQ3Xb0thke
f/gA4mkryRFQ1qFCt5Zr854SLmm1YzZOL0C8nDXPH+poLVbnlWG0IPywgRWYUKPg
YYnEklCzX1rvZ70ZPXLQ+ufKsTDubJIy3bY2rpsMWEgRY+tfzITFsEWcoTxrLqy8
esCV5+IpDdVu9FumEG3P1VkIVHYB9gSAdh1LcA+1OPqFeNdRsTn3I+qV00e5tok7
py2RgV5T9dNi008H63kaCl5UlgFZklUjKZimLiFNSaN/+FfIi3Vto8fcy405jFz5
PYQLCggyGGo+t0t6u4jyp0dj6RLyEVmDjnvWAn4yAygP5VaElOBoxrrehcHr1tuZ
l66kmuoTOFGdnfFkJXT+I/wZYIG+DC/ICl2iiO8GK8/KaQNtWpQTvL3P5U73/w60
sPsa9i5Q+YC8xVGLijK/hlDnKDZaDOeQxCHtuHfs1INpEh3eeGUlUWbG9JsgGv9t
c7QdaN+jXLN7yeZenSjsaZsV68lSupsAg8bRla7wpYvAqnOzlqIoX/wQbvwdYNoI
favY/iONaOgS8Qy9jqZp8f3MHU9k4oHzcRcEXDKOblLAdWqScQX89RdgL1fPADLe
pPcfcHHp9s4tmiXKVfD51YZFE6FVEqLLSTEgt3fxrQwXMMon+1KM7n6+cTFKUQAm
F6BoB2glKvMc8nzLgivghcsJqEer87vhNp0b/9/1KOrVWdSdhsSN1BJ1jLDcTHS8
pcwgw3euysWSaIxgsOzxEmKz3P1t2jslrxAtnLxKYiTqC+ooLohtcKxX5bgpgRlc
CAhwe7iYfE/GaEDXUcLPn7km3p7hds7aUY9C5gDMrrQh1MpDtzCsPqr0CRqKh8CA
SnLTChqC48EYJdBLijJ4HvdKuYwS1zpggg7H+jbSWn4yysXgEWMau6i5rF3vK+u+
ELF2gDlVS08F+g1Fe0gbMZqrzZ9Wq4SN35mKygXWOnZQ2tlXYBxGb9ya+fIsCoEh
0sLIGm7U2QccBPwBaDTy4JVvwhtdpYoZxxsfWc1N3svrotAqQaWn6JI8h7qRv+cB
DX1rsHrOTFbsVconGNtHP1j4Zs/JMZTkQIej5YK6wq/RLGD/rFLiU4BLALsjmCxP
qyKoS1KcjfyfCtummG7tdmYb3hqmR35Fu3TVaCFya7qkeCMm9q2WGy/SVU2hPsBw
a7iUex5aTSDffYimdV2BMTmqXQRbg+TNODScgNGsn9C2rKc0GhHASks3WiDQMVAQ
vZu2gfJx9nvdjf61hWw3xecS+F+4g7TwEhsEd33xO/aFpU/VlmHXlx4PzrIjYpHl
uzJtP3bWRsV83/3jnGWeNVZ+P/JlbjGfz18PEarFoydmEjE7e7Kozg/cyLJSGY17
M/H3KOZ8SeuxMRT5bZf1QzFpZl7GfGzK6ZkfU99Du0gRAkgb25YZ/s/0PrKkZllG
OpXGVVYKGJ34BTBTH+4qmD/fYdLpVFUGjvJU+ujOl3p2SQAnqtODZrJj/+4jP0hE
f23x92R/MFbxF8pPk+YlsVm72fEqnskaP9jUHvOXCuxS+BTcyfbkH65t12zdBPgJ
Wdq70GCuB0nIw7AvljmDtXYTPnKfbyBVfnO0oVlstIjydyJmK+S3JDKJP4NpSO3k
N39skGZY1n352UQ8+g8D1G7K/PojMghicR9PWOHYRF48Yu0HkuaAmboyDTI/vPKu
Y906W5Q1GJ9tLbuXrJgPCicoXYM8zi4CkMjPM0yH80yHPZ7p464RPxIO41vsb4ov
5sdMzqSRkxdH/SQTyMCMtltbE9xn6jmNPzGuD40F5nd6G14qDfvibUovAXUnVOgx
1rJdV9jupfiWKXmsjFZ1ONED5ls6tx2WgKIKHC50WvYzYtmbTikBbpPh5DqHGNcP
DOW48OSzcR5AAPqbpikNCA8vbkTPZ4vtKI5u25i4dUVY0vkwEPppa7HlNGhztDRY
D4WEi0ovHbtKr2l+QZc+vRDGLgEwB9ZOo1S9qo/FG98bpWeVL4MYfhQuDvr2UsQJ
ufdHXuBxNBXJkpKZNIfzevYQ/fbtho7gEGKohzbh5CO3cf9gnOclW/AF1qHvPxnQ
ZiQULo7+M1jCH+srUFt8sFxgCohEcqXEr0PMbYGhS4eDXmKgN1W0s5pepjQWZ/7T
sSTQq/nAa08NMG9Ip8VT8Pu9FXYrVIW+cIyqcDUnkRWFmwLQjmpkl0T2HYSmTMXO
kX1I2EvLn5PUUTSDY706MXvZqij5OAuiNdsdp9gDwQe1VAliRYzVutIvfcvJcd50
N0KVdvBZtGVrIlM6vDb9+4TbcvrCuVQ4IycUGAaWxTZTWXMvBsxk3TFBsAvzkf0T
Iha5ZA+vnQaiBg0vjxNAXUVrSEvR9B+uZS3Fpmc7//RRpOPTqoSR+Bnl6lwcyqxz
4hFqjIc8NuIZfSwFXIH9/Elw/jffL9eQu+Ov+tqFsIKP0dEtRJEDrZT4FmZKSy6z
LaXhlw9B0xAoXrSfSgzxPIDcnE9zU6ycQ52vMJHIP3QyS36vbkAZ6IEjSeKmkkKo
JgNRaaglkwGwLu0NXOT10gaVtC2at/DhHMgJL7WsuVRwIZfoHawt0H1sv98CpmzG
8hdtVVy5V619ep7t5uxL//AY5zMnP3jidZ5lFg0zn5Ya7wfrbp7zGXhqKhQOecXX
YGTOOj3+AGt3AvKwlDpbC+aV2jHd1IQC3vddSKkK7kaNjOwhsH08fY1Tu9ShZGtF
B98aokjNudOOLNkF7BFzgvsruiIPwxLxHQQcuU5XQb39DYfxmDidHkj8ER3i8LFT
4sS76nL9FFdhvf4rRaQt8fmxOWWD072sfXoqMdpAhocnjCBKLBK5HkMhNcH4SUJ+
8CbaX9KwENRsdZbhbbP6OXgG3gZdC5WUOq0RzwPNTfI1Sg7IDoqZMAEGWg8uQjpb
R5YHoKaiYmv/weooPn4cwzIE7oMdilh5liJUkgmuN89Cnp9qwyP4tHRd9Hb43wO6
wrf59qsFY2H+AU8HFBsypRCsG5AzJcEc5Omzz548g65DprmtJ2IAj+UJ+W6lu2iT
GzEnyWc40j+g0dWgj761G+yVP8+SzjrKexTWszxSoqT0f1QIU9ZdTOI+cwmauMpG
PTGzcA293ACkLoWnCROIBnNdX+GRMTDZtTJRhVDubb8CYRFdZaKmQmvI2wsVCD5H
4LtfRKl/iCcFPo2aPmzZw2ZUm1vyiyv7rfxNoT4nHWTwvaz6huC0pCAxBx0osIfJ
n5jPF4QBtbEzjIdiJ18obhqKF0tu2OnsuEmBmDLC1F65Ekwe1K8q8WzWMkFU7m8D
M6pUJWS7+lwVoIJySe2IU5MUwJ987VDADNsyKbKQppVw4qOYu/wHKw77cZfHqX3e
jnYo7PqKBQefZfxgUBi7GUMsE81nSBxxejQO2szg9N3A6R1zi59pPFRPgCGjRzc+
jS5qpIeoAfQu9Le3MT+bzQR7hkHLi+gt3VCnkRtE3nPX4uQnIHVRIm6dpIoe1EWi
By11kUOUyqprMsYYClLD/CdGR4rQvsX5t5WLVnzN5DZ3JhmyIzbLvCTcf4Tg4gUS
hx1ro9SESP3k3s8+mbjSS6Hv0rDuGIkuMILw21xtSlZ3rczsHby7vE47qblce2gB
xtRTxHGL+tbUgEEjY8f2xEY3aZ6A84wlnwEDCIsIVzfcjRX0eaC5nKw/jZVxyy4F
9lmkHgHo6ePSkeDXzu5yL4GfzgUVIz5OQdfU2GBB18jZKpQTYT1mDqNC2QD+MS7O
ZnYM3BVcbelT93aeI3suxE5jT1acFJGQ/cyute1wAQYV9KPyNyNqdWEcxBT3S/NA
e9Vikkf5IUpEZHHHrB/F38lKld/RiYQZZzDhIRvQa1u7AOgg73z67mCASLTqmz7D
KGjDR5P6m+qC0xvc4piW6/z+ii8Nc8cj5T71nIlH4vWK45nRYLcaBR3UllEemfki
HPAjD8ElUmJ2ix79Gm/+GC8X0rZWl5u1TtMdcTAHjasNou7B3IcXomAfPKKWX5me
Yh7gA2ywDX0236vsaxVVqvfItRSL3v0cj328gItfCazEC79X/j5qxgWn1rg4tkIm
I2n0II2aR5G64295iMZFNnRlZzip6nQ8GH0lXjR5be2fhTP0+0ErVIqYHvid3/vq
2W4b/AfkZXwWzrWbdbQmbm7F2Xn9OHL6M2x7c+xPzqEgjAMsWoOaXpxQ0b11KWsK
b4VSilbV/96wCKye/iIH5p+cGF2TPDWW8K8tk1KDR22w1WZqmR40uIeIeW/+qroj
o8xJr/n2cluyB7x6VBh4B72JC1Zi0baqmUVUFZz1bK1NWgFqPO/0MOIguicAc2Cw
wn80qcmg9EoBcBnDLi9V8q6Nk7dPRiTD3LB+OytIZfweVnbVRg9b5sBs/KSiMMMv
ySZtVOG97vCsVmeokG1slthZPWoz/vr93Eyc4NB2IcmptD8q4ccJ4Yov1EyqVmN+
pRZH/AQWyzqTk1z+r9xuamcKiw7i/XkTiL+bL8rl7ft8HALuROn4hMIHfNryZPuT
fsd06SgSKJmkjDGc5fuzlODzxeTrmvGkScPkMasIwuHgD1z6cGl6c7qEEOLbBVAu
1jXtHg7PZOCSNGgconj3JR2OJlN4M6caD+1nadMa2snr6vTCbeGOuX/HtFPwaXaU
UdNmPICvvjL291P5jsJ8H+djbkpYAcobvl4dfYbwmFRCU9F4J5wVwPWI3ciH8ElG
IexDKFtOoGRdvoOYaS/rXHUpoBlSs8A5jACbwI70LEcVlrr86QsJyAyv6Hf6r5SZ
lPNM0Doc7h7nKJQCqyh/D427OdtPMJ+xES35MuRZMhVcKKp3pc/HWxdLX98zI8vx
GTYQlHY2UvlCw+8fDVEzpEfTp0WtHQ1y8SqlQDLSIqfjspMIThXAIMBanaCNQXiU
ZKZ3zpmEqc7jgMmpx4xQyAJ6rQoXNQ0tS5kcn3Dkrajf1kD+WFanodii2ApCuXt0
KbkBpc5tyRhqERLuFuHkY31Y92bQGIYl5k7GH2af2u1Zh/Vypbyk37nY8jUJbxiR
f290Q+PTyLufNL87k1oyUFXfXumu7jbH358G6aA4IXbNzinT7O2D7yfH6QAH7v8D
d9f+qEK69212N4kK+bipYd+IItuSVgDGfXZL4vJgoxBnk94AdFXBR+xS6od2ez5D
ZX7mNZYUblYW8xVQaK38jrrbXMWTp35rDpv/LN+bNT1U+cDw7Y2d+o9zL1iC1lX0
nMpUUFmN3XOI4aKvM34b6L15axyAxfWr2ZFLXXJHPoHPXVipm2y+QsnZpeJeO+3r
bd8FickCGUb+B+Useo/wbPP7seVsGnD7t1dJ673dmfFRzs95V90YzRv8zi53Mkna
UlAbnVkGucJLLjAK0j+SNXW/KHis49CTsBhhYohmlLVrKUNvTAV3l183wADGf7Xe
LcgNESRy96ogp9AWQPpuSXo+r+XmrFJJKFh+fSkifvXP0CHs/mWmJEOl+2EBQiiU
/WsM4XpZQuLO8c1NQTpZIbrUhFafmCppm+GouPG00DeO1Q8F6WJrgu4CejaghqsY
DjRu3lAyeQT8itWVBUQE6jEzsOaCYHNqDLfW+zMSVCRoljAfaLXKqsgxyYEaZVX8
mC7AF8fMTJ6HHZfnuKbh/bVSPbDyIBhT8RhZxCzN5ChbEDOMN4VEIDH6rJto/gcP
WW1+0PHLJ/HbBj6vSlwidBEkN6v8S0U6G4U0RCDfJbeEBeiAtttBkA8zN3cMO1bv
NA5I2HH8XvD89QdieBY+8TE2jaf6bJggxW/QNU5LJCcqkBFr1Iy1dGkNSFXTRRyj
rjDfw7uWfWl+kS63w81tIEWdeLsOTeTmIT7o/xVhIh3JOP4CSTgyJrrG1m1SG8sH
54Ub9EbmiapmnuZAwqasUeeY4l5PiUgb+Up9mBAzEevwY9a2DsyP3eEXPH5Q5td6
4ngbm/3j7zl45S0S3FQeoztMC348xulaOJP7OVUPPLfosdFwsFqjEs6XlIz0VoNE
q2RnJn8h7UdjqEyhEXLnAPW6KVjUuOM50PJGA80dBKrBaM0xOI5FDYtcshfbJrs+
lzvhQmbqUPq+JNvfvuv4Ay4mgzjw82ug05Te1ZQ1WWFRXYATBJax18SwgpKt7Fy1
+o+L6QV/8d6HMIduMd3sjqKxf+uSgG6W3oDb8Pw9gVeoGKRZ8cX/JeI6mtUg/bt1
KOh85zrFEaF0Sjx0F0HBtad1QgyC1ELkrXlNjgbueej3yIBWrtAskrlV/Btwril2
BPDRlX3WRmYfYKAMqiBDvKsqMDW1KqhI9JZyYMBz3+Xnz3fJzpyvB7LA/KA68XwU
BeE01/bE3GJ8xHFXUsJkms6HvQYk24FeodkL7Wbw+ZAg8VtcxptYOXIhKDTE9z/6
naSpl4jMqM2AI70IGe/colBxShW+ECzKGy5nJFv9lz+iFoLHSujzD+T7JKO2/qDH
zr1lNICkILimnGlVWEmcBE0W2u0E5uS4R0eGXI73pZ6SfYOvRI9Rw27xiLyD5Y51
gTxpZoA+nJsWnGfZOHijf3GnUH99TlA81LQumOZxqT+oIuCBJ4ECLa+pU1v3Ux2w
00vBF/ZgMY//qU2cXMQqhC2/oxYToti0rUxNUDWosQ0oYU44b59MqHPP1BoHiLDy
OLpDYK59Ng1bXm4ZYrbMgpv6mzkUa+fD/dI4H5AScj4tISjxtfonrppUIqZWJ3a5
plywgd6vVLv0XLLhdVIDnJp20hfCWuVogj5KPIDrhJYa/Glyv1OeMJ2+6Vc2f1ae
D9GB3pNLheE5mSTTHBRphzPfoFiVp8r+O2YhiKE2JZzckclATLY9HAl79j1wL5ii
jPb0N7nWYIvLKAv+0tyVdaRv/xLm3+bmQ/9iENvF7cAmvE6WVqMplQ0+lSMc5Rpn
W+nH3BdyayI6pg6akfd7SaTTLsK7nXgDoDQzLtkmhiMv+aKhLUNpHEhG66G7+fru
22GMkgcf70VQdtgBMG5acql2el7ZAttext4RCKBGINrV8orfvh7JexRGpuUyt/iE
yb8++0jijYI+IoA1GcUKcsYFjvuVzTqMS07wJM11SiNneUWzufNUAciHFp+pgBAS
p0TUbTSdA9SnTQyGsKlxxQ0lnD3MHjgyrW4phB57ZALmherYBqI1yrrvkcDFQ42p
XwSuZy+sHyeS6dxmSpDrqme+tWmxMOfRNmWeGgNw8xg4CCZvNGiAxXYgfb9t+wm9
68yftACJVm49BZGS6gCaKuMnMJ4bs0T/eyu7sDczCzRo2wPsw/15KZKD7o4mUlAI
UyTZ3yI6rC/C+P+Y0mkSYreANUikFCz7hTKP63epE77dPmsc6cVW+H9tA128EVTc
TeEGvA6gjpDGfaOkMOk4pkHmT7DaoVRHAdRLqEg3KCJrbFoJU9Rjquo3z+lp3MQV
ETTHr1u+p/kfALHZHkzkV2YFotr0xEc8x7uKkr07XWvDHY6DRZdHPnACnWehXHBo
mnMI/eO6D+9Rh0rXMYF5Z+rPLBlIXPLr95vvVoNVznKnidYLL2T7nkCXcbzmoaac
ZOFuiNY2IyJnCSLjzBSZQuK8eWUUYUn79dho4OZtrqJI+pO9nzE0+yjEcyNQt10o
6YUVOCo6Jy0rHPgH5yhFMzpg+/d/VKUd2oOiXN8nRe/i1LRFMv9w9q0gggFTWLM4
LtR7/DdSZTvPTe1Fmv+5de6WYARmJvZv1/wRD+ObQY80GZLktfpMTiNNhZAWS0hj
MEbGTQ12khpc6Ic7HK46UODeaVZk2ulBiqwlcIMHjPrS2nccMLrmTpD+gif2NNc/
pKes6GLzdgAqLeABcAvaWu9xm3w+l0iRat9pZLscAhClu7Tv16LpVlLQ9jhBamXa
qMw1f5ATswQG8s2WwHmcnLd04E7BThkp57Bx9N8ZerF5lf69xgiw+QGYYryi4i8X
1BGUErfvTq2vBKTMpFzBBjQRDNrgeDl3k3ELFZ5lr60Wf3MpkNN5Ta4mr8Lty0ee
ydozJfQzGdiW/CJomu19yrteag7KYslzp/K9fSDGZwbgoyqWDR5pSvXRFgDmiggO
76Haa7wODFWNmABUwya2VzPnfx5kuNHqOcdMUcwraAy1PbhI/JCtwfxwlUDde4PP
og7NSXTHyOglwuUrHHLK8uMoMsWXUhMA3+R5JUL6a7GD50sAQZkv2XviAmlZF1Ax
z2O4udW3XvNovFRheEd5Eku5xYigpXeYa7doSWASHzQxJrcMiNaOVbNbibWzyFNb
LTVGIKHfgf1HreaRTY2NpEldhxmZiE7lrfaZJq7wOUVZ0XrFRjKlIjhoZRSOIKip
mMxf/SUBtFzVf9IzAvlFDuius6VtWan3+ltLjC1urOnn8OFsu1exyPzQej/3v5+I
ELWbU0T17EMYP3df9cDUArqntI9PCyz9ERBoQ6cS2B9QQ5BO2E5dRiPqihV/f3fw
IO5/fco3SH6/jj05yExvVwqhxbnDkJbPt88hK6uwKDM2xcaaYf9GGqcqGxXMnzml
HoKKKf7h8w5+OcErIfpRb9rb+ZUQoUAuhkxR6QLm/Z+gjtaLRITUWJ5go393pP7L
3sI4jYr3lj3vouc67b0A93kEdAm4fb8roQAlIcOjhNMK8aVsu1yN1vqHdv5Sxd/z
fVu/fPaItat4KUGUcnSN0ZE2M9LGyFz7jj/7ESQf2d27FtYRgFsOfQWeuhGIE+1f
BCZExzWZXSb2+V0SYO6Aj3IUgKwZxLIaX6bHEV88RaJaLyUoaEQgwUQXhg9a4Nma
VxbLDjI+roHsyAloTrsQOg9uFryYpG7FJEI6GbEQIGQkgn5xrxYzapLuAvVGjsWD
J5qPVihOK5mOWkahRZZm01eND16eIMLXEW4KPqcV3Gm+vQxUxRYdzzQL81MF9X6w
Y2MwecqxIbhJ7J43yJymzilw5ysgWny40NJVAseorZzrWEbareNCEVh9/6d0NULw
yOtmJsJeiV2Q7d3GSJ5ALq0FFz9y/wHdbT8Re+UGR8CNXBJCRN073AJoRqy/4W4d
RgDuBqVRj7koEsM9gOYBaRxdCkgX76OYuTR69cg0KPk3B9Q7s5+gAHZ4QyApvbr7
OfAi9EEc0qn/jNTDW+uQMmr4mDNVw2AiXJPIqFINRTJmcMWAga9AAx+1GbiULxN6
BkAb/1MECBxTdA8Dnvg2hBFd+PzU3SUHfN/h5mrAir1MnhZJ55A1emofxsP5PNnK
jEaeWjRZqQNK1I/nt6KtN54B/4Ni1PBwIGgL198w2Fhm3kVxnNbrcdheSDoDA1jZ
ZsXcYRcW2CffYG+yUl8O05LUg6LCtnlkya5WwyZ4bNPy8gnRaVpthvPVnpg5mNuF
VYjCzfYiO9kgDphBYUwLRqlsFfb6SBWbmU587jz77uTzIgyN52pyTXkZRanHkv2V
9exmelH73/IMRWLNSKj/fajPwysbFqpfoIj3E4SdNWjZSm6idWYU3wozkMbDrv0n
sT1Pag0Mbd1b0Y/4kAo7JWKqHJKFsFsKGlwvR9cN4RjGgUKzm0DXpxTBBQTPT1uU
kgHFGdeBJBvpvmAJ5XJASLGBJaHHP8fBcFaJt37OHzRqLLV/NFMvBNMijB5SnHPO
NAtDAycxONI1s1i+Qy5JMOGu2UwSjmKO3Lm+y20HcQ91WrszPeON4HfOcdQV9JiG
35b3/akaFzMn2PzugWWsS8wKHCOIHIlPnA3GhuXVgKCCO3KdbeTdHNpjAJ3oeudd
iVCXiPMsjmlhwsVV4V25fZ/J9IjeBQI5JnqHZ9KexJvt0NQOG8uCDKjEvJuKICdk
/oqX+STZfwRLe+bSXhRw+PsC6U0+CDTQGMCJgRzLKXLETkDJuhRInpX3QeIzxgEo
5IG8t1PTbjGleMl9u4PD4n+CSEiw53oN3zolzhOb8RabNZ2frriiaB4KO66cDDFE
joVf3oCsblQ3X5A2y2gh/sgwct1kBvW4n9xPKsfD0+bSKPLkNBOKWH8lGbMusXYc
IiNAzE+CSeMk46DCcNi89o1nRmLCQ7GudjvUtL+x8XUlRctjRoyDsB98OTTNpTSd
P6m2/g76cnt798sTRoGaUeR31ledw+lMxyopx+t3Qo4O+V+bcKBcsqb3PF253K9e
UnLyBgi45L6LAgLRtnQD1pGbnCCF2RviDALelRduCXpZz24A2GZ+iYtJ1z2sQwTw
V9FaXQzhaG/8SP8tOhts6AaFp6nnP7fxLabrNw/r7X1vZyqGz65BB9/tbw2Xr+iJ
av6T9HyQpygagUjWMKUzeV8AW+Tyn1MPh/P5kS/zEq0nwhWkGVagmtmksYQ1wq9B
6guJnWUiOirSBtZKj69tCEWmSDgDvoLblMkZuu+YKmZAmHgJZuppwG/FkN4s7gsh
nz6nj75WpTcfrGMmgpZHRYs8Agrh/+PL3gIGUQj+NCdoowGCXYuhgqG0NFcumzw5
5U3c+/iKPLCNuz0R7OnS47LWZnfc/F2xvGoRKA1t64QU4f6my0H+d5hSmzcZToMj
gTLVugn25KpR1aYwoIzD1t7xkxouT+hgL9SNYElDt1cijn6ojfBDYtgGEYxO9pio
dnoENr+ZWp7c09j1o84ImXt2m/aqyMbDkhywy/1mEY6pE41jUu5Sx2Nz8qMIVrJ1
1Jl8fAEk9HKgykkobGrvtms3H/C7L/SAqHA+uQqo8qkwCYitEu1+/jLYzsfrsf6/
8xI4ytfXB0/OtaO8rARVRcQqSAufuZQ9rpXPA3C05yNLdHo3kByYCExdeI2N9utr
wucjg1EpIVjSaIcGYLeYna2BSwklcTJwxiTqTEOM0n1E+lTJUMZteHYd1E1GPh5x
XA3mQELpVPw9XYxwmIiVDp0X3sNFpW+NCvAddmVYLoC0kOSD6SIOcnWTcxkkEgin
5grQ2GPhCwl93ecfPPbxoCX3gpxyLB1DSAItPIWQHX99RFxSX4SkDv1h7iP5/jql
1MPlabmE6pXw/toLtS2zswjZXYyl2UoDYu3c9CROq6vwjseRXhIpV3buWWb/l8KU
sgHNkhaJzX5PTGu6NCjY9p2ds0P6P9KgcCQhnbgZ/UN/Q/RnJnRAXCCvKO7iffm6
p3VaufCQPetQFYI/NZw8yE8qJ1aj2ZUORqMftAAJ0C887U1Pf6eAr1l+/nGCdvT5
5EcyZGCdmgQMSO3i4BW1glEa7hdJu+mctHak70uzgs8GTOKwzWVHGT7kIQP6d6CZ
f/8ltmiwpxzfyoXKDOM4rGLQPog+P5JuM4O2AyS++03U+OAS+vE50rf9o+v2KtkX
MjSiPXx/qvblexDnOFXT1sMMkzOhFuRF2fmQa+Lx+nXbOypGIATHCAxTUGxi9PCZ
ukFAsURWbrlXrEF6dkwHzrpls8FrargMtW9xhKidJqpQPGYmEpfpc3r6VxpVN39w
y2hzam3oKfhEACOYeLf0h4LlI8JndUAQy4QJEuMDYX77oB9DlZXvQhnb7wYUJOiW
d159mE/mXor4QfyRrurWrDKi45r6U11yd47qgmVjbjYGixmt7RsE2kwlGrtqOZSh
KTR9I0bFp1Lf84D/Gcs75/tXF5yxyP1Gb7WJ/X0t9dkld0JCGuS5Ug2qxOGkFZ3r
44LhrHY71LyD0ENGQrHUjiHs3djLJc2Ffj/XkdEK8L5eIIwG96M5R6Liv8vsbkSM
cH5naNo39RNRxY59CP4prfB2caB8DRISEqUxS+Ht0VC192lqNEbk8X31ddP0tqpx
zdNp9NCMVxFlvGdbpIzfUJLhYRmiQEVx66fsgaFcnkjM1PAA/X5M/fywmMyHgo+C
P/VhKojdmPVIcHHUNuv92iWjRWlgIfGOHiYUYuTj7cLXd57gVDlyD2/rMV2UEyOT
P4o/FG6UCKYBK4nf1uW1COqWgwipN58SvcUtFjRgB/ZytNtkfG7W424Z/TXG1bNP
jvtSmUSlBFYfOXTS9FycAo5fBuvuS0ePAZwMhGkEjKJ8WqyvGfy6WlRmSQrbCrUW
VhIn4xaaABV//PDHvPKTKDNLCLAlGR+kcsG/zH7KLfrpU2tGRDrSOMXsePEcYN+y
0J9ZIirXNUM8ONnTL/s8SLEu3sLTwdIe+VF3aS5SD4e2za6y1MCYnBsvXVKt/xw0
rT/wr9/vSbCs4B+gA4IX84t3jPCpQzhwjmdeQDpjaKG4oGFBpUs9u+2BsWjI1IoU
ngYe1/U4t4p2wSIXSHkRFDMZet9UZsVdFnB7yvzhjsNAI0xkTPPvUSX/PQ4ToGnI
/mTwFwSO+KKjHXALm+6gxN/jMrBPeSP728QubH+WzMQKD49UHV6En+mnqvizq0ZV
LXUeSMZCdKq+uKoldTkGuFGpBRc/Pu4beuRFqwYUgIEbpEm18t4AYGawblIZBfxK
0md5QtU08Hot20PR7T5zkubH9ftN3Oqlfnjxa9L4uPCw3hy1PO6Ww+cXUGwFBQI+
X7Ugya0Za1AGJeMsLCqFTmFy+lwxtiTAhbty0RTXaGz8BZzk2g5KAIqqC4dgqk83
DFmSoJHhucZ02johRh7WNEqLuYQC3RSUul2e0BxmAnLskW1Fz50Vw3boe+8OLHUv
Z2IIVHSBpUAGgw1MfTm9WOj3WQ+ZFR9sQt+ANR0faHtqo4ACVOWHgLEgaZwM3E4D
823dGwwg28tnsxHOZwc4fuz2P3ftMj2L457wfx6vHqhrn4HBtMDGwP3RhxmV80O3
s8O9kSsvK6E4sUtNLvwbMzhYj+FJfwXrjcrvEaoIfkEv6F70Plc9EFpQ1jNnRlsU
yKkw/GRP60G/uzsUI9Btumt8R46AeOEGAG03Rx2R/FZj7Gq98SUcIFuD8d+A1LvE
XNbnljmMCtPfqYKtjDkwvSefr09FaW57PxP42E9nNKSCJWy2QBqzxNYyyKLArTUW
CoEO4Ppn6uPrxiXyFVI+WMMXRqwsO6HXsBrPkGeGAfKmhUchJc4wGNYcMx0mVsJC
IM/aYPCfVB/BCDZp7hzaAlfJEAQXv1YD6BK890Ouqdgb6xFqT9kk93qgRN4TXMpL
XSYi4LuaIKZ5GXXJr3JRfPadCLNA4E0xg0aN/hlI4DuDVAh71PQtHMoK7UQszvHy
n8w8tdnISkiPDpuGrNr4VxLCIbfWo1enSmEgMjZhW1q4r0miVQD1b0bsBkzCs9jT
58P8pXKdq8vq0I6s5RtMMtHcH+4JFAfs6nA26QyO2SQ7fPKFuYKuYDardWY7NKCk
K2GOiTjrGc1rKrya9KLa/8N5PAsRo0E4GpOw9ABH5hZLkkGC6tbPSnLZ43wmT9yF
5zR6A7GW6RWmJ4OgwIU3yg+44NF3L/PsJM9zhj9lTCL+mQH3TIOyYh713iYDlaHu
WNCmW6eht273l6OUrIWY4ExQKn4k9QbIXgQO3aUaaX73JP/KIBV4tcnpT4kY8OPL
mMO8+C58tSJBVdi/aDEUdxSKpFRGam+jmoMWLzxDDm4LjUqUFQz5bDS7x80YhzXF
+FEDMeRwLNFAEHcYn3wKgUKRnEjs9vjDH1OkLeg5gmuWCaYs4ERthAMOPp3syqfa
9zfyO7Oibp1a6Y9pM2xoCnWPhKsDfyGneWp4Cx8pgGCK07lvhwpvE7cUGgmQ+EDN
tRgd9XmcC8shDyypKoQmCwQOm20hXfGdPRo4p4UE+1y8F9Pdi0JDP8V4KkIc+lL1
9c9xL9ONuFYDiedYwhoiOTWazJt5ScgH4m46zVxMdL0i3hkCoAYgw8vDE+SIUuuA
T+r4ABU+Mqy0M6ewAWQbouubJHoTLGRd0KWfKoBqSRWIYaipZ53S0W88TjtrIDSH
35T3UGxS/xXHrSLJBeTEVWaVh1riqMjLb9cFOgldm7LpXraZSl/sUuuD0V/StuCy
bD9VYl3qyIi7vjomjzwalbo1IkXlBIQS1F2ILAvf3M6nmLooRvKzZU0DfbXjcrUf
IZ1k9o0M1NsjhKD6xQpDQckTkmmGABOk1Z4nPHjmuh0FjnnFW3MbGk7HdddT00x5
mLd5NpeqyOdXNCNiQO/HVvz4PKVMVmoRcMghjzZqInCZsoHA1DU3USNXx3MaCBDF
qOjHgJk9fuFtHgIy3MnvoP6OFePJ1skQlxpDLSBoEqhg+v/g/kLvJkep6e9GCrvj
wDpACsU5NhSV3gowGSi+GdcMssSDSBQxSKgmIITPdt47mB3Ma+r1w2NkK3pcQqPP
T0Xny0o/pdmi4b35nPmmgPTS7ybtSLBWUkHt5Glou3nNS9JdBAZTxxDug0gVryH6
/zq4GIVeamF17cF+Tp74J48Cuat0K53Sl69gU0MJgi0ukfyiAvASnTglJtPYqpgH
84322HRY/d9mDx4pmXKbKTPdYdaEB8FkfG7Xnml2IwtDW8ZMJioQXa+uIztDDm55
oEPg1hnO2IGT2wwLGHbC8YmqWFa3G6tcmdLwMdTx+ouceZ9N1+O8YvRH4lhiXHe4
uKLGNjj/+qt1dZ1hG6kqI8aMmMkGatit7SB/bnp5tMt1yHOQNvhnoacWw6u/2Xqz
F7L7Ezhfwkn3oIH+zi+iH2viRRL/iVPtdSCX2QTXdSxmrgxOFXtZdu0bKdpJjLwy
zY9GCnOOm3nC7uhwmTsLvCu5IwyYGRngHd4mTPzuYvICz0xCHSL9ApHAgrH5pBlg
Ge35iU1v4RSEc5bS2uSpvsJ4W2YfweJygVStiB+Xx6qqtMdtcU2XUBuLuyKdf+Q0
WV/EPxCMiZ6avG/d4IdC+rNWt/Mnc47NRhHiQtn5Jpj2EAmihFM8PeFU2padwc2+
QF2bQb2M9poi78XScD5KtN6plMrWPZFrd3i5Xqf8ifPgPrXxAXTx9F6D6CE7IADd
N5Iyy7pyCT8PoXaquOcEPEsWqE93jSmpQUJK8Rf4WBFk/2PwSfJvpIH6gm6Lc0Jf
T05gcUF6MfO4qX6Tyww4XUOnIhcfUfitjoU9Nchj6Xz9Xo9fXNtVJ0wGaNZPa2L9
8CXZnkikmXt2mt+hkRYFmN09EEQ5M+RJZ7zNTt0560T4PPmmVPretbmA8DWEyop0
pukh7VgV6jKLPc0H81kgEOf6pqI9shBMeDpPo9IkrUm7bEpuGtn0pqM0J5QmQC6k
BBMu136CkR/vSRFM242oW7+phOvHtiGmXN8H4XHX4Mu73Znbq0q20Uf4zUBXe66Q
4NveZaCJvm5vJAHCEv9geuQtBmHkVV+W+YuFSXJb6KQafAZBqiZbcqEuexZmar0j
khoWN3XWAqS7ZqHRscwUdscEhrreEgiRLB4HWUMiVQ3mylra3A8xEsb00A/+VvYJ
naClNrphp0jgsxhq9hRjAy+hMYPCmUKDjMxwANQCn5NI63FJzrkwpzn4+CnWxJY9
DVc59DDfHRuCKjbVDKylYRoKLq3dZXoiF2X3dylQbaZ2DVDgKRxTilPiMuPqRhVS
whYkkW2gbgFM6ll7J3ETjt2xn7UCSNnzg/5DwNgx1WT9/g6wA4qQC7Vu6KuQSS8k
L64//DOsqRVdt+wjNM/0K+MJAomqEc/KSyVRAd6LXk8j03ahN7uCRvbAwCk7EGts
PHLR9W8/gBK05Vk4NXrHwU5XhC1RrjVxVtE8vYoTIDYhvr5RDwQHktgqhMpluQN2
jmfSU60DqEhRKeprZPdo0ymKz2gtws66mdJAMYwBzPl9iFVYCOAAv5+wYtUZo+wO
N532PbzPAg8/U1sStVerAKcaMCPMEajUW6CHVVu/uTlORXcqhrUVHZ/Kh0/LKhD1
6uRfr+TdcW4O0axYXsy7iCwb3tghod6BOdsCBF2xxUcA823H2l760YkUpJW9bgUt
do5Ju19E5JgWMkav/hoLgD7DiB7/TEkoIaLa7Ykdj2b+6h5NRKearQOCFP+iYtK1
Ob7sqCvfruzh75GJeAnMUSzoaBM1/sAL/71qzV/YgrLwgoaeKh7JcR/QMA67OWMI
ZOMfZwMOztMHa9P8+7IrbJQrYMk2uZCObc9Zh7OhkIylUYfLsJNFfxqayaZczi0H
1RDw4GmgDtD1rzeTmnC3EYs8bYWnohdV/7I14PVb51RI1KY3WmEv80whsecxAEHt
R4E4mB9GLiWWorxt+KZXuttPQjWRuwtdkwNFAy6AHRjEa92b4Lf+hqAxz3CRb15Y
rDszA1LDT9SoFUe09ltjecW7iMOjr/A3DF51iDjKT7T4kvKgmMAcDXi1ejaeOebP
sjMOLaRBEqk3HPcxrKkD8ZQg8kKXVwSAGhq/faxIud0hDpjaQzJ1u+RxYPYsBZRp
MjWKaPsL8W1KpPU7ZVQ7wk+zTG20WGJjdVolhVZYsqI+2Z7693wWG2aTdCZVOiM9
BmBtugEBvxr7Sgk1MuinvcZbe8kWDWBIlafbXE3CufKrmnxXIXXVUW7WMw9JJG5f
iAz0Lz4MnrwMIdlBIYylTURNY7Clyn6xCIMjk3oB6nZQDAf5+4H/+0ekU1fNX6sU
sZyfBESLz7gnaDuJA5aU/wbASsztRQsAoYU6lz0gLRakfrqJloxYx0xbJ54VXLlG
3DdDAb0JFCgEPwRBTmlC7aXrSA2hWXAVuhLoC/vQt4JOXO6Qiqo0vcE+5VzTb/x1
EJ4fS6Pf5zPgQCxdo9ZAVDQk3rUT8G2dDpRqGOvm5bUTQC0e2fgnUt8WU3anwdrE
D+2Hk+nL3POAnXzU/ExkKhBNMZg/sJPmBadK1Czh1nTqHGDtNrkwlOy3PTDQp/4T
R3V/Grtwq2l2cUnJD+RJZWxTxgKRWNL/H+UY3sg8TRpG6QGEAFBTNbEiRIaN2Ms/
nyYuQ72Yu/TyF17GDOmBUNAfXhx8Az/uzb3OISX4GSqnSMEF8mMsPrHu4vPY3VPF
NtEYw9IAES7XT1hjLeXXRfuOe26PMaG6w/pm7EosY9miW3lSc8oPkXVjBlDSIwsM
Mstu0H+7M3bD3sUIxEDQD9qOiZYHsgmoAGeHGV3Y6tZRxdFRkN2Nowua2H7i4wX8
DO7yu100IB+qa7twrmQtjTRvMXrM20ai83alzZbwJF+UDIem2y4RmNouCKMPJ+3c
923N8uXNckZlNtFmbiYUsIkC265mA/Qsl8extrexHv0ytwza6WFw07Ef28sQzdjE
FVUsC7Hi1w69KEPKJoE8Ft3ZbytoetTHpnYKNBhBFZWk0sbP1grwGCVEAqz13+49
qVKYkmlEkz3kz/Ms0apypnZ6NWk6oun71i08UKjQMYIyaYiRSMRm8w/IcfgQlPhc
VFf172iWbrA8B938AZPwzBZoQzJ6FEziGtp3VJka5+xsGOhhP3noMv+XhF2PYN/i
iMAJmBIn6HS69boA4VHqGp/pbn4FrQSGCPKE1oAM8LDZjfJKjamKgZ2rKS4KyezP
exXQlLLDjE8tmL8uwBreKzvzsmlmp0sE4qRUf2oQEqaIvPqzTnyIh5bjaMnQ9uCu
XxFbbzV2FtWCEJFYJwyAFLd/8flysuul+FJpPyE1bH4RuHqIT7wi5UW96trZc6XR
aQpya4KKyF5zP8JTGv5qFLz6tTyOrsfltFWRgV66F5dE86xlvIbUavkv0VhQtsV9
LC7vHwXOMBnMYExiGV9YQHJL7nbQJ0IsvdnFPwV/qaUn1v59Fib+bzC3IP9LeyFh
1V0hHq8zMM9ofqwztgADP8szBmTia7wVAvIwXcddX8mzITiS0QiE3T7dOgikp1uW
8G4XTYP+SGxpGXlXHZb8nF+fJuGSMUJRQk9DL8fq6l1nj8jSkmeKoyHHmMjy4QqK
egTpWCWfziWa/6p8N+KbxDbNxG88eDcWnAtjzV/FFcwG7fQYQkzg6Q4m4d8jAPR9
eg7c/LM4NC4YO3nIsgxIZ+cHbQhCBiwjLqsLuaBSB9Kq47l/4Kwd6fPz1qo33VVf
ehXbdRGHe02ZkZ715YZPYmW8gPsYTqoVM7jgO7OgiRCYFhUVXbHLHEGOsyjDgraW
5c1teZdQvww0IX0Moz/2xWNqBP1i7sTh3OdYRxh+c5x6SsQpAOpa3nTx2faqg40k
BH5oAMJykeYJ8RcwW5QaxeEUmb+kbiXJ37NAcJqocTJ+i4cP35pY+WQKa/9REfQS
6QjIKh36Pc8feRbbYQAT0nw5QzvGH5bEps7E+4s/YC5UO58b6opGfmWhFrtXBFiD
5bJQQoTNs0zjRgzBH2UQo+aUn7gGY/dJ1M274uiUV6x8KSDu69Uzpm2Fd/bsBVYs
GOqVV4rLsLVaB3LRTJwFntpCiPzRqcs6YjCtG/SJhYcrWpf8MKte9ErEOmgEA54f
PfSe6gZgM+xVdZvJ+5qq7yAtGA6PNKiWP8cX3IHMBvqLrdC97KyLyvMVR/8gpbAo
ejLU0WwpQ79yXIRqGIPzkRAEU7isOidde/WnkD+yhUAcnuYIHhCwdpjIDjj5KG69
fnDcyFv150A1dMS9YjD/6gu/mVhBGOPphaGwbuvBsJ9bGfbvCrk5y+13pFhH652c
ThqXwLuFTHfs5AJPFDvjQRkH1hxKA24prPk0bAAPt/2TQXnVYNpQugGjzuMWLu7x
/oPFN2SPtcgL2EzKkQk20itiugihEJTmC1cGoMcgO4LuiA2gsZBdMGBCCIJohJ5P
BUijZCzRAgNyve0tDqRLadsVfw/E3WuFKw7X+w8fS6NB50rijf5tnGWwuxbJNX4T
/ev3DCwMNvJEeEgtD9KVG5Q3qwwIAxeomx30ADzYL96vHVKhTff7YLNkv0Y4bhgm
aneLN/nkuA2bhgzBOi7nm4XNaM6ZomIJasmlk2VQf5zh4NcIjpMM1OM0cl+ztkyk
dpJoj+LYx1lAhXIsSqFrjQ/XWaqhz2BOx2vLv3/MrnCXnlDqdl8Hnb3ysXS03TBi
yQ6OKAl+Rnhle1J07u/knjndV0dU4lL4ZSmDe91NrGk7MN0kcI6phpwCJgRUMXv6
H5Qi4DveQcyJ4kZA6/95qJwYfw+HIG0IjJWC/VG/f3KnenM33yGa9BxSD4X13BcW
kzRKT7+lHCLMaCpoKUNwYmXXC06uY21G1tXaQdnD+2OyXSckvRsun+F6HK8dmPMq
SzVfEJdsg64KbbBfGacu940zvv5tNwTtcjY52u0+NnNPImIj0SvblTwI/UCdCxJP
NVr1fibsa0++ZcEAFfIQ8/FziGpWQ7KZLj0W2n/Hv2OdcnS81MEawGtg3XMHvTXP
bj2XHCIp1dpHTP9cM022SRlihVTcwvh1Rdc7KauWVUF4dRJYoBzWci2vjPf4X2L6
oEoO/3K13wSl4fJgrYvXwQQ2cjYcq1yDCQgNaDnY5lKwjaeJqeePjBGU/asgBqUd
IuK9M0nlJs5og6YsQjGWNEUS+W6gEeze1GS/RJzWmGf4vhmwazm/Qz3v8Z+K+sp9
9HW6F6fpWEPk8Wuenjo0O5oL1Uw7XtBNJSJTtFrSSi8LZkkvtiC++D/HJuGXaOSZ
fDns3lVk3sENdoihtApx8qNNBWu7XvWOAdakVYGqBezmo3r4hzs4ghB2q/94hCaS
UquQpi/QCKglod0itH9okX8mLzEWTVQh0ljiQxqE6tRAXyi9DSsfpLF6hd8TJs03
eVDHdv03N0dtRb/3BlPwouM5dibrj5TuSiOjut2LPfEsbozrC0W1FZJlDHCaGPzt
MeqfBaXpcFp1yNxhBat1ZSYTQHez58z66qh0nKq2lAHqon2P/VeuFqlvR1jAJzi7
XM+CZHtmEn0vfvJf0CcjURhj6uoyXx311vpY0zEY7wpyVccI6EzkurOCiNR6gqQ6
Y6S+0A4Vl+87NzmSbt+5sjgZOvTboKe1qE9Fvcyt0pxQyp5F6OBeddQNvbzfn/UK
anGSJqyGQ8DsT+fhVX4gBpfubvTyv6vIUQABWmnv+N5/fAHM2ne9CyBuMYmE7cgM
+h7eEZcDJELGRWf4fEZgwD8YmxrFxYyCtMu+jb1RMbrBq10uYQ9gpPZ17oxVJqjs
2G2HKqdsIRqmmVzqjNOp9dRAcmjOvdXY9azEby8voqZq65FJ50TDT+RClNUnRK/1
uY8h7mA8uXOFazhAYQuhNvbFFOQkbdKr1fDSAIO2nGWkJGxuVVAbuugWNd3FCIKV
CbnUBbWvvWf4g8nY9ImF8km8UDool4WOH1o1AJ6gIqyEDdpWJ/kN7mzD/hDCwMw3
j3zPR/i31qbg4TO3+28zPjy1+MP5UZJzAQUVLal+b5kAEqdNtTVgX1fcJr/y8d8b
+F0HtncjHzLTltlMDlwyCeAFeZBCgm5ifF+fWE94rwOdQH0MdMDa7RZ34vL+2jQT
TsA2kB68QGHtzh6mELxBG7o7kM1K/mx+dDSlRvw5kKoK5wc5eNMtGXubh8bjnv4R
mFKm2t+iK2KKdG60QlD0xmsFprNZmY5sS57KPyRdVzRTRgukIy/5Lxn72vwePqp/
ExwxScWqzRo7hgDcNQZApxh7PPiWMhZU+BYYtDjgFknti8FjVv/JWb/5UhkekqpW
AInsnKSg/HHN0O4L9itcSW9dlwryDzOo+GF3ZbMI6a1XKOH0muRs6NThsT8iaFAw
RTiedBvUnETgRNNDDc3T0rJB9BwnA8oR5V+Xaewrhkb8bgyDrm8URgqvX4i33I2C
bXu/tB1cAqpU4xLh3369ge6suv+zP2pZcntidkVJwPB9QgREV7Y3zJ5HUQk/3pyn
hgVK8KRsNoU/z+oUafpRmoVPdeiiYokvAiua54462LnvY5M6ulDrST0Xyoy+jggL
OUsLGm+xKpNrpKEn7nsPnJYhacWLcXNWItMMyuyUTDmbAk2MIbah1LT+NWtroQR3
QX4OeWBJusdur41i4MZcFjogmlZfePgEGo2Es1olA91OI67e3lk1I7rKvrmac2lc
dLPQRtMlDAOt168MX4VgsiL3vKiBGbyET299w27D5LG6EToA8ndWqzBh2C93uxdh
a4w/9qJEfdbR/q59TJIzqrT610IWIVCj4UI6V8uShQlCtc+LHeV1s816XXtcsspC
UxCPnY/22ZDaOaxSRxuP0x2Aoi41KCs7nw4s/BUwT4ZIt+SpK+ZLmpZffuSp3g2V
vlviL29ZFI/aLpbPfDLyEiOWj/oDXYl1+4lQaJuFQsvMFd9Q2q8TIHCiZklhoIBi
EilMa+KqIvj2ZrAMDz6eIqb5KTeEDp8IIuM78s6hZSwVWS/kT820TgnlBFk+pGyR
RsvCXmu2sR26nS92x93DbJiuiYqRM528W4CzXf5WHv/hTVLfa4Bs6i+JJ4LFt+Zq
XA04HS3VTyC5gJnsZOoP4ugVyGACZLSYJ6diD4fkCOX8DJRK6DiSBDPt+rP5YYZ1
PKkFsl49CnaloAylaP8hqvT+xIwWWKy+JEc/GoqOdvE21dUCqLt9kfV/UV5irKA5
LYtTXMTiHYpuR6ATNgReoOVDAR1OTeR0muT9GKGLRxPAihbXIfgIdh/60pEH5xUZ
/MWyA6tiyKBVDcC1l/pcyOIoew/VDMgGaa0OOH9MLXo9ibMZ331Mi488vMymBGIX
AgDy9Lku+AAXyPslba+SelOE2mKXHECCZnadzeDaxUTT2idSTXHDnqIR7buBMhqT
Sc66R1uaSVSZXjLoD8+Dk+PCc6qTjECaoEAyIaE8cpKZ+3mgx6cckKbB88YLKIae
V+Ta2WM0xlD4CzZhYnXJS2Wmn12lQjEUcxJV7a04jmZylNTfeGMqGR1pDH2K8QBp
F796SSXywaZFXa2Q7YeacytY6nfXzsUkEc7et+4G6hJzd/6mNVfCn1buGNBB63Gz
EgCmBmVe1NUiXFs579QDL3zvLK9cpD9PKY9mL7LLYxbjsfu/hk+Injt3Llwl4bBY
938aKG6QIHUn7ubPBBJa7kXbssoTM3NnwcVCtRUVvjxJvgA1Gy6lz8dNl9uh+PMi
+i6m3earRICmI2DarCeviX1LKVaAedf0S00gaQpb71/r8ZKw3cFU7N2VAw5657+V
eaBBLT/rhl5hGXAxuh+SmmsXTYnpOOX59qOwKW0j2eAIL6tePKN92OCZMSzZyHG6
Q2/VqEX0x0Yz24kmHWwcHlcx70Lq9qRiBTD7TCAg+zX/k14yWh2U63BIMWQyFU9t
M9GL1MmWPbjmmGBTaY8TQmMQzvmuax60NsGGgOEDp65Wmeewoou/T9PlaF0nAthF
4ByYbBGhEWNb8bMQtdEVIZmIh1gukmYDwviWnexppPvby/nlo3YiP+BYrg9Ski7h
vkq+NvFwNv0oUXe1lsNv5ZehAJWC2hfJgbizCs1yyx2NG1KLj+izhXkx2nuoXgVv
LNSxBxwgztJN0eL2n6XYmSRC5UgwjbbiUH9ApCU/ukht3qpyhGrOzygDToADAVTs
2fPi9/Wx70ACpmUBbAxDlzZ/eTyeAHpZqXt46woHvGQMUdwKIZwm3bRvjz1YwOEy
lMTk5qGtXC1gvoV6Q2DuzFWRoU3mHoCcTMnzKPb8RcQg7PgYMvMFMskTDoYHSGzh
kPfwIgWoTwaJqyGzjuJJVpFZdzoxm5iL3D1pmwr3tZdeU2zwQrx4hTs6c3yDvxH0
qX0cRwrAzKZffnX5RgzC9J3xM/D8hhIBQRuN/0mzn0hGzQU7jdz/n4w62FqNb48f
Jkrf6gJ2Cd1+USoQVhQ3AQwK+wSOabastzcSw39HvouORq6kp6VkN0FJWBxD8tBw
fWydHlynmEJOGXJE6o6m7VMRbZ+RkyLu1qkF+HZBbFQtQkfqLJnILELSZmECfYeC
kuwQQ5h1pkXYYkBSuPX0sYRblAwvqmyjJryMMp0vIfpVRvKSjVrnC2WhYoNUmdIq
33loiHFhbPps0dhUrQUcqO+3fbElNWkEov53cz8A/nMBjqY8SV6RGMWS97jjyZLB
LhOt2xqfKSiu4eAhewLp7kMz6++YYGuS1OLqEpZ56PuJTQWX3CB2lDyVH76TBKnm
S6vL64JBrd54ciKX/0EHx/GBL/S7YymrXCfc7xvLGrFdUWw5ADO8ohLw5x6tYCsy
wl14sh9svulkhTNoXTDnTidRJe49X9yS+1AZAuFYil+yK77urZXhyCrPE3IThTiE
78OigwZOcv4SzD9mqI7fwMIsivfSAmJXYSus06uNlCBORU9tudQOy8ZBhGA8gWAG
XtNQULs697JF7xlzSejOpqn69v/b1mcx9kvQ99DdoIy0X5+2uD4hhJlL2BdMhx9n
EDzemO8uVFAGANnrH68yIhR3Mlj5RzQW/UunesB65rGq6MzZlhu4OqTCwQ3dzTEO
FzwWktyqWl3xVmcvUdToa6BdBZCqp9K4yeffEnbeltU1R0oTKIUP2EnLVfQ0h4S7
YD+SSWj0vlb6+37j0/1/raFPSuNCOJ7nXAhrCG/AnkCsPkSKGH8MCaayYpVfUd7E
6vjgNrNme+H+3c8IDmqwkL20H0vk/JsC8oyV3aReAN3vCmSow1yRCjzuB2MTDZf3
8ujSKONQ7YwNkosupL6b6mOAg1ZjX/xhfYbXjjJyN+gmdP1x7og+4YQEKE5EBA2T
P6LlriyQYttMY3jU5nQiOPy92tgRxui0gktLQkCNgNAp3DIgnC6W5dMPXK3VhyVn
tlE6JD7nKuLWaptM3CH4a6u8/jnzPOA6TfJb009Qnh84zARxxag6F5yS5oWmJ7HT
HJcmx/FfoASjyq23d0C2zMxCqqlUCXmLBWoUjwJghFzHR0nijq0+nzjyO0QLS6+A
difFOt+bUh7sRmMyYdO5uSdj29zvsmsjAn9KZIjQeHdaH/r1S/gwfjzhZaZBLDSy
jFDjDcWc7MaMFbRMrRlPN0BSMKiOAYyLx1zoG5oJusKy9xFl9BUEk1aoeasXfvb+
p74+SXdMBgxc6Lv+nNx9NNllEpNpGbjXiSJ4knc3Rr3Iij1Y3BZEIpgMQ6QEq4CN
Zi7lh+poi8IXCedwP0eEvn6ot6PXdlBVEhobG3g9bi/eQiOeLAqzmbngPC39LqRw
suYieDQSA3603t+xq13KKh/ofzwGSqHu/k6pWHx+WqaKjqQyPksemUbAtZp34R3X
+aldLXLpIRq1ICRhZww8wY+20OttOEhWJmmuj5lgPwkRgr07OUEcCkZkg+V65zZD
D+UBeEwNs5M7sfhZqkl3n7TnP49yb64FGsC+r3xqffQIaPEMpTz5vpAXlHiTJbBT
BOcdzT3IX2RmIlnnULgBd1HS7UD7OoOurAYOhT5reJi4vDX+5kIIS/ALnJrM8O8g
3bngGKiJqyrO7HZBxT88LE0NddxA0ckZBUA8j4ldaMngcF5AUqlsZWf9PyVO3q6g
xIecHilizoSp9VJgwIAwTvAQPTwSdzEKqGKmXzr+1ZaqMt5BGsSsu+7KQC60nogK
gC1tPhMmHentybqY0aePnfhawAdTlRi/FriDB8zSbMsRzW7flg4CMtQpUHK03kwa
wNsL26tn4eDh8VbBBHEbQEpfFcbT9gKNKO6p1KBq7HGfHvaWaZZKdJf28xPMvhuD
Ixeq2r3p62yV5y3F3fuxLpLET+t27W+DfKWcohXjuaIeDHI3nOGZK5VqBur0G94l
GmiKNomgTkTAoVp6poJAZAueAhfKtHsytCa6GVLOABRLgFHHilFmlr9O3mSz6NST
KUO2iWizkg7v9QyKCELB5earfcQP8Sa4xTmHE9rwarcifswB87JZ2SWmHhyzQKw9
QPGDAYgj8QKx+XSh8dxhOy098MoXIaEnZuvevoQ8WkSh33MW3ppXvncA3krSVXTI
8/A766/njXHrOrCxO/3DVq/xc/igQZWDmROIlrUIWL+X5RsofZbeEbHkx8l1yyRd
ksqru2fxm8IPYi/cdu8tY3w9K4YhlNGZmgO7XvQWwygbYQvImipsT8Y11MAkrIwJ
36oLuDD9FI4hqmuwjYYk+hKs/rYXnNenuiSJj2YUA0eyZcEKsipG/g44G0n8UXZw
vzsOstXc2vCuU4UTXsGexoxVquGDyp8GpkaSDMrlS2fL44vxSIjaryKJJvu7ygcz
nfeEYlCx+gHRn3KO80fOKbiVN325gj6PKiLPK+5TiDK1nZA6lxgQF3PnI5/OQHMI
/QMUusAQHdGg9DsQChuOIzL0t/xMyT1BucjxD1k/HC/5dNaNHA8lhfSExmb1rhPm
n7afGtwMQSlj3UKX8HK9Asq56GPuR2F9hiQRliuDWjpOO/HTCQBNRaUrCkBwob65
DfdWojkCVtGvOXp2zJPrce7UOvgXw05kzMxPXC9y2LnGzeZGI8fobhOCmoDXCp9H
niWDPq6IRSqI1inRV6e+ZE8dZecXzdLcnlcqW6nIyVauYvPl72QJtnL5d3IJ5nbU
5cauXxDkC8qGl42+Z2oFuxySX1tKb6PzXr0bRh0UawkU/q/shMSfsgR4CYITMhnW
h0/nrwAtnaz0BdefkPpzkw9u60gilY0VHdS0IRq+r+wUynpsWr8tMWnYm/Jv9TBf
8x+srhS0GpF3/Cim6c8lkqAtTNHwOnGPe62mDuAWBmErCWCUOg2J8v6pp5SKo1F9
TJjGLpw3IRV0roCZ/NC4/qWaJ3qOjpKB57eXVyCSghCoEldmzLdMLpRwK8lNnI3y
JtyPVTVZEwrgN589+MX4d3SHeSSKDLFoT81hKxQwIOlCVugqL6WAbsnzuyB7bvl7
2m1uz4yfbRR23ZgAA6RxWlqQwvur/VVQyCO2UBugAZgXkKjwZA+MKAgEtnTefekO
99H5kbMSWw5motNGyDIcS0pGVbNnbn6EnjiQtby/uOUasta7g3fX7pV/bWBPLbnH
UiNku/StTP4nemuoIYX0elHkn9GlLQVLdQ2VsvvoRGacWvu8/KXFPbyHKSHYngZD
/I0JUhjYXciTqyiL+5jdhwLGOHG/+bO0BWF1Sj0w/pdb3fX3BwkJAYBif2dwAXrS
ZB/pZVu7qVFTbeFXD4UE8Cfo4xkai5H/rO3sI4MXRT864X+JtZnUGq7xbw/ox3PW
gMz1t7LPoINLt6QbvQq5yOzftxyiNnPc46spsEN9KIAlcXuS2WTAj3cnKzFwKtfK
ceOcGL2bPKH8wEuUR0NkiVDKumLWCHpIRnG3d3DsmpxYSGrFNRHR2JKjetl79fH/
dIpQ+uH7i4+rmFDl0W1Vi1+/X3f+CiargtHNiWjasYJaDRqdbY5+ImZuwRfu34fy
m/HV3+RatmUMjRphOWiPZLBb3jGBf/Wfge7oMzBhSUbdc/byb6cmONP6r31PrcRA
x9T+Q8PwHY82yKzzBeoowxw8doPj4gZuwiEoWLp5t7kpeI3VVET0SeMm1RVyAf+Q
IenmHWLl4ic2j2NsGBEmDGg5zSqZj0QGRoJrDlQHodx7GH2GCbZj7p8FbxerNFQD
FHUyqc6gb5yq3ymf5QVHsjZt0e9nXbSFMn/wyifGLxleHOq/jxAJ0Ebz6QrxBCLU
XWpnHkI52qY9No96Qtf4+zg3ULZLJNykLT+AWGUJYf46699J3gvFAFB7bHOQfPQ3
ktJG/InQLiTnu3kh9TNSiQlXwMp1e7okew0Kc8iXmJLYWr8K4VhQfaHmOdaazCwr
bQgcKa1G649RQOZqsIV4Ga6QOwv/4Fzswk+T3l2cdCoDxywp5VYTEnvIVQRz7sr8
t/Dibp9Ir2mWi20Jl24+A3e5jwYDc38wO1pm74lt7Pw+dcS6iRo3fBDT+j5rxGQL
uCZLI4ftoacLgoqV9TbND8Hps4dpinLRAvJFhjhL/d/N6u2pGMVmyS+pwpJ3sYYv
H0Sm1xA+m9LEjjEmsB2I18ppNqjlqF101OuPtx+iqbShXkdiAcQ/xS1GYSdK2NRI
kNrml9LGV7qmoqrSKEkiwWvJ+uACyvDHHT1lEFH4dTdXQqXpH9HTTcpkt/agbXFo
EA5jHaQb42Nvr+Qyfn0vpJVsalezMbU7hVeVa5YNHAujzmr41lXrzqJq+akX6ghu
gvWPlyUrDwFl8xyvl1i/lJlvUaD6w7zzrihbFpfvAyilCeVg9qlww7/KRJK2cZoK
JfDBTj2BJwBNXFJgjLZvNNITQXzuIfGc9BdgBO3PQce2kKvXD99Nnv3iqIpB+zVA
tFgawx+W8qaDHKMiwylPykQeYxy5iborItfYHPzld5zZ/rgSZmbU2VLcGqcepdMV
XIEQ1EM2C2fgvJldul6zYJzN+wHUoT1HSrZqnde28OIlk7UwD60qtpeRZtjdTA/W
k+CcgYYX/8YjTGcZXrQ28hJKR0PG2b00kpgnKEvE/QFCygzXknJmBdO8/vP+Wx11
V5amQKqVkT6S6Ym88+6OR76XkvSkl/+QBdBKIb9ATcLETpULx0lfJtvEFClOHjtd
Jg3gvc4iZaI27Kyqu+Kr9tB/1G/ooSBaWfdCmhxHtf49TDff5Y1skMbZsknYN334
0JPp8Bxsqtrw2X3DTH5w/wjXAmCk3Bv66/aTr7bRKmvG1+gJVl/Nnk/FOtlq3uq+
z0INKviaJwG7prQqBqjJFsb/CysY05lAIgvNBHKSpeKCr8nUF9GxIN0hrXE0WEQU
OW1HEEchnZl3dr8M0DdJ+bu0LfcqVtRayr4xPXKHtgAVDZOUCjeFdcH/aUCm9K3j
lv3n6tbSZ1XC4rBRJ/ueHzlOU2gudWBaLa23zA4gnYmMC2/ApQwj2YHgKTpMyNok
S3aBy2LIsqCKuz3FP2QiasY9i/Va5omUl7fzpJUiQB6Gfr2PjtuEqGXsCuxPYCTv
FrvTZRwdbobIuJwcX6VoxeSkKRooTQI2FIgXKXbLDsb9u79eZnpKlsIlSiFwaKkE
lkSQZCBe2tAKkRsxLraaY9j4Tqlx2OwkHn+yoP5mUr5MDWSXwv99dPOLO4BHXbag
CY8+zAQExtz64Y6xH7oVr03GV3LYl8Kq4io1KxJAmSWbvmr1XIv5UiqvxXSatSL8
8M7l4LTDG8SNdH1b7lWq3c59WI2qMomBmVv2XK9zuibxz+nEF/AdxHYkUpcsmM1w
mS4PJTx00WypuqUiPTbVsmncZoPuumNfb9xH+GRvkwb4tDwKzPpz7gXZWBKiAJIq
ZWLglhAt76ilZR7vU6gcjC7Hph1KIIqKAF43Jj0RPWF2OYYa1DhEEWBGilELAg7O
giICWWFu+C3b7P5hnBf8wuABtudvh0NFm48XNX+HKZLjI5kmwBIn7yDWdzlbYII0
gYyrzyBncOfl4lMalC383dOu7pvBqQ4HQGAkj4vs3xVbp4lcbUJlJdCQ5ItkHT8I
lRZcmWVPIstEcSL0KCWOUJZQR70Df3m9QReLVlBlV6dNo0kP7SG4Ynk1vuhOr4QI
8vuWTJiLcfIjXWYXOeE4bf7xQW9S4rLoFh7OGNru/vkiVNRdVnkUxe8g+Hq/bIHF
NVdq49+fpVOJiN+ict80f1A6vp53VxVK8QJ+6Di3AvffbGsOmq3s9XPLQ1KWm6fr
Q+ex0MAhDoXxJeSBMgQqNk4TAC/an/MinLValk3M03ImvCPwkuSBTUmH9x7NENQG
XJ1zw+wVw/VOGXfCa2TKxFtPxp7Uzw8vhrYhZa/byEQ91CMvHbHvJAjU3jlOM+M4
Wu9hrqyI2RTi3SGSRKb3McMt8QF3hsMZFLIgjdqI1ttQ0g567i+kNtP2QGtS8M7O
i+RmBU89rt+gZ7kabE/RmR837BnkgTs2oKA4WcpBC6nrbwC7LH3P1zfmDcI0ckeQ
3YWTvohvyYBzG6EIoUJcM1HuhkWYy3ap+kmITnlTP3vZiRYluVIl/hjB1mSQftQp
HDax874w8YIMu/9q0N7PbPbRj3HF89uw2r/o0qDomxZHAGPP4bavewChgz32arX1
+H0k/76EAM2KT7EwIOwze74ue6JAs6ClwfAsIfRtUkxCAIZFAp5dR0SPqYl3Svqr
Mjz14tkdhrehw446dbTE1zYBQh+ccM2pg4x0elxxO9pIfh8N1Z2J+4yEH50i+OLU
LY9rxrzla66xte3Gqs7HrYNh+UGpqQoVUeuS4r1AV0V1TcaFpU8gmk0g4HKqWZnU
feWFf5JRilwb3rXr9SMbfRPm8Ydx9k6GDOr7U0bd42WUIKMWBBUWq2C5jBz3rqsf
8ESJ4t6jObGHIykNoEV3zyh4qaSGMGJwaZU1kgyTU4V9T8Dancl+iPH8+sHZ2SeA
fV6kMX+olrUFynZKuqz7yugeK8o8UJ1GkVko0CutSm82fgikO0oZCBv4brRbR0Kg
y/BxhPe2AqXFjQ7aBD7wwjNQu/tj8wUd1NpzByS0BRgGGpj85w0fXkSXIZYCwZrq
xf6bEf6KA1LKA/5W+MqlLADJDZ9xbB+hla8UUZlQ5zs4+yphgE5BeSwLZXqIz6oF
oIiOXnqjykzHD1GBb1NgpRLveM66sCsvmW53AlEsPIDDWJLpmL18bkRzBd0m79vp
0S0r0CaHH4fQsLGZ9ELZvjAXARs5/Gc8kR0Hsf+OMqTZz4DEKM+mtNkwBerF7Cbb
vXScmlgwFN3EhHjO61iThP9f2KtbxDqtrqIYX5eUKYepvMb1SUUUXbjjql3ezSTp
+C6U7dC6TEBTX186VwD/aWveMHwgdh1JVu7i9sDbVjRKLDaKOnfBBfUQHGq0zrMC
4JlwQYm4RW53O1bp4h98oCOsZrykeoP8Z2mWrKCodXtHR+cKGg861nt1U2NZAUlu
uWLdyygK9vj2QC6Bb3nzjt+a/xvr+bfFb9FGNXyaVPN9CSkBsZDiF2K+NTrvkR4d
iMMPrswxD3ye75IoZkySkm7TJ7WFMkxHEqQOZenX1dkLEYN0Ez5we02qZNGVwXp2
H5LsezdCsPg2Oa1ix2BTtedqM4fpoITx1NyfQGECJ5wXgwmByCgm2R526MZhMCxI
ad1MlSaN7wx+RNRabKsuH+paZEgI6Aj4udUWS61thk+BceMM08dbljP+36thkl6P
Jlf4CyU4QvDaVuPt7+eEmzJSia69eD+qsZu5NXUVAxXsgqeEL6O/h5QeaUhBzYBR
fuYCMIN/7WzMOLY03GOENyNchCJ450UVvgyXHYTDllkCjAkO7274q5JGvQTvC18w
9EImnVWYwDxcxpOghegtIdp2eanh9RVV5yJSVm8t0ESKyDSf1EraXWYR6uNFVHuH
ymF+O4gx15ryJ/c4yIKR+hJIpSJYtzur6O7s3jjlTEZlTnXGV5fcH1l3LOwh250+
vzIGfFcxzM4l3CQJyKgosnqjrCZhTcrZUM+sAx1BDfH+cQWP0IBRpJnI8ZC09XQI
+2e7p3x1eySsBCtvv6cJt0Gi37/4gr2N54JbEa164dp1lc7KFPnnMf1YINqrj35J
qFRXcQ6RrT1+1tjg0OopGH+53j2OBe7E9RUdMPKn0gWwt0vev6At0APXFnHDCg2R
7xeYHCieTPS/v/IVT0w5wnThtREVv9o8Vr2ZgDuPYnLaXX+R9Qq/gDgkaVgBMxtG
CCt64gzmyhDzuiJNNGYBPNr8jrH6R4FEr8PlKjh61VqjoXDP1fJqF801QGmALv0M
9i1jrw0TbPX9a7NIQ40uLDxlfX3nr2Q34IQPgBKoVRTsY3E6XjZiCbIZFYrhJPlv
5sJtZF/CfGH7ZccBz6hL4F6Q8WlS85z9eTslBQYR9ZYZJe5puRnXiefz1AMBxqNX
0v2GZSLSi76musL/qsn1rA/s+F5T5TFYZfMvUUvibKOnqk9qIZsyLi/L/Em/9QQi
1la3be9RVuKEXEhXitQzuHZ4YQUN2tNeNdkVqbnxFXUmFOfQvBwSEXHIdBFnjIOt
Vw/KFgIzr/1Oh47NfMGVGqeB+cEu4gbMRhRsAAoOO6P/st50/2AC8gVtgM9P+jPZ
nLZNsoFEWOg6a9MrToPyBlnkyJDeOxgvk779xOnwzqYuQZL/x09mF+utvYyTW00Z
lIQSpUFopf8BkrKBQfrV8Um8PCeG5u85lbxwVOvcgqt9lDijPHPLvuSR73VjoMD5
bDkgJ/IjWYFqCkcSYo2jxglwftgxY2OHrX7UDl2X47zxKsX9NPOFdw5XMdURcTu7
+ZRiUiOeBSfGuRz/jEq00IE0x8VmGKJQHnL3VOXNJnF12eU9/ba70VtMZ3EKUaYe
LTKslfOgBW2aN70uCGZvDEn1YTsIl7LI2WMR4rMgPqtwxiLjUcDlQsWIaLcKMmgQ
/3zyZfsXBhJErGu4I33ozICdpzeV6sjehchzSiaKmXxLqoDFNinzsQH+D9UtOgIx
cchDjtW86bDE1GIGj0AAtuHuefJY46GzCUXR6JHI1i7YxMuVydRYDu6PBZTjUBZp
gsv8C8iKADCZJANvqLAgM7kCHw6H2KQHBuqtdk8Sd5hJqQewNeltqYgplGc34vre
ArVrMo3l4JTpoJ8mzJqbjWRdEr2Y1zVUn6uCboOFxRJbDIBZEzYis50hxos7Mq8h
ugX2m8ooSNKfs+JOg7aJ+LSsy+j6s/ZXpcavzqKBCuagohdXiiFWJcPUgk38WACF
0uAfVtOwelxLZH9rBFNRDZGAERzOOq5aDScx0l8vR+sD9sBGHfFceqzz3EdKX+fT
/En5uDMNhy1WlZgA/iJP32hJWqQ7E7d5RfMnx8gXBGQ0UkgM0kNr/AOQpieiA+2E
LBtPfIOr948rwk61geASxf42UAPyK/3cvpBw1FxT1SWCE+14+tKXk1d/QlN/BxwA
D80UqK/jWNh4Ywiuttez6nRoky+tO7FWLttgzVwzD72i9pQhUu3+VYHV4ePmgYbf
JOx8MxriZniwzMcISCmE/ACKqYah/0o1IlovZ8PVWtKEevluMQboa6m5Cw7Yd6DV
0vdvQm1GC1DYKwKPPgFYz1C0pRHX4cDqan259dppqBOawhFk0MAy0Qsi8oL1Y1am
Qb/tTEmZhy6CGAOEfvWSHYZ49eyQ4/uKNLiJiLZW4wMrFryy5ru70d0PbRdvc3fd
GqDC1PSnV2UMRWsrLaADolGtLE9dt6v5AlUK1pf9NgJnJfLhsUcEs2uyoq7/f4aA
33XYydmFwNMf/0wnNmonUCAngAe3i0mk9AG/Ds/izC9tI3ps364t+YIaeCf/Gra1
dc6oSbbwZ55fLwI2OItZF7VEpaA+ZeKe0ompvDliNj3FJcWK8a9zlSH9SytanVFI
ioe3gzD1eDRDnJUfgPx121pkIMdjCuumvAGP49x7wujXeyozkyPNJyER+QGSP5YX
qzYgc3vswU7ivOI90m2SHDj3HGSWtoLRajPvuDSe5xmAEyvsnfZSqQLAOkkicUf3
5AXRCtcdRST5q6uasDEO10X79dwv2iP2cKlHdkJYgx3WZsW1ApRGJVC9qG32VQnw
2A6Q0x+82y9jntuFyRFWXOTxjpEsk5xrPwi04WHTBGt5F1XkzZobK1QwOsWBPavP
hch3C0N7OLPAb4nr5hpJQs/S/o+ETG48o9Uzq9ddRa6IcMoXS7fPonclOfthXk6Q
3yEuE+Xwjolinh6iEXfFFWrAVS9m/nD7p23uA+E/S79yY+XxUOxMl52f2NOiroBc
fGoFGTh3wLjlbnuZIUGGW6PxqeIAKoSsVq1wjseWjbj6IwoV4NAqsG23hnetmeAC
3WojMOMqeccWcaY9eqDZRFRcwy+vgTHilsYFtdYC1a2C4NcBWlT+vKnwCvzP5HmN
aWEQmt/p10uX6PpaE61nn9rKYGhHAqS2/C0OBX7VJ+91RfHwK0/lSfNHEkdjIzq2
aakkmM/xADvRxlp2jb9uI9rLXrD5jaK08bTXQTWKCIWUKnyswWxHBsSLsJwVPX7N
zpB/87lbfiHVc5Bv95WjVky+DfugeXTVNealIvBhpDuFhsRlYmw8adaoEb+lPLgp
W3509z2c+Hpj5uVGhZb6BTPpoIypNq0uTPgC52Y1I7eL16B6rUgOkb0L+UPcgly1
HtQyk+Eyj4hqK+MLUvkYQ6JNIqgPrPgdwE/5NnUjg2DwvfVFYQAaBX6qIgu/fMR3
PuEWH+Q0A+1LN+fl2SSFsh+SO1bUgFRcnGNwUdgDwh5NRLu4jx86rF5W9zP2Dial
AWyNtT7+72AJ4Cc3F7DvhVozCeM4unP2FsxMZBHj1Z0AJFgpl8vjfCIxO0dp6Nxd
TR3NppelCULRuz6npFX7w+5GtcEXHW7OWHu6vSmK7j83YF/9UH5ZKo+l58sgFNHP
MwbO7Md0d4BIOtpGVufF0488e59Xz51xHWyeR72LlCFo+0zmUs6+8oWYlpC+gOl2
7/+FES6SmBReVC4aEHTX9UnpXfcZagbL99I4+AogF1dT9qpawWpm4nylKs3Z7MaA
a/i/+yjqOPXD5FLO+vbzCaxOw+gScXllHRnkVSkyPRl1FxLKXVTVWna84xIEyRJx
FcInaogZu/9hRZEiVrALvV8xmttKufNbT5KCW0yl7kkUKyi82ijS9gxRISjmWv3f
cDx63tfEgorr3A0a95cUH74E4OXWb3L09GfPfOIHxniK7wefHkECu8rmCgwXFwE7
0BHe3Pw93CCRLHgNLJiL65sfrnR4m7REJBMQxc3muOWzXZF+kNvDXvNpCtcCRXsn
PlOKmG9fz7gBllVa+1nOeXSjE7zDiu9ENJOmLkKWzDDt9svc0tAROYJU3WTv+gES
6V3pEP6Max43M91czuNYnF05uIETU2j221oNI9I9uR8wpcdi8+DUdDrvXOXjweo5
9ryIxlO17wccQ3IagTJ1LAs37thCXKevKefaQF0Lp5Li2G0O6aJWtjITeq0zhK4q
v07jqFVVlSQaZFEH/eblVTT/3Sz1a4+q0jBWnhGN88uHu2L7LJacAMcTw28wbcA0
AEzaX/XdrNA9jltMa3ttHzgjGUWnWCN4QLS0wuYa5ZhKNDejLsLFp44HwHADmDjs
0Fk2pBcDaTjxnTOYxCLIb2bk3e6uBdNflHt0P6FzzXXZx2a62MoP19D51MXLAPc0
EEAtAfFXEk5WqszVkcogw/SZ9CQoRd68OREqWQ3kTlufe9IrwBMxrv1q6CecmYAT
o500A/mNYJPq63GFvPXEQdDGKrGsL3QVc9wwuAJ1gxJ+5MdaDrExVGNXlvBU2ABy
HaJhyBhuJL/ylidRKk+INbNYuV7XI00MwgKM2aXAKuAuqMwXssYQkPHmEP9DkATy
4z6Qg8Cjid1WwThtUAaEgJ8PB3qaRSNVV2nyYd4WU/hRdPJxj2pqZ59x3cai5TM+
b6c6UE3kNdOP3fn/XZNB65Xpp5tUMMIa3ahwdIBBnz/hCHak4vI9betESYbJ4JD/
0X/Zx14KPYiKV6mZ3jSvLGzmGFivBqu47Hb319iUzQIlSMngsoe5k2xQYNBLyVhg
N3G6Et/hvIArqxb6t7oAa0GfD2dXv6fTS87wHEIZ/bugCpPNjHPhgDq6KITNeG4j
6W92ZHz3cp8cvrmS5eDuLIhe4yWovoLiMlh+NRTt0LlnpS3uF+/7xpmgwWSKWxQk
TcdoozaHwlr7OvlCterdshkKENWz6KKY7Y5BVgOJBx6RouDgcGFLYYcECMf6/Ig1
Dt0WUbZCgL44+OqN2L5w01bgvPHOy8irWM0DrtTm5rUsIIv6LStxfSYNSDVDQgJM
0gt6KAv29o8lMg18YzbyQV9zbl5VmLurjnYbX1BhkKrKMu3GL2I09rXghe+w77Ic
rlWaKoEb2V4aHo94EbC5f7unr3DDkKr6qByltJX6jbqPopY5jlWWf5nMo6OGvUF5
CaPe3svpF+Q6kyxJxG7Newz/ZjQhFN0a2gQOcmWpZqE5ls9vgWk6Q0FpxKq8l2aQ
udm2y61hrcrRvS5aiDbN8qXFV6TEIfS2wTp27TKEQYp9ZAAqmF9q+wgwJ+FGsFbA
6yxyQHiOmwY7UtcBtP4BT/ARdFVnuh0Usw3o7Ms6PgdNLgWakW+inBl4oR1q+Gx+
RxUipDk3yazpitmH4VF2RxHAvlpiqkqoHiB/3CP7w1T+9lw1ihGCkOtyA2WYv7Qf
Lk/vb92DjBraO2tQgBazn/QXXmjPammwel0+NnICKXjUbegz14NOCqCS4v+9rcTh
Vt9GDNU56T8a0vXH6u13X6KMDAxpQO+xtzq3FhDjhSFMJrjATdv9v/90epoh1tgO
Ov1BM7Ey9H/Ll2OZQ+3um/1TR73TCju9zQH7acUXlWtw3/CcCiPAzF0ldTv4scaA
d7Y/dx6UzK0mCvyrZ8ScLRHSgq1HHLmNWr9vNDBA+PgZs/Ii5XntsLfoYt/Tl8mg
vc8Vvx7GlGHAeiHdvaWIqZqxt/KYDN+Ar665IbkHRcLHez3QfXPPHmH5asPMn/t1
JD0setK76r0+2jn1A4eAoYTFFrzkohWMKBo/47APgKQKPDiYxQGmuJgU1YQnbS1Y
SRoQfFeB0uHb/rBWSnjuzvq62D6TBAEIUuNdmYERU0LpIqGSpXAhl25W0W8GqXm1
lHfW8vaFrssv5ygn7bkuLW785apczset9YiqKTWQmhk2Re74gG46boUTcdQdnjIp
FS4zumiY2qDma4NGjYH6vVfdMlR9kcxn75k1UdH4B0mLnSGho449okSs7Jy+zjga
NEsuSCPtbMez+5T52/oZDApyiuBNPnNjgsDfcU3L8c+5SO0PibX6m8CfOyU43zvd
JBaH3uIfmMj81ZoRPXFz6/AKnye21LC99jmdD0dZDtDS3yZrOQKxkjjBBBrjlDna
DWf5AxyC2gEw0KIPRg9IqAD09j8iRj4LtKHoYSxc39cZ8nc+1N6ERIvYtbosvxFH
nQuoiFgtMLhZVGHvDZzhEVOR1Kgz6+fRpj+Yjgu8bxSgQDs9r3rRFNDXLgepoVv0
woykYbp8BRA7mVNVu8sSYpB31eysaKBqIVAjNyfD39jdxqqY7P0gOpMurLlc2caf
3xQNYB2J1OXGcDTHLY1ej0GayQHRBeSLfBypfhOz7FInd/mbeFh9RO47D65byGyA
eAS/K6xJ1PALeY0dbn7KbDyH3JiVUCVxqoAVlU2n2ABfjoHhPtzqtx93HTKtfQSX
7a7anmp1kOSPkov+G6bXypwxi+Bxh9LJXY+l8CAOxGqiHLnlujld0I4V7trP62SI
ek7s2jqRqt/eqP4du5p0yAm3Wq0my3XVQ/kUbpg87LE6eS5umX/f7butJZuurqgZ
uE3qYw4L4kpPec15ddN7l58TCADl78XZSVLeK04B1lpFzgPiojE4NOHJe91Fx4iY
kHyIRucAqd3UtAnBXlvqoatjx9mkAbZ86JT4iawsalvZThwA9gZAjtKkhG57pzAZ
BNoODvv2cz5S3f5Ox2mb8fPBx5HuGoKHnbaRcRs4QJhc2ihWhFMVnTUngJjLpi64
Cra6GiZPyPEs6cJvlvBiUedw1gw22hQkAv14tXz9FKHQYm3zKHiXMHAQybT+fEGt
LQrTkSw9Dg4OqtYRUhI6iQOaTGz7zs3+surrRFlIxBYxRi/1Ugna5c+yGsxXKBrm
kELGdq5N3YoIuY9KrKHOuMbfdIWYOTIxWbmZtls/XCVwyylaROe4LScExIP043eJ
o1oj1J5PV5RzICrOXjbyIKEsHD/KbUcB3l2NDFrv9lVSbSBFA2qfgoA1v5OA5Crm
e4mjslGg82k6iS9pcn2b2j7XdXkV2iHRDdPfhExQiEwxBHC8iHdeRix/GWWwVmzL
m4XrvAiAVS9cE2QtIn3a4VxSPZ5SODW/C/NhgR1FH1s+qOg7Nue5rrZ31AfZJ2Yq
1/eVZ5UQwzFSi2Hr9L152JB0PhUA9jHtoQnHPQXsj2BZCzvBQFwMxKhmOESua1yp
Jn+DWzsfnlzXKlG4z+cpMwK05DOvI2La0vAw2q4S+rOVC5k+JxmvPHx20mudZyXR
/P+taXykraQEV1J1p513TJeEiL9mQuUuuxZieMQfjSKx2wgn9mmCObH6emWF8XlD
vPOUaMrV6l+zpTfgetcQp7Ne1TO2aOBAw+hix78aX6fR1vhvV3xJK9gPiJqoo6wR
PfEsmvyXojR4ansG865iwAX7OkILlb2az/tLPaMwIt+RsiK/3R9NH4f7qBcsSQVd
ZWL10tlNaf/sgs9t7wuvzidw6a6lo3uGoyWtBh63Wf/CfMvNC+oSh0PDf+RzfyEL
b4vysjPozdP01Ko1bYUaKGBO7+90WBWRqIl6r/bsLbOP39NNZYEOx7TbkucfNYat
VJFMoKgyk5OSM5lu+NOV7F7THmSu5pN9Sa2O/usGMNjXiF4OSFNPwEfB8L6CHlVg
nyJ6ew5RBm7lmAPTRZ3XeGtZ1Avia8pja/HZ+euwEvV0UucLBN5fZLZ6/RPJFU3C
jqUq++2EbF5NeIUjCKLVOcVl0PQSfSCIfec9AbPle1UjBUPgfIRw7iQ72J8Aeuyi
BbeB7/F60AX9yBcNkOV8aJUGuR1lvGVv/SOCZ74vSTU9M4zkcTcwjY+D0nlyqw/g
+I7n8hpyyOrlzu20vPCTsQgGWTHvpcDPjtzHUjffgn2OhEpr6izwJqjJfpYdhRl3
b5A9CPnAHVgIlvIrvsG9A0hi/AuI3vsvFK1lkY9WHxDNsZOd2iGtvd7LKFSMpitF
WAfGjpt5GLKd8DVwUecpp1qSWF67X2NjgRzUw5qKysK+fnG9VqrTNJXxNiiU51uB
sni+LSp+NiUZTLzLFpm27125bZCC0yr/35ORoLU/6P5UEvlHIDiZ//9gAtqWISZ9
FWIOgqaqaDNFnLZ30nloI+EXeLBqkRZaT9A0KDOPYrE3JrCCe8kP5b8TPxrvff5N
2QYIZsVfb23rGpqVYViOnOZ+lBOpdmExavR0fc0D9VIgE9CUZmO0z2oY19xZyKpC
B1DrWTCVTsaFtKwTpqH0zX7aLcmYEbsr6oPflNvUL4it5czyV2Jqnbj73toZ3SEM
agz/uT5amMoU2IMxisnCKa2UfvsySTkup5xNCjrCD5B2IoujaXqY4SjqawYlpf87
/BdQc9btGTsiXtk1i/8lIQN+ASFrrGKUjJtZ58aHJwtBmz1CgkBV7LwsiNNS8ymm
NSyie/BE7or7n9ndTw0vqAZfufGA1DmVi9upq6yBQ8jQciobiHl22R67No3ZVYFv
oWfsrdQl2uBot41c+N+2pS65iIe8hM8NyP+V7P0uz775wosXl4SZtT0cGgSRvrD3
yhalSR54mQm1MvtHjzhuuTq8VKo7Vam2l2igqM4W4038CloAV1/ItybFhdzQg+ff
q1TOiuMx6nzYhy3vSjBUAWg+EMcdhi0XGn7mj6FIncxElmQ1KUHc72ju020efLU1
CRwjd3VezlMdwf/cDviH1XuupEGCuuIFOt3H5cTvUKx4bc4NFfoHEfR1RN8/Tkf3
VaK5INew5hJR9DjFjI21dmrBEMJPcxTA0636Mi+oSFHkWMwu4WroJ9nfyq/dvQmm
8kQgdzf5U0ia0VZj9t45zF1+sOj9gAj9tJ0/XLVqXCw9+k4OrffAd5GpaNUiQSB4
LeQwjg9CnCMfl1G+wKpufFAeFDptqduMyVAJEfW1O10OhnL3E2EfVmXGMDI6mVEF
hMkhu+tYkF4aMPg/p+EMc+aDJ0Ss+CNvD8m2OfJs4Kht/O300/AP17LnMeH4RzkB
dHR3Qh9+WHhzE3m5SGxxIn4o/FN+2zKRyoE3nEo7vNq5jBvUGmOU8l202w5jDMK/
/cot6VoKxGZ9vKvVqmXtuODftybFH/BAWn0+A7MWbBs029PxfyRww02oQF3Hx7mZ
uczkAPX1dFMvPzFQ1cmCFsMYbm7P/WKdXt73CT1y2GzSTUcXDHwS7XWtDktztAFd
0pXHYgx6jX3RTymZvVjVu/DoGbhZMtycT68QGoXh5eCrUg0oj4nWahD+uEhS7zVA
wu10cp2PqtR8mn9GoOceiwufozoLU7Er+GOBA5F6Q6l/EVqpi5zVR1vlzhHwpQc1
9te2pJg6Z5S8fJ3X3rtefMyE2EOJrY8pRzUw6q6lWTPmiTDYyenKDl0UQE8aQ7/7
q7ati7Gd/pdGxOmvB+vfhWHSnZSJZZKaObfRJ+6wMky1x6UcKTiXtI0eYLz4+n/m
hIfg0GHjPX/BazGuEI2I4W7sEiDFykcnMkVu0avGNA0H8xs+N6dOfDdZjTF4WhKW
AakVOFVIDSpiLnroYUzgjRLFDKTKDRVoSPY3L1uzpqRczwPGQJzEjzFqicEqcsFk
PAE4ujzwC1ysPZA7SXZTVZLbqx3cWjhxZRSbTactShk0/GpiijevtXa8y786WHt7
R8SxDi50d0RKEaY+vnPcpHAiL7tAYaRHD6feG0C28azurM+/jjgEBj9Xws+7u0NB
Wd0wvtXIogGksbeJu2ZXX1B8CYwUyrfA8aJf8pLjU+5lHapJiZyLd6kz5kj0/3ct
9i6JuqPhNLVMEEKxqbwwXDaL7m4pGY02rMCb5/tiLa4MaD5W+Xnrf1BGuffDD/it
+HmC7Nf6bfYMADMPA8vibAP/acql6Nf+8Ik2O+6+2Ry+2xLM3tLeUVK7TjJd3HEY
tmGnK/mUz1y3omvUC+kztYmNJCsotmzXHTVv9zD+rXhpTrcd9q70YCjK3ru4rsj+
r7oky26Q4Eicr5MR8HeJpXMkCwYsbswApLg4yzgmrWBF2D3pnJE1053CzF3QS4CC
tIXy6LwzgseqnlM3Qz4+8V5GWQk195qXzZu8K47dWtpfBJcc57wxic7Tbc0SiYQo
Lj+Ed1VAfjHdFH5dWjXeZnDbiSppTGVpPV0v36xAvFBLEkMWsIIP7BKNLDzAK3+h
53LM8ffGpLCIIg0/IWbDJtHTtbQ4w4lmXKanzerMtgwNu3Xa1KJP4ina0IoCV2bl
L7PYencUrn3XyGYxI6Ly30FpQ4HxdKNOemVsr518Dju3RUSRiTmgmf9rc6pFjR+b
6TGjOf6wMhMDdM9QT7demrDDCeOr+AVxhr3V2D4zLVdmLIcmIw9zO1JqtJAe/Hpa
ERohYHEF8Q5jQyeyXWw7D8yiAzVp9Jh4HUjyJOH8jyNH+UAX33bTsuTgLHew+Rda
wwRxkEQNUSlNWtVPYnhPsLI+9IY8BpW+KDpOiMi4Bc8AV3L+Cp0eSregsH79Uxqs
fGx5LNBdh78rzcRyWyU9yz2F1YqXhQ65PIfJRs1+pNk7ClZaYkTOOr4/6DtV7MS9
loUVLU8UloM+9pAv3OvgGQhZKYf2pPmZI+8qnwc69Wm+oage49inkcop1oApyud0
rlqnLNbkSxi0cmNofZ/nioDb2J+fZotoRphohk4UZkwbzA5a/0bsrpnmmsz89K6S
IXDMB2DQmUlJlkbNTbkU5StBu+RdMqJqS9mhkuk5tkKtx17rCHnmrdCNpusOy25W
OeBoMWVqNZX89ZpCI0NTCuBCYS/4c0uQkviMGjMScAbuGafP61llyV5KevzaEBfi
hfrh4KrxyZf9skJhL51qisOCHytweZrKfeGzBLviUDBomvImYPuSL5sg8Ml3tTh8
HYMGyGuZIuEciI3BVMhW2i9rTtfu5j5DN4CduMrVTgOSnnUJ2faWTAB4or0a9VUm
xYUEp164+AyihXbQ00bm0kSuvaflC3fh1i3hDHs4oWX7ImHgZfEv46rCDDK658AO
/0Pgftv7a/4q7t2vxPSnxUmT1LiY8eadNRI+nkpYDRIBiZGemDnCD8UZeqJA5I5T
OWjtapSpqsZzMRTLUcFx7CO3lU3kNEothI43htqUC+Kt2OvfkQRksRvzMK5urfH3
e34YD+mN6XWKE/GoHu+1cY1hRYh/+5noBFgGXnVasL768yhkQGdW9eE0/fO4t0Km
DhhTiJ8mFjH5NUYB5fTKyltfbaQzmKID9kKwnyLg9UipwzyioZnU2owWhYKVfuXU
T19+Fbm2Jsgvla6XR5Bmxk95+j0CMkU2HaRrYJ3rWYe6xcngjjpidr4jUEw2PzIP
XgFCZn6iMM5hJ59p+4htAe96SFi2eQCcNmLxtvKtEXM=
`pragma protect end_protected
