// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:32:40 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
FX7BVUqxzMDEhWW2IpiBBA2QF10ryF1MXyibYCFEhRvxCZhN0qw3UnSrGK1vHEXZ
1yLpc4iNAytsBtzXw2m8GDDLLsJr+TjDcqSS73l247SyYpVMu40yBtmxcSbpNC6b
ijCTGs51oU9P7+JNhgMDF99pn48L6//zaIeKQ9Yimpw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7696)
/R8dlqOxLIwqmVYDMGZurTHpyBovPHYl6Z3FPSTzs9ExvmGjSugGUVreom5havcv
16q2qfFtJsekoHtrztEfHRvRaQjrtKjgWUWhSXrtgOJnhjAWM4GYevVWc/EZvGBY
m9PiMj7k0DdyF2moYQJyMeDOAE0QKvPK94F47++8LnqBeTgb/WekYKiZJRTJ/xSU
pvtKX7VXtWB3WBh7Mdnxl9PPELbsKcgst3wrgtSjHB14kFx3A4anE4ggL9TUqzUq
oSKgOAglM+4lZQotdGuWsL+RK4z2LQuQLM0nDW/jDxCf4vPPR7ntifWu5uf29bak
VfinG21nY2TrZgLMoX3eRQBaqemKIP+jeV2p1zrS39lTR43ADmeifzfD8Jc8R1LP
O9YLq5iOfA/5WEGO61AzFBbN96LrMYbqNmetAM2gOovVJzSU4/6/EGohqUFOi+Ga
xpUW+V/n+o6OECxX+qvkM1xy4AgMui8vFO7ZtG+S8iWhxHIJT9ZtUu9LNWoxAS2X
VWct/lK+GLae8zW0DtmsGwSh+88YxBWVQ6jS3Wa+L7l1yElKkCapErD7xVPYhAr/
Ezi46pXuxXNaAR5JHr0PM9sZe02/peHirY/8Nq5VmQ207j4KSpSmtKBQGSeXsME+
JqseBfsN8kv9iSwkIpPyVIVZMImpD492BnkXtBvIZ/7CQbwrRELCFFeYljmSniVK
T43zXweoLmGq2Ye2ooihsYZpUztrol1BLDJDUEkSHt2u1wWULglczklpt7mAG5OW
xP/hWeJtWX+9/fCU0dxSXwHDg5SNJo3tI6ISvpqcYY1acyTo6I2tihzTxJ/C3J92
HOYDOeq4NB5pAguQJAr1ogOQp9d6EAGHvERgSmYDx1ZraFI9DdWj9jLiLEpoDekr
NsSUG+rRCC4Y/olOpPD82D3rct2O0gCap1xPgnCbmZRhZ/jTPzaM6DZ3mRdW53fV
mkQE1CjGSyzMJFxs2SGR7bkUWaT04j479+X/A85IX2Fbqgc6Lyv7RBO5qT1wa4O3
pV+J55rBk9WntOt67yEYVJgEWnvY9Nwrf/T2VwYKragjU5gl4KaUJn3sV3FJKqdO
4CamVURFf94F7txCgXdq7T1SdEwWPSnkkvPovBLAzhPr0o1yh0oBP3PZwbN9cPHk
v8lY+iuh2/dt7EmRPQTFf54jeMmailhwmC5ZmnFOkXDhD5oSczCpM9YMqoAeVswI
4xD5V2ClJzyI9l6jRMX1Zd7zOjZI26Ynztfpopv8h1doDXYrORnX/rKTuNdJFbdm
9MTSx555+ePuXoXyDVsDrCFfEfJufvTivdFJWxJlBv9NTEZflQUbi8cJeHExjwdO
27x2Uh9aCCJiaDYNRZUt4uTx5JKLgqmtdLOS0AjpHyYcCxQAxpn2VoCeb47lUKFq
VQqxAPogMOffQ2eUZ+zaHG8tOkjgkWmYNyv2e272Wa+jYIgX/wGzA+xpR+aoRyXq
G/1tkAqmowR0Cf/6mNarBelSewuAeyDihleY/OxNaR8TS1cDWIaQ1buGjbpYU5d6
0QqJIgg6AHrOBNJMXJTbV9bHZ7fRAshEROpDYpiPaKQw91xm6uMmFungYbKykPbU
n/b1cJ5B0Y/VKnALlKXE8xBtXOWRbyv3NtJOrlV2vNPt0o1SkUKYhzvJmcDDunNI
GPu/yhC/HgLmEDsmvqaAEssGiIMHa8dT+vBvuoDUV3qZZe1imPHBvmO8VXjWFlUc
GMJVKy88nFIgwvtntgLFAPcisXUALPhg7py1BDVIyCbhhHRnhCO8gcUulUizTvgM
m7kbgzW7uyqOvVXxXR6sVzBmINgYzN715M6DyKeNm1iNHt5EdEoHqj3XulzfJyTj
t2NegwTVBtgyu9DHA1cX6h6QxY9IewNG1jT8QL+ZSgnMFOh3vuucOTyDALvgFY6G
7l54F5h+pMDZPr96eJ+N0iWFEd1osB6pJsblsYlzQ8yJzhq/dxqjxNQ+h7TuKCE7
jVdr8JJ9wendmCOtosj6d7Xux+Jcc3PRUORAJaYtwBb0HizhNfq4HtylwEYm/I51
GWxR7WiiIQuliFiKN2j1s2jJJKhpC4k7EImAgMgyj/vfRvpHLatDuSSzRgpm3C/K
Hl1h4T+ghJpkBwMXhjfxIEgG3PrrFKv+L5x2uLOFw/Z1wEsrRzJuJFuMCrwUDmn4
BS9EOqwXubZ2B7ovKODE/cJXnNjFu455TmJHaI1yr7wtyI7YlMZlESPHIZLLHykJ
Ra2qIx3BQBtMUKGlLLYpmW8QWjfGq3hpdVLzuimSWCeMuKB3xWuZ5uBM+h/3rm2N
mjdAa6HQwJpOd/cWAM1PhbGqUX8V2zFuxgMrxNp80A1fhlwZzXzH6lOroJZwkX04
ZfzsJnVr9VnOPFRuMFo6yX8Q/LM4TqhZ1Pe1NTMB25FGbYnJUtLDcavxe0/Ym9HN
p6kfJQrDHd8hb6ereSxx0D3LxEstCcOxS252P0i+0b4BG+6umHyFKodCVdHqWsDz
yVzQnqiRzs9pJ8kjHqKKk8vYIXEHwJ+AHa7y0QKlpXhqMF3imB8U2xWh5BvdEv+j
VSv99ey9RQuqJWMYnjODKLeWYTFaKD13rfNoiseisfhIKqBrW13pQ/g2TAgU7FhE
N7D8pmgC+xZYwN0RbJALI6Mz1AjM11GBtQS/sVeJT46/kY4Gd482O7api1DbfS8g
dtw4En7PyRcQm9/TUFbVJwytzMwYW3Le2wwMDhiIv6DsxRuUPq2NAFvAhXngm8oq
XGrIcILG7iIrX4Bta8+vL41rjtPdepWcb4DhMkyWqNIERYHWeeecSCxdNTuAo+aj
fK2LrqLOoidlvCrTaGeCeJDbi7eiDtf7DaNpEmrgPFosqIyLdbihzPR/tzDqvl13
3b9Zex5FHb3BxLnQTdjT6RFJEXF84nyYG53koBa7UN0oBAIVsnv6JkdFO6aUK49I
pYy3NeXc315Qy94O4WIDuXNq18bSGEttlGTADp/1Of4sGRj9zzjglVuSWceEXDxX
/BIpIPQ24DKquvyqP3l3VXOLxxNo6reE9I/V9yIdNzuxwdud1nUPX40dWsSebfCf
e4UqWBsCRMX5+Eg+OTm4MTijQAVQp3QMKjKpEpQgtxRaZcdb+HMLLcH91PBWuIig
8N6rmBu1AgpTXp6BThHmSZp7pS+o9B2YXYqNXZVKqTqPWlI7bNoR9Z2wTBh+N4pU
MDs3r2mnUOSTmyRqytYe5y2hijy5ONttkADvM2xeKh2QVPWG01B/e4PcNqXAIACJ
J3Rjhw3YXdk2plUPq9UbrXe2RFiUQNE92U50QgZRtqSnLIjyaf7+6iD6tJfWOSMC
dVMJWjbs2YNHiiMP2lGd57f5CrwF3J1y4OfY7R54JcihDRR2cke5DTl67mjota1T
ZuYhNqicxNUJeO7pip8psfw8CRGKlgnAAhJHoMUL3J69tO7EkUoIA1iXU7baOMGV
Lnkftd5Dp/UZcYOsIPgtL2hOUt6JF8DcU0rjo67SWHoGIyF2bANTwMoeekDGIBvj
0uAqGoo9Oy8WWzNygPTGHoPiZKO/6es6pDw2yrasy7w6DG1w0nc0NvB3Xlm1N2rB
QWlLrUANOHo286Xg1vI5Shl1Sbzx3frJuuWTMQiMaS+tHC0aca0H7CbeL3MTtKrU
smNiP/b7ROzA1r5FvAeHsIE9J658/aa+rUpqJ8urdCZa5cUCeM7SFWtYJwCxGnpn
TzsesBS0NO9EGxNT73/piLLCSOGt4aEGLKrwv1znxIaA6wPLArCidzuTQ68i+8cZ
9p7360HG4gZ7z38qX3jTH/xbP7LwymWXs9IGerqGNjH2W2NjWti6JIQLoOX3U9SI
tLJTFicneqHRTRmJftQaQ+FNtIFfFjFp01V8srzx6Ew4NVHNyzsUcgxzBYJOH2mJ
RQ+YcCU0leW0oeI83V8W67JeUl16Un4vfzaZHQXGh3uJwJb7bA5sDonHFqtC0wcC
ZsisWltLToWr1bX7QiLyMFJPO70o2YQZc60Y3f95ISCwi61TfSmiWKi1e8zVA/AE
ibaciUUd8lT55Boj26JF7fYW9gcKvMMrtXip8JEGJaMJZ3khGCqC97ibUbSbRmwR
B37cmaujAos6YA/bHgWYoYDAtCx7IjBrFd5MveMKxSFsk4nLHqjL+bOywfEsIkrb
rWed4LQuZggnGyHnLA51BcX14r/kL42/kNVrFrO2atIJlp5WbsHNHYTwVQa6BHnA
PRovITwdDtYL0Ggl8uEInj7gy6GuayB9gpgr9Cx7Ht+6KP/EAS4r9jgn3Q9HiNxL
RXX6MnApDRajtx1sZesBDYuhYQ+9S4TOZptDsP/HKt3+EPeEWTuObjQfqE0zVUbt
leoynPSB6FNM2K65sflVgrwGmRXpgXpvMToj3aXtyBpo7YN8RlRp3OzCwPPCIPzT
1LlYZnrhVmEuZl10TsfalKZ0sedwEg5xj56rx9zUZ6eXSFfopBcf6SL22KBKjA4C
gs374obnLR2x4QlWPNoNf6uij+LyuDGgmK3frfCNdyQQHi12ypMUNUOuwrqcu026
woK9u1w63EAy6zZWBYxd2cEXEbSqVLvRMoeVVnT464/gXYZyFQw+J3o/iwO8woAd
BrwKltPAyYG6IYj/BTna8PW6TnMTwhmXpUWy6ISQLB8f6CPGf42Xz2Uvj+jB9Ndn
YKfPIIHpSbEfbUkrWWpwmYKPvn5MYmvDfkaCAqJpyHob99gW9vwDtWe5jAQ241II
GReBCSdixIcnqZ9EjYLAT+n9UAJKtlcAcrrwOMf908egmdT2kTBDsMQSJzgjHLSp
jwSd8pgmJPxLe9x4+GjeL25nnBu32VJP2rHn/kZBWTdFwcvJQYSKkmXynLn34cc0
oIrA9eKdgV1ygoMeXJK+kuKwRqcSMFPFl6kqZLQU5E7FZb9zy1TWFJoRGQuums0V
PBMhp+Qk1tkbhw92UVTywhfGMuWOjG06ERyHaVUS0wehM9z0PECssr1afmCf9Ju2
C9Mc09oscwIvVU2rHl313OcKrUJ5NW6tlixTy4DMURdgTrIS0rFlgYMvsr5xoxoF
cDz0fD1wjEsjsQ35hlLi1w30g4oqdl/QlYk3IJdvrhjNhssxNOSMe/9Rb7hCRwSX
8LWE9T3GNhIuDq4Z7Zn0LgcGEjd447pP8D/by62jGCFDy2o1MM/VaoBW7mpavmwH
999VO69DhMJgAXf5ABHg0yAICukbwXBqWEgFgRnxJPr0Cqrx9kEOl11X7qqVgYkf
gTQ+DqhmDyXr218aI3skUNpSuE19QlOfppJi7Y38Krj5ORCrtf9Qce8LvMtWgsW6
0Oq54RGT3qKnM9Dxw4eSrJlCB4OrhrnfKAgxDWfNtq4AKg04pOcw5CZAIAlEXJem
RKW1dYQCog4AeeMAzYcKsUldpNuFOnzwCCg4GegQwiYibrALRWJqpTs6KqR+ddV6
ZrAse+lnF7hBoB/HkabQcvmJxKIqE7zWdwB1hFbjmN1Bs7ESMS/3XZKpSVgd/wP1
DT1Qus5zPdq5YxgLiJ2eiZ9sBJCFhLPko4slSoCU85iE/wHw2OEqaBTSHwpas/th
7cIv7j/zwiBfVpL+kballcOqwI4Yb0bYwY9kPIhM7zqb9oOQh198vNu20Cwn/vkQ
zjjZWr9ie2ZKY4WR0snvXxoyoYJ7gBHQ92dOLtivPbsMlbPQZfVp4xOHmluXEXhT
39dy4GN1Ce+267T2P8hCmI1NmX2km4uuGkcVL1c5Gx+ftGYFSgIWL3Nf65M1bbjw
mojzTbeC6XNFkA6pinhzUnisXz26x3pzTjMOKa9YK5U/KCJRyWbeeTXliwMtCvgG
aPs00DBuFSVrpMCqohmYPq8BjO7q0MDW280Ynpdaetl3zCP4ScZdBsj4ai6im5dX
9336IQ7CcIvH2dq/6vuRNBKkm6AVi5tQkxmGASTVrfEkI/fUCEIrsSBUWOuUQHRX
q8wbbRSvhAYch6wDMe0EJWXlghgbkBiauYvRhXWW24m4uM414/nlIR5Re+SIAAUE
UpxJv4M056jBUxcg+plwa0dCyDVMj2UYm2/9oOwJ+ioSSm6GT10YYrOggH4mAnvd
AQjwDzs8aYY35zbU2WdGl7U5Li2UpFaUbZ2HfzkLHRHeIl8hqSS1UbII6C/5p5KT
X1+uXkSazcmzFK1MkpREQmC7q3Hl6c2BRD7LoI3Wd3tg87nR9MUZBopTvWKMNKF1
8ssMI/y9mY2kiAaL1o/jzEnIr0m0InS06y4+r9kXdhlNHwE2xYnA1/DhYcDqU0Xq
ZLycCShzX2ZSYX8v/YjSE8s26391PD5cAPLryejARm59kN9yFqlxv9Xt2nWSJNnN
zNSE+6p4WrHA/BR7Xfqalv5jk1koZqKZaaYjTYbTmqkNjnRpWN2wBgInZIjoklzb
MiujqAcWuo7o60MyZE2m+IfeEXCv7w9hdeW7AEXW9PUPS4qaUTL4bOM4QTlg3D5r
FaaUEcHtz9x6gpAp5eaPIofytoWxEQ32Msvdcg9nIyB3GgHCVB7CqW/2LeJX100Q
rpCFUBSn2bEICFkYW61SaK4zVjIUFVF2umS17KbrrbjaMHVrR+Pq6IOBVLtoWLFA
+uMildU/UfmVKocX+18HgAcoRiVZEXBplErRvxkHLo/Lw+lxNGU6SasxapyhWf3A
EqrJCeVbdlO//7Jnrwg2K92/UuxV/ORz3NTmc2gK1Xw9gM/MkFzMDoNGUkMtUgpB
oKHvLkpwsc0guCGlYXVHZ/2TZyTkVng6FdKYiBBx/vFcneocq6R926JugUS82UtW
umj25bKp77xW0SBr/FCepX/We4ZqZzSJZfpKMY3yRts/wy/+S9z/1QYseUZGZerl
r3BvsYhGhjc55r9BHp08IqZmN6wME8ITtj+0+4YHF5Wr91ulrN+HqkHbCdk6VBLy
FRunIm3ANUEhcKHz2V4vD+fJx+EUzjWBh+CwqOkvsXeEVaIRSnCwtsuJcsJzzbiR
oPdlxmx0JEpoy6KYfULuhWNx2nRK5MQXxw6iSjphNexkqf9SKc9hVPsjG5qHym+L
BPn/ObWhQjD0PAydhzgVO16yZuifcptUiUtJOMvVRoUjQ4LG5MYmxQFAer98jXEr
RMCUkU8Ure/Vap2Ir2AqTFQ7cNbRRLYsoY8vILvZ02FpoyaOqiil3FUrMl6r3gbr
KMtsiGyByYRX36zq5vT8nttggvXV83pHq+YDSjb3QBZhq2lETgkwjuL2ewqV7v7F
pzmSaILOIA8U54OBiM9k4rQjzp2ENQeruMJE9aHuGNGtjDWMvxHYKqnTT2sh+SPs
tI/xTbIARpddhmcfX3Fdkrq0X69M+TU7vrR9B3dhloX9zS4fgWNKtU2+fCqyTR6O
fsemecvUkjiUCluNmPcP+Ah8+HGGMOUSxEPX0LjZcqrmtZggFrEcTFoHW9fiyk6L
E+rMeB7vsjZnqX3v6E0Cv0oQIFxqOnfrDlBZ3tlEdGTOUmweTbKEQEIDJSWH7fKu
B7vvtKaL+a8OWVfazCg9JA7dO9AtnxJeEidkosN4qU+dMWHE/UJMYC6oFTTqSguW
+LrGfGzslzfcBwNAnoCI7ufJsNdN0tFjwXL2jdh5HqYTFSSqcymA07qQR8JOblMM
xfO24hJwH7UWTQPZR1Qo8O6/0iExkAMCHPBR2WsrCf3iTT7Ac7ND/5S6cUUmJ1jr
BuM1fgji0YItaHNFUjxuGKKOnKqINParZDqxdFDLi2YhsfF8nRORAns765c85n2c
/l7vKgLhgJnR3rv+wTVNcHFVT6nIj1wMI/egUUoCaRTwZuXIMR6Rgmm0bml0nNCd
UhuXH3j8+d7+YDOa6lIPU6F63zOG3P9w096dN13aL0wl9hddIJwNKXpA7YKnoXu/
qR5yD+1SVJotomnhS2CHVFP95XebqUqhx7uiPVMVbnYm+Bl4isOt/nDX2Q2jh3lp
0wPt9KlN28t6thnSdY8K5+4vtmY47zXhHVzsN5FDeI9wHJ1EO8N0Lh92QAguOHg7
9hRjXNTwdV38boxoiFXUlWuejZj3hGvwpQaR2++0Wl8K8gqE3meAPZc0F0VDVTFQ
B/h5zUGcTvx+NEKB9+zB2iufTevMXesQsSxVSIinHtuV7f0qgqMnf0a1PDajTU6v
gwdvbLps6/2KiP+YEYuLPyy4dJP/uWtaWIQELOhi3hQm/7bhW96viVU8Ec9DBaTL
1ZFVdx/lLZPm6pgjZPjpQywNNJxgzBY0p3b/+b3pIhorCqWnfnUHEZorQ8WI0IbW
Xdb5DdkeRImyNjrQMpCmsgduqau4tjv514IXahN/2hAsG+wQVSP00fams6Ey3CpY
gmmFpkXshtDgBeac1CT677/AReTydI3W5wZGD2lo3lVxuUVZX9qV5kHpG+3FjOYW
HuFDxTjuCwOgs19pTLeoRha0rGWaFSxNrYZS/e4e8uinygnMD98TnGr65E8CLUkw
2ZSyfB+MMIZ/KpOHMpLgczw2wLqTdJbgyWw4zzOHx5DLe4dxPehjsuymodHCjEno
CorcOokADqmWJtZzLQ1/nM49CunrTPf40Mh2uF4iKqsIy+x+Mu/whI+J9GudKsQI
78iZEbKzVTzoqLNaNoV92W0QkPbjqZ7ulxyy/iFRjv7ivb2nXiCSWLHd14Q6fnAd
gkA45SdUXMPWEBmfgRwiJuwDYkR9gF/BQaT+ll4pyCQER/2AuHg3LizH9kqNFJ/9
2QTW97A7pwih1CHUzmSeeQYILFTQbNPtCryfaimsFFPiKzM4Q3Guc5hTlcfVgvmM
ni/jPJt8HxSg5Elm6otuwMNR97+97g+hCLKTY/3m2dOS0U7tEDexJdwcpyyxeWQo
76McZp9eB9Hf7/JPtVumrEhMpyCzHWFkOPcntP0u6dm+8e4GNJlqWnjoI5LJN+KG
h61TkIZ/6+onblIhFlH4pNS+JBism7hnijM6v2b1e0MO3wEqlMMtFyNQxdNXjQtQ
hJNqw9vXSBc6rlsbXDSw81OzxjeANpo1a8jS4sTbHUOQLPStu+WMcgpuPyFeGkeh
KQnbC/KQDt1kMLkUokILKWdxv1TZ3tgRNKfkqwvdPhtI9lZjtW/o+uSCFpe7XLBU
z+hxQccwNIcs4om/gsPwqhXv25jahxgTqMNNgS8NTg6w7RvYTubhyfPQ7Qdww6lx
EkjhrJCXND/p0E6sQo+DWgkRA9CFSk4eRBSXVyuaYbEWMm5jttbaWiwVArpLD1Z5
5GoL4yNkQTKW/ObJ2JqBd9j6B2wiaMbz8xy+S85iE6kpXZinCZyOMvCIpSR8jgMk
nmSIMHSl2QCGsPKF1yPdkOxRXxefk7QWu8EJRNBeHzSdHxhpYbNOUX9Yz9VCOIYU
Ig05wyVF/g+FW4Px1UOs2824imZUFefeNgyrG1RKtfb3s2IfHTfqn84j0m38VR9z
E6fnm/GPkYn9zIafU7TQSskL7y3nbDsw9FXGdJk2S2eGYd4bJ3zQ7WyXDX8f3CvV
0G4qcLycyaYN0rn16VXUaPDOydUTR16HLTCpTzdzRtGCJXq7k3cc9nHzkAWHZ+Qy
bUQgu9CZJ5SELLzbs6iAh22+TFJMy7ixcEuDeyMoFweagKpWnAn7WN3jRvEI+lG9
zWFNqhf5s+proTvj/RZumEK5tI7ShfNfOa0bvuMqa/mSrdgkbm+i576TW3IzHaqC
U4qORUn4cylXGnyzrbhWhEDQsIu4nSz+1Ci9TbXxngbUJra+PdcaH0EXi05dUQn+
2OcUN0TtzSsl2qDMY4BDgBcffMxLFHydSxNoJcEwbrTzo4tTKVTB1pX566BnWmTs
qwNpYvixYmxIFoJRd0C2V7CMnlKnOvMPrBz+46RIpUHYmz+MO4zehFabyEhkK8D2
+XfdEMAQYdC6Z3xEQAoQhjXvxoHJC467OIdLHIy+63ewPUKSRCFPSfsKcAtk+Exa
00KVpUxA3+5BC/TF6Tr+OfWWzpaU9uckRFzZCwWNPs7mOKfZVc00iM2PTxPB9AGQ
wWz2zkq/wJ5SAWC6Hm8uCaIkiJqJFYzdDGIjUzG9lmc5y2lt2MZnMbozS5k5Cgqx
Vaq2YBjNVi1I7hYjXXuQIDZy4vmea7vCaFZyF0AhRhCopVOIRKBYdM0awc7Z0NS4
H6c5IXnaeLrcssigBhKNxbW6fEMa7sIcayjyOBddjGK1HT/RKhSg3FkbuwvqS6TM
kgCK6vxMMQCKfn9Z00DobnfqFyGooGT2UKhZZ3ljEO7Gte5krIDJinTjc8YQpElD
4uDXzOPw6y9H3gWc5Gagvw==
`pragma protect end_protected
