-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
H82Ye86hSV3KdmG9yQlu69ij3fOZzTp6YzPiOAjZjqmlZtdInVLG9xwUuDqDHL+cNHtwdQvUNBp1
Urz/1/jffZ214s+XDNSazd2AzbKu4fJsgnFuiA/S+96eHujfIttcNnRa7MA7h3V6l7DBm4Z0ikAE
HawVba8E1at0ugMKlzjdPgNouQTFikVovugu3AXotYAo5KILtmUdEI4dro1srHf9+oNxiKm9NCJi
+15cY/hIa9fI1TFeDJNCdnMM49h28g3XUA0jujkvEfQq+R9ncbqYq0SlylbGj4pWqQFZN28w9GvG
0WjClZmMYO3/40k3OBYvtH9r4T9Qlm4JkcHSvw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 5328)
`protect data_block
d6Vh//y/WBkfydO0unU6Ss3Bw2Gcy7MSviebR8Ygggep9LefZFyYvj/O+4vE3f70eIkHwBKZVXc2
JJ84gd/tOU3VCI8sspQYoBHI8xpw8K9AbpBZnSYCtNfEvamGPEYt1Lm5pNAp46IvVDSqCU0h4khK
KWRcSxz3Lc5P9AI7wFRohEMs8Cze//M6BAPb7yMO5b/tI9nw/96kAPkIm3hcrgx9LNNvlxzSozIj
2lJOPOdomOUGye85mqRupOPDGsZCslr9/pgo9hlsjRoAx5CJtvNoV1D/pqWt2PpWvcqQzUTL18HR
o19xva8RWy4AoDTsT4o/wJq+X/F2z4YaNduskRlqWYj8soMxJKpM2MSfHSuRQJcjuiBQHostzAUn
RJ3x9TUmzOrnJTkIEvRe+KsT/setlQvuLr5THcZk19f+Fc1PnxomIHNLpdX8AS91gK3lZDK6vIY0
Hdh+IqtHFLnljwPM6zwdipBZsSJvL0xBUsiUEz5x35q1DXsXlq04FqF0cT7xjI4KeFZu9hWoLlt2
mvifxVqi+tCYigDQptIHVY8555YAoBCU97QRdigJGdNw04NcjpcSNomDZt6nWdiSOV150zvZpSjZ
fhobvtlTuNvlKBQR4AQ07ReXlBqD2M6Qru6psLGuHGWu+qZ40bnYL7+KtEv0TwngH/EkPUdOxkRP
+8lVQZU1k0kiZ6bb2/5i3ZcSMo8+X6RwQ6fSG2xhfdGqPfgUCQkb9dK4ahn+aWgqsdAfH9Mqzl8A
DZGpcXwyEvKUdWlld7709l6TAhnqX8N3FQG+r8yBq7ZDteHOj7PbwVeIB9eNGW1fLBTUBM9fcoGj
RDc+dV3Ydzf7meVMuDH2uu8N1fzBl81gJcPNNg2llgd7CprQPCyK4LSJZ8XgP6dHWHLPVP0Y6fy6
rv55zcIZZJv/JA+uqwrB6Cw2vziiMDufbE79ZnvZRv89xdROqPFxTcJ48Q9rZdzz1fPvZSVx15J/
BkEnE6jkBJeJ+gRYfk9svzXnjzVY4s1Bchjch2Smxgf+gdWGOL06MgChr0ytVHKmbKcg+ZNZ3F0V
2uEwWfgnNRQGlbnlfTK5PSOU49EzvbRPR9cSYucs7I9w4nP/zRLZLAuNN6voA3mxpJw9Mk+6HH4y
kEImT9QVosN06itDcvxCPE/jJ3lUeQ51REWTGMOr3OscuRb/QEm9iKzvcXrjLpflDmuwh5K0Ks35
o/Jt9FimOVIqVLLHu8VoWp5gJOcdRBsUVMElMaVeSRKXxqQ/LYwimd962viWKxE0zWd8x4c6Vdwn
TZONGbCtTMZqsXoFLyc70pq8UkFu/G5TjNJHCQi1b7uFOKVvyfW5SfBPpP+roUHUAoYkmhCdHykt
fGVw4MkyjLF0DlQWe0rx9Ao55nW/gxvScJnTFiBwCo3unnigYP5IKRjCLzi/TlFwd5yRJ7w0nAPK
ZHOIUmO8YJOWYmSqyd190NUjopCQ++aJ9NzQw1i36R8YmpPy8LASzw0aefWGF+ow8ookccPxVD8d
z2Invb+PAdEzZeUY+lfFCDtMy2m5nzuychKE4yuYZExCjyvug+SqoHSyRATclf1fvgZ8984MCE0M
wU8nP11pOZt/vXTfv0E3qHRQtjOvPcVLSohfvK1i2vtQ0mfa/bSJoZG+Tx07QRJ4v0Ls+vDW+rhu
RSCB032yvChF1sgGB+r5LQHqA4J8DKersy8luQbMzp2FmvvEeqFlNr0BpLhG5YY8swp0D7k8YKuJ
GiO+1eh0cvis9XHnUzPiMs9rb7YhAAleMs4mEuujTwoHHThkqx0MVByNWKJaNj9VLf1o7Vsc0Om2
EsJKkRPpdwiSZsc22c+xpVDCM+wc14ac7ykTY5OmNasbefeW42UcBzynVz98vVn12VDcjalGC81U
UFw0UNY4NF8rtfWrGhTksMn0zToGtN5kQpHFdEWNWxXWZVclgcswURJVZDURkTcGYfOhWPAbTzSY
DKQlbgaTFcbKDtnZsezsxWIfwnBWK0+nrUnPBIYgYXQsUzFMwMxlHOUAVF+p6lGaiDxc5/G1AJUw
4XozseI93BkqF9Nt34X8Rpi0mQL8yaOPGGrzD5SGSGP6vo728YS/YDtMs6/UzEaZL9i3S74672yn
puzV/hGJP7uqwcq/NDB8KvLS9RwIAWovTucVrpdn9Z0WBpR1nyDZYXrGvwAvQfznkbeJxu9yFA8F
U4JPfVaHlWbH4L2HoSSw+cnGDdBCXpES4yIo2W66mhCbmlEyNMZxuMOJmHibYLfotZNH61sAkUNX
KhabiKrKgsMsbhZGF8HUhF2SFA25vE88TF613d1e7hbITObWNBmuIi7xAw+/pMjIKmpvNbkFjQoq
F82+NTcEUuxfUj8cxA03bSpp/deVItr6YCvn/jIKyr7Zu4TZTD/jjViTE+ALboQIk7BWYvXA3xBb
Udz11Ebn36gOAJVPfKFZoIZqfFCLlO8vhKrorg5fn9ZgskezMoMU2oq5oJawwp09Vw3+B7Mf41Eq
MCiYosI3iCxe0ymKNwcdxMERAotH4X/KgWA05KaBSJj0tSNQB3ZpDJO6LTspY60Cuoale5uXTPwA
S7YJAMuBEewVLvwlBVnZJM8DA1uF89JB9GLwvVpJkBVmuZNrgtpDVsd9TgRPVa/TzJw7Aa6o5F0J
fQz1fREypNStqfngYIkQ5OfamtMUR2SCjnIJaQ49dQj8L0uhn5GNDO4dCpe/DvFuwvdBD79qKSpI
XjUYMOHiWt0y55NRk5UsQBrmo9iFbzQAxTWecc+5a4bKnlynQUADSZhMqEp9h2Rt9DkKDre6O9J/
dWtViwS17uXrWAyTu0f13Mrzxxr4SMaxIH4l++ewcQj1xO1GgwpCSvDQshwkw0nDqqfolc+XA/o6
X/dGcmFoBb0Beok8tTjxnfUMYSAo6x36utYKHlHFyfpvViYbXdSLiaHQopS8BjHs7jFYyh41NCYN
iU60ORnRH17It/xY7g/gi1C+Lm/ld8ccybH/46FUYdQQ4ILZmY2pzyFpX6YfJWxlgynTO708sFig
BI3FNZkCjrZoA9WXXKASdmGBRGPJhtBnfe/kjPoJvC3IddZ0ZhWIvSdKBvUw8gLVR1yGk+A5zcf2
k+1jv8l4TZkqG6Y9ApoioFnWXiHimamW+kl5kPDSG4P2ECL5Pdut9H5D9615/EIeci7dG7rT8Mcn
kKag0GJqFC4IytVar02XN718Amk0gaH5XBHiGJLrABcJmKPurQXxKP9zBhdmM5VnfZNLIHXBKSiO
N1In8k3l7svyoecRSwYg0gyy6HI285pi/EIsRGRsci+FFeETNqAUe5DxhH+xjbYkBxWVdBzJGNNz
cR0etLhJtQCy0V743k2peyVlAKPe2QiwrLUDeIgdF8kxBk4PG7HCBDAAzwiFak72+fe/7Xp0r3wG
nC8/2bIQgeY+Kd4zmUO3WZXfgFCGpSQLMiA1fPby85eq7DWDBWLfEGOGs/sPMKkyJPLiPb8IFymq
4yThZLdnARngeNUpjQ1G1v8tuL9Y0U3xxwaJWrKpWD3VW5Tl/JcGOOim5dlBselLHqXtOj+T5wWn
jzUBTyHCZGBbDLvp2DbtH/2DhHI0E4AGMuUxkct0kDeMVm0DLGnbESqbnVlHK3bUZ6kLiZguYE+e
xx6r4bzjUqDgYaoQmBf9U2AwBn1XsBCbF9rUC5MF4qmpXodKfQoLxsGmRQcq6rVVmlN/J7ds5g4Q
Itl3tXFwpA/dHykyFWvo1/p2tkCDMEorHMqqlJZgIEuuvoqd98tWjWH4Muzv1tOOD3eV5OiwbDwh
8PpjSla473vgEOOtZKWl8M32XFd14D3Y7HPxWoxytzn1+nwdcFBIrEBoXHkwsKTzi6PLQGyOYIVU
bN3S3XO4iozej0LjWz0j+Q4eZ1xF5iApZPU9/kL7QlWehL1VScw89rGB6LrfJ9jPifY/Seg7Q4VD
TyOfm4kFO4xpuDAGf+lGzkQq1fnKbZ3NsY56rMmld8NsANyMo55OGrPEC2mi5EfVQ/11TEvA0z9K
v5L6Z5X0KbDVIUzF+pzzt8Ml5TF6Qelxz1TJZY/ID9msONFdBLKYx4h/CLJK0FOq6Rn739kqzaFx
dCM0fyeGqDUYdq4MgCt0e+rD8aejPBWDZRvhhqwmz4Mxo/YRGKFIdk/HFYlGdrznTbsleZd5tOwq
Vrur5dj51v8INpeDokTbkduttT2igFpRkpDsSL5x5cYeexNwjePYmgjN5h4cXZw0tQNbKxa33RSj
xXZhkwpTJ5d6xcm+J6pneLNomVltE5KI/eQfrWex0QSDDi4nHf+LakeqJ2wTPCAwUHRcIJ1209r4
T23VTy2s1Dl6ami2rSsThtqRu/Dtxr6qpJuIhyoVfL+peoJGgtCnJjLH1W0ybb9KohvjdpBe7gZi
2mTYAl/uGiJR+/MW5+oXuKNQlprxbHKLbuaKj5IArqr2OptKgBaA8X3Y4xbSw+X9owQdK/rH2vdc
XdIu9n3qsohP9aDCuDHK/L3/7r/OmtI2bY8iTejXlpgBFLqTm+iRzYjCgDjqh0LPwyHYzoOYXp5O
m89uEAdEePnIvNs0M1uFeqkk+lUB8n8vqMxdRyMzJv/gZesoN+SgMu82EsKRekGiRqp7dSzmKlvj
kKOB12lf+jymKZI2X8Sr0ohpkz5LtI29J8dlVjQGL4imakBpGdH8KuJvMlY+8tlPlONB0MubELaa
llye/HL4OytHM+nK8eGCtBXO8m5ge2TjRlRQDspMLU1z5DN5e81scBApdFJpbAXzoZhiT2832rIs
WfY2uemJM9rCxpaBzhxdtxdPUzOjgMugjGUvmlUU3v32Nxgyr885+39cLaSoA2T2+rD7uTUDtc4e
DJpBo5ZnYy8thj7PpPPlehpdgylKf6m5pEkr0uFXW1JB7OQxrMj0MH7CTc37+dNldSp1q1UFAJcv
ghN289uKq0R8Hy1UATClg0sHzuTdgaeW1C86yzrNS+eouQ+cGrwjCdOp6kfK87x9N7Dn3y+rKy7C
muP2HUjytZR+p84OS4cEIQnzuvxvyCTT43vTMlZReRSbxMQ6PyGyZexjjiBhrb4n0OPuIBEsurZF
P1SrlBlE5gsQn4LHz01uszpHZRSFLVxsQklZew5gfNkddOKEwQ4TuMABaCNV9CbSuKpPgPSSXYQF
5aOXZj7LvPgKKsenxP9zAJlu0TsytfAembPCXC6xtPbVC1GuOHS/jPi+6A4T3RxjseiQFDUN+roM
csu78fzeFmr3e7GTzBsAOMDSoHrmzdIL23crFXf6p3AI+v3I3tZ5mm9Q9KDh12P9i9ibAYefioUj
a+Vckat8nyr82S8egEf+fUWMqrikRCa8BFYeFL1dxsFFTmGRVAvF1qWOkV03OnOWpmxLF3Iwnf+P
sOTuK6x6iM97tEpwNyHNic+PebW9r1N2v1cwXFiDI5S1tqd3tK2n6nEFjQ1r5JuKVfsJVkENmvh/
y2JbxXJ1OR7hvZOTvu1UMj8kq4m9985ggWVHroP/trYzyrkAmh7KI4J1xRJSbfoBz8aqcU3WoOH9
2dtctP8vZiDbiRVAOXwpjnRrm5rEt3JDNBNYlh3b4SclXjCZsB07RdsHUCAUz8HzxvTfhwlE7VcA
PSRQsEuL67vpfQVAc5qOOmBrSqsXiVVhKcIRcSEJExLbM2goHkxair8KpBmctj5BMeneySqZzMMN
3Up4SFP8jANKs+rtsBHtOhiXN5mxQyMcssmH0cE9nGZcjhhd5q51tTRMP0qPUlgRvF9qjGO0BeK7
GCp/6t3E6LXT+5aaVQaAa++4/I8Uc84MbxeWIMghzLOaMWb7McOMy9H9eq+oSTSnatanFs81gN2l
V9fwmLkhQzkIXMh9fTD3ufEnaQLae45yK6TvPcC9P6Utve3n2cqNTXHPwbj2B3iDocPGtm3hBs1h
z/g5yBhzCZScgJZAtVDQiK/e3P+mhtDen4AL8nKjxKkaDd6MbwrnbRQ9chDq9pLY+QeYBIwzKAGD
jnbYkDKjdMGxrl5XAHHEDy7CoLV/WAp+gTZA0G9u+pDMj+yirLm5cyiihIADsG4L1V4bPdmjXktt
oRVM/wwekbNJUT+7Brv9ncgLzBhEwpj8zrr2EJ/2T6uzAwbdZqRXGGxm8dBHI2YFH1jJzq4h70oU
fn8TQ8wdPmTL4sVP7+TYKlB8qDNYfrCsxdf9DjyYNUS05uedWcM8vnb4Uy7cW7ywQ9hC13P8Xu82
K/yCYK5EhuaxJ7h01MsCGdnyLk7jXmqg+w1E/xr6kbXPwOfHD4lUIazocOOARoCnZYVVXICQit8A
7Xbn3GpBjb4afc5nhD9qgnxQaU/WemYY3r9B5p/tOmpUeZSmnqMvEq0m9ItVm4nsvTbGl3mgYupm
jy0tr5F58y6URUP0XCeVzTupxhVEF4YuZCCgkb2JFIpOr9xF3gh8oCM1AcmTxLfyTvSjQm/lJkDH
Lzzd8nkBZpzmFQyZE402TiF6XWnMyDc4rLCqsLfb9E4J9WezJSomwNhbC9snBZu5nH7RWcUEpVDV
mdvgFwlGYmiAubVANMD0BoqqV2DHUEeenVP0Paa3JS4XxWC4+YvPQk6B24CvaLt0RRkzabyq/yGl
T1hHSIxguKIStxIuS/nUkN8yH3ulrRqHCimsrXSnNcejDggXA+PgcLTSilAPZ/TRCbZjvQVue7e3
fVbOM9+u1qREUocl15ahx6Wcs6QSXgO+vXAwSJ4LLjE7U30cyF+HXiBoST9NTP1RyKzIRqTVvhNG
KKl8StNWuXNozaUSXpw52sid0c1xDUQO2WEWGK1PO3UI8/i3SPEEMdn2nNXxKbc3vvcwtqCKD4bJ
yZ9+hf11yQaYlW6a8mX47lfjY74n/3aGQNtbRTsIaYIb5EFDxn7QhqH2+5FwpEO3PRN67U078tbD
8bT0wP/3k46w+FlAmRXonZnIfEo1zuXuVp2f7fQspG7x8t2+H6eqIS5Jm49LfONP3KUAYK3zlwYW
s/IJ1FEMirFG7G2trUMENco22IhluWWz+KZzM8SXNsfjR0TVKD1lti0PXgIK/xZ5NFdC7WR0Jbdk
7YlNwBZhulAxcxxDZh9jsUeaCX2iiEQRxoqn
`protect end_protected
