// megafunction wizard: %FIR II v18.1%
// GENERATION: XML
// fir_v2.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module fir_v2 (
		input  wire        clk,              //                     clk.clk
		input  wire        reset_n,          //                     rst.reset_n
		input  wire [27:0] ast_sink_data,    //   avalon_streaming_sink.data
		input  wire        ast_sink_valid,   //                        .valid
		input  wire [1:0]  ast_sink_error,   //                        .error
		output wire [19:0] ast_source_data,  // avalon_streaming_source.data
		output wire        ast_source_valid, //                        .valid
		output wire [1:0]  ast_source_error  //                        .error
	);

	fir_v2_0002 fir_v2_inst (
		.clk              (clk),              //                     clk.clk
		.reset_n          (reset_n),          //                     rst.reset_n
		.ast_sink_data    (ast_sink_data),    //   avalon_streaming_sink.data
		.ast_sink_valid   (ast_sink_valid),   //                        .valid
		.ast_sink_error   (ast_sink_error),   //                        .error
		.ast_source_data  (ast_source_data),  // avalon_streaming_source.data
		.ast_source_valid (ast_source_valid), //                        .valid
		.ast_source_error (ast_source_error)  //                        .error
	);

endmodule
// Retrieval info: <?xml version="1.0"?>
//<!--
//	Generated by Altera MegaWizard Launcher Utility version 1.0
//	************************************************************
//	THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//	************************************************************
//	Copyright (C) 1991-2019 Altera Corporation
//	Any megafunction design, and related net list (encrypted or decrypted),
//	support information, device programming or simulation file, and any other
//	associated documentation or information provided by Altera or a partner
//	under Altera's Megafunction Partnership Program may be used only to
//	program PLD devices (but not masked PLD devices) from Altera.  Any other
//	use of such megafunction design, net list, support information, device
//	programming or simulation file, or any other related documentation or
//	information is prohibited for any other purpose, including, but not
//	limited to modification, reverse engineering, de-compiling, or use with
//	any other silicon devices, unless such use is explicitly licensed under
//	a separate agreement with Altera or a megafunction partner.  Title to
//	the intellectual property, including patents, copyrights, trademarks,
//	trade secrets, or maskworks, embodied in any such megafunction design,
//	net list, support information, device programming or simulation file, or
//	any other related documentation or information provided by Altera or a
//	megafunction partner, remains with Altera, the megafunction partner, or
//	their respective licensors.  No other licenses, including any licenses
//	needed under any third party's intellectual property, are provided herein.
//-->
// Retrieval info: <instance entity-name="altera_fir_compiler_ii" version="18.1" >
// Retrieval info: 	<generic name="filterType" value="single" />
// Retrieval info: 	<generic name="interpFactor" value="1" />
// Retrieval info: 	<generic name="decimFactor" value="1" />
// Retrieval info: 	<generic name="symmetryMode" value="sym" />
// Retrieval info: 	<generic name="L_bandsFilter" value="1" />
// Retrieval info: 	<generic name="inputChannelNum" value="1" />
// Retrieval info: 	<generic name="clockRate" value="240" />
// Retrieval info: 	<generic name="clockSlack" value="0" />
// Retrieval info: 	<generic name="inputRate" value="24" />
// Retrieval info: 	<generic name="coeffReload" value="false" />
// Retrieval info: 	<generic name="baseAddress" value="0" />
// Retrieval info: 	<generic name="readWriteMode" value="read_write" />
// Retrieval info: 	<generic name="backPressure" value="false" />
// Retrieval info: 	<generic name="deviceFamily" value="Arria V" />
// Retrieval info: 	<generic name="speedGrade" value="medium" />
// Retrieval info: 	<generic name="delayRAMBlockThreshold" value="20" />
// Retrieval info: 	<generic name="dualMemDistRAMThreshold" value="1280" />
// Retrieval info: 	<generic name="mRAMThreshold" value="1000000" />
// Retrieval info: 	<generic name="hardMultiplierThreshold" value="-1" />
// Retrieval info: 	<generic name="reconfigurable" value="false" />
// Retrieval info: 	<generic name="num_modes" value="2" />
// Retrieval info: 	<generic name="reconfigurable_list" value="0" />
// Retrieval info: 	<generic name="MODE_STRING" value="None Set" />
// Retrieval info: 	<generic name="channelModes" value="0,1,2,3" />
// Retrieval info: 	<generic name="inputType" value="int" />
// Retrieval info: 	<generic name="inputBitWidth" value="28" />
// Retrieval info: 	<generic name="inputFracBitWidth" value="0" />
// Retrieval info: 	<generic name="coeffSetRealValue" value="489.0,876.0,-70.0,-2692.0,-4749.0,-3398.0,555.0,2463.0,-170.0,-3341.0,-1651.0,3095.0,3463.0,-2093.0,-5255.0,-34.0,6339.0,3092.0,-6151.0,-6637.0,4218.0,9891.0,-396.0,-11899.0,-5023.0,11705.0,11244.0,-8596.0,-17023.0,2344.0,20835.0,6597.0,-21160.0,-17006.0,16843.0,26969.0,-7462.0,-34141.0,-6396.0,36149.0,23002.0,-31106.0,-39563.0,18157.0,52580.0,2100.0,-58413.0,-27395.0,54005.0,53847.0,-37664.0,-76409.0,9709.0,89627.0,27145.0,-88625.0,-67787.0,70207.0,105197.0,-33845.0,-131396.0,-17662.0,138758.0,78005.0,-121521.0,-137805.0,77247.0,185706.0,-7947.0,-209996.0,-79344.0,200625.0,172776.0,-151266.0,-256696.0,61154.0,313452.0,63640.0,-325790.0,-209760.0,279512.0,356995.0,-166075.0,-479596.0,-15262.0,548125.0,256015.0,-531263.0,-537738.0,396490.0,831504.0,-107394.0,-1095361.0,-387855.0,1261530.0,1194690.0,-1171615.0,-2607191.0,146187.0,5583607.0,8388607.0,5583607.0,146187.0,-2607191.0,-1171615.0,1194690.0,1261530.0,-387855.0,-1095361.0,-107394.0,831504.0,396490.0,-537738.0,-531263.0,256015.0,548125.0,-15262.0,-479596.0,-166075.0,356995.0,279512.0,-209760.0,-325790.0,63640.0,313452.0,61154.0,-256696.0,-151266.0,172776.0,200625.0,-79344.0,-209996.0,-7947.0,185706.0,77247.0,-137805.0,-121521.0,78005.0,138758.0,-17662.0,-131396.0,-33845.0,105197.0,70207.0,-67787.0,-88625.0,27145.0,89627.0,9709.0,-76409.0,-37664.0,53847.0,54005.0,-27395.0,-58413.0,2100.0,52580.0,18157.0,-39563.0,-31106.0,23002.0,36149.0,-6396.0,-34141.0,-7462.0,26969.0,16843.0,-17006.0,-21160.0,6597.0,20835.0,2344.0,-17023.0,-8596.0,11244.0,11705.0,-5023.0,-11899.0,-396.0,9891.0,4218.0,-6637.0,-6151.0,3092.0,6339.0,-34.0,-5255.0,-2093.0,3463.0,3095.0,-1651.0,-3341.0,-170.0,2463.0,555.0,-3398.0,-4749.0,-2692.0,-70.0,876.0,489.0" />
// Retrieval info: 	<generic name="coeffSetRealValueImag" value="0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, -0.0530093, -0.04498, 0.0, 0.0749693, 0.159034, 0.224907, 0.249809, 0.224907, 0.159034, 0.0749693, 0.0, -0.04498, -0.0530093, -0.0321283, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0" />
// Retrieval info: 	<generic name="coeffScaling" value="auto" />
// Retrieval info: 	<generic name="coeffType" value="int" />
// Retrieval info: 	<generic name="coeffBitWidth" value="20" />
// Retrieval info: 	<generic name="coeffFracBitWidth" value="0" />
// Retrieval info: 	<generic name="coeffComplex" value="false" />
// Retrieval info: 	<generic name="karatsuba" value="false" />
// Retrieval info: 	<generic name="outType" value="int" />
// Retrieval info: 	<generic name="outMSBRound" value="trunc" />
// Retrieval info: 	<generic name="outMsbBitRem" value="12" />
// Retrieval info: 	<generic name="outLSBRound" value="trunc" />
// Retrieval info: 	<generic name="outLsbBitRem" value="24" />
// Retrieval info: 	<generic name="bankCount" value="1" />
// Retrieval info: 	<generic name="bankDisplay" value="0" />
// Retrieval info: </instance>
// IPFS_FILES : fir_v2.vo
// RELATED_FILES: fir_v2.v, dspba_library_package.vhd, dspba_library.vhd, auk_dspip_math_pkg_hpfir.vhd, auk_dspip_lib_pkg_hpfir.vhd, auk_dspip_avalon_streaming_controller_hpfir.vhd, auk_dspip_avalon_streaming_sink_hpfir.vhd, auk_dspip_avalon_streaming_source_hpfir.vhd, auk_dspip_roundsat_hpfir.vhd, altera_avalon_sc_fifo.v, fir_v2_0002_rtl_core.vhd, fir_v2_0002_ast.vhd, fir_v2_0002.vhd
