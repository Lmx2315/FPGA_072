// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:36:47 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
n/R/49UhU4ZozsOG242NByEEZKDr7LuLtAMZqdx2LyV7YSaXjQX/qeE0HibDUNdF
3+la6Vvzl8EIUVhNU32DgLx8/oZBUigkY+H3aT2f4ZFAjuoKk2KlaRToj8dXPhVM
1ECQ4cSbWLuOn2jgVN04XB4kqWePoDehVQ3cVuPEH8Y=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5552)
Oixq7jmypAajhEJ37IWDlLI6xZFYyx+qqfWs/nu2BbCVSl5i8Lwh4GC9IvIj3stM
v9aMgUijMURalO8FMIoTAHlploZI6aoGs2RWwSBNOYFnXJZ1wsO0z0gOUaD1JAiA
3RypauLOvSuvMGA1O6vqNR0qBghZ6VKIHE8c121frYP69ky0EJljNKdWroamEzAk
svFx+vPZThyGhi1g6Jaf0XMD08uN9OByPFXzykYDH3c1wjfolohjKQeEw0gllsBM
YOX5A8dSsSHNI4qKqJU8C32u78IaGkWL5pUPdALX+Kz5sv2f5FBVcCTbNiHM4pHI
kVKQkClm4hNSW/GPf7skAZa3RYExiGKEMU+cVaZ+qfRaUQtTaZDHt9eJkfXh2OwX
LdnUxyAlIFD/neu9Ksw3gjzyXuxbGduOzPuLr+zImszjWVaRogl+r0CEtHsr/rvW
8S10lwM7yNOgh+be0FZyOl50Lml4MWAy+e8QFdTjK9A48D2D0l6vIO3psj+DTuih
Y/XD3Q4J0FhRBh+QPUWY11X4RdXVOfiMtfPoVSIsawyoOM6dvbgNXZuQmR8qmLwE
q+dR14XmCQXqPwdNKC8LsnRoa9s/5i6R9nemGiIxN6Hp8uu9VwEdojPkL+/+iFbd
t7nol0IGZkxHO1CVyS3Rcy3gEGu7UJNQ/cl8LPp9a/+qbJu7p0MjtESODOFw83Iz
fz1zoiSIX59aIWUj5gJyCqSJ/WrZgq0OKz7PsDwiVAlg9lSRdKYoHqB90M0Gl8AZ
8/dXq66niPAON81+myVpHt3JSzcELw6OvRkvpf+kw1xOssccgPO4/bYEaq+kIdmD
qeIr9jLz7gkHIjp++j1BRrySisfLYrF0sf/leR+Y8ekAPBXrQJQaq+h8p7Tipi1b
JdvG7gooqNcGkw8FE9uKmPU81uPRjKgqUnTpBXZqarfCog4YKiUMyDqW5o9YWvqv
5810pUB1bBXbdT/JRs9EW2o8Y5Yo3T1VHWJznr7nNGf2JAImybI93spSt9dxBEvM
rl7U3dlAI7sl17L35uTmUlCA9R5zF2lCr+WNHVacUdZj8+h66/0RowNfI/pqvWPD
boqgcKbWcJXzExtP7uf4KfZAa32ABviHJA2if4T3YpuBXh5OnjA4RHBs6/2T/ktA
PND+8YbygwmU2lmNoMB4TpqbKt7gMvox23WnJtUBWWZ6wz5ylZFINVCv7CGMyxzy
ClrQYgcCxMcpYIVBHnfhxiSR2c+xCAU+LDkKwCJ80GbNv7KO1/pOtffMzNPgriI0
NGbVKdqks7Wp/lgs/jETuTJy7o1a4va0FCm+fQAKfFAbifWnVtVaTejLcmLa+cVr
jmZX+bxC43Y1HBx/Vzd8u2b6X+eED7DXia+nnsuVJ92OOqSDdfreK0W9MbQAEOAx
74TPY+n44syfk6Bno/EppDmvb8bbTqTtBKTK/kVgeKi9+MVYESMHnZKdvq2HceT9
zXd0ZEbt4m5biGTw3K/+dbCrp/B14JXIu+q0m8hCwtwEhy58jwU4mogf/xRNz695
boiVk80bdDFNazNEB3y/dn6ET71Cw05TVJty6EuuJAasKOM84CeyOTexoR1Pa7j5
XJclmN3srzUVUkZC2RkbF04GMU1VuaeT5PxLp9W1gqGyyfP5Squ+BIt2NE9m+73b
lSXoAWgsXj+GK4gs3GBVwInJtM4Bp0IRbUAonm5mnPK2A7sLBWOlBl6cwWqtPVCR
RGHFIhAS7i+5e64HsQIvt+c48hKVm97BxF5Ab0lkOdgNLhqatn6lUDoQQtLJwA/7
s4QzChwqq5hk3J96sE6k+VWN+5MGiUPRjw7Z4tOl9HTZownogXgTYGHGQXwhxLJd
+qq6NIa5i+CFZcF+7RMrMYOKquEs4CqKLKH6Vd74VYGpjIw+nPK6yukG9DA1KbNI
eD1dAfRmZxIWzC8eT0tUhKdruf/q49QAF8JgSuj1u5MNoXPQ5h+w/75La9QOv3eu
/u28qCekoGVBAX7x6FbwFzpjNcViRuA153MXl5pYM9RuyePVcNc3WdWbz9TB4KNx
8n9hbJnEHeGA+evHkHH8UAQaKy3Aka7rbSFW/PodW5EBb9TAr1fTk56UVLBtX4Tx
t9a4YwC5Rby/J5UR4IDZOQIjRaonacLrMoNadJ9wy1PbS4RJGcSKhDQ7lwDKbnt8
egcqc6QAwIVUPjv8KH15NUJ+j59NYhqf/hpzJCCnpylcnWd5q4pts2F4FcARQlN0
IWb8UXmEfXsXMmwIwOTdMBLRxNgCDjkU5Wp/LBiOSw6nvyVYk9QwA6Y6XGIN8EYD
bdAdVyUy6xyGJW5mOVmxJ6R4lg9W056XmA77ho4rHWvSjhNlRFhe08otJBwQfpK7
5RyG1gH3JX+SvOZECN1JXuVF21FAtprIzJiAVuKgaMqeG3yN3+0l1G2dLNDE8cN9
KQS9u/BD0lBUTfoiWaVgrF4DKvao7ThopMvz2JsnxpORr+7yG3b5EGr9YcsR2tBM
8kjpWAm8x7s+zVH2VXv5ipPT4l7G8SzNugMKkRvC07Q9K9MrpkmkJEM9lB1zhJcI
+BP767nf1DJoiOP78qo+ULsjCNC06rtSehT72WqeyZcUBLcLDcG5psa8JGNS//S5
8Nzd5ZanshOC2GlffigS/U1LIL4KOdFr07zjBnm07hjfcSPSHtRF2jifaoI9CDKK
EGBo3ScMPxGA0z8HMODks1ZW8EcJZsoMYm2mo/hcaDv1Gk7cKMnXffSDsN9/5xrT
TEXAF4DTN0QRMejezw2oa7lvmIbJdTREfxZTxZh3jL7AW3jBR4dj5YXqe7yvF86j
L36rWW94wXGMjrGOsAJ7shSx2viJsNWCt0E4mVvdio/nKNLOvapcinyO4uG2eLEg
mxSqbSYP+9B5VYdgxMDFhWE/RLxLN8SrlSZnsUVtUe7ANVBFEI0hWR4xA2trSUAt
FiwybUpBriarISaEBbiz5ykRzs4u6rF1LI9mDfGdMQqZPlZgmmnjEelhe9+VWrkz
4krnavs/OsTg/7LFcafiz7tcTdTd75hbp1MEXu1Ggu9dfNnCEL5wp9LAV3nZSb6A
YPjVFeAbk03W19ALiAI0L/F4nqaCh+zkRWionXw6EmEmOSxPmOXXlTQJZegm80ma
W9T2soRmw/cPVI+3Sk61+Ng2/FYD+Y8+bbiSgH/7tFGyog5Gw8FU/vkQp1wOqJ3B
PbwN8NtyGVppHOtS4lb58rqBcIVLsUcevB8B8u+6YzjzArGvKs8xj88Wao0pjxFI
Cw/q9+S/ixlpt1IiYx2FbUL4zvvHyuAXlfpQC4dXfr51lWVwz29W4aLZRDCzpixA
yIqkQbISckFoOcTkWC/n+EioaxI+cZdGgWU7wdCOiUakZ/1SH77lUQiqqwEQ0B84
S1w/dbZfvngbkwIxiTQbv0Zxe9ruFJQHs83FnaWMOnLg6f7O6C9XC54G6i9Qk6gF
9CBr7CkSv8TgA4noqacq7fqOW0Z+WNW8dGQEQrOkr0GFBpUPjvqLNPso99sq2BmE
pLu2bwShmwEri4LqaTpA4mlufXD9npHGmnJT6zxbxyt550CIIh6395ssKf85dsyB
0r0mLxC2eG1HyA8xJ7cljdumI+mk663N2dbdlfWiP0x1QX5AVyHjm57l4HKMRe2b
HbqM/dHXpmpQNPPi1dzzYNQmLMMXTueQUY2Xog0xi9pjGept1YcqRF13+pk8JGeY
JbY4+G7HtwYOBMtx2NYGniLI/S7ZOFkzU0ovin1FU1kf6ON3WR07ry67YMu+Brip
inDOK9aRYbq+/01r1aQXxBnnrZbYe4Yp3zRSs4oItBduWpAQH93t0d5NrZI6qymM
6ZZxWZt3BQPzgBbz1TiLKzAG5uviPEvVosprCJKSGem0UGkaXEfL/VQKbdBn2juc
M7NLTC1OkSkXaZuDMCDLtbF9ASTU+NnN8z/BzbWdUL5w+RayBWh9BTWAL8qFsjMn
sWETXGmjPT7j5cBLc8HhhMiED/6o8DqQhkjxcVkaMWhxqgBXuktPzYimEORJoAcr
q1/Y4lDXGS/VYLgMRW1L6hPG3q6z1zzlyBWHzNI3cwzu2DIcjUfVqIvaP4CEnoR7
i0fjaLs428tHj4jHXG3yYPWMl9/X3+SuSc2rCGmFJKjPu4jKSy3HDY7k5wMvtibs
YAKfoKi4l49d05LjoFUMoKIP1PPzdqb0BiJlnFgM/8eUSVV9KjZkZc2X2rYMr5sL
A/zgMkURaCJTiT1lGBrxTgn9vCpHjG6pckz447K8ZD2zKSjsYK5ANgry/UofQh0q
y+S/D3mVHvgcgRz51+zY/KCjCZd8SIt6H9rkQm04Ay0YSXpuJZ5khRSyeaxLXJUR
s8zsQgWYVFzhYzPxrTglcwz8bmEzhIX5vjTBaMph1ZxqiiCnNjLmS5bg79jHuCmu
6I3sgZyZB3lpGUl4/SQKlXoBy+sEmLfj+noW3tFfNA9hZbFD7Q7JdPppt8JaPpJK
uKzOYlYRo+bK3BgGN+v3Yrqvzt93dGkew4dXHe4PCR8pHDOhqhfHQJG/sYc/G029
8TfJvuKM937/VBCFnJ37OfQeUXj1l7bSkKKwndBM+Kabj3dOKULu9jv8+QVqM/sP
LSv1I2ip8Sk3Vl83LmPD5VP3xgq2fAWczl1SxSYtw4gGZ1Ge80tRiSQhTXKr+/VN
ic7gLaw9zI4RGIIPjuh3pCYtbh+v1Wf2o5k6SkCxxbBbPUFHtI+ySOOyQY0hTqhB
c6Rfu3CUWpqbQK5mpvQnAWKr4dshdPyCSDgMXq7QajcEDovWw0xddisU8yo1NVMW
4Em8iHyvOpaP6hBQgbOj3b7SvsvqVW7l5u/GDX1md3DAaUEHSwbWPfVwjeEksYIe
8/+aWjMSVGeoACEUSQWirMxv3wlxjyOvmbxR32mhun4wL0Ra720nuin4iyyQKXSE
YuyoGpWdTVcplvjXWtlPvX7m1YEJX39RcfNxXe8/U8pM8DzgihTWKjgf3zvIEtIi
cOYJ3Demrmawk8KvayPWAWmV9dalRYviutUk6Ezsp1itCdaDGFwV9ELMJO9TPnDS
2m27aRhOw9RW6wdUPMc3BlP8LPDgAnMmgrAB6B8A8G1fY6O7o/MPyGMziSf3dmz8
z4NMT/ddPEg8X/1klK7wPx47zTwh5DziJxrcPAlkuiEFL3riZF2cUNSOcOeczVvY
UgFbvMg1luQfbesEnvuUqtZxffC8VsIg93tgS7QBCdX2ijR9dGOSizjR7dFOsCRy
cew0jnS/Xgh3njCSlg/aepbLFQpjks6SYdTwm9T3RcQNdhA141xq4IxRH1YREdxy
ICAbE/QheFH8JCRogWIkPtA/qp7ItF/D3Vbmhsv2UslinGb/NPNcOIcNaqwBVCq6
2Hel/fbRk4gNJosKq6r3gG9cv6OMTrNJPWaWlewJRghYFuLTIzaK+6QFvs/Wk9eW
oH6CE+NxYAWVonSjR0LZvd4F0Qmp4AaU66FMvhTWPxJbsq+PeMNpwl+g/U6SRPQa
CtqnhDDMeLqqwLs65xNkks243jD57qfGdPisYWRKS8hhkmeqGJ/a9pzQDA1FWya+
pH/YJ2dKH/pt2e8E2tXoOvAlY6C/LWkFz+ZzDA/8nO+aBYvUX99ZboV2onJkNbaE
BmBgsf8WwPKqfWMd9GLBMo2KRCXEUvSg9H7jkn8yOSeMOk5w8CFav5mw8mttVVL2
sLLJPJBsFI19xdo+P5bZ7qZrxc/CDXe/zjfTRKoyTYaDyRvDUau9ragUBP5wcEnJ
Ov1FWBtq4XLPD1yzKxCBedQYB69Pwo68B/Hv7FmxtzWKJDRFpLFCs0Je0ciWO8dm
2Hvzji0N002btQN6VypHWl7IZgejaHcKTTxRjpBKoQpAlmRxYcx3V5dRlXG9PsjO
1Lo2yAcW4gNCFbLcgnM7/zhwwDgVaXaBVlLpXy/HMitBXUhWphQDIPnt6JQyKzqz
Ps51t3opUd6pRuuwPdYU+uh74Xxtt3TF5LmISVwt2e6S0oQluHI1sxF74T+tUAPg
4Nt5NUCmcgaQe1lOm/tWn1GJaI53wzSxl5ctvjezneEN7bteI38ioxFnmVu78XJy
JXPDVLdBuLbi4wK7yIISkry5h0h9TqnHPOIxxOB6JD2N1CsVgX9PCpqIVfQvDyFh
8fLPX2q+BZSVRvjxw1XiKNgoW4qN3rzvi5SyuYjMrCjLxkL4LAJCXUXTIb3AASvd
o1Ci7W8XYmBi9QO2G18FQRb5GuYcjjmZXV8cPfMM3Dh5qXQCZyd3CE6WG7HaRqrE
HbicUC+PDxDuKhlKCFuk/R5QyxqGieIlt10Wv6zGfnG8fthwEXoz6j2Z6JJTi5lm
TnjQRC2xd1n1lk16xRwOFcr3JX9DSXM+zA41ph+y4Y8C9JR7Cj+pPoiDOrXrIQ7C
oiSd0PZ+lCKFzlcs1MQZsfNDN4AqJjNaA6A9zE12MIyvHvZnAxNg0F96a7RwhnxX
9T2NL7MAkEfu5AaqXPTHjrsT0gw3li5+V/hbrgXE5/mq6wFfsbBh1aEE4ftZkzK/
Crhb1fOVwm6fpni6z00Kj2gWBcuMpbXnvbh3vwXYaQws2wdqwfIgzIZGV5WHpZcU
ZMPOrGi6l2Jr8gUItKol3QRwG5C5QZz8UxTMMp2/6FzWe8g8W+Ry2KfHyDvfWA7b
ZbOdKFQwvjvP5Kj7N/f8Y7MZjpjByL9az0R1lQT4iBR3AELdCrDn/exNc7NDcY8Q
Wdz/AizZWcDeYdVdP2ZcOPP08/MwxHqMAvWJslq8cVZsxzLydQrIjlDoq6zPcDjS
uuKYBJCnS7nrJfupyfy1IU23PWdCeoSf9f3VXXwTp9YrALuDMSKEMjtCJBnSeUFt
W8Atp4bqTgXIn2UvMuFuVpLVNKdKlG9GVZ6AvBfz7v/KI67fV0oUNPrRQH30gdt7
XbS6ikGn7vKurJHDTX2FzgTNdsxtHa33NV6qUJLNIxq4H3zcGIMwD7a/vxGlwqux
nP9fhOhaeQ+MABTJXTTDiW6Biczyx7UbWt9fY5z7uzkU0lJUpG4O5K1g3VqB3Qnz
5cITKvNMiiS3Zow27FZ1ggOjp0wjgeOB0fyHjq1a4jzV8kzG4kYxZzg+ekjvTNCa
Z7iQQoM07AF4cOwZwS7yKSFfSusfxWZ4Pyizp03G/KgxFfPNgLhMAsgQ/Dx1LMdQ
OMPSexV9nMQFd2zJUNUBnCU8vKhkB3EM0+LH0ogbYWUn2KPYOI5//oNrgtEgLOyE
9CSirAsesdpMb0o+AUyyYtplbOYeMLr5N0fsqmGhlXOcZ3tjKBUoWX5rRZT/8L26
4bBZF/ifeKFKc09smz6bo856tOsyTeTcQJ5JDnbaN5lAGGCycbmVoBOIv61fEp1O
ezfPRjmtaXrEttIHCBD3LFVN8I2DuH3sMFun4Maj/cg=
`pragma protect end_protected
