// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:32:37 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
rrJ9DovKDZRhKm0+ovNU7wTT593sYfGQQ1ECyVumQmR8AesYS97l5/G+YVrzxkt4
4cqj92bXtijokgBUSp/9s4z17mAzgaYA1cDoxe3xmryDD6xYrHvzcoILzQ5fsSZT
R+8dmHQ6ZfSUWQwWAQl0DKXVJHs4zPW/EYPLQSRlKLg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 35376)
YoPhphC+syuNFpKRS7vgu3pFAcCAqX4OMgz+M0oIJd6EoYDByewlGomf4NziNc3a
fcLnVvDUPXqtQhQ128rJhwRKnf+NVScvcSA0RzbxT/NG4013bvvBm27vtgncvO3J
sZdtTqfBBBt7IrV7HMSBSr1SWKZQEMpjjqkrbBK9h90lLjQO0lbRd9lOSpxoSR/1
cct0hBTpgeBC42517O6amusBtctm+uqRT8T3wVBcqxEzsqpFEjJ33NwZ2IzSp/qR
/YmZb1RlzlKHyvA+7y1mk/iCAosTHIFfzdSj5v/5SjRinMLCHwJox8Mn3RKWgYA9
4TC/qUVoxqLz8zUmLEg1Qy8dvoi7ThgcWlpVfW462XeA4S6BpIpiiryuuCSSrmUx
8h2T6SYrU3Ia3FrxdkxsH4SWBaYtSwnmxaKBGaVazI5hrp7k50q9TaIq3AdDn8Tn
4JneWkH/OYRJoj1gbB/ZTlWchO9w1f8HKq/jixYlZ3XYK1ugbm7p8+s92e3p2piY
A+A6fpJeM8kDufTj/Uw/L5hydjSFgXmuqrYDrxa6B1GLaxdCp7B9QVah9dgylHxg
sXBDuwYmAB5X+1esdwp7j3wXu5asaHHX0F1q8Wa8pFFgfqvph89ZadLgsjRBoXTI
HqJPbIrrBmCNv6V/UEiK3qsdxA+v746WfbBWGasoy7yA1rY5RfKLYEr2pukA8HY4
2yUwzHKifbRaw3w72cx3/VG5O96h760Un9qsf/CSWd+IJ0woJ+7JmIH2Yy217Zrj
uC2xU+P9lSl5bpl6UKQAuSxmuhY5u+VhzAeMAGFRacfOnXaBFF3twVjZ1SiBQxs4
MKYAFXsx27lOYD8sjkXxr65e1XjWShz6M3XsvklQXEhkQxQe5KaOfAN6KRBXTR8i
mBeSPoYYjdjbEFmSrKjqqXCievo6K0LZRCaHX2llT7gFhbc0xiDoay0wb1ABMApF
M5/GjTXp1ss3x2Fq4vmIBEuYadAiLRO/CPe/cqeNxHLYw42Mud9P81v90hyVyFD4
MZ1cIYVBEuhtFo/DtCepACLqIKDzExeWwdkD0bcVAkbTVsJnp4csjzvKVEK/JRlM
Tt3zqx+eqDKhEbONp4hV76RqSiJ6+FIl90k+b20Lia79vhF0xZb5GSIANbPtc4co
PHe1nz1cY2g7Cph3eF9sJHIi2a/ld7exblcz4ho7fTK8mY0XAefVOowS0/C3Nm5e
hBrG2TrbB6QYBKycn9azwHJ1N0uKVBMQTtY5y4o/RcQ/6/BJfisX8tiKD7Iau2j6
K4NkBBl3pWoB9lYgaTVWKG2irnLD0wUZBp6V8Y8D8THE+m693SXA/Rc9zCeWSkC2
fJ+89kKO6RpfsAKvPuz0W62Jj0QxadT1/C9bClUE0guY3xJaurCuOianO9n1RrlP
flxDEYTxRrOarLXRBMrVb1NSp8cooHzprCZhmMeCiahric9MymSve0fEO2Ege1bg
Rqa7bnl9FiFjPLcssDDF4VQAbG5B/YJWTSbOZoj41mBbCggA7lgAUVgHYPRitWRw
7NHNTdb1dr/0Toic1fVIiOMHdNzP7zfVM9P1+DtfgCpKc2ETjrsD1/B19yNbTvow
cK/3PUHMn1jxxIcTk0yArV57+EL4oUVB0yy+MNzRIRojonXZEzhnwQjXI54B1Pc/
WdtbHKKpGCUar4xlUCZTlLDb04aUsRcZ3ckH2kHrR2bsEGv9ZeIt/omkIUys/wv7
f2hSSbqhbVL2dI1WHPK78nc9EpJumrq3p4Q75wZk5GRY/kvICSkHOdoWFK+RuGmF
oufF3iYNISY2Nnfz5aRT8HeP+MqkMMZvW6tlIn8vB8HVFlFCZu2BpX88RstACx0N
BI2sq3lOsJnDGc7TOtmjDfY0LNniFaHrYLXGDPguO5f7P4G763QGtno3q/g1CbDF
XjpvKpI8GgpoUA9k3iVDf9wG0O3mhcwPokUwfxLUXz8rMGuPSqi86bqVC5rU/iY9
XWCxX5/c/rUMI5h2jtSA6d8IUtNSTrc9odN5ptvaUszGG9hkNIhXV7g3wKWt5NC5
pVDc89zQF+iV39cEGNiyC0BzbPtbVx2+QvBaIXeWOlAl3nMYgJWNrK7c0CmFCS0S
ziu8TuAz0kPKxDIAFq5I5qRC1JxPbba1Ai8WsQrw4OtFVfe4YINuTMLJkCraWyht
tmPtZH09tdAF9q1eeQlErruy1LlXxPzlne+vHHu+CHnYvZDNpMQnFKzPt1rsePUt
jyhgxfkNILBlfQ9+t1Dpt7ioLfMe9UV0eNXp/f6XqwSNYWhXWH+aXIswMtOl7Euf
bJe99qWkCMK4L0kh1IfsJBC5zZNxsdmBP+NGSK5DFQrZBzpA/O1hPu+aX3HM3VV9
FWv9Mx7bDsoaco04DxLhCpXasWbQ3ySen/mzgA71f0E0687IAXIBm+lP9xxRi1hk
phdsjTMPXYtxJNE8a0dlzRdXCUMcIwbjJFkw+p7afpn7XjKlp4FVxFWJnUWPRvNy
klZCHgnJjkUKX3T3Hq7kh11e1Eg2WxYvIgO9ey2tv/FRp8px0Tl/l19ETKSaJS5d
FBKDWy6a+MEaVfYNn2uPq4jjOW5BQPVcOJfkgWPKiq5DzPeRRtfac+HxDfcCvU/i
s5cQphnat3146vCMEB9XAXnaVtPtfOlCYtPeCVaBKv9iSJB8UkUQxmq82Yl3bLCZ
LO7Kl3jWCGJntZ49QUgM+ic+eEQ9J6KvEUbdLE7lCPve7BDjOIOdvgOkQlUc141W
nhSZ/1ryLAjZ+yRB4Td67ZzpOw5jNwzpXwecQ+ob+9e9F9svQXWUENyUcX8JYsp3
XH0csMV9yQ+sAzIAwO2We89DuYH4rFWd6oj0eKcIYNT1kQHsvaU/wEiDXJbeZVyN
dDAhTTHZRuyQlwunLi9GVRUC/Os0OYd2+YG+MSD52RVSVI1IkZPJlQujHmBWx9Cz
g0C3jBvkNKtMulIySs3VeZ+CebsVIlMOzayMUdkJqXqMrZRKqQn+b8hOSDa/gJZn
wiQ1BddEhgIRUx1UMPAEykdfkYlC2mkcJXuNYvxAPbOwJLTPhuMFOfugMh3xppom
OvyEzcuTq1I1s48N0hylL0uMK9QqtFJplEhYoH/VibLj7wVxdPxaQhnVs5Jg+dIC
XCP9ngwjEvI35exYeLR7pa2D+ol2FIUJF/qrsUs7ENIphgXpWud4AbyId1cm760M
8f9vISwevtQVzufW+bDarN1ia/nYhm3CtF4GFXk2ilpPk5Wvnk4mVxkTZr1YlZOa
b9RJ3MBUW6uS9DYZKpbbkrkGJ8Wm3SioYj6vubxnn3y9jCLptGjCLVHGarVztxSC
VNFCj+h+i4m8lvy4lLeyj6qjooK2DzrSaNMGqLyfB9I7aoFezyBSY3y+INE+63BB
V73JITzbbGhzD+Z1opyWWagP3Ua8y3uOkeAHHeslJpAmfJoTFXK3XaG1iZgjB2m2
AToVEUFbWXPcMGxqOjU/YGCW2o1T1QVaSdDGYVZ53RzQQq6RJ0Q2E60vNZGmOfka
63mrh6NJAZrpMfeyigm4Wf8REZL/6GQSRSFOvHegBSNvZjqGHjkLDTlaVShme05V
Ppt5E2g+xB16mRWLFcTLKXv8rFEO8ur+cL0S22CspP2qpkXpZIeeIMQkUialJ4gJ
4nEofxYBn2nh2Q1waZ1Jz1UMckg7JJ1E6CneCjuQg2FbRlvTHIB/Msdw3yHhY7jj
h+9YRKc3Bn04cftD6BfLxYCPeU1cT6N66pnrus6qY85n0/z8XUemJEeEoOYc6eaB
Wpcsrb2kKp1F6XzZAORaxm0kPM/QkrmwooftJv4nioYwIxc87f1qz++b20LtgCC5
Az8Sl0uW4J3Pdqgy+VmHwDJZ/Ogliq2/Oca2Irx8YbDXoS7MTLIanPmIRaPPpmmL
VaPC7gdVEM36CReXCtepMZEbCnY7PasZN9p1/ecpSCZu2CLBum4yTKqs/ENltvEz
QP+SSfvgqN//MqQ751AvfHjSTwY8Ka9ABRrMi4U6RnMhlzPDtlB5BLWC/7FNU9HH
bRd/B2N1sEpUOWW+nDw5QkOMks+ng2RKOvdccGIXlT8jWnRKWsmEUWlFGO5Ivngk
ZISdisSQXMY2SJ0xMP2cWctqZChhfODiS/wO4akGfQHnLmroKDFQ4tjuxmj/VI4m
JYT2mJXwY3OPTWrI7EZICRBcmNbESu6PRhLnz4WWg2uVJaiP71z1b4ZX4VWEFS3f
/o4skT1qgGGGFwSIGV2cXZZ+cv2fYvlHQbPZoZvphe/TXGvwt4DO6/uIuZ8y0x4Z
aVBe/uNptwKXPd3VC4Grud829rppvTILw5miIraFuYqQIimmxSixOofUHzacGaxt
JsCIXWZxa6Y7KCKrVcEQpiwgSA43snCCyIXPRfP80zpgJwGOsGFWEC6l3jFjeLFA
5qbhZ3t6NqP5Vfu2e+QuWNbm6bp/Q3pHPLma4kfs9bYLI86wPSGiuPsMTnGL80a0
EDYzMGvGHLjctuzvMb6fzfiAB5HbM9USdQnBES/fY3h/0TacXUJ+qEuA1yfz9JMa
3aZvu/0ZGTjWTWActARylA/0qx01qEFOX/c/t9BYWfDh+EEMfMX7wZxkPBt3qAOs
O67pFDh0loJ6+xy2gvQb8cMNXOb13Nk2z/R2XzhMzQ8hDTK5hBwKuzPCS/xczPpZ
sdPF0MfTpQ/OR9oT9ch3/dtpRP6P1dPbOSWfdAuR+8AOt4cZjxyZgZ1z6hUlp3VQ
8eWBh6tH6zZImuze7U46eC5wS6mkc7o1oDRByO+B1B5QvKM3/9c7IOvkh3WTZ73B
LIoJB9yj+CBS4o61fcrfdEk3lXU/jn3EWdif/weNOmDfuWgAlxSXxgTuNrAuMUcl
3DuIfm6+rBe5RdpyJCuqdgCday9n560Umwwcijqm35QJzuPvBxaCwKQoTW1JkfZH
29H4YD7wTrf1LNV/R7/kUaF0ZLJvvVyAgExAC7bZYCi7FxDogYs7ALMxWhxlG40v
hraJrrNaddo1QKW+6PbN2ijVry/lD9N8+IERaykOFOnvq7t8SjWOmXmsLT390k0a
ASGnyWYbbFC23doO5efQOGmNExXm+VUB1G1v5edLDSDuUxoQPILXvoztk76hHENb
6U3f/vdgRori8aB1Ms6nQkemuIXP6qe6xRKA2XRg7DWBuICrYJKIFPPZXKuopknk
MadAW4WsVS1wcjtjw3T4NJ0Pcd+RDUUvNpBHJQiO4Gz5/DLkvOQTc0TVX+g8aWfa
p6+Eh1Pn6S18YX/kcUmdkdCN0U5jkoZjYEv8xvbVp9ay7R145KCc8vNfUc//Nl9A
68MPLAWyFwZVCJeoAAwirfrFNUYk51ekCEZuxa3DcoN9IvILpVJkeJ3OXvpqm2k4
l75rjgx414xSYag6BzO/YhqRzRGOyvdJAxmQSmzQwjU9NzZro+rZ6Dw9yL0mDyTF
wJE5Tt6yWXH/26KRiMDZi3xpSY4FTwOIiZd5RupKFyJDUp/qG80cv5LI2/aiSxLr
js+fUEEicqUmpaY7j+2pNQz3LSkn+c6d/C3klWNKhYQmuWo68wk+INVc5ZtMFv17
CnBuZIbh/G+vgCWHI05fefwhtreStD7KemXPms5jEMewLmCBJbx0YFjxfyVj3B2+
cI+36zfEkYj3NGB1lOrm6zRcR2TVq5G+DbRvukRQ3XzHNxHvc//hsEsBzNVtiDcq
pp7OmXPcmiRMU+G5LHZn95n0M5ZClu0y/so89WJ9bPM636+LlWD/denlVgmvNnxS
Q53WIq1Rczu2zslvblT5TIi026Td7A9ThBCWQ39oUN9TCp7UNm0HFSxl2abd1S5y
quf4plLDZilP4cWAHkckt2JIoOvYChO3DPPnMQpnHV9QZy6zRUi71vFSf9Py7mjW
uj8cc7hmf5ls8RoJrn0MOvio9JeB6XbVflJvkrJHJFFb/e6zg4dCnzAuEQS072jA
NViiRCrnvqu1G1wuBAI/qGWIeHfVnyMSYB3/JRIYsL6LkK75Y6r2n/plIxH3vWh8
glRz59PAaKeyNkzl+oPWWEf0Ak5byRWdkWYdyMd5RIpMY6GiwjSGywheRZOcDdEH
6u5aCJjZJVLhodEf9AeqheI/eL0UHFpVNaKEKRgPOcwyG8oP1WhyoxnM0ZaWhS1e
OX5MCLecjW1VkwUPuYThdFOjNNe8MAv7ffKnmBm2rc2AWKY73rl1M/KBZFSXcKHr
ZfTSratnSZI4Yu2GDThnYK8dHyYKihgX7Sljm0032DvfM5EdKTu8qCrWScvQ/XbE
SpKaOgj7b+JB6YGFF29aphmD6ndgRP/mi3mcxoip3RGfvYuElIYvmuHLZ1woLHnM
WohDgEFp5QzkvzOfXO1C4ok8oNnDxPo9H/r8GSCDToD8q1RslRgp3SPwkSU1aKSi
wNwU1tEHcmELhhqIV7X0BKA//963fBYRas7rVhOdKOl4XfNNGOjz7Nk3fbmYBTSd
YEVMmET3dWrcX3bIaAOgFYJYGxEUGhNFzbDQru5uokygZ+Fc3S/TR7TPg0FpgkQ3
vo6W6709eMGxwJQZKnNnRIpUV+3jC7djfqHb3C8dgpXxAzM6ZQTbVTQ4IaK3f5Oa
gZcO8Pqg/mnhaEQ7/dcFwsgnkKkcpk/uBm59WMPfgfhzV4nKC88jiaLHyHNh6uEu
DJUSqJSdw1EMBZ0ngvNRZFAOPR8B1e/IYwOgNuGq13blpzbz0zVh3rUe65iy0Rix
Dh2zWsg0iWmX9vxPPv//KRvLw8qTlk6Dnd4LYG02iyYU0bGPTkD5Wx++vc0VYdBR
A9RQwvCHgf0WA48Broe9kSQ/Wg4wSls879QKrYSMFytYAZYHdZWrx4rZ9j24AWmh
F3R97zFr/qXjGsH5nxIEU1bhdnOiiCmGQiz/Y9IZgmnGtCQZWHohKwXT+Xeta2xJ
YtZq32aZhrtuuhIEqmiC7gLQKdZzq2eGqNxom64kQOnvZdS76Qcdtzec6m0NLWCk
OxZX9ec0htoOGSBFjso9DpfYsIY891HFP53di+dByo2mCgGH6YL5nhlWa+xEMsmz
fRZT5C/CQ5FEY6I6HAC1jrAM0rzr0Nw8a+9kdaqMULas8hXJrYfIBGvTikdMIlhP
bcneS6t3ZuIIi5IESc5ejRUPAna1/27UVl90J0TEacqHxwKsd9iz1pCgXnaUzU/A
m+5vLxIEbsDV8unRWD7Y3rE1bNlHMrKmshuTGC8Q/YDHhoQewBNZm+CicS4K5CCf
KPba1GVpInZPAe0tO0vJRW8WnohqM6JgD6fvZkchwF2BFzvc5w2pIhpxBXiul0Up
n0p40vYwCZW/GjF/CeAiHLTEbW9d0ng+soI/iwG0f/eH3FI/t9b5xiEeyM0qh8gm
RQA/1a6HHObX32Rog9STwIWvXLpec0VSAMLTnHMf3ZhIY5xIbNsswZqnm3u3GUwk
Ploag4z6Cx11pBeo2VR0UsPDtAi5v7/ooOJwaA9QXEXsbLhDfLQHo3aT880kjtcP
D05TislVLmpNXKMsYVk+KuoQelu0NOPmT6G01o5NE8zlv+D0XEi1HzcRhzHqb+1M
sS10OINsEZzS+xcVRfm3N+i/kJ3aJzhpLxIGCU2ToTvtbateegkwG4hF5GRyu1XU
yqIFPBy1b65bs9vhPhCvPW5k1Ze7V/Gnm7oR+FwWBbfiBvJYGRTRmFHI+cyxBx1v
8Oh64Astu1IUZFkU8K5B5MUuaylKMHiF9v98CCBdLmgUvfjxQ+z2bpZpHmbPk6/E
L7txVc8VMyNUFvWwAB4KGtkAXs7Clk9u/JxhVaUtYfrDGQLRHeM4I32tFgr58LCH
ZpEPKtlWH/FT661t7IWZ4YDbOfmd0b6cIYq/0Tna3RPmDZegBk92XM+lCndE/EOm
jJBJIS2qbwMYZoaw8V2e9hn40WXlb0zzfBhy2eG2gi9nASNmz30YjPVKMIPqWhP7
b2Z66QrZM4Ns9W1EYe5Y1b4mGKlkOmOS/cvDiXKPZhQ/RFtCso/ueESGxEEdEeTr
CuIaDINBEXpbgUEoW9Clhkam2IgoyMNyfcNtFUo/n4wtlINpVNgezCkXe4LFOz18
59Ty6PZe12oaJe7D6kE38wwiy2LqFktA4SBIVc2EqPI6ThQbXI2SEUA14Exd3ZlY
3N3KbsMwXyQ+d6VmNtLOQ7COn2sfNuEKG6HceKXYVA/SR4u+cSu2VBVKqkVmNxFz
DZp1oZl3NMbvpg1VL57hEFr7HTXpSOhk0TWJS0WbLKLtRAQq7nR6I6Uk+imLHkAI
qBRjGwEhSFk3LwOquRdUqvms/SiCNw1bbvgX4ekIgnZXr+PZ/57s01xvY313LDIu
d5ZalSVj4bgn42v3msrzkpRxVnoISuY83yjLTdsI1g+K5gYrGuCR3FE3w4WRKcXk
E7E1iFLr6PZRg8jRXmN/1NvWqQw7/hjWRZvjmuoBYguM8tXKL7Gu7o+E89iCrVgM
+QZS35iN4PfXnHIibpRkZzfH9PqsmyUJPbzM8NTTNH7Y7QWKessUudQoo6k28zgP
ySdkjRF0m6nrWQmIMvIrY46luJZ4Wh43gM6vc9F/vRrjZfIIjI1ZFEqX3xVASmlf
NGb+IrzLNpQ9d1i+81DO9+AZmV44niAswIIZ34poihMy8kjESPqcr9HRbpQAVYDP
dMqVYUY1WhRU6zCQcJ428cyTX4SxfV8X7SqsWlwd8WjgpoDYcZwdCnMpv+2uSxKA
wioW+6T7LcK0zUW6ea19GVdeU2ZL2JWYxsvEcbtb/oGzZk4BqKvwI+9atTrJD9QW
VzL/iIAMCW+VJ8EQdLmOP1AhTtCkC3px8DwZQFh7b7BvTqhOPcSmt1Mo/i1ON4Bs
rRjYU2H1lHJIyHveI5cvHLfu+6r2IW5aF88wjbbc+tNHIXqyba33RQrGWxssN0Yz
zEpqKGv2YP0SfYxjrlZpDq9+euZv62tjmeqImxAkQNZHGQgHndpoH5PGXSllh8wJ
SYyBIwxLHd88JmDB/IaW+4H+0jmkjx6ZWT9Z6XtM+WtBujl0fHOKVaPXVCaYH5Ya
d0fmr957Jt/RzVN4AOVyfBCy3/JKgu6HDBSNt+scBX7kggaSL173MdWMGecEmMVr
AA+6pknAVzcbJLo33ahNTbuCafvl6HNjeDTxVVuXNUKYsBXRZlw22fa1mIfeNYxI
TtUyjbWqEJJmT6+tK9Kotz41UTzs6qnsYs3rSC26OYTi6qAF+dOy/r4S//NtCaDe
QeOAKWeChbrgkErwAZdS+iJaaJ2qffkNh9PB2C2+fc27m6Htr+KA9iVuiNVsRnsi
Zy0Ha7ktdGq87trTGaH8IQZaFVmczb9eSKYUAx0MCc5dYnHiKdrTwWnHKsWqv8wu
hbbE+p993OR+qv4qrkTlL6KVgaO6QvvFZq28h56PTbXJLhj17OwU+FcFD356iVzh
+btO8CfYuvVebiya3X4ugbyuXWKKZYShrrgaHPiBbgbXb6lqbCVj/i+PsstOkr+n
lquBZ3o21hb2LUTUULSyw1OkZqeybCjAdmeW6Mny2I7ILFZXwN65juvOgpmT+D0O
xBm6Q9U94JWwbuuq4j67OWNQ3cYYvL8rhMmHte1zQ+z3he1DDwuhZ+nVm5cwllMF
++cIGDA+U77pfirUOfOLrv/Urnd5U4MYLvqGmHxLfpg5/ySUpBTbdxpthU8kUpIn
Lm8QHVHpgi40o+djn4ePgPuAeBoSd4SbPzqzMNINQ/Kdk5men6nhgGUr/fih6vNL
m4OGZJG1sJrkFJSi3JyJufUxK5u5Zowtqfinz2THVieCV+IgtVnDJODbOOhXqgTM
NfPL8ygcPvV8hl1UHkJKKspjFucz4AJqOBXgq1pyALFUTUKRFyE4SmCpzgpo7XK1
E2Za//VEzAWG4FiZLHQGK77P56gPiIRt/llIUE/30gU7lkHlRZ6VVP02yhP3Onfg
jdrJ672Nxpp4PBUppkJabLXK5GLcRfjHK555Y1dmUiGGSmsjxLeSsgU0xetr6UTo
sNr7hGiBT0WlUWzzItMKzc2BmBT2NJa9R5BK5+/2xvZ11+gJSnycYyqwYGraqS4r
X3yVtZzxKOi+8UfLVaJclsxkUShjwfalEfENHazWvbxEoMBBEvy730MzC4fpIZYC
YwbyvfP0F4jMWOf022/tMnORkkup5C778ozIUn0LcgTyTzvLVTtsDBm5zpYvh7ir
I2VgwFPM/Eb9zxFokHX4yeVEyDWeax3F0y6A5J+9KrhjTC3uXzT4K5JkaG+12Ck6
k1P6B8MjZY2MJrK+8hCXXmoDX89zwxfvzRCeTcOBw+a6q0yYEv/bVpfwHS4oy5N1
ZKY/+1DE+gshjWMTx/z1mgbPIR2HjlJIrY3sGpXiLcMsJX54aGCxXtr5248iGXOA
MGyuy/pl/djSMFHB5/7J71X/kY2+JjBN5Cc+U7H3PcbagrFb1Oi05Mb1Xyf1qMnf
lK3B6W6Iv+zAVEg1KAp/CsQfC/ukl+iGK2T1AEGlNEI3Hf+K32ILbQ2ewNuhkWWr
sakHONvdzFDbiUSn9S1jhF9OGtWrc0llcP4YlojO9Qeb4NzmoUwbBcQT6xE9kjV4
S+Mz+Q7lGE9wKs4ZneGOXQ9FIx85vTAstao3A8RWjIGjyyueSR1zoUCXGw7XZmvH
5Ev6OvI7Fp+iqrM1TuwHanAg+QUznQgWvkdgatmEkQsxAfsKGmWk/ziJTEYDnUMF
wosNzIjEpp3VzvbDlLBdmheEcvClvSZAvQfI9TPzupqU05cBGncNETxnlE9DXnQM
dig3FKGT3hMGTJHt7N5w7R/WRt5WPmdGrirk2GROqba8YnEO6VL0lemTsU8JaVuS
bE11jUPicEDXHTy4nQCBUYXAOC7eT6LuF8aVQPRvBPfww0NkFYN4PL0UdsqO/9ox
qId2JYhfSV2OkES4TlX/uPOSeJ0uZPIHisBPlXIl8te2f3vxiPdLjqbDrpnUHSUp
YWp/ncKl+P5Oa1Qqbc7tx0E0ZqmrybLst2okOQwlPN+A7w5GzR64Xkj/rXNcoh2+
4lVEwI7vUdBKeCZgVPdrgqMl0NH8gJwIXSp/BeIsrg2+0mkh9nsmHvyLEikEYMD2
RHanUXWys9nNSNZcVt4wY5nwiO+KNkOLbioAsxbTxpNwQbYBFE9ea68AqRnxXjtR
5Jf/aGKEVZYAL71Vw32UwEWLnc9wOOgMlut73FuI8BrXKkR0J+tEHmb5Zpxo7wYa
8CvmNEPbd4P735BIwyJo6LIP07KBqzkjgspDbkwRgvMozcWlTVFKsTsWS2ZN1RZx
NdNo+kg9F3SUpPtG0JznPt6Tu5tf3qCHzWc1ArZ062H5Zcr0BjDnL3wQYBaacDLt
juj6t5Mrl0o694jGZiXvtWAW+NUVg88pxey4efej8+RCRtZNTOizFqQZPyefjLaU
CyKCW92eIIufVz+nJAeCziRkbNVgopp91OrDXEvIGjBI5Rabk8rGydajEoDSOBrT
sw3l59fMuhpK77K7+BmqmnkKtjqpC2f7Ege6W1SOUcGYEYXL39v09v3IGlQ6PD+y
k9Hr2AMa1j1RmTGROPYHygIrsfPbuL0NALRCD2WjH8xEKe+f0nZ5dK6+5EXcD1vR
Iw8IJZKPNqAd/HpyenG3nKPjscksHx9Fr8lbA8V2i1rjyMMV+3ixv1PTTPYGW6jd
xV2tnEOyYrtCmFPMm43eDVtSrn9zlI5LXVnY59rtdjvaSNN8dHPtAMS9femueZVd
KRH1XVDDz54n7ky90ajZPWQWVFDMMi0IGfQQ3UefDE/EEgUNzjZuMKveuPMdLkMg
HkWu8dxVd9QZrVXibwBMRK1w81bvrSRpDESkeS4QU1WrOrZJc7dKTaih6/Xtwxmq
4BxLmid9+3LYiTR4JzFrw0DP8JIczCM01eH8x/FHt0rJFU+dPb8+tCviHsEihkE5
I/sIIgoBtBbXKZYCKkdnTcLdmO//7ws/jlUSAdhGKYgW7KKIcZStIDvwv5hsC40R
+dQThy3xfe8lSI90He+Wh5hO3VkWTkGYFAmsPu/1V2L3+DGznzbgYoXyHeKJU6xO
BgY8SWVB3+9H4fIjzXhavqx5CcG9XRo36HTukYegh3rJ4RPTgu7sTVHJdDPyGNN1
EG1hiqKZpXMGGs5kQzTT88geJ3j7CoLqOckU96wB9QC2tavbnU+JJMZY6XgRwkWO
9Y0/BfWKTVTp/cqGrWtbW29B2zMxxtNeyssFAPtDfvJTRX24ckjy+qPfmuZAx+si
9oheQLB6uiVkDPkJQkpxbnCi33bqMXWlmlat6jQiVICoDCKiNdGQExTqJdpgY7nf
lUOOwzCzpClxMOgDof8VYqjHAw6DKNR75linW658Cfkk8RvBgh4d1Bs86aWBGiwX
3PofIyhsLDuIw4FjpUT6yIc7zu3FBm8bZiqGoTiYSl+thkYq6naymNWBicog4yeK
iHk+fit1wP77WAhlcQz2UD9FWzhi7YCtj5JAhX6Jh+Zp17RUUoku8MQZGhzBL2pU
7OJsSpCTYpdg79BV2qa2poE49+nHk5Xq7zCLWfVeqjagyBGL4Gera+r345/QUFUw
OkHVep6rNqzivUzA7LKLK+qCn8thRyZqWcqeopURxAkUZDgI3snftwBBALxMYGAt
gp31XAwTbes+kWpsWZGKa/DtFO75jrpyLYIqw5wVlNsAT9EvCG+7baYbArVt+4T2
BbKz6A3z849rc+OIVPObI6G1HDCuxIMkgdDpfdhL8scvaDF6YbKkaFuB4L3r+e1v
ZbSk01JZ2VhlMMgz/OU007HO8QDJy084HL/AL8dfVb2ddPVQ3f0937MzBPsk7yVp
ltQ2fRM2SZ1hrzN0VOzoGKLUreXfuvQC3tYrs7nhFzXMRgm4AWzOWC1KN1RTCux2
MhXjl1lC/9H8QFE8hPXH/5os1ztRW881Yg3ifoHr1IJ6nizubmxQU0L5WC5UsnpG
p1C0NfwZWgZId+RmRIQ0hxhCNt+IMqO770V8nb3hupOFI37xqBQwu6ZmqzrCapJ9
Ojxg9TCq8MpeGTGcnYHH1AzO/0xT+57ElDSYKkAtpeR4WvXfnX0dEFKvuwarNZEb
WjhUq0fuKkiFrg2VlEBxAQQKbV91BhNCVfM2p9BpdRGdNE1rhuELVvT7CeK4jP4O
N+sF29huP/ToSfqPSkfHQGdwDt4dv0KjhaAz9isO1ZrJSV3MUX0SSy3b1BJKqtO3
ehYNnryW71CBroZIdjiglA1J+m8k/EiFfDh7hms3yOfjAXQ0BoUyiM8QzcPGGNES
14QWvVVfJDkPyO/f9iVq6SxNfzNfq3ozpyckQcMwijeAsBt0biIe5gZ55swXPz2f
3kC1sgKZFxW76SKes3A/qzFP9LEvW0zl/Z7I3d+9abhM83wOyOj1y3ZtcWrEJcXE
oQ2rcHr+QONJISn+AEDjp0G34PbEZJGhpbtV1O7vamQH+gKmMXy/SmAeMbFvo36r
MeFFz53I3QUl/pd97QTOY3DiQIl75siJHi5A2FcMfNRaAckfS2cl7CuP9WH/6hwS
93/bC45oAw8dMTBS+1o3lvy9HSJbqwSSVvunMAmZEgyKGlrdLHSNASwznLg+zVsB
a4wfZIeg/IOKWg0WRs28Jj6QukPwdVUmrFbSUQ27QxYHtzSo5/x6LLMqaybceFJe
DIIpDvalB3lOz+8TaOgY2huALihHByNp0ii71l6oxQJXrEqGZS3PF0vDAt+ZpvkK
HEO4U+klobHiVc6RzOKNUeXG6asO5sSsrBErsm1hHj8VVtK3lIiwADZhC2P2wS6Z
zQUF37FpJoDQ8kYjXJv0xLAuXaPlGHmSYBC4irBTZgkAGJFYVa6KUb0WjbH8tG3S
Yv1otfvh3HajJMwr6GdWp/oC7sZV8arH2baR7Wv6GdhZ2tx5/5uDQ9ZDdSq5KOEs
JvQe+m0ZxUvJi7towEkLg9F7IvFzeKvjWwxO/M9d7Is6CFVNlWmJata4hQnp5Hxm
JAwEubVPGOr1cRuWmORNb0SkoHvLnU8+Ro/khDDO0NISjyZMnb+6QwvEANxRuevd
hUp3oDg4n45H+KtWPrcmqn139cwZEoIk6Rssn/5pyp5REhG9amLrMvYa/2iJb/wb
4hs1dVupjeHv+pCFwux6faPE9/c5Cr4PMKM7+sNVft6gghkMa98y2Xzolv/R9vk8
X7ZZjvDBDFr6oKBpoIgBl+CdhCJqO+pXwDQCuTG8qAXINbqZBRcfBHrpQZ0i1NYe
gvb2i2qh+tRFm5GH4dEg9r8G0hiLuVHREpszUlXnXVVlyah5fJ+5BZks+hIG4CHS
hv+eNpGpN+fK1LUET46uuSnRys4RArnK0sGqTao0zl9+8Bv60jxuNmeLS51MpI3e
ocV7uDcIHIh2rDyygwqdjfGzjVxzJj0qwStMFouA62/MDI3FKIu4MlhlDLaOebHE
1IEkXQpnTJzEBDnovoEfboroC7XyJeV/DDHcO49wzMKhgrRCoQXp9dHcbgBXAAff
+bXRTK6PAjOFQ9OX7fvU4utw61IcEEUvbgzUizNgo5SvW2+RpFJewN4WwPa7fy0e
8revLaab2cOGcgZ6NeOWFIsNs5BKP3INVwHRm4VN5P4RoAeumPGgANrRC/48jxJb
FEkxbJS+7Gkf1KcFnk3rIcrZn3ObKVYY+E0aiNwCJ+l5tyPs7wuMvXbNxlQTVgKn
Q9ke17cihPGJ7p7lGKVWXp0svWDKhECdsBU8c4r8EyeWi89qZwcyoQFzg5Dt7MFN
WZJDFgoCXzoyvpdZSWf94poxGo+0VMiTkifr+6n2L/KaPzk5TGjlqXmA8PwIWvY8
qbFZ1N4fb06L24WKkU+CUy2M/Jn4VPrqVjcSFsN7tuiTcpCtJTWNIfQZ8j/5SQ1e
Qd3NlwOzMDKFQOgLZNpiWsbUNTSo6OfvL5EiILclqdOeNx3CItMiLDapeSz4URlh
Y/8BDuuQe6Wy3u+FHxOomujELV8+xHUidSJGLiLKO5yR6g/viRlfN9nS9xLhSN1x
Yt4HbJIhKMl0JRP9ypalox5ezOzL8smMLEmg4jgWOcWw7/hpxt6fzOTMeT0lue8X
FwV/CHmsTVKhoIv8jGbvHRIkwexz18HH9RC6cggvMPhLchJToWpRTBg0RUaQ8ZRF
0gKzq4C03uUJfcBFh/h2bJrPSbs+K4K+B9Mq/STiIJ/YCGm1A6sB1qa4b38KkdPW
USks7HKXunpv/o2Cqr775UzVtqjTbtqTmWiA0pyQj0nijIwrR1vXeUK7/6A25dIw
Mue7jcqUNQZPWtPFcec5czlFEHKWkIMUFsmh2Ine7RBLh1fuBLZJE/HlG6vCYCEO
kEsiCRAMT8gLEIIXpQcmU66MXKdGmbO9OJ/qX2/BT44lGQsp9OLvxTj7ROeAvzI1
8bRYseBfJmXXCjSM1ri9FU0LSIQGvwkwcWdSwhZYP0EuuXAsAlL6kt09k/4UUwIK
N0hVucWUOYX5en6JX7DDcibuB5IHx/NKWgcu+dpLomotcNV6Bys0qkAYLiyplXmZ
actOqp0L0V7bLNBpsKxiYQZ2c1nJ4K26OvYK4Vcms8VDr/K53R2LGj1gR8gtooJa
YOjBpcG8DZcjKu5tjEYf/i04GpzYp9KeBHS4ePLwrTDHf2srh3q64pDaSXN1QWkH
SWQYIMgEXPdQWg0jsxRgY/usrGx4cZCslGZx4p7FJ+Lhgwmwlo+j9UzgeqUy1u/l
JweOdAAhVSRjhi+eERfiEkwMH1LPXUR1Hf0Ul1TOPJ/e5y3MHi7CINfojO/TBwhs
Pq70P4kvB/G12s5Bu4agpCuJCYqzoJDxT5oJNSbHwt+oHW/MimH8EFb878JNEzUC
3F8tGCme8vMLAq5lzoYW7P+I28tW30KgbSYWCNaBhGXVDi6t50eH/GoaAHmzGHyN
aDVWL+z/mBtRugbrenO2jJo42o/esXNJ0ddKKFqYDnfv9LmeY5J744VL4/kFdCgz
j0kRQRSBIkwgLcWRtbKtSz8oy8ps1DOmfJJYFdyTs5qyBqbzXOYgFsDPqZEuGQKN
LlUgfvyRfaaYIzq1Ufv7FrL7PHc9NKG/J5CVnFdbP5ns5GQTgwfi3vwbBzP3sSTx
trE2/40+xuCNc5z9pQrig9evmxSWxBasxWROdFuGVAva6M2eDwZ6X5qTo/aVKAKw
kzS7Alw5i+XVj1bUGSv5v7mg/rE+FecM6ymqDvSP00MMyac99wofO+z+Mwu4HIjq
7XocQjolcJSobEjWJqtkpbBex2l0nKQNDZ6CIRmpXxoDBk1kp9X1jkE+QZVRG+6I
uCv3AuZ/pMKJ1u3ZsnjUc3qMAC2BfDgr97jQ9mlhZjEmiikQIz/g4ueUyMCyiHzC
tIZOKDtWqmCmK8QkYeu/W7gFlImALbzbsWxOxznyX7pGsdzgViXkjdOtFD1MH9w4
RDIPS1LwadW54Tfx1sG8u6fwQW2oeeNqtDjlXU7mRdMKlkjLJ1x6u6Kera7wGGkL
TnPDxJn50tY58B7eFlBQARbl9bfRCn2Tyqi/tym4zwmC2ns7mml8v3CojEzltQ3T
5QQ49EQ9RwEqGORTPb/dklYskpj4Q3dtntvodDGcyCAZ13A7W97Au4k34GKelM/o
SIDk6eINNT3ljkYnDMfBn8e8aalunif8IQl3gjTMf7VJTciP0UmyWCL2WEQP4zb3
+8A/5OdUlRoFuswK9fVnn5PH5CpuU2vPGLAM3kWXUoiwxRMkqkDKmdd6ZWdIVNCP
ZQRsbo6ewA0AMWgXeuWQo849RJPpKziUOmMXjfrmIbLeJknF6+nQwUGYwdRfZX3M
19Y5N82p0aXuLeG5C2dawupy9Y5Cu+BALBshzfN5qtqGoKNwv4qzdsHT/AimLdnF
/c3ylWelsQ3ifgp5he5ML7X9/b6D00s00yV5j1Ftph5FRVZqj56y8NZNTn4j1ZK8
BgaqoJCQeUD82ybnvB6MSpxY5Avmcw7r5cwrTqWsNXWrFa1ZZ69RHl28PYyxJt/G
69dhxWsSsfw+XoZw3VBeWVCgN9kQFiBVdcOGdVzf/CXZUvNocH1bxORN9xvCaS02
5UBp1SgeR7gRyim/3qe7t5BVNc2gUZqdi2XxILm1HGTCvddtAptQeVUIYdsOgGju
wSfwQev3v15iEFjTvcTzC4/zQo3DYoFexVdcwTKAjwnlOtdZI4BM1J3KEPdQ83gt
M5bBrry8gK6PPunzJko/LabMN7TKZPAbhNn49iQUd5XcctUTs4I9As2hdUFUKjQb
1ECUEwoR29O3GkN96M3oBATrvNkAT3jnAQE9eImqpxmhe3pfcKzZVxb3Zj/NErOM
/MkoLNPukF+qWaqIOCzABafXvk9iDiHHdBZBGmvcnDJxpy1PNaEB8LcyMsTr3oa5
I0wcVmX82YhJWSHIlumBpBXtA3S5mNETtf696XODTmlU3SjSUOFN82wBl50p1MTS
k8t2k3xbA7yNjh9qdU0D1XUFMWVaulhC6omeXsYRhEeU5ilZzgs2qJdlquqIpYY2
MllQtF08TbLrPeqMDW6OqJWmRdhVwRAQJJuJXW9nBIQ7RsOrMqDcBBS3SlGVVpfF
plQRSksgZSVamnf23+1D6lrovxfo7azxNT4/xUEGEACSAX//oZJ+F3PWPEMjS87V
HckHElA+PQju8UMC422fXco4Xx9JF6lU/C8TdAeZa0ZBCt/t1mdNdaMElNqq4BSy
2wHww6i4LVp3rjjOrXaT9J4I6dv3qhaF9gYqz2Pkx6lR/IxfZhtcFoUbgSJfOzPB
sK9aUb7kufYJ3VUQAFJQJEElcjiLbE+Ol4bpeKr/pyP7EGGzBRvMviKu/6KOeBrH
TRyOUFidofa3LPtQyA1zqzy/S+vj7FNiOonAIWcVxXRDzjQmOfoGJl7ef5nAfG+h
691WX9Ldb4fKvoUipkCAG2CrzcjXreJqI147aAQuxIy4KWUVX7iRCho2koyTc45E
3AINQgOQB8VTRcfWW/nxCBzvNqRHkwa/Pnm0QPNLbREI7EHLC1gyjil315NNlopg
PalYNooA95lCs8TcRW+z6WzpPeHC9v+L7TjhQnNHECN1V8SFGsSgvQnZ0aS064nX
6KF4HU/ZskJv9TMPcZOwGOMeBSxEmjX22bim8gnt2QfbecqezK+Y2xuZqQF7SjPp
esfuozS8c/6jIJsgO+jcc28XOHSZ8b40Yymc6cnJkv3sXg8b+Ap7AmGpSmsfDaAj
L2L6WvuwXl3Ms4YHCUC5hAQiEy93QldOnoCNEmujLdbA5f8YIKq/fCCc0ElAxrwz
xFhd4zjhpzKKFlBubfKisxuUBAt5ViKq2plBEiTUSyNshyBKXEV0Rp8pZcitBDmZ
VsXSvJ8+z2+OJXHIIjhR2Xon1qIPJHYUnnxg3yuUlgLo8eQu0sObBD8vASTMgoe/
oD+PvyLfboIUt4XKnpIDIV76ny0aJvBPV1XE0ogytJzwaDB8sHvDk/U3SpJufeoA
GcxKWj5oPeoXjl8pOFnyIBFeHua00YsdSc7QG3eOxNuC3MeIL595VO0M0wPRUtgB
kyQNv9JFsLLpa4X4BgV8V9yAZw4Sg6r6J72llwxlA0pnFRmwUuFS5Swsfot21EUn
mno5B3o0XFofGMEYCIOV9clUuQ27Fg/g6q2PSXeeDIrU8wYEZp7NSu/EVOoAHsGD
o187wjDHuzW2Eg3L24Gsm/x1vGndlOecmot9nP7vnWzy+2LSTMcvY4162DBJt77U
Aq/JRNghsNFPVhQb0tRhFGgkJ7oRz8quSVaSOKs2TxhNthP1DSgc5rBzVD49iLfG
6Puh+9tyqdI2xZ+iCIq95linwSJYGy3gKKOM7TbotIfoGEV22G3v+mujEaNGF/nf
JSHC4sMonuNjAOimoB/5W1oFp5fd84nEOIRJWb8+yNOY5LlwXfhIt2t3X/qAfHDr
EM707dMvBpS6hSXWtoEQGgJofQUcPFEBil5XJZCEm3mA4Jwnw4HlNy6hwqNxgIwD
35cqRU7RX/LdW/3mjNMuYlIVCber0L0qRdobujoOl3ZS1HWgKbBjoDVjQd8MChjf
n87siWIYHpLMfKVsCvbh9MD8BZFVr+JC8nlk1RTlSmYnWVLtnSsMefzVwElijsRC
h0dWSDkh9UzHTjGRVZnexw/IGv5+iC8BpMojpoZXUBLh17auD/B83pzhiSCiaf9z
y7ykK150w1gOqj/ISQnlgUSj0vDztxZqBnppBOjuChhM4qly2qPd2UIK3cictb8H
GI3A4+Tso+dTcCsey2W0aPLotJ6A4UYvuSkQ/zy02phy+NgmNJX8JG0sFWXNFg6v
yZCO9fUJI2VaZRNIdEJM+zKGHAAZ9cbC2jsNoe88GVa7cHdRccE1Qk8VBdsrgyy4
fwlN+ii1GR56eFNQls839xURZqbWFWjwO2zu6k2JLcyuPpU9XarJoO+HzNQ7JNvr
oLdRcfw8xhtctDeQw/ZE/hHl9OskopyZ5kYurGor61iadmrluOqkDzLFz2RKnI16
TsIyzTX+KJtY7O6Aw/eGA6QtVOMjDgetHEgVLN9xFWlMTu1zds2QWwirxv2fAMU3
3MMFoCi/4Ej5DdIVn7hOLWsYem6nQfYavspW7WyC+5mgbG0oBzipC54yjQzg3LnJ
ufU4KhJcHHWafG9LYGBI3wx2GclGfFlaIne1S7ftzK8uq4YOEq3lhueUou4YhEUu
Y+B7htA0XTVwW7iTfKjV2h+/fkoqxM91tJ8d5VnySrfH8Ajivsl+GEjpHn2FZTq9
/A+OIDwqpd1uRCTiJHYiZXASgCFKGBzODZ3PPcIaGoq/dKc2n/rU5yTy3OyZh4Lt
s+3CGBPczyfmAmXg8PVEJV6UuXe0eJ51ePS/6TIrsIqvP+3rxXJT3BOG3+s+UJDa
lhAMS9rV6QJgtMODp+nmr+J7Jda7J+uYNOG3MhMfE0svnSyAnyjN4OKwMUVksB2t
WkrxwRsfo8kbVxZPTVyrjohPlwdIAyR4b3arbPnanuBAmEXkuy5hQxA5oPbnG6SC
iwM6JtTnVL4K2IjdW//Y56AnZSew3pJPn0Vk4d1zGWIUHAlzlBOOcGz4Qvo249qY
Pa7wbdzaWj5jS5oCT31lE4vhjBaqzAXB6ZYSVn8YMUo/KKMxnQWrO1PXbSA7RBHp
FibVcoxgt2ynJmxmqtFJRs5BTR/lHtfrIJ1uSeb6R72fkJMETBK5czZY9wSvhhRL
sg3QgjAmjJBO5TIt7dJZpHHgjUl/qkM+vcN0WdKk+yeteEwT7jv8q5aG8oxO5Nvo
08zo5f5WeD9HfYS2yD54zCJJrpg1ZrC/Wv04bhwlL2yybg0gH1EweVrMCclPurCG
HgsgG+GC3MvnkDo8CiE3DFTuNOtUBCaK50D4mlR7Eo8j8nRWooQKJh3ovDPQQK17
HBicCdx8Nz2gq0jCCqaABHhblnljHqv0hfYbBP0fI8seh4rnDE+UHa16qGQH9WFS
YDA+JVTwniQN7rvGi1MCiS6WwejPeAN1XVOALS+9nn3QR/7IvtqtuZ4ASXeXtZ6M
uM7WKPp1v9ERB5olGh8G6gnUWCYV3qbadgfrFjV2dQY4q1wkU/AksIRLkzPJGKA8
uItT1sBXMPYY0yLZWtAC17a/IQAyRfSP85OjikI5F2booGX61xuy8ASmxoRgkIgW
cE0YquyuPRlDL8f6sumRak0H4FXtI7fr3FH2VBMNNt7fcHsj2vBChvCl963RBTy3
fPhuCFuLqs2RcrjCYkTFJoDHB9ccekY3CXBbJxCIaLA0ugzQU+71IFgntfQ9Hf0h
iyGc9ZALHcbXgaAAZiWebAkYLjfKFXkCGRvuynpN+zoYwdlDIG9V5jGnZJ6VyYyq
tIc5SYTv+AsxW/YZkA+NOnLW2E1EIr2xzBTSkKS7cDKCYq6uPuotV3NqpVLxnJSB
X/TwJZV19q+l6KXqBNUV/SiK9XNOiD2IcR83bmgY89Ks3outkMRuYruJT4hhTih+
3JKC8mtDqiGHOaHfNuALRT/OjG6rgoaadfsd9Et56m9o0mXGp3FN8AsM1jBunbim
sF5qTqhP1AzxkN3xrOM/q3qNy17jvgiLZFAH7LrZB4Enlzctm2NzeMgsHNg8X5cp
2gul3Xacgu+s8WoaoeTOeQUzdMuZmHWpScAZzIIq2htts6hx19PLaFVUl/+/p4EO
b7SWYyBndHl3m856hafiTnfJRCY3LssCZTl+yuhE4LbtKCSswDN2oeMwYqxcH/By
Hc4hbxqVDkrkXVb8OLpWQTQ0CYPTasV/wu6voJS9DKdniM0EhTJYTQUNyhJoAbJe
EzVDy5ZY+0RDfovGmBongXun47RXh1ftrKSAFWm+Xd/jb/Dy8y4ae8WLz/hg+43t
Rlj0fGA5aXa7KvEWULlTqH+gwWgK8bNh6F4qBtLWXl5fiOj8UCmUfPX0rMERKPj1
H1PVkW1EBjgTMC5vnR7pHBQFYodka4YtGcC4X0LTIVRTorLY2R0fYeT2ea7Kp9jV
9Joi/Lk3WvEEGgA4edTlz+/OdlX9pK0hDsx37opqxFQPoKBt+R9TTX2Y5NwmKoRf
C5aShGERhLsmgMFWHhuDn0i3SsrdEWNwl6+K3LTKbRmVB0LEYRi0DKMo+zu7fFL6
rAj74H+kGhEAxE05n1U5e/31csKDQ3avJEoHke392apP86q0bofMFFRwUPrwpWOI
l7AB57GcHqjY9jSGzznDJwB2BuaI/udDsPujMK0Z+dFcmmF06LNFbFzxZkgpYs1l
RfkpXolFsI33PjD342Chr8YzBjkffIw6n1fPExrGFHS50CoXPK8o8hdmdNULJBZw
3AsVE7OYHZlXvAmsFyUzVY31NzA6idtW5gwQ40ZIIJKql3cYVsiIPdf3dA3YKs0K
RKIseU6NrYm78kQplWW6VTNspU26sLgoqxWKAvdw6ZI5iykMGCOGHdfyzVe2bYHx
XBEBf+g/ejKC9LwFtkWovFJP6Yz8hf6uO0b7WnPZDL4YgQGVYOvbP37BczCd7qQ7
D7WBgBDRssErIuF3NO3hACw+mnGBldKsNAPnp5jYWZRLM02TdTnsMqL62uhQItrR
KGY4q+Grcqc46H0q5I6mXWT1mw2wxHWmJUxhAUnjO52h6r0igQTFT8Dwqbm9rE2m
afjMDuX3+Y/Eo6IiCOKMVRJq0zYOO/KkatxAAZtE+SeHQl9qgzJjay3JoznWH+pQ
Ylx4OU4AmQP0xeh3Rk7BY9K1lo1HdIwFG9Z5Jvb67KiV1GrlLAOlFY4+efsvmIIn
tF0OmF/KO+7bGqLnIDDQ6Qg0oUq4jSSrJQCrbB9690tsa3MjdpdxamqS250YKtZi
zr7Bqk8BzkbFxnUFvX5Fc3rrYpdF/qivSFDnrJqiB/MP16ItGTdL2IxcgEe/e8xQ
e+ppXb8xU/9OfXCXDmnRf85uSCwEG6GVoe/Da3Wlk6xcUT3/UIf8QNNWWlDcIZgz
Tf5hnyEl3Fa85pcfhYP1hgL0C1v6cWZUTsH7akBH7USEXhDTE72ke7y1k6J77ICT
Mf9pcHM8J6PyfBXEBiEUTnMJGYdddlavlXA4K9GhJ3C6lozx7FI0cIMrUzTdvy+n
9Exz0awBIybMtWW5MYD9ZDbSmpZbfqsWft7mnMQbxhjX24e7hsxbUq7poII4qD3t
6XsGR5CX7CsZKzy59r1EyhfFOKH447GpM0yKFKRIQ5PtA5aKKLAnbFq8YKmKWFRp
yy/l/8L9LXnIFsBvOqFv0YdGeLFjiuYYOMpWCrLo8JSsXLPejKYkJ2Dv7Inkjmnz
Wf7ljJh/CdwS9/esrtrW7Aa4PSogv0drsHSi8iUv63ojIM+XJf2CzAP+I0mo61Sn
P0WuV1RWguEbiF3dCuThplM1PKoOcyndpGfalQPRYyQ9nwI+IjldwGt1T6CqPGVD
IounF/MyRHweEc4wThN3JaksMi7lzv1mpOSIhhFShQ55nC+2iTofMVR5dp5LYOvO
MdZi6PI1s0S5tb5aa9jnYc5b2EE5wCplWyuh1LuDuVK3dhCk89WiUhqf4yPXeCZb
8+qFssgZb9Ex01mufn7DDAeB1yIHJfA9mdXTUOhSrZrPwamYiTqZBN+wcHqUKJnL
WA7K//rN9zn0mBcafhaN3G+MlE/EgDGkZhpKBU4Uef9je3zT1XLdxp/E1zRA6ETU
bw2FteSZ2/Y7LaJGAH33BvSQVPWSdbycBqgaUmtjDYfWL9tmDofNychJwdfDadL1
evmm4AOKTryJI6mMcP/W586Gw4ArN6Erj+3e0BgbI8aTv69m6neFL9xjuE0Em4mZ
fcyigpn89+L5o6ILz6fSSmSGybl8Nrhj56B85AZys92I6UISzEDwIsHyuhi3u1Xj
RhBR8So3IUFoHNIrt8SB/1uq7I3MKtEbYv25U97/srO0HrAWD8k2Y9UjIupWiB9c
I6zGV5fUp54Us1eLXLlDrblNF6UBcI95S8tEFVVUDpsUwX6bFBCkLJFU/dZIL5r1
SPevraMebHjYT0WYSnxfiIyQ3/H1jHTg5BLqKgBq/xlbYEkWWM3A3U11wXDbj4O1
BBf3meNS/lcBVo+rnXckAt1mrscj7371XPLjRUnIizArfuyN2PoEcnsFkFYrmhTw
UDsyhNFadFlnRewgBZ6rPTIz2Z0B/sPn5koPJrhGJz3I9dNQfjkk3uux1aHRQlGz
WAvZy8I88UYGNcygWL9T1tBkahjkr0UcuPjzlxahsBa+8dzlJn7ddFY81gRKtE4O
xc1GE8Pgywz22jEeKf7JcaXezMBjAA2/DvehIdkJU7O/1hC8wzFeMwiWsSBIULxl
+WBN1IYX+vRGEA+l9KlX6cpP+DcXbz/ocXmeQg3Sj/honR/BYtFB8n3b8RuZOk5/
zDLLqddRQCKaDTos63jPQv5pbos7ueEiiDQtEz6gcUZhiokwiqrMglSWSE/byo79
NbM7gnkrgJiLjqIN/KyLWGOAJqMFygw9YO5ZmIMBzNmYXbieVrzY3zFDirjaUZiF
mPDRiOiLWqxCmD2XY8xIW7NrhpTioDtl6nEw5s8I0ObXQ8PZ093ODqjFIJ70Yz4i
XxlJvAwQE+Xew9x6e0MjluMuvJXTnG7mIWO37Asn0/X5A0G4I8TSDHn6QzT72XCJ
uJYCQyV3F23riIM+WnckG+S9e0NcOM3pNyjrgFlk3SxF9AuGZPpIPbgzOaFbonYX
xCoq02RrKeuSZx6B0sKOkWcQwE1btPMmWfRJc1o5vUWAJrBg6dorMT158t/A4sWV
Taxx6VM6rfySitPcFxgoZrRYuOCru+Ds8EDWVi6gBQcnD1H+fCBKOOZTq3PPyrcV
Mt4b3sGifVdvRCF7k9j3aBw0QEMJEzSOzKf7NpQYMgzpzaKujU20r4u5NMLNRfef
UyXgg4i55nTi9LofDWm9Fno1MD9NvC5mlT7Xj6c7+Ng0ho2NLa1EvUnuCHm892SF
HHvPzW6u/OLxH828nirEs+xLazSWJdEC14DsBmu4So607GsewpDhFSULt/x066lC
ToAZZ1brmdaMaJH39DE8hJ9jyyOU5RImIJH1jQd2xQTPpm7b/fFuaXJWRdK+I0kX
jgrHven2JpoWYBoYy9h4LH6ggbo6g6yWEWy8pPjp04Bua4YIAS2C4q/8LyulzNr7
j62JscpZ9G7Y4Q2pyFUQMXI7dZ1qRPZnuphQW4q1oGK7faX3sHOEPGXzwMuTU+Mi
QvMTeoA47Fqt6keAWdkv1ixuUQNLXOtB4vMTPODO+hFoDz44mqW4VohL6IdUTeDI
YSjscDuV+eMy/70H8JBKIl8LBFle5j2FgSh9pwST+41b+lAuY+wLqT4fYuqI8cNI
3zWTxg+aNUObHhLD6bH71P06J1Qv1o04D0f37y6t2Ce5/4lnBn7YnyzKC1J1OA49
qpv85b1eH5oKrfAEuEf5bMbjqhlvGNM0SRW8ja7W5BauE9QoICD0FXF9nVkQsr5t
RU35qD2eREikVSL3utDErwbU3dMrV9PTH7MHLFrcPeKW4XjRbW/EI4vT3C/Vfo4q
mmToDtmkcWPQ/GscVV7vXERdZb6V5KJFQzjq479K2WZkfGv+FYSlZ3H4M44FfwZ2
LqW/7hZgFCg6B7xAcVfspU/RW8fnC+jHp5p+XfYVoCln4g+uIr9JKWQOEIZv2sIr
Sa7nezDQZ339ENXAvLfQImAj6k99a+zrsfHYjCU2t2rr+ZdZFL1TtvdZvaaWWm5M
KuOgaRWzGPodSJsjhVJ0Y6znRV/4o+ML5OlZZATBrq0PsJEzgD+3qI8eZQPkP2q0
tl3TN0mdhUZBTAdGccCA7NSbEabJbW1cobvskovvEnYLU65d145QrGRtoOqMTJHx
l2bHD3SmRzMscm99FWMAKda4NaJA+gI/SQsNSTwwOS04ckDE2bXYRtpEBft9JKCn
vdEbpqXa/3XVFa/HQSfGjzb9FqCYnPRVbKZ+nKRB7ISrRILAsLP7zOFTIbrkrcNk
FsMBh/nEEOSQEVdq5AEk0T3UAJiRY7eCmtVHZ5x4eJonu2WiUTvbmzxAoGsomiSc
w5gahxS9C7JHrEln3EzzO0Ut0BkdOZecwWL2VUs0sEwRoyNoy51837Diu822PBuh
N52dZVbkNtP+bmDib5bapDPv2PGKkAUpNVPNnsCABNUNNTKpOSGVpyj7PQ0thsB7
uLLso7hBNfyOLhdhh1GRM0VRAJXC6i7cDcO8e54KrYDwoDrFsuOwSwQLvLmYZx9r
VObDMmAt0RNf9vs5XWMX2P4cB4tZ0AfeyoHaw3o0ZuxmQkbo+8Ula/zbdmXGFQ3l
NlQ/0wJxXNsPW7op34nMlkWDrdK1keIGlMyzBJE/265UyX1bNYyvkFOy6/VxuDHy
N+/MK6W9JKHc6yGNqwRWLEZd038M2I3tiZgHLRiKZgDfHhWA9ymN6rtcWakuUYV4
E2DIQgJPzOAa+NFgJSd8Mnkw0qMoTYt91tnH3Twk5MxKZ3QeiD2Ir1rT7/sPqSC3
jKxYDltFTyNDbI7vPObIMeU4VLp2zgUKTYTpeqEaeGiLb2vWyAkAoHfxgkkNXgec
mqb2h3gFuFyI6C+ekUcKHlqCloULPacVbhIvQGHjFzFC/q1r+iVTp0SNLtsE2YFo
8XUHx8pQxrWyXkuqOdBmN3TurfjX1E09Ec1daSPZAsSpmP7J2HEzo5RSH6/41+Rn
HSq7CIl31GvKepbIn4stn/mn4hvM+NBQBjGgEZTd3gn7W8t3gNZZ088lSJXzLFjU
eoNJJAjc0lm5VuMXRO/ChFkXN7Uiv0Lg+u1PGjOCAHjCzd5M5JnzK7lcrNnionCt
zCKZ0cW2FdJIsD1eOSaOX/Br7qjZJSmVBp1lG+4tdmuLX9HEK0Y3i1xGaFJMrgog
/q2Bui8m+HIL2sLiitQEbudv9yU5AmUQNaIZqgarcCmutniRxF0UMA5KLuZfZU5T
mrA5vtm4ba9Iw3zdN7IyMkv/BQ3a/ukXrU3g/WLSH0cArbOT8GkYD3YqQ2wD8iP8
X5SRU7WhwAP6ipzWqbw2IYG4zHMzMNgMUqBOoFGdjelfP2z1/8JnlxwVchuDaReq
kOEGcTd+4NGzKmzSne26u5glUcqsHCxYI+ksVRFw/ASAhCipRLzX4vogYEvxcWyh
hhzfJ6teUiKCVW1BslCNSnjn+W3H0y45fV6WuLSgKeLY6BlefHoLhnCE/aVjBQYY
LDMkefpvGKPU3MoK0OgVa4iygyNjVsqUWQt5NX5gREyBX6+xd8rsFX0aN7cOLeOz
wFwM3nMo1Dr5nMb3Xwt+b7i8Tkz4Y9bEgxZFz9kBhxu+lKwGyF7kX4A3bti0nK18
APe9zZRBqqyZu1DsxDE+7zgmVHMVvWkH/WCf+QJeA9m16efhkShUAIcZRvQQYJBs
z3KejJqMPm46c9a+34CS3QQRf0qZSmuJmr1+qqASernvQjsMZBZXt3Zx1Kwf2BVC
sm0vALlre5pXbD1zLq7FfkWK+Hcp+P/pKZegunOj9YnP/szDNq6cm24MCqmFoBxq
Uy0fPWiIHZhPYdcXoSLCO4ayjSqMohYB8Bg7QDIcHgAMOyUtuMonLmORA80Z1euN
URHk0mLyoDqSpB19YDl3FdE34CxQYM4P49m7uUsvtov9RrBxLGjWvnHBoQfw/m45
q8AId4fDvIxuM9Pv5BXgVncgrRyideyyoS2nbYqsqlStYomcs6VySl7Wt9FOgXQu
yX7RLGytrT+QXgXSfQ6pOQShzO8GIFaLqDEVnRWJIij+Mh74ebjVpHOTcMPejFUz
Bvv6r+fInJhETfwIC552Jxvb+G9Z8nsnvGG8e/leaYVtEXinYMCnq7u+USv2YS+Z
EM0OyPJ8o9/4juKDAkypjTmdV43zxnpBKDL5mUFvaGVaRPCIbxd0rqO/KL5keVnc
VpHcGyV67B0909pPm8NpM5tOmvOhhawyiRa5lCghRviRQFD5H3Dfbm0tOWLZ8e2s
blO4Pio8LtBMKmUq1+gAtL+V7Sbbe2f8kpUPStR8mdwjjYAL5B+pMBpdaVIr+ZEu
Y8+ojzraXg3XzY8TxuRNNTiCUU9bxtP9+N41H3tTSMjKPjZsqgSPE4TnDVQAdruN
XX7yzNMjxXxJmXQCPDG12JEGe+i9ceecT7J8Ugqg6QuqUUm5jccO8sSGPUjD19Pz
WrNrDBAZQUOKhssASroOS29Cug+p0R/wNkBG+2EWy9Xa3Se0lZ3J5b1fTYYX5W3f
/jVcoOFXdbv/yD9xauKqzMin+ONUrBjY9wYj/Vhj4qPlx6ZvaQGxQvKdiOeSYCZR
dbgjqbM0IU2aL+P09qJ37VdC2IT9aGXUXFEN6VESzp9S/MLJIeKPTXpKTEf4mlZm
yqUlWnrGIMT8Mk2DbWcYIps7mI7njuNYnH/8RNE6AI5ehfbNaaBTkzIECkUyUmab
Dwc3CtZ0wAABHnsXiIOp/rES9RGWxMkHv2A3fFx5+7ylPwI5402g/7CPTzN0WGpl
Rn20GN63vpkyjifBoPBLXeAa/UipeXPv+wmcahXS082oG7sEG21IwXCm6pFq0k9y
4xvJ7Y7P89tAhLchavoHcCYCv+usMkdsihh+kLfLw8ACdWnVVuCpgAj4vCkksVSp
8i4HtDykddNjwjx95w8nLjw75iRGJ0ENK1+DmPVCW8fPu3z3vqyGZvZqJuRlNuJ+
yhpLBtEvBlz1cyUhFh9SUMo90MnhoyO+MHRlokerkALFIOMPGLpIqkE2Vw4K/Wo0
Czy0lNNtV3/hOayuS0oWNcYIkgZ1lFXiaUWuHx4oW/jDn78avr+JB8ijdDLJM5hx
UU026pPjXGusyBDNzCq0CAs4yx7mXm1yJzGdGQXItFSO2Mfxc+Pk2ENAsvsCVmDJ
Fwhyvf+8CRAWDhZlJSW1EZIeRmEQuemc9mOI7ajK8u1Of6gvZy3zKI/2xXubm+uG
hIeslGljO2Jbg37iEsv86XsYyQ9jplNTGDRaEK9I+XVYDFH5Nt5PD98SWtVo0CZU
zio0C0q4hv5nkvzxVPknb55dHYGCd7mM5KpEDzqIs9UkheTMjHlIPHOCFf+KxV8p
Yedns2cmyNn0Tji17U3FQinVjG8Sw/v6jPxL0XgOU3eHqOa3SB/fl+yj7hbIJ3vw
P809HdICNdSb0A8T1S0gQmhp29L3VGpOyF9Zlc5XaRrdPzx6fncnoD2t7mEezcgN
coxf0sZqbqnZcfrL+tihk//9nSJeAOWcJllvoji0Whs/EI7wojVnkFpqM9l8u3bo
DDknJGLpsjPJcJIVqQtwKhPqkBdowNRso8fa5rpyHDVmQUwPOHfv305k1/hLj7PG
4A8wek4P51FgXSzm8iI9R4AeDdt1mzocdu9kjSPj6ykXJEOADSEZUTRmnCQ/gOa2
QAdx8xVEXR75Sp0B8Trs5z1JvdqhZ6L82BIV6smgVyMLIFgVWollkxEkNbW6E1a1
Y2oCslKMIOyHz8CYEGPij1SrFy6wXRhEwtA8bW8TTKdnMQXgdzPfG1N+PJ59zyay
2wcbGaD9zi3a6bV+RoLigdtHdWKAdt0QApuD3pbyxpEbuzSq4JCJ/6TzY9Dg4qsB
pd0DOkiYm0AhwYdKuq2Ixwlt+s1peBGM3ZQ1gbGmwWexEaLdDlpQC5GkYOJglHTz
N4WhrVW4ZG6PZ2bWWFiGL9mv8bC62hGOt64/e68fQecXerCUai2dXp3/UXnCF3XU
qZvtYC7HrtJCeO1UU8oVZ/cf4m8IO2nGBd6OJlZJxu+WE9QaamqJrglsgesHFNzY
DV4JIxCW+qc4wXQYMRlk4XCpn5D/03KuOei2Pg7bOgJSV15MfiIY+pBgn1kwHxBu
mCTdXR/7SaM/08m6U3fYbilhNGlkFr9apjr2IvWfkCpqVppDASruz/f0zvbQB7iW
kRcB4rADTZb3V/lSZvvkCx3XVR1/d1YaZzEilaTQlqsAJ88X7C5LW8+kHGmFz85+
tkOwatFgOrL4rcA4wvpTovr/sDMcV5R6APhg6odB5J72O2JOSEwaBOk6k/p+/NI7
nMGE9UaMASsXT6P/XOOsMBhUpjphPHzIUN734vf+JzaC3ahTfGqsKU2TzMUleQBH
bmrK9h+jy4RMR7J1+nzuX1W23IIdygBWs3+yyd2YGPnA/7DTem6XOd3nKo7ofZ/v
AYtV+0Rq9FoBBtcHpn48sQR3ovBaPDV3+8Q0TIi64+AAF7+T5ObkEiyx28LDGYiL
rlduk5pG/3s7aGjqpMYu79VDviKRUJDJme120hhF0itBFv959Wbw3SNU9kFFVlFz
ZkaOuCmY6VMwqUHacMi+9qOQrHZCm7to6GszQh17Rzn4XcD3lrAUuCaHIghg3eP/
xLF/j43zZ5HKMsLurvZhHyj+1uxt94SFm7195fKDiYu0szbxQC3pbyyHK+p7/qWK
ZEP1LEgg9VKhOSjseDF/zyTvl3ySj0auXCTPYyeVbBCPgRNUEZpVul8fYXmJjOhH
zDYQ8V+8RTpPBgPCvQu1D2MvVbbeCw5AZ0zwBWq7IB0JbzVHRsPaaaoE4qQ+MEQP
bvNJ/ACE/mR+uizfDJ3TvIFpcMKJQOUqjCNLPMxYZ35hBr5fgKwKjuhkkAlzsc+E
Q9+MVPhGk9bkOdK9ucGawHHYfaHOaIxKHOGgUsZR0GU0ZFx+I8J8+6Fqq5iN9ok/
FNdy15bL/htXaKQnjImwNyU8c7vpYumjPZ6YOwuPCVdmAB6Ti5a5OkKzfEJMB/g9
jsWusszpNEvCC6CAb6oSkIBAFWhRHQuC5H9qmxMF0vxWmZzSUdNolxRt0OK9zpNQ
RGgBwjVRAKM6RY+b4RXjU1/W+kD5FynMp8T413JW9P4vFlnNxaG24Az+y9B5iS1u
RZCwaEQMotFuJlK52mhwhuosUPMbJP5Bvx++FhqwuXdeIdSSCVlCsC0AltkAWxJN
gno9Bd8QmFh9knMQq6GbnO1eF+VTyCPf6Iu7ITOZr9pKTwAsfjZcLRdRyA0T78Rf
QQb0dixGXuyZhE/81w7J++lp2LFgGnUe/8U0a5m0VieB/818TszfoQYBEEL6c68p
zOoK7iQ58xTsWACJ7qTOWaFACAFXPQuel3Hq+Te01CJcTkOhLxQKOkTOBsYYww7Y
v5yYKIKYczpoB6sfpJNSxeJNn4MNt3pVXZh+/KGYF8rDWByQoK3cALl2fUPOtnsA
jMQhqlBmNBPXFnuMgKF7oqS9S7UbDud0aJylLENraoCNO+tfraAsXNOwhhN4CarY
XVzwLoq+Yqt3tFpPlcEBt/xYtduKaKFck4+kkH4lXz/miAel3EVmThrcs4YBavuA
1EqP9JTJmb+Q57hWvYOWUFQe+XqBGvMUBMjHkzhfCbZrwpd/+Nkf9UWLC+p0v2Ev
I2BsMy/koRyEAsiVSZ8W3oXpwSqcI4Si5b47WLCsu684wNxY0oiF9Q0nQVFCudXr
5N4wWAVjPrJqN0PNDDx3wwxoniVrXIdtYw7Ojcpa4cP/9odE/KtVVwrVkffPSsTG
je3bqV1dmH25gGt6Ys4XnV9ZvSrs4jDxZmipmen65nMsLMZi9tW728uk1E9i34P3
QNAgh5bI6q5xUl68RJ7lecsQR57QW/EcecVKrben2ng76lYGqR9+H8Rqva9T0N+N
s7V2+zYuogyp4Vf2i+mIwVTn/gEVlKc9mddGwtZLrSDLoNRCY+ff+lJHt4rRl9lq
nArQjD4Qb1y5ubG++oFWq7ocKUj6l+yY1FceBCHzbqORoF1eCzMI2xxtPXjl+qk3
FIGMMr0pJFN3T2Q5zdlKPo44gy2/NudcpHOwAd+vDwE82IkfH9ag4wfeHkhLo3fk
GlWZCWfkez0xDLK44eS54Q1KcYegHKwkklBdB4qmFWgiYP85ECVWQBOKqz+sX/c0
uI01kjlWZXZh3IhSUr8oY+0KT6rLausZr/fcC25pEToQl3yC2tIwptVgyUN9suy0
CZPF782ICHflKVqeZlr1OpEdfvoR85BnC9W0NEdu2zEEXdfOi9Cg9Bx7QO7vECnH
O+k33C85KQ2I6y7kjbK9r5vfG/0+jbKbW3YsdwAY5G1kc3962bCjRKAhJxqdoPp4
VfE6Ozl652GrqnQrEtHShEAf3GGz+de+TEU3btMILuDjENvtrpQfOGtUmzUzwsdo
YpO0NPvh00bbTOJV5DRwq8so/7xfIb3DvjfeI5hTC3PYwcfase3FEb1OJU5r+sDl
PvihxT3E31Ao1mh5UlhYsHTWKSRJNwgnXYjl1jIzXj+Zps36g/I7YFFY0nj91qQC
emLki6FtiGUg4uB9P5VCS50K78MJIylazcBoarUrDGON4GdSh6EB1Y9tAAxYZaAP
9wwvU9ookmcOBdKQtFY2yYGqFjkyd1kebL9MVSr0iw6XFsZto2fn9u88wx9GY5N1
P7OuR2mN5de7XCbxUjGFz1t8holARHLRFknL2wRtOe5lH2Wpio7QAsIMcG0pSkVB
BLTNGH3uEkH2+U2D06r3tVOmocFgYieCewRGRSb4JGaNoZ+CdVwap9y9WVZtiU97
r3722/BSV8chIUhA6P4E3LEOLHNBTJRSCRhmT4i9jfmfXqoEHy0SqfKb+bcj+1as
GZdh0ULECnl6boWkZvi4wEWZTUXhbCJzfTmKYP8WXCPEiEcAK9sNOf4ONw8jHkhT
Fwi65AZMF7Mt3ApdADWk5idtUgel+pJ6k22xecLmlL/EQNfRC6VPDT6AxqolhfMb
KzmgS+ba+pxIh+9hOz6eRn15a2j/wFPhq8mMWc+K3AXgp6xzmLOy/pHVwtJLgKaB
BNfjJZsnNxkkAt0BZ1bTLWaGZXHBgcu47U8W7VKewwYfuDlf2f5lEW3ZO584ENva
rk5egpKuLZ93XJRkf+HOJwb36FnabKgIyUtj9C2aCTZ4HXS2Z8NxDgIpjXX0SCJS
8fe8enTryUtSKeQK0Gmklpfpj7qKvfQGRzT6si4A1OatBF/LqA+A+dG1TFpImidO
QjWso6RNz1UtQyoEvAYFcEMKOcEsFYJlehmMr6g09v3NYXQ/QdIcnUJ4xFxcQ7ET
PmASQRQzSaIgdzeNKKZrrtr612P38/m8BrUAxkRIjfX37UchwR1kZXItnaMkQqLl
bheAJPtkoOwunjn4+ofL/aLizCH55xg6VYLEJS4R5dLd4oJL1YGIAII5HCtvbCBx
++f2JlbC1oCfFQ/RnbnbtjVzLpHRGbf5inUJkEXMolBvdfobkVNb8Zuhtk/iqmN8
rMniuRkxVz9cYcrHNvRhavsPQ5popywlCESZEjO7he6Jf8hLOyMRGVkoN4k6P60/
oDjZy7wLLY85b6+wLIe+/mWs8x8xcdDMTlqexiAiAiLjn+owVeDyflQERJEqxIEo
QEUzhagkIm++oxs7wL3dOyDVIbUBLiz3+bMKOtCjRVZaTL9Hd1fpc7R560OCV8Fi
ZvxKXncW4kRG1LKoEuMlVQQtkppiSSbUqkRV2hBdXpg84XS6ydwP77ly+q49d3Zb
ok5QeKGI1LtdNbDsLvlGV06biSZ9yQc2b5uyp1TQe/na9bRBV3M32pURi3nyJNy8
dEYaG0VKmJkguPLzMIXRC4z/fDU04JzINf+5KAyUBpnArGKZNXF160H+Mv4mE2CG
/ViTM6F8rMqOI1E8dUj6uH1p2DVRdDw/h4Sl8JYLRnQRHdxf3pFEAoncfvu9P6SI
Rxk+Pxx3DzxfwWPiTkzj3MMZMQ3i4exo5WFVUgum5GZdHT3LTFV143Xp2aRnz8lI
qxsaiRzwpUPJ17+gUMRBZg1mWE4CfIepXvlKj2CT1/ZH0aKp/dGOQ/O231p74T8d
m7DXnj8mRolhEjD0aOjpYO873UyJfmDYyWRjOQEVwASSoW/a8LUwJOcUrZzmpH1J
97Q8K5Cvj4AMRFKQb4YRACnC07ZerOBEj/etxWngf/jt+IV20aTWwbA+RIvop5+s
rPFlcmvbcyhhQoTTbOIsz/GacnWqTYvMTuvu+MKX4SdXYB0O2hcGtih2Nz3LyLd6
1yMg3xbB2r6kWZefxWkfLqIS5AzJ4VDD5LPAXTmfrObwq/HPO8JIYQ0EhdCJXvGA
UDBpG/wTe19k/qZoq/7z/7SRDTNxmrCES6Nu8LHC/wnOTU3ho+NgjmzYXmg9tRNy
z2HmOu63XfIstrnmZWSBc185lJ5vY+1CJV1jluFzqdD4ju4qRu+pnsTW0PRgNEI9
pIWQGspt8SKV3WTBM8qMDA57AIQCa/WirpRrLIqDrSaTZ9SR3IxQAIS3YctUKZ/e
pAJtW7AzFo9+Agkr79WU3Zl0TcRZr1UmB36TToApLEu9vVeB14ZAgOQTORSxvR4t
N9ufmpOpWe3F7Lbab7X88L+tri8BC3HeN9xRhwowDt8L5dsnLUsvep2HRr48HuHG
l6K/BnYS73XKJjxaxcWcImNa/vo7mrUl3Lk334mqMxVhuePmJeOFktpOFtp9zA/q
tEUAZiHtdxOxGTenLvqoNHORJEFXti0Zm/9R5ferH0+ZogFg/cOc/CGgZI8w/oOh
qSQ6tZccse7FcRWG8Cxjbn6at5vY4BFNOvMN5Fe7bKURYZ76627SPG9T3C6XqQxA
7Fi1ctW3sevyCgIDRxjyD1MpdDYjcDA3yVhxDGiEwcHpD/ZZ6KRTzxihyZ/3AGCx
wjBubhZaG5c4+FzPHT5U16GbOKTR8RCmKp2FgOPJEgdQBBe70mUW6FpYKhELN3fn
SliPcJ2aCMQwRa63tLUtVLUflBuJ9XmSftkDBmFxvwi16wenb4fUPU88rVrK0gWc
prUxx+z/oKDdXXyza7B9032EWw9HArj49P8BF6wRPDvUeU6RVEnYwjTlDtvXsPyP
SyzCR7Vg4YleJd6NEDP8qh/Qj22z4klWW47j2ZOXg/CueOt49OmDon4is5nvVnLH
hyOP5L08RoegKxk8jHB+2vCSq+TErULq+CDxomvgDfv5EZn2HVE4vnpv0XMyo37r
xtnoblWA/xlbdzQsbvVWrZDr6Fjictpd8VXZ3nNDs2kqpsJWACiRXehhUDC5UAfw
lO64MK2EkkPoiE2Ld2PG7DxLxpbIIcdXtnZ3/LRrX2cfzUzk/gIf08FTIGYV+D04
3rbkMdX3EbEaiuuBEC6XNo+kKD10cm/JrXVEfcPmWa1neyPvyipyfEs0wizB3D2g
NeyQNIKCffXJcIFf9KODiW2d+9gUB8+QrG89/o6YYOdbwWv40zbdLT4BXsNqILgu
UM9RNTh9N06x8dX8UPuwUj58coeniEP7xF7+qoxRaoB9e1knFa0QfA7dTj59Gj/4
AZvTY/cWv8YZduK2FFC1GXtHJerIU0R1L+atW3EcNZtdw8kgmWOXmYaYtDLxsuW7
O3ZgqAnyKnpaRYTMagxV5flpaU/t/84hULUMFQNnqJxYEmWe4pMYobjSA5O4Ec/h
G3b3YhaabUbVn/fyjho2yVtxPJhfj3dDMsKWQXmlQjvuWQNKJIJUEEnZaPlsdHHK
thsOKKDIvrh/khuBhrnwWzYnqjSDzmNi0l4xoM7ooh+8P22esRJnTzI1+QPQWJha
/Tj9XK7DsMGDX+EsdxdB8uXyxjpbPOheJO3RTlWvZp2iiWWNowXYgBymHmFxwmbH
TnSvjMIiRvR/f2MaoP5Xvlj0jG0Kz9QP2lsBPLmeRjWeBNcTCwgcJr8NWj7vAdsu
j6jKLqvg/LdWOM3sUObBfwsw4jm8+phdOI/iZ4BBbUJrjH5wn/r6x5lwZhWEiWKf
QPmGEcrRv1WkqX+kOCYdUN3vo7aTu9yYYIuGk/u8Q5PpvbO0sELt8yTwjFq1i8pT
J6HPfctlwQYXStesIvYwBRRHV7U86CvqVK57+GdLZUZ6dDmyFl6rbvQ6uvamZfmz
lTSDOTzcgMze8PvLvBJWTDJZ41f594+8TDWLTwrwQ09rxL7D+ockiqimHSLq2rtk
Ejz8+M6GmAYS5NMumzZ4Oof0IuOey7+2JCg5ptwkp3IgkuHrfBhB9aJXquVey/fd
8dMNSedpo9ko+hfuvoz1ZGRsIjEZybgYiAJbjlw/5/hYu1sC4tjNKF6WHlQWmx5T
nISaMsc7QjtCIzrFt7d1HsYbT6R7/n4pVGw1bjlLQdL/eBv3CQPpg+7XlO40+Ks9
VZYfm7GrNHjdF+nARR+F/0T/1bkkBJLX6qsfV6mYXwZ9kF+Pm8PaYAZfwnm502MH
SNREIRPGzhi+Y7fWqmT7vl6bgA2GtT4A5fsDaMHThSuqNzmVJiRxmUFuOL0qf9ip
CSoqFJkut5durrdi5103XM0C6h2t0+lKRgcpmI9gDP47QdIswOAoM2FqNK9DyXeT
s0ND2pbqBuheew9mjX5QQDPBa/ol6NT0846yg909rKBFvCtbrWBQkDG02AQtcmZ+
DkiuzIsQLBpdi8z/mBPi+XWtTLFIXGZaGB1IaYSDvWhDFCgFshlP4M0rkTEnc3Eb
PxGdcDp6x97WSrHrFchtB5XuBdxaIQXmCYR+9y3CZ64RFv4PjEJenMsHQOOCNtEb
V7l4le6XeEbpq2WnqrLlDy2LGfZAgHMw+oFVoldKiybOg605HlmKMYAlBs+cNAmA
QxnTqlbpAqSq4Y1CwMJWhzqZk1MHduHhwMOZGZ6aMJGQxvyOJXaH3EPuxOLYtjK5
niEYapm5ILBeSEn4BlKTGnyj0ivviLh+/dxM52wpD1nqOqbWqVOGI2JMau9uIOhQ
M7FNeEUpLylSq5nNf+gxZK9vuqUyIYZcLci0IcsGb3o5Kp1gu41iyWBZ0f7G4cL0
O6ORtuZ5ysVVwEi9K+5md10/WVJ67GpSvBlNyJLN8KhKTvKSHhPPno+FE7lJYMCT
zRlg2Fx6lSGXfGj74R8Ir9Op6MJ5/9FZviAasqQltO/d7JJNNZKJ5dWHkHzKCKtF
Ynaij++nVfcPmXTkbjV8Jpzh+ymWy3cOKXRYSCj02Abasd32Pl5yhZqwIF4axUH9
81jRfNPioD91yVeuyPij8TTBQLw++4IMYix8EK7vwKo3pQBec55GQDfJLQUeAOoo
YgQ92D1HRXf/HjkPQXJ2XdwyMN76SXuA9CrF66tZgAVYMvm3KvJ17cTZXAB7btwY
eGDx7pP4I+BHKK6bM5ymcP+qkwfDc+5R+ND08f4mX+8aGoLj7TB6fcS03KaFlelY
xdCiSeGpZm8CUEOn9xQRIAoL0Chd2X1KItgmIzmlz7JC9aRRhgN5cGbfFG/lRmrD
2LMJx7dy7iIVB4O+C+ewPRGaGHTo43sB+tr1QQ66L7V5eiWItjKWG6Io6m0RjYbn
LVCm+qVsQLK1asJI/JiXxwPzAw7pG21utePuswUnrhaJyBI8HE4Uios5+TYmt3gI
Aygbngiiu52IrehMoeMrvme34am+4ePo7KN2/+J9F7mbQ86qF7/xkRf0BgYTTiXt
DdqvGkacZG0AoB2ABjcxb9+Tj3YWdMBUFdBNqRetW1v+CMbzcyb6Ifdwp21fCY6C
cfuxVX+zPA57rROYF9ns6wPTcVOMNgoslgS0A7IlYybfmoGfp35x55XvMhABl6y+
9Ui7vssOrWKmelUGO56GCZ3zdtrBNuF6dMmPZLa2Ry74wBnn/evtDKfsyD5Zo5+Z
9ZQFIM+nTCKdJwuxuPsIfrR/eLJ8OWQFvlaJmcEbfahVY1XYnOuN7vhKkRsYZkYP
k9Sy08Qmx7KsMLxfcruvpaABB8gmQ4y2EScjqfbPxfVGPvgVsHOcE8+120YGEa8P
vWyAZ8Tk/PZox7XLxGEs9FJeI3Ax8LbgTtEoWFiohtExVQnbAm83Ay6WAJw5fV8m
7Ge7uiDCKZ79GLSrxZAYcM4R6IaBzl68a6rvf8CbvAIz/tePTJaGulATp7z1+w8H
uEiL58NT+U/VE6aLooIljpKoc5yC4v7ZR4x+8yBalgoYZPE52wT3tRLmyryB6z/f
BGUCgGBxKkaEJX/TtxxbmLbEx8VN5rqOitELFf469BImGd3GrkCmJbUt1g+BSAHM
ujfRemdaPrzr2T+t8tcUtvh9To/EcUA54b5GWes/W/tfox13mG58WnILKVrtCAS/
Ey5ETgfHq1maUeIodR5rCAXfGZkraxUKXE6pFpMuRQDs2h5t0d6eKqbisUrkuBlV
8nz+Kn28tFM7bBkYmlpGtLUqEKHt0UHgJ5nEmW7E6l2h6MHXFlra2TtsVTDaluxJ
tPZIKQjc7icHj2l3fsSMfA9Sf0DvfUyMTDWl3Ut9lQ4OP+0RNcUGbZcE490sT9Ey
VPn+ruah7AkgN2SQt47rDP5wNsj3NoaxjpDH+OmHY9dje3GWbRoYKubF5fn/ZwBN
qx4+HAJeT9r6YqG4dfft5z7EbSJW5pLWfzSb9Ev59Yw+SwgDvmX0S5FJfZf4+Knu
QOvQIY15zQlMTbWDrWqWn9tzcG3hv2zZsM3TjSdMOJDPoB3bAiQEgVkjUNSKH1a7
6Dl+0YWSI/aMiSxRJ9U7DvuWtlegWPMYXOTDczPFU6MbFTf7osrnAU4BYFi/MMVj
kZaBRnn1pTnAKYnBxkVDU2HNzmmVeaOlImBPjzjulu/bb0ObYXbRJSQs1tQgRBok
5yAzpHPEboC3x9wQdgpqc1bZAtyIahYi2xfFd4NYVXIAhBOlVwdUvHOpIsn0btly
Bfb3h2gr9Qvg596h4ieUUwB7eLN7JLHU0v0rsd+A169G7Rbag7Cu+Fxdm5oz+E4v
br/e9oWO8LHdgbV0KpkKP6IgZG6ehxsRfr6oU13rFbPWxptBFK6OivUjV9jOTCCa
r2Cn40ub1NTcAoux9bc23GA3nV48Fai9F1727yH/SPgnTzoe2K2eHI0nhppjasgv
ehcYgs/Rkqckm2YZycfVee77DatP3vzQdmPkpR3RJ0AYgDe31+VlupV2ltaJ/qQm
bCoiToGEf1+N4DPd8C/J0Ty9flAPo/jVQHIbttKulSZRylY2xpLxFIzwaXftj9Es
aR+2uOnJsJFP27LNH/cv+Aa/ROkTTL7t/PUlZ9QWmy4CGPmzAlV9oypOYQUhFKai
1V+KgVlKGuDpAXIBlFTmOPFDjsHB6SArOqFolIukLL4KU1lgUQ4r2CCa5XLT9yeA
M8hE57OUYQjsWmJSUGDZrgi7ypupiacl4EEBo0Y2oXo8G+Rt8N0mFxBp3/KaIP2c
OroAlwwp5KBjkzoHE9IaR9/3w/1NgXVpesvFAnCHkdh8+T3lh9vm2//+ygrzFDJh
CUysnz8AUAegEj5w2Q/on/vNzgXvWg7Y5ZLedSBuCpNyERpIayXQbLp501CBbstC
xSdLv8sxIgEUmY5ETuOuzHL4ovMzMuRDSX9j59wWYcrIL2GinV3q8D9XuJIpnvj1
vLS+jxAYX9zgpZaGJq9K6o9zPLiU++h17RPNr+0dcby5SNDHr9tr8SNl6J2+pcJJ
pa3SDSGXI8NLh/V7eoC3ajbLhwcfRrNHCwLEkPqJfz/lP/gB1xZHWDOq6klfq2jO
fYjDxaGskH+vrQx3lTgDvwPjb6UoEA2AADwxymds6pO2B8NgOf6PFobqBr4l04CN
mlHD29YLrAOuogKMs10YeQlG2qdd1Lco+aJABm3GnOrWhjwSRanpjN2Qtu+u4LHe
nvDx+khKrs9+bA+e1oQ33k0wYz9TmebRg6ePFdvdaQKTmoU8aF2P8vwSdkz9jb3K
ydl55aoJe54ct6/ozTVNOWqRbVAgf3gRFDqjCLBMwefWb+jyK4AlLnKcjeHU/w5F
75R5/wdCUu7kU0tfL2sgzbCKhhPeepkLdhhjS9itMnyDmAtBVwsWIr6U30Hl/Ig+
qBXU5BQPb2UMjgkCA7WXV4qIKpVUOGgCVOtyEwV2zeN6qboFWGbn2wPsd9ZX+yl+
h7z862hI+MnhZA2/cMPvNOPS0qXaPOvLnO4HNsOStYqvS7mDK7NU1ho3ElescREW
mIn3hodd62OofIluBZ4pVzIuoL1EhL5KOCE9WaWa/zhUImQ558y1ZYXU55C6uTqe
Fs0p7BaxPWb7yM0rULnIpq58JlDO69D63Svo+vYsyzdNxiF6K9xtIY3qIQrOxPL4
tdWwiA7r0zCHdAiIl5PVyuAZcfcWdn8bjG90Gt7jZHO89HepJowjvZQTgoVZcPHN
/ajFVhtqNXEuXmwxi3CJDPaoKd5bAvtm73M+zVa5kvjTVEMEvvbpvu/V2lTMkhxc
TXk0XQHJlXvefuIwlK5eJyQ5Uj7dFGbzSmTquwVZ4AhhIcaOpOKXtTuNGZOj9o9c
bGBddRMkwiqbbQqd+d9rypxyItxgrgCcuPRWqk9ZgRD6AEA9CcDf3aR6NtnhxWiY
HuMXOladS1xQaUQK0O8rC53ik5560JVFLhgyudHv/gRMEDPSyTFGhJLYwCBPwYCk
1zNdq2eGm+aFdyqFocz3GKZwB3xJZtoV4qmVMmMvCzEKtg0GUB94LL5fgvA0t/n+
J9hGrw7sA8sQI+4ydaahO+cV7ADMKCA5AhVdLeyJMLsi7XWedkd3hjYxv4V0opdj
5NB/63psTzwhbfR43CAI0SBL2aq1LcEY4cDjxKNU1iAnX8Wzkon0w2Ylqlv88+X0
3fDIVcCn4EA89/uTPe2cDSGsfby0Ql3HLBHOA4NmR+i6qfJKdZyQxjMpbxE4/cFE
JyMrx3IgAHmvrGOlNN/ahttqIkPzCdUvlcadencmLOjzCyJNAwwsycL/qTsTbrSo
Yi0v3kICrGqGCo8xle0QsIjjzG8xKqUJRAV7JGZ7OSLBzJkXY879aTddR6Vwp5+P
aovxvdyxIDR2fsXrIBrU6ZteAWh7dgmuhpQq9tRUB59qTEterYZ/1ztgWlS1djAr
cc404DNj5Pd1Q63Jnlsz8AzzH08RvDarJZfR4licWaQMG1/EsMBItZuvByza9GI4
KROya5jviVVRtKwAj56qCPpnUA3jNAPPFRs2ZilXofHnsSuQRj7jgCWSx9LxnM2a
YlrWUV8vRDtAnakiqWsiQuLCf1HlA3Q2SAhro+PcRYplINxtnvge2m37TJXhoW4V
7tUud96yzocjwmh50mZTzDC0i3cgCh1mdd/7ikXWfbQWzI24d4+EGY/vCtidUHBf
w533g5hnnquEfmazpylZ9eDCT8NM52n9a4hNmNo1a4aO06QccyqFH1OJUJebukTp
UvRBGydxNoH9bpoZQP9scEy9Hi9j6qIvPJP/r8UC2ilq3qEOW+lDO5GpXP9Gewys
Kz1NM6TlsFiTMkkgfVaOgKbytVVf4xGw6XuQz3HuMJnISxBjxciQmYeHn3NssD4/
rX4GOkxEG9iJ5iYztDqoFvX6oak3EE5L4+6/Y7ZV64J5BnEFuNCe9Yr6b5jNHpLE
t284kBKu6a2oreSjp8okJxhb1V9OZt/R0r8Aq184PLA1zYmkp3f/uM7uGIGj0rXt
3/BTl+9IEN0/aE9ynqmPUavj/JgakJ8bVnJkSiuYJ09bxcMMFq+u1+Sov+PqiuHM
dzWTfT7MDTR50iMlPgVIU/B730yxAVMTA4WXDVbPdhRF9BzQdwDLQrqcXsUX8X3f
a8wqEM1Op+KAPPesjKpyffQxrUI3AQdKdCTnnbpJXxuQhxNTsNzHR3ON5K4LTO8j
/p7cmqYeFD5oshcKwZROrvGvYWzC6HBlW7E1n1Q/RR7AkikXSSZD7gWrm3trF/S6
7nhGfsMBKRXPVnf7N8mBsuzQSSV5UUG5ocWKFp3mj/PahumAtV2wX76Yes253wNq
PY5UZpdUcCITyQINHK7qB26JzANYuCEwfUSxFMoLyQW2+0QUbEjaSOpAedAGJVgP
+YUSB8zEDap/YIXYbPIYixUA/euNiFk6ClqFEoT8dMO8Npbo5x0tvLsn53D9KNhX
wVLuuROCqSKDXlnMH/6njvFr30J6/3YUj3IQDe26VKexA2HdOL0FA5ukaVyrvgsb
Wisy75SXFAs2knt34XEWScTg2DxX+SNIYqiYZfAC54WAxO60f+ebpI5wGJr61u/+
JkLqtO3Jrhm015EYnI2ahaNBK+dA4W2rjTsw4yqdomTTQFMBlkN9bX/HveYQ/4zH
s2HZg98a3Zm/egZz3HpOEQQuZN1VlbpiCPNuNtxGAz46MoRzaTXnrer0aIPF83/0
8vqueRWDXfPasrcB6sPIx3RS8y89mGgeg7XuXAS6kmHACYOGs29nwx35YRTLUldn
Val22KpETFXR1L4DsKpR4j7OwzlS6MIzPqQ3Ix9oNIu0TEsRH4jleyCRi6LwE9nx
IJ6QtZnSLMDL/cjUzpllJ9LIIGxU0FGpnOOntryNOAWok8YuXpgyikfK2npUzc3B
aswjdk0iL8H3VOJCb6/jEk65et9sreS/cqC42Ag7HEbjQy7k40mp+Uc49NI1Ilpo
FVbiVPYe6cWcouD42UtBayC8ITXaDK693DBtoeVujnGfhD6b6p/TrtEcxGAKlkI5
G81vOT5dB1jn1ZUcaPFBxkJXEW88I1fId1e/WX6TqgteCuyjRzhwYF+md7G8JnaW
5rboC+Ur91V2KnoctVzMlEsXt+FJJ9I5k39MB+J1y4+ByzddZVRKUNw2/Uro8aoL
+k0o/CkMsBGYoyZCZGpr84zXG+YAJa6FPh1ytnEGlujdWWN4eap693hVwKMJYqjt
KFlTXv+7mn/nJswBEh2+kvj3mrNgJPCQxt8nSawMaCCiQekIOznsPpMjy6QpPPCf
TQy+NUT3iIpmHdKPk2scmv4VoIjofgyHFG2FyEQ7jSaATLCIDdNTz4kY2k0/KNAv
4WeKJnNdUYedgw7VJdm5VIsMT8wRhVffGM8sjJmLqY47jbk11EbZ9iG9/ZSyzWuE
ttYMf3wgotgbJDy3oWh0pAOysLZS2hPc2sgZ/CxFVNzx7SZ2KqRPWYU28BMHBq/W
BoR2cZvF2v0lOgaUBWfjUkIOSTC6Gbk5Pj6d/9gySo1Z1SfOAuHLNCFv5KVZq3Ki
Tp2mMecW626c7r93cccWqQJuB+fysI/qzJZI9sj2UUFydTkJIbL7paVtOcn5Nf/x
TPClN+yflL6e6XYycP/LA00JDUMfJ0POb6HnMThTkAHxEZ6O64khvsLdhQE9gfex
AQ3qZi4sZmt9TYFJfs02lVJtLAES0vkOU8aQvOhOL7eIcGtiLi59y3Hr+xlVU5Wu
MfHo0GkTPuoelq33mf7KfxN4bkYub+U9bTk08wpmSPOukWXj+l9PC4OMcrMWcA9o
gs7kC3Q29z7sZi9NliqsF23OwzaJMaLIj59a+slJrRhYUmbKcE6prbzc+wCKDsNA
bZUmvnBfPlm/y8VCGgFKV5Dl57Chr3ujQD24y886FTgJTiRJHPtQwoNxHxL7h9ys
bSlXg6atum6PpiXMQa8fnkBWQbRm2gleUzRQFURjpreyuCaeHJ7W0R0M3fLF1ek6
KpAzQwU5jHJh0fTPYmkoRQcS4a3DW3NvaAJqgyiKotw50/ITkX7uNagrIPpnQZJu
zS8WZawb95YPhSADTOTpzv/TaX4fJD87YyMhiHAIcOG8LSITmqSaHeP/13LMDc4B
9np1zzSJyJnqJPdn5ayqCKLoDmryCHEjUK5g+DYhJj+fR0AsdQ2USxUgQtcOeXMo
gbuPFIra2ishnSaIujr5sjjKT9kyPMzvQp1gqxH4qAHfz2iLoiVEztsGmAQS5SyI
8z2SWQJV5xXN6TKYh3lLy1q1qrwtw3dUb/oN6PVWlp6S09MixJ2hX2uJNNAP97LV
pWvhFGm+6PeHPc9lnDA6kOlTrD7pLrnYIDWgwvLrXHlEFw0Rcf7a9BmljVYm5ZUA
y0XB1HSNsxNWB6jU4VA/VF/w12IWNx59D3zNIJCS1v63DToa8tJEgPyKtYCCli7Z
LnQbthXmzUnN+qzFekPWpwXSasYPY4IpPeRLP/cGdeBTorFf06Zqqzb3dxjFloxr
hOlUERVg98mEn/zUSwWX0hPrkGsjAfat0L7syqsIsy528i3Rg3sOpYesWvrl9KtC
Dr0lW+RTtDlts9pV8WtFT2NB6Bq9ZypUYY+A18PGHWc5lH66gswelFJp6rFa6WEc
l/Qe+ut3PMH4kYv250E7t7+FxhoOG8cxUhiW0L+vjj8lLUiKlN1554yRIoKZN0tu
DJD7xWg0UqG/sSGghSyrJKcEjEuK9DXiJw0700aJsgC8Pu7PYYm7rLjtn/tTI8HW
m1zJk6grKx3dRwjAZ5twUkkwRSM1qtv5wfZjIW507b1P9lnUukD668kkTkNERGff
yfkACLWeo+YtRKE+yCxHVPl+C9ZKlHj5iHLai2tUPxPeIpmqhcskRC+sLzZU81dn
Ai+6nrr+txq3vyNvm+c5yG/73vklfUgD+HSy8A8zfCU8xaJUht5kpvv8/qCjvIzs
zA9lfCU/CftxzhwMzCzLPDcJ/NDKxZsFbOGKTwYKiQjeQVo+g0O5PMmsjsyYsGJZ
UyDd/d9MYpolpd9jfiu23L2LEoz2AUEEb0/vgyxVNVPf++AHM5u9MFuoOwPiQMV6
XiVySDLmeJdiuuhuCmNCDJPA534zDkZoGEjX4rLFo1RuiSETeaS9ulY6TjXgGotX
R/W5fx//wLMsogYez2DDXXxhOh99SsqdZNn42m6vyNBdKoU9y13Ya9UWEBUI0+0v
zRAmMoGPNBDJykVBCHUKQ8dvhfsaP120YpuS9VcmPKaosrh/IihHI5RwT5qDQHt8
QElPpQEtr7glQLaJFq0252ki9tI6sq/lX+JedHWXUu5gdu6or6N6iAk4rJVdKKav
1pcnNzYJg3vMU+1+e/UWzrXSWpa16+a0l2qgQRnu97SLZCR0fE5IvE+hIoN7TPDz
JtSHzscpLr8Os901hg1gCD8kJWa3Gm3EqRx2bMCsnAdV7xFHnlTetQjpZ7OX44nq
/+Lrp1vi0N5nPVM8admeqgq2bRm5ATiIjx9sGMSeLOXzUxxsg/g/eXR0PqJGzv1O
nTu0h3pFkdVHjN/RMWi8ldSlV8IulNPzoNumRRP0PRvLfHANeXLp9+F1GWXy8xwG
wAfoiaCtYm/5yi0gbXszlq58l28rwvpybeRrbmciDdUZzAQRFJNUjXNhqkKU74Jb
4HRicez0rzV03xafvxAtxiB9L/fLcdxgp7t/HXXJmrQMEaUS6SMHDN6/gb+CoK3l
tROVzRhgy5/LcvvGyuhPnC+6BP1wHcGVRmOm9V5SjIQY/cK4xTdrcz2y9zMtSeNF
fePWa4qYW8VDcww/TtMb0GsWEXpLC9VspZCAxPERGIanJjFDjZ4icg1cZQQwn5jN
MfttVFgsTeUDsipDNAgcmRoDXafq3HXgSzhIZZiQr5czgewRSEUfU2OqpFWgyU2j
OgM6dVlLbwEu+V2cxNbXnkgGdBWOfrpqhVb5jvBAlpeqwglde10zisftDXd3xh7D
I3VroPtDZCCjMF+kA2SIRsBCipXFVhrpPKqPYs4mIVeFTEOvGJFPV80NLjPMdknj
23ly3xVGLRXV5pJYD//fTxRQu5NZ0SSIZdYX+5fhMGOcFBGakD2Zjo1j9vFvGyIJ
1QQl+elrEacdtqXdCwm3tURTM2M1LmpkFTURQggBMII/s5vvjR53suFcE07Eztma
WmAfFB2SGVV9C8UE9M5qZLg0fPVEy9ehLErvxGPAgCNxQNoFJIOgUfXtCn8azCqZ
V899TVSPhdh31HBsuZzcVznrjCiLFT0kLyvTDW1cnVr91t5tQtsVRfAaukrenKXN
cC9T5JS3ux0IzYfCBdDO46p8I3LgPdC4gRJrvi8f6QGJxUUHjYD2dcm2PXOEBQhY
aGentemYUH4YTb0XC2W/ccPsg3ppe+vTeaLPjJkaI9VOew1NBkVVrfhTcH4hwl0P
U24fqW+JKPsWr6hblZG+Vtvr6HXpp89yj5EwecD1TFDJcHvADr+xA/uU+jWfrlp4
WbshXBCn47L6YLVQHz/RG2d60FGaXS+KCoIL2hduMKc7juztGeUpTGclhSSu/Kb5
5De5H64vsPT/0Eq3jPv1POc3S4bBQ2P9Z+nzCbeIWVOp5cGXeUlRBXusCf4JAOVb
dpARRPPIs0M7liEISMIYiTek5WMPubTUgZtQGUSwoy6YhN/gaXvXQaO/1dzTRk0j
J1QM69aYka5FEPS1h33odU+dYRjq2eO9h+bIblIGrGZZ3mEoN5ZWERIPuxPRvCH1
eEsUGmk6FRwoHt4TyXkvTLb2tnsraXl7g9wEo4mmS1aHpwfM6gnfuBPoek28hIvD
iwskt98FAysV/hX+tA9r5ic5NKs+mFmfbgJ4rUROpTL463krw4XEl1Z03cXqPo3b
DK3kr1p3q6HYdyqeg+S2x44YXlwQfOtycxdxbB92i2aVM9IO41lpGxVKMEGPOWjG
h85ctrFIKBMjuY54TjtYaLefa4Sm2QWlje2/KBVzkHHQBaDBP/Lv7Rf+ijqRjp4w
KnNZ5/X7YNN04CVdgVglLfqicr+IedwlQ4sn0Pj/XbfYnhCcajO0vVY6u3qPIvgI
PNkdlr+vkXgzIujDy7tUyRIJhwo2WpQCSLA2ahVWovLmR8wym3rg5EEliz80NCMC
lME+tD/NuBofG5d8qihrnWuYTkM1utHs34jfOyD5ov16U0Rr/2IDM12Ku02Hjyhh
W7XgYGSSd0d1h8aWbzaw1W5DPYEtMHLjFv/LSXiKbG8mLc5lgBeAyedun9b3SKhL
N5T/8sLhTRInXkvyaPFfdC/zbFIWQcXDyovkmPFvwSq/AzzJvVHjYunkfBIt6G32
hMOT7RIugfw5UI+MdO0zqXUNLBe9hypvRuAPGF1CIh0B17kx10pMOfkGCxjQb5Nw
s3aVJw8NsT6g4t7ST+ZwDUfKJWBPHQ5X4ng1VBbR1GSv0PCFwFcSKGeVr5lkGrzf
ILLC4wNMYtRKnNL3RN6isliUWCpj9Ty/H+cPzdIgbzP9DBPi1YpM+aVPrkeutKSd
cTZP9+pvOj0xYbXN9v3LTYuOPoYaIOvr3+KxDjiHWiFbDi79tzLNC9FGGn7NHBiP
CHqYcgif7jYN1Xq+54Mw5BrfzNZtSnOt4B613qw5yh+dIStR9aJ268/nmz4aDraR
9g47kdp8kZH3VjkptkHc/DX4Y3BINNQ4zwgTTTrW8QR1/Pisej4Zc1jIajUduTuF
1Jhs4z1d2yJf1l4D8golCTsI8G6ogaVGRlTW3+RgAVtbOrKrI2DpgY+BPjHNvJwu
OV3hm+4TMpd6xVcOrFzgqtrTe0IbDEbuVshRbJbiUsfN/JVwMxy1nsi+BIGZPKUc
ajLoJVzYqx5jLjsmlUMn+zczyCbwJHpFe2sic0+iQ9Cfg+8MmIdv11CFvb0VyrPq
DsisUAryOXB966sn5p+uQhcPEUlW2uamp0T5JzAZw7u1fIQjMVwGZ0SIw+lWQbxA
eMGeRNI6gIS4H9OMijt0Lrhxkf6nfC38hRwl1WOjSUt4r6pjukxxbMb4PIdep3JW
rycFVtvsUS+GqHqhCntPvV5aZw5kOoG0MqOY6VMk1Cz63GcO3g6V84FAz07F89eZ
7ob6uF7NdCLb/W/vsHCrPGxnABsf9kNGwTMNTaj3gBRY1FRYgopo6fST21ciSkQF
Lusq2neLNoYJHLfUnmUVEp2DpzDln+vyD5rNcgXGhVYeJCjZTtJTcGQjvgf3eXBR
K20MHIMbT07kq97Fvs2S/a2aDvx2Lvyc2p+gC+Wtze2HjfLw1WfrIw3dhe/rmgBk
2SmArctxyTKG7F2QIPnfHgjK0Uouw+7ySzlxn/5n8n+lE+82v26ivSU25yjDxojI
V6p4ZOhx3b0Jbd24ZraNMlg8+UlAb5naCG1jYGuWdXsfbSm4EWpT/nQKormRn7It
`pragma protect end_protected
