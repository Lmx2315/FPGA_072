// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.0std
// ALTERA_TIMESTAMP:Wed Apr 26 13:33:37 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
SrJzsVEEZIH2M4uVjABj5PuNnMTINjX4HO4JK5wGmmXlHVKftLPY8uN60kQEFBUs
OL6/6I+n73q39fB0tNY+nGmkbl+//u6Yc26DsOWQoutxtqtJUAb0r0kKT63Felhy
BvjzOdamQFQHtRiJhOqZ2Vs1iPtUxWN5iGTG/Uw5eCc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 18368)
n2eb15vN7e5wAZ+MYU8ZtKFVnTH7JloYxYlBWkj0kF3djWB2lp+KwoYERIxOTGpL
xZMLJ+VVm5piKxI8NxC/m8Autv3ja204Rh78WFxHAJcWFLuJ278rurMaGoEA/ldW
mhrHF1YoY10WlqgyBcgIa4Zfj/q3L3veUFgkgbSJIVFq8XqJWRx3q02CZkT+eylq
S+vpDtic3oTxeqp/1v6cpXnhQzpDlgDBbx522AxoC4rInEWVsnJ9hAepc4FOcLvI
PYmg8XNWYljSwN5bdviNw9dBIdKbzqr/u0XncGi6qLZeIaaKRG3hiJHpvYxtbab5
oQehjeKsu9Hh2aNZRN14b0KsjBfNesDMYD40hpqO5IX9zdEututKJAb1Slf9WA1d
BV2PjAAAiI19jF9jjYcL/R0mhHY9O2qLYEjWkMP/1naDUdQIKr19wCtWDxyFlIEd
wisp+qrY2wikHSRtqslfUQLfUplRWzmfWrYUXtyO7RN9j0JfSC51zJDjm4w2NuUC
5XXm5/hkI99QSt+6XkiAmJXF8qnkszzbsL1GGWm6ksuxD9Brw//umC2uKEWWfzog
hr5sKfgOH0s9h6+5ngxVL5d8DldMc/dJWOgeVkuXI3RIaX6M2X3BrZ3e126pFk/2
8zoiOgU+xnzdPWknHD6xiOoAQx4AF6SNjkRsXF15L78/dexhiX5lqvBg4sQQ0lpf
7fIi15rA9WCLyRVMz9gi3O/UtQP6PqxI7x88iOKdP/lvTSfv/I9KTAyMbJgc5l8i
rsGRbGiOh1A4AUh+IAPVG3z7zInRKBEXZu+3nBqIDYtr/+g3MWV3idbHN+kvnNnE
MevB8y7bIfyUr0iCxOnBnCdYEXUAdWI83QCbL2bnm1+T1sQF8zElEJWVwL+xo/05
1x2NHvGmR8kvLEVD+c1emFQX3aW+K8appZxQdLiR67kgJQlojVqF4l26ECKJZJpX
L904Hv1xW3z99idtE7qLdrVgmea7Az4GxRU5lDE0jWgx3FrY56QY8yf1fu+HPcEo
FEW1eJQV5vxyQkfE2/GGMRx7oVJ4EisT0Gx/nUfZxLA4s/EIhNkVBtvzmYAPApss
9dwiCbp/stxwpYQ6PuQNQlHv/tJNXhfstYLOMRhDW7H+yBIYP+2yv202ANS//yMY
RYs6YgPkLMAe4yxATRai1UPu7RFBEOQdKOBJzoiEa8B0KQ/SeW9cQ8tZlC/nmhds
1tq6Uev/35KukR64DqqvlTiHDMqyw4QMzgq8IjMSGQd5JXxY+3fCijeLvxBHukz9
bS+nooCsttjk2OFf4JMF6GCj4SO/erJzGzwclQQslTwTBIz+ZthM2QlqGKLM7C/a
4ssK3AZIPuU/l/sYET5OyIq48hkjMRa6FbynCKeB0FPPPv2tvn6WcUtnvMjSl8FM
ThT2HVojbuoY+BAgLlF5B8i0FWsabIDKBJRZTaeG9MMYG/8T624xbQ9sPK6oA/Yy
7rjJnB6gNWwdHaGsACGsW53ydAgZMo3U6Biq7rbzcoTOagin6SwQWoLV3PxoL5ck
lq9OudJQewQArXKYwUbPsgt4YcDCeUgZ7JBvjguQqGET1IVx0CXcdePp3v0OGaiG
7QGoZ/q0sTGSP/l7HNu4ZOZgUdOZmJ755yHJmtYR1IWObbLivEhM2qr7h9ab5BE/
1i++Se4Uhkhg02Iz27W/vayPfZaLZqaFM9pecQnwrtE+oQiZK5/7X9wBIi8uq9jq
UdjBb2AI5hhijSimaNUvvgZ9lgwx4DWKezTsY+9+3PCvutaBLHfBKcTcK+H25WGH
XS8vfMZfo90T5c02alWMroh2TJ14I4IUj8FelRdyKvS6wjHI7p1YA62v8nLs3X99
x67D9bkaTq890LRfu4fIlR2HNXqt8qRszMTfKpDXhXgF9FPoeLh5mZQ3AX/Y0+nA
QtlJX93KOjfPWWd5/E0yPzorQB0tN2oBtmvRgWjWqMz5rfWaPSuSio5xXLLRtWSD
BaC6gIVVK/e/gU9E+rCEpuRGqzRNQD9F3z5YBId6FOS6QgUEmNWhHnTRAdQwXDCJ
GXsvoHr21NZtykhm+YpwWGSdiFjNaE+4OQAup7M1Rj/m9XUT91MAsMlE/beBENaT
CWD2TIzYXGxkSSQb36DmLO5P8PHImDc8uXi5oK+iipHRDfQb8QJIta4vMcaPEqaQ
Y5Qy7hLniYKTjI3pX9fUVVKspqVjdBEO8JJq8Qc/krXRgGgb2/buGaRdEVHUfNKg
HURgAuIo6R9zxo+KaSBnmooFOp+U9Xyk5egh92FNq87+bIFD30p4FWoX6nCo9hTM
5PHnfoKEQYehzs/ohAovBxXBs+uX54vTd+tHJrbely5XGCHe7PpQIFLRuJqHFph4
CSHSQDZQkjxsMcZ3LBHYHWX9vTFT+t6L6NVwskgrfMHpk/1zCr3AsedajrnuN+8K
+SHkPitdNTZlmw35v3BSbIOq7SHp3yidc0tNCOqVPCGhwjmZUMqRsPEfGBY+tnJ4
Ixyxp/GDDzJ/xYX5UXV5BEFq01ZgJ2F9wAO+3PR5A2fgCkq8Zi69C9hZMLSx38CD
50D53R0AQ0B8hTLO6jlmid6XbdjkH6VBpwOiLNR4R+vFC+YSogy+woEQpnri4G5f
KqVAk3sPM0o8Oo7jHmV8siLg84PiANS5v43KJCRNleGizCLjOJMThNu9bJSOdQQV
W7AVua6I1qNGnjiSUzqiABA+RqGYM/S4Lg3kdL7Zq5aENfkKYUUaUom3R/i7Kwx7
tDH34odkPr1cGRP4cS504zWwDLorWoR1WPSbf6SxcHx2pu399NJv3FOIefM86nn2
KePSRZdMdnNwV0usIX2V6TRPO9cF4TaeLmyV4Vtc8mvzoctbL6lxlOFyIpEKIe4z
7VxZXNu0DybLB8/IFl9Ya82nI1vp0vVoCkL/mzkg9jFSnvfM+/kttR129d6hxUti
mSOsy0HYxvthJ9pOrmLvH8aerHdmWitjPVCIwCPdLErr+R8pVBB8GvIX169fAw3h
ollA8dlU5ynwyi8ma6nKdgD24+jdJk6q37EfnSNfqy08MhMiEgq79t60+MjFuneV
kbhAqDvrinaNAHqZD980NaComRIp14R7utD+bgG3Pfztbf8fXbpstcwTPtjQIijh
9Ga6A/AuCEoTogWCMNP6nTL25t6oNyz29yO3idqSvjxKGA8BBNp9cpUWJ6UtI1dp
3TfTVUtBiRq+CCYpTmSWgLlm64XwMjBIdWSa/yZMHXy1tz+07Z+vQHL2BVNdcnsz
s/bnzBdc+V/fMRbKSZlXNO2TnqDbsYwcB681NhkReJl3Dp5djGJjjTO5M0tEZcEE
sy+0CT/oH94QxYSLELdFubepukF1Bvp/87697D898LiRrWeSdRhjigsL/u00ZzZ+
0T6t51dlF1aowE7iXu+sSj77ymat49pcX8SXG+txQZWBLAko8C9zgMyZ5tCX/Cxw
6Q2iX08rSfUwQMFOD0Mng1GDTKS1L5Hb2mtBa8ofSCoDgPx5tWeUTHB+43ByoJOb
xcM7xO1j4C8kwq3c6kQesbIYJXRVAZ2c6Xzy4M7abc0ewxuRBDTBqZcgrQJ/wY2I
89p6BdPG8MVNZZ4zRjCXAOX1jeVbB+R7wk/jaUsUBfEJQ5dUvzBq5qbsQAODgGyQ
jnhvcnm1/58bqR17q2ahiGXyuQNbs6Wz6CuD0OoYrzYOVoL+PZl/uZ4gl1otGL/+
9iL0BR8v2hXyZRfWZuwNU0AIwCMSp7ebC53jmF59bG5hvY00TIOhg/n4d1c0OUCW
+Qgg2tj3eQzm52P2+vduy4fgM3S6H81JnEW2xvic14AI+SPrdZlixMyrIRxoDTRb
mOEll9MuDohFS8PzIjsAkeolCH/StmWrOi3j+wr2vP6Jrb0qq1E93eB8YfXtO+OM
nlfUA30WPwVqXmSoCO9H/i17aRXdnl2NmJRBxtBTVSt1808M2lhO/jQZKSgW/wtc
gd9U290xSxSKg+tKOz5LWOJ9W24P/imp/kYTusSvwxrQo9tDvg/Ea1wYkniD7OM/
DGMhv8tKOgweM3BghR3gQiFq37P8bTWHUzqWy5yVRmhzSVNhTxARgyI8/iBiI6aw
7TBkLYP8wS2vqI6KOfRL8DfbzmN6d0AgZb7IQ5hVXthZ3nk49cjauWFpmPTPsJm4
K1CQYj2fuhiTlvA83gurGIgo2rlLy/TQSRwO7Thp216afTNHFKAlYmtJp+B1ibKR
2z9Q7/Q50GoUmYF/Lu07Gb5s41Vlj7mb6nRZ9UwStSoe60QWYz42bV3eJXQsL3/F
HH7McxdUUwl2LrfgaCiUTD4mQ8nZ3wpxOjGi9wLVQyEk+ZuWjEy4mvj1j3gKfiNf
/V49c3aVT2ZgBwth9veIP8aKHrf3B3LgCsgX4TrIFSW1j+nurHgoverxcZBm/NTD
GyMfuyAoixUgyEn8U5GxIrlRQcX77F+f9lXNf3ONuVkjfmBcs6n2cR1mgBXWuPM1
qRIJUaMiHIP9OjkGfwqWg98wiIIu5wPhYirjEi0UZm/k0youccsiQE5x7ErISkTi
dWiWA037aTxSm/7Cuw1pBjk0d1symocy7zNK5JvPdX+8tPvtNVZ1uxQoubLgVWMz
4KIA7IcqfOp3KBAVX58wjMGiE0LV7KMv0rnf5kvkyiZ/2iwl8gVQM92Mz+4gpjzO
TlbKnpxGdV68QyKFsd/j8ilI5pRaOe4JKejqcWsDvzvPINtMrsQWsYfd5od3Elis
WFavIu6uq9q4JM2uDDYAetG1UJQo3RvS+HB1BycwK+nm7NbvJ7JbxcAZ5veQ1GeI
kBTGMaJLZKh43kSovby8AssLr7NDl0wIrEfDF6mDi7TBA6FQahF3GvlarISTDnYT
S4VDcn8G3PX1ZRzv5sKgBAvJ0qS6uuUmss3uVQbC4FUg9Cj9/Tiib11G3zfBBVxc
16UwcxZHVf5xCA/UWAXOJtdOb9kJ2HVPwxq0zT5kcJgNKcJ9IYn9OhjzOaFhGvqr
9+MwDVQehCf+9z2J4hfo987UUaWuuGxxgoj3TUyDgZQIKKkNmUoKgrSRzGL/v3mm
AKHgI2WExqfsz6v48M88F/uT+veaC43c84dv3lEbzzAiU1PxJWcq9jnafAusBxK5
M+WfyM8jkHSHZyJcvGl9gl72N7nr5Iu5wAhib2269HuPOU3oyGAli8tI5CHeV2BY
10lAXvFxMqfAIc/RA7THsKiNMR2IkgSbWIkVsMdz7kClOzz2YfJzWBE65fIdI+tR
SgUfNTxZSYESdfccBvBUhybs1VKLgum8PCF67PsMai7pIJOkrWpXdJpA4rVginYQ
UcsTPciBE+HV4X5oyEBeOT+HC4bmLTQFJQRgzTkirVEgNESnVAna+9MzB/p610YE
s8zD56CoIZEGedQ4Pn+gleo1k5R/1FCCtAe0RgjRCq0LdlguGDIR0u9WOHvrHFMB
ercftq2fPPmRC02xyWy1M8hrGXSC4X3a+5YVYbpv3KLsL7TJkciVoeUx0s8Jjas9
8oxGTFEsuNbPxqyX3uyvGvqgKPRIl+dh79zVXKMI36rDQ2MHZ2EmhzN2Oq4IR+39
zzhS8aHJ0yIrs92vGc48DkomsZkKJyuCT+mTk/s4GjFZDrM9G0O3ZNKb8DkEJ4J1
bzLBXo1Nj6GRW0QQC3qDS4DpY5L+3ZpBtdFbP2jR/bDWT2R2So9+B/HkRmVzGyKR
4bJmLKWKkAPc5nD72VV2iUUAH8NZ56x6b8LGyllYYY+I1RcktN2PvJ0mnwTcphKz
FE3GAkYoLqtlGUV6rXUerTS1479zMEnxqjAZUR86khxVABlG3SlR7AjbKB7D3kYs
BKiWr9l9yyvlcPc37ASVKKFyqQ3KDAp9Am+5VMGcqWWLwcWwBdgAeYgxyVbzvi1U
Nh/4LVLublyAGGqUF1BQA8hPJPLt212ibkeCqi9L7A/uWYnPnLUUpCmZmffnXlAm
9XQUvjngIzeXtMwLF9K+d46DTy3BGGNx921C2yjbjze9KumXn5+q1nbyOIUPIFzb
sSdTMcw1Y60DfWk3it96Cz2/r1hZqzbmp5GrBITkAcQpPLCmE7PpewcPhyyZrtoT
sA7EafP/ql9d2lJvbKidvn8dzRinwBcFeSrdzoP5MR2NJRqYCoMGRGzyS2QWZrK5
eSnk7zwLuvM62PvKDzB5emvwUj46zgaCrGPe1vqJ+s6qTi4esVoDwkHcaw0akUrF
BvV+6MKh0WHCgV0qRwslbnU+mIhhLz4mUafMZBbggA3bRbUQEuN9GLEHUYZjl+AA
mqQAkruspTgJ9kkDmE9xqy/P9yvR7G6ZFAGSgBP4WT6hQwp+CY5x5fjLYv3W4clJ
t5Z6IQZPxttIUly505uCcAKZjWxregREsXSxE3Li3B/8bQ4W2uqUrdNmfJDh8hAn
GI8y8NYQOAKvgTQQrDmvBW7EyzVDWRGWwsbeJ2/O/7cUhNPWjygXfojU+VzL1N6y
5XqNN72VMiIyqpNR+dZ0t5Wde6q+dJYlDdpEfkemMypJoKwfwFbs/FaCqs6XSZ9J
vTBCg1QwubGjcZyGx4Pvm0LiNtdelDMMcM+hB+75mZB/lZBVlSgRbiieEI/SVGDk
dVi+/GsW81pnMPSLblKm3NJQk4I1oFfCTEMg5wmhav1ESqi23CzRlYp+O4tpGlLz
ln2JxqE9PChTczr6oiAafp9OSLrJs/sIOk0japRpjjmU3MVwS1gP1hNHEFKbVVeY
ZpgBAisWNfXGriSfBjv2r2vyotImJnExf+F+TLmTl4Q4BLdFnbPHGhaQ+n6EInKi
BhQ+6W1nMCb6ng/jTADl/G/ZFILDeAr11u5uVpP/ZL7tQKDIJfVN355O4rF+XLPt
1rINTeTnxJbkowLfspqADJZmaFFxXw4RfoK8jWNaVNfaDfLWGYViqwxICunPp23g
ZsIXqgrs2PHJQQaK6zO3+KRqCN+YvdyvzXIvN/eIQhjXKvPuOqM6oDo5gP2fq+ln
pHLqUXqlqS+PZYRAuaRfOWDcPaQLCYaTYd8KOCpFKxdM77JM3JjfaO68fkKYHZZl
5k3sSCjD+sKcH5an93Zrc0cHXVPD3XBwqPgqXvlVE29nqwW/eTWHKnLmAWLsCYHF
szppllA/9OExa2VGX22/378e3HBpxC5CaFoHuZ9cegrGMu3THoK5m7KrN6YK367B
6OZ01xBvsfbgSKTjxoDUQ7qxPGA/ufM7EsBY8iDfNCeE+CNvL80q8BC77HwagSak
NeaUhaag+1OPxqnkw0TeJdUBruvPwx4Z1wQG6Iui3rkGpPJ+CTdaTGJ4J0Ij6dcE
UJmmQUulEcsa/bXBmHJzOZejcPxuJrk1GC1YGtcG2Pj4YHoMtlaruQWLiwoj67Nf
WC5VKlMz1sxSgRyziCU8TXNIc5Xk5iKvDX5OZT30a4Nu48h0NEKN13BbQ38vdodu
62cu0PxqQX4sNSpNj8fZ1j/t3/6labjmi535e4UFebjbyygdhe57DbaWek24CeLJ
Y/wYtJmNfbysEIcztR0f1AGh2InUumk8RhAZZlCZPazYlHZxY9RD4T0m4hEAgMHN
lrmN32sIvswPMeOZ3yapliIeHdNXdWUfNXL9jaku8DLBAqdG1TfrW8+eDzx3Lfk8
AUB4DTYUMiXl5fIB9JLJi8H7+EhHoaO1ca8vi+JxxLDu5XtIKskAy8TKER68cXYK
m0PqCk9sSgOWe1npKdl5TZwy9ft0vwMAPGVj08Kv8QBu5GkrtDMT/Vg3FZdIKfpN
i/MaSQkCYaoS/Y4gFe6i77kJBBpLTNf/vutBeef5mE0AZDQNhP1GLSruJ8aEf9Ac
h9mbUXzooYfrh1OUS4saniioAq+wxYNg+FXx5vr0j/zIrNDtkFpGUJ8oChbOdy0T
44A4PE5tSu4Cf7beLFMYpUhQ07yuFBYSKe2qUhXpcfvz/YapXhqaa2DnYTQVnaeZ
cfuDVR8SIBc3wW6qxjoYKr3rUXlEQLBhT/5hnCXLwa06DR6rk3Zt2Vils0ikA1kO
xs25jVMRnb7PZ4vqKTmvoGETWvDbNFSlSk7NvpxQyrh3d+XL18sEX0vNP8DkHLuR
cauSyjpW4okss7DR2dC7J8rGkdzTRlo9ATo58g+bLBHA7RNm0SIn5AvPyV3smeFG
Rd7wkHDI97GE1EwnzmrKCQsQWnd4jaFk5ZIam87BC2OSNriNxOhI0obgcRwzfmTr
iTB1xf4BKukKhQu3Xb9lk3yfMQwPM+f30h6J+PHKLl+5fsfR+ylUwPL7Gua0BkM3
7mmvNNDAJnx1nIvVAkxokCMfazBVXbO0Dqmg7E8hyqeaSJY0UwYugB2BoVgkqI0y
7ZjnSX0vLncVtBi9UED9Ge98/7IaWIJFxjbmB/k0JQx0z292La3yChBA5mdb04Ho
otMv1Ty4STwvF+dztS/aqWwPXlLeBDEsmAux9hHcDwHVaVF7Joy+acaW930uuPx1
RZKZIWCq+268m4CraR9AZcJVXDJZw9+1hrg+QT5f6U1lf0TL1ltqEzgb7TdUXiLp
uj91i7V+fnGrJQd47/x8otghqe7ld3jgwuc6jbab/fFAX09StnDwoC9A/9xZp7NU
oah4J4FN0dnwvcjVZ+AFb48pRG/RZtTRKP+Qknh8Ec4WQOfb0bbGnmQYQW1t/JBR
ozuhsQ8cPbP5SnQuipZz473rPMYvwDZW3TLIUEq1SPdlrQvEbTqzPLK+3ciHTCzo
P8LbU4OlDjPl2iQ4JIcS4tZT/EHWYR8ftB2upZVE4Miej/m4ihgOPpx4K7kdA6xo
pTn4j5IAAxGWUMNEoYIRAQTKkAS1wSn51T/Fu6c1Z+GWqs5swd+wKhnplkm3bL18
ivPlEwcxn63KBQqBPFUTlU4fMtvQoK39tJeafZu/Arqs3OYiaClpwrrck76NLYa0
i058dM056ZhBzR7SsDXy2z9UTyQkGbmlZKCMPwLNUC+dAREhKKiGHLMhgwl3vvbH
hVRh2m0deuw4o/GfE9mKRNbvbSQAUpHNEsHJ40XjZiOxJTMEPL2qpyiULRZX1odY
53QErvGBBVAwPh1cff/w+mAVHE1nAssE2DMw3Hl48MF/8tVLSGRMAeV/6oe1JJCA
Kaqr/pxw8g8i7tpHIvoRI3HBZ2IzohDYSNciSvW9Rn8sg9M5L5LcMwlaheHA2q9J
iA7zZNzpwf47YIGOT2oMK45Mm0rUghjTjD7naMZkfDpUnWK63FeH9WrP+7ylTa43
4QFESKfH8L/nrg3e8zO3R+2FkkEEAtg8lZuGT+I14PSJ90hALkhx8afEHRCXRw9c
l8ds0ADLrL8YOwFkOE3GPLgTlx2WKnqnGmCdKMdInQSO75Np6ydU1X3rMtfg9bcV
olwhQNmXu85nZbYyxfBCnkpkaGSlZEyZ7ERUBl47+dPTk4Vam5XsvXLV5kDoZSUi
j0Sd19c3z8TBNwuX0pmDevXQGk4MYQCdWyURsLTHdpB5PO0NeZ3rrx5J3810IFM7
E/R/1MNICHzFbkA0a9tr5M3ecoBu6aklLOJVbVJmjlSqIxv+BM4FrpjsTcSFSjsI
uuEHivazU0+hJ88pG+l3oQeZaExaM2hno7Qa8PiVqcyV/y2dxf0XLurB1HlbesQ+
hd1HwuOThgRA7ZGTzvvyh7gN+0/VPNGZiu34cWAAtqIVSxAWo0MAuCNTUh8k64E5
HhXXWH3TVcLH1btVTVjH8v3pzjYSDgAPWZY4Dj01sOSCefGHPqh9WDcIOn0mq4mL
6uVXyfFMumU7o1UpnK8RdVY9XEUQG1WiYHbErjc2HUUnFSPtJi718ftfuYmEOWbA
ZuC8nWUHxyX7g0jxIuZzhV2cYovae/imTxz6mpAMdSGXRaxkRJWdIsSdd887a+Qh
gHx716HA8tImXtTOziG8A+PBajFYKAB2suN026hMGkhTPigXVSuzzX9kptQvvbq0
qpXWJ+nFM6Hdd2C5UOTx697f17EZKWUPSsZ0wUR4KtCCGL+Ahwo8iu/1h2uG7CrX
z3e8f/kHNizqUhvoXNpRpv7fAh5erFW3PMbGzrxLz5r6E9n4hpfMr5dxZUps/dqD
Jmr+v1es37FdMf3ldznu92hy5GtBK+MW++07u4HvM38oOuTqpR1nymhMZmnpFlfD
OHEoCknbcNoI3nnHNKBDx+vjpZAFgb6YbSIr9BXESIjlQrhKd+YJzy8yAINy9Gir
1YRPOTrhi93EReQYEvhcNrAI0vQbrLvxup8WbsEKqSKLGEcQiMSnNUgdI7cX4DSB
BwbibE1qRSIXzvnqCFbshhr1WzYzHy3etfNB1BgHEFU8aaCjjhRuBQBrCjLg0hYE
Umn5fFIPodZXJ59Dw2G7NhNQCnb2rPkLzIFMzdkFoOeVkN4BQNfXUZEh5Ag6kOpn
THXqs5FhLCriqeBhbuKSjAO7XDncK0CIxecIc9fdt4Cm7/GCrtwclI5cWBTL57Oo
BgiVmS1R/I1gh/Ad/ZV2rDD8a4EvRwhJ/4WC9IO5x/NZIcKEdr80lBIZmw7NjLuc
VEhEqPRuJ3MsF19Q5huH+BW1Z2ksBkbbvGri6Q//JkdXJj07qeYn/FBZqFOqdELY
m7nJ/XOVrkSM3uMCPPznPpIYK2RWWg6CgEqkzxNOYZoUooZxl8v0sXOhXO8ZAtbs
beA/FJM8FWAZx8+CItScjuduxWsx8APc/92dNxmhwm/wbqC9WvlIFP3ODJSoCOV7
/2JalzLelH30cRUEnpwOEWqO90GsA/DM7vkV7mcWThqb2bLp0v92HC78AoG4oc71
uq01KY+J85ygULcg70gpwneFIHnbVv0toiKk+va/CDUZNPdacYBQQ6BaOUkz8T0y
CG9QYDpmkms6ZgF2oJrrsEux4OEms5UolWmhU3E0SLzc0nZ10bW3Wz8QTaCvnma8
1VHR+OVGDIih0sIbJR2+mg8eCTReopHyBbKvKDjhJeQXhvISeiFKnEt9Dy+NWkr5
iLUQSvmzPSq4tXglG4F/0Axv+oKJeD8XxWQop0Wb45aKvlA1PO7Xcla7VRuqpZ8T
VImi+hgv/N8KMssXmnEFtMKkpCs1YwIJfhiUQaIHXKPm3q40SiYVoarllZF2AD6R
6obpLEqySRDdFCECazIZ9OGkfC/bN5Qaxag480xE6t0QNPv52OXJBKJaac9DPHPD
AlLKF6EmaJ6UrWsy1RdluJy1VF7fhiMqRO16456ZNc1VCW/3hPgmRSpba3ywNzyZ
NCVhOQ/RtuT2YgSkSnr2v3QMnwAwcI1zU1IxocRo9zzajz4hJhL68Dey7/XnwV5M
wP6BtSLTmujzwbXAChtzNakvi+0Vq7ZuJnnkBPcuf8lv+0U69W9kzudqqd66ZByR
iWEOiPXMfCMSiN2/LgDqMleUh0Dzx1B/KUj9G8QaHKEo4nCiifyin3hweyeptgRw
3cDELFfuUEhRO8plRx4Wkq+xVdXHJVaDkd9EL6Eeoqj+9E4EYlPoC/fbJb6r2/uS
dJM7+iF9Ci2+6J7LVyOqAB+KBitaQyFinru8KOvVQaI0j1Htjei8HCWbFiwLh6mJ
tco8eP28kt0Ml2LAg5B074qQf0ccANMLB4eBU7cj8TxGZZloRmtGjYh3A2o4x035
EPl8Hg5pQNE70fDyaY6DIG4njzms6kydWjhKbdr1KNKxSp9t04yl93+qYp1+OCgg
3MrRrjXGkFeNd/WL+03BpCS8idG7bKblP9nGewnwegPwvsHKoMzJAWXn5Ky/aFUo
GGDT7jangRGfriOUUix+oKZp5RafFP88+FmiSQcNolFF93WoTYVLSCWvGA+Q/Xg7
BTt2JpkkIcIR+mTIlPtPsvnAvwxZOoIyGl54QVsyWLJi5WKCNhXBIMZtywJsv1t2
Nj4jLNXPdg3+JusM3ezLwuVr47D9d+c3J1QiquHLAPT7bTW48oTNZdnVaG4ZQuzp
KLNHMb5V1AqIxFmFyXOxSRwJbRKpRnBIJlQPzqr8ZB+u6lhsXS1eG/eW5MJiDxij
VU4Xrp9i28A7Hy99mSoZ1EOX7Oed+gpL1kUz+vkezY47gE1MvIkCyf39cvgKv8LW
WoKwkYDWE81jWNgqlnMCXp0D1iua4WXG5VNi0/68IKnpMtoeGWBfmPc0xl1Jql/S
pBrnmDVZnAJcwNd3FRubFvuy7EPXEgSXT0bgyCBQ72DJKbryWZtH6lnWJHyhqFpS
vcfY4DNC5V/8lgD5FAbFpUxT5qXadUIb8VRFb6csrXR2Jjo9zvJTocCzLpJIY9YD
TQ6mur+GuKHErKgfMkR1S9rPgTsaLHh/3X2nfhNEeQVjhybixsc3dNrolXZpFy/6
oe7sFsSi3l5I90yZob8D8pwSnxLMqI4muKZP3JHw9vw1avhHqAg5C2rAbsQCJ2bp
j+pNSilosdoq+7sih+5Qq7MR6l5z3NxpqilXxdLHeEKXp/pMeGNSKX8vdKfrWEat
c+unrk49q1o8+0Gr/Cenp5OBpAZwJ3UG7wJqkJwDHR4/qORj1DfcG0/i+EQjZY5X
02ur6RGQEh8G9G8D4kR0tES+sLaxMmKCKTcfb2lhdjskhxTN+tyMqepI/kuazT79
KCO9s6h9BCMXqXveibw0ircTLf8gzpOAW/knu620OfQpI8IX9gWmL/c6aCQgRhkT
pOmA0hebc6B7otlZlTOacj+M0WrQceRNv9Ez9cUsyhP/dLHAEWqYzjV2YpyuZSQ6
tQd5pSfq2VaVUBsslqtWTgK2cfiwwhz3zT10/zXBjUXTnBJN6BcVq6KQCJ7sBMsk
EWzinWQuK7h0XUyKE9A4zA0bY7rYI7oLW529ZZ5rGBQdkQBsji05aLOVFeJh/OoG
gRzBd6RE9lxLMU/iJ6T7CSTuH7p5ZKqCsRe1K2CQStQJtaBuwb2XXhwii+3nkiD+
ooEkfc7uWceWWhEhz1l6QLX+3WkYahGMpJk7iPamwKCxDntCmmklrNoyS0LEWazR
mhUfaRkg5vUmNugN5qvcDyXFSHhEIwiugNFkSmgXWeSSmiqBca68JQjYxKYb6V4f
NOSAzpUGPxZP6FgXLV18Eg4ekTi3RVqoA9Nnh62TxJzcfUJLY/kEvJq3WMGc+dLv
CzSS/sAkSzRpiiD4ijVGi6hTRJs1pyHgBDUeZoyyvp1g+54bZh8UcjZS05mxaqM/
5S/14+sEWOh0pVUwIUnKM8xHnqWdHWTlAk5m/I8tjKo1/qrVvUCriJWN3DrlVNUt
dHlz7mHc60kxMpQVqs6/N8cZYBi103a2V9l4aRRpaw1/Tiy1+Do1wWjVvKYMBxPw
mw7LO3bO1PzYB3OSvfopiOcrl+peFL93ZpHKTlM1cWlb3tCIP7FD7XuAXaxn1l/u
bRidzABAqJzqM22z81KuUX9yS2Hx6ErK6mW7ORPbPcTmEuM+1uYpDtN+0nS1ZY75
GHi42c4uI5xzem583/tGcBzJ0HiDcW5KSru12vdYLJz3BtLFYDW0e+a2ZPw7CkKn
C8h9AP58uNVf722x8zMYMAr3ZDEdMKeGti4kv0cML+ksOyCWZJuKGYx7CEw7rZ/z
GRxe62sMyDZrZ77Rvx8o6DAkhe2rdywmQfW3so1x5KkWRyi+zQo2DI6MRD4Q4zfS
6npOkZ1hN1HY8M/Av1CUZBsBKfCzXIAK1y1qUp3gZArJEtORI75/jp3kXlaxc+dY
lrBWixXjn4TYdCF1/pWolKuk2awNrHMtFJoqUjTQ3ppfmYccw7Wk+1pajqLbFxCS
Z9bDXxNG3WkzS03P7EShvkiSbQSK86ElVA8V4fCAu4PQY/WbAmmtSCal1HN41X/i
qfaFizJ86fgPPQL5A76JGttk5iSjD8nw63gcB0tV5+w9SGTvD3W3sM+pbbnoMvxR
7JrLWxZfwuqvUxNXmep94d07LzwkecU35R2ISrhVcT8UJUde1JTw7fW2ygOG5pju
UzZM5HmdtnNHg1JSTyhc6Z+BFZard4Yiyty5/Nl3n9Tvgd6OT4omf5jTTjBimK1K
TYu3rIjKK/BxmzfL88ohNRJQUUQ6wtXjVGxLsd2oMWgTQaleQYHhnKld0bdTFglI
VHtknEkTJZZ8FXx43Rq7q9iT9uhZcOcR5uY3+ENlrj5qv8CXngvsmLx/W7DKQVah
5+bnm1B7McFv42kjs57iqCm03yGkXNjPl0B/B+7qbyHOvuUquP5+CWC/UDeZvrEN
eff1w+Vx0/On5tuPP+gFcQiQb7Gtt1Opm9Ow8F13HUXv+oUmB0REe4ieAN3F/q9N
vOxrS38/hzaSdfKemeWiTH70CoTPN3pQoOZAe/wKYCKq2jAsXN2qItS5AbzKf4oM
gbtsGMY6tQXAlSv3DosCFdijHpXot4vtQNfIsVWxRxzZWYlByR8pGuo1sU05raBa
X2O7qdPvbVjQF2nAzETjPQk0m2IdA0aXp1b5FTUB0YUn1dP6Tc0uTd51sl7kYE6n
sDokeqb+HzvrJug76gTqgnRQUaBDvU9A04G6YTGvIQfg5m7uO4yDU4hY0fr1aUJD
++4+24YCEf3bCdnelAobsT7WiJLd6O6r6XrrvCLLhrUdT7QfCtqSjRtYIh6NFvLP
W3gvZb1HIE3kpeqAHjJro+F+Q0+z1wW0ktaJh2xk31HDGUzdXp/yOb6A2KDEV4ED
pnbtYM69sv2N9OLZi/eFoc3czHoyf/6Db8eoilFQ5IkoootIFsPdjTtTgndQ7q/R
bUnwPmamlIvXF8tjfMJoyzS60+1vyspKtSimRfQCFDOSFtT9DbtUCuio6R28vZ50
3feia8IUphxMeeLrowtHZAWxoK+Fq1DAXA/egEiXgoY6DKq1BIohs/PfqXXnAg5+
RSTloTjp2wNUNoNgGuwFK4vE2bmYmu5Y9gQEUFHfKl5qw82PmnI/48GrpFR+B75q
D4/ugu3OrYoqtWF6UdPAO8YEyveyiNJh9lsC8UF25GMbyndDf0xV48ooK1y0330e
AZIrYXYdg/Y5INen9ikvJab8P8lSB5vz+FOa6Fo7IXeSW2wF2NRStMneCoGDbACd
1Aoe4DGgTLhr3KmB14BSq6m6Fqq0+838DcRtTa7FpnGQ4irUd1WXzJmJ35kK2+z7
0nk00UqVW6xSuiKoRFK7dKZOxEb2t/Xbk5qtNvP74e0i0gDvAWhX/DSz3xNZC0Y5
ImUrD9sAMo9j9jGPCVZi1pW94louk8UAzJwCE2dfa9etAwT7470R4Xv3HWdOo1rf
xn+EHKFPm2+Z38IEhvyKx6yyfNeB1RsWHDpyGUsaklMFYHirg+qYX9Dul6YzSGP9
BY+qxCiMmxkjCK/C5IPnnDXaiHcX55MZoaHa6cOJzKp5p5tFoOIvwvgoS0oQJ6+I
+MFUUuhmjRkgI728VvLc62ijBf4upnt2t2ZmimjVX/jRa3m/X2T0iq5DWCyx199P
qlGymdbYSgjSnQPB7spAbNWuiLKeHhuMdUyTQNLPon8te0lZ5N9jn/vlmAYO6J9e
ob1Zr4RpeslKetDabv9FFMLD4JsCBzOm8nNLIC29cytK9eSgGrhZNZruHSzsI1S5
ReiBewTnwW8I1byYSE5cbGA5dbSwNbnmkuOrfCT7pyTL9et9CsIWdwKa28r8vPvO
2HeSwFQ+v7vlUZf/hjsP5KoUNiPFrzGOmzrT1sKTi5/wzJDr0IPUddslDn0E9oac
e0iQ20BdYYNjbQJsLfIou56YZ52WqxYB1SmJE+0M5hOzCFzfaJmjGVvjCJZL/TFP
npTq2YllpJT8ZsJIy/17cLHM8gyf6ZfiY5TKVfdaLrKAwBGBSONu8AO5EFFPo3Oc
Uq0lFTEcW17KUDwNU2vpRGwlu3A2eZIicPqCe4xu/qBACZpQfHIfazQHKdZzRMyU
Ul93ZQk2dhm9TEiIf3Ozjc7/3WZS71y5pkMcVwDVqWjHbRuifsBNBw+xvFovSVYv
ibW7hoioyJyCygHjAMB8uobZQwE6EGW/FNBQqECk2KugHrt0kLp6CtYJrSQ9kvbF
aoObv+3JNCDfKVk2VRCdHjGq5NBE8cF8UbpxnzfPXIA6o8bjltFmx9I75iYoekxZ
QNnt84dSSib0RbmcIm2jg+x8JjAmZh4zmAyA9qHHIiZogaZDIfI8suLk8t/K6JIs
J8/hM4n57fLZgHd86uIZL+xg5BTld3kkGiwVdzg2AHu6wTVSARkIKdsWsvbbaLTD
dXF5vC+o9eY5XI5LEdyRHy1CqxfSfVK1P4VBKnI3Unf5eM5fybhKFGkJ6dIofJTi
/R7tTJ3ehsi3Irop4qA9ZYLSCNCsjHgRyXt/lH5MxpfIFhJiyEnLVQzGmfvkqwuh
uIgHiHbsV9Jcb7147a4cfGlG7RRJhsiA3T2sitXtBqzGSlKYx6LUciTrNk9Ntq/8
D1NT46FyK0AR8oPvTepbFPIt7+8qj20g7TlUfSd6qkhn1agvSpOj9nlZ+JJLT9CX
tb27jWVZ3svyyHcejRkUa9+z+432Cyf2YRxH2oixkmGrbAITc4VIIwka9XrZLFuq
ov0wuXgPL5MUkBIQsZwAmY0pFz4FIPuwXuqR/CXXbKAhrkwPY3yE+hoX3/F1rKQV
QhZEUprQK6SHVb5SZa1AG4zoJOL7nMRBqoworZBSTJXL2pQH6tExe+C+aoLUBUv5
t6ZCUw2wPVh70/9tdnHgKsd/3g3JM0RPevjcqADP949nJq1O8tC+CSLxjwBJTVJV
UMPNeC86Q40wCcXz3OgcBmW39ZYiF7swQZ3XknmPS1Ifhl7ffUqdyEfXLDUA0wLC
6smve/rTaxDePmof2lfkpNisC1xUFVe+wP0OtvmS2p5ETKayYRCbsV7kP677IB07
KXCb+rlIQ5FIwKL92W9/WKII4xvL9Yue/PrqyiDPCK4vJQyOd9WSZCwq/b94CF5+
wHSMq+HwmIp88ZiieRI7VApW0sL1xZ2nsvYfhinQA/b9MDFH/jWo8YWyxz/re7sg
Q/PWlhsvPMAaDGK5NJufdklQfZyuvflLVSfEOGRI46MiYRx9EstUEYvTA9SzR99f
H8msu2Zc60zddmicMsQOfvFWDXwL9XPCH8s9f2FGPA9XCeyPJasmfAQKs9foz+ze
+cmr0CLdd8JgA/tyMvgsKGnG08hnQ/Y60yRKuchMCF07SU5WHX07S4ZqpGejzflX
NGhxvIa6e3MV0ltMxlC6288LBgHHj4q5pp0/uCAUtsjRvo8zc8Y6LTxDlrSsEhn3
3u2IImp1yuzkSdtTv50hyRCV/zCnmNe3PZP6XyGUKQ0oZ1ttiqrEb0ba+n+0Nr5N
WFM3iPDuHZU7EVlj4MT9DiRD05nfMMcBfrxBVzNesXksnlRaUYQbUmyK04QYAHh9
5zMGwBsdJKWtEt+TVVBUDWGNKlBGPYi20vYYupEUjMkygrvUr038Pck+HtjW2U7W
QyCcyN18qEkQPFAODwYCoI9NP+wuY797wEvSF8Vy99MtScCo6Or3GY7F8Z9hEWVE
54fT5Wi99f1U2vSnIbqn+RO5bdzkQXLan51oD24WA6+L7A2x7iVHGSnuC8mFKlbp
aY/4Wn7F7rUuSR91s388Q0FF0cg4C56j6vYhUvafJWJuvdGhZaqHgoQG4H7+/K3r
UVjihYm37DfxLzer/dp4LHtGJLJGs6rNWny1vnuZLC9U1kBDjOwo28yLp/J2lWCh
cafh8mqaOyT8uqdQlkpxa+bJZDXUQTCpkBAc9d857CcP5Uh9MVpKZbxSSo4d+6IT
MvPxiNg12T/tDIAYd705f2XmXkju3aepPo6J/+T/8BhelIHxF8CNCDuJddWJkdWi
NFLD3i8P7V+7vAPDjTSgh7UHQ2Ex4T/8JrbTISAQ6nrgCBKgPpWGYJ+m1L8nM9NH
4n3BFsvQGBBYcwQAO50izv3FgQP+5FqVNpXq7exZGyQc5OamFIWT1c8pyx+tzjWL
wSIvtqTxb9jP3YH43yBSO4IeXEAeA7nG6Ggut4M/o/YDV4tSICMtos5M8yxFuC0i
fmeQ8l4AjuEZPQSrtQAzKFn3XW5gg+NKOaqUJXrJ9GySS5hqk81ZtOsvzF0uYnOi
AZ7jIaAhdaiilyP4VOJ4sc94CV22eTF1A72NN31+HVXsaX+38/She0Hlw6dA5fFZ
k4XgZ9g2+AGQmwBBqSOZUUlRpXyFBJYzCBZHP82Q4cTt4lnWA19CUMduNxwruu7F
i79HEmQKQVZEinUwk9cpC7Woug4sBsZv1sgw/xUDRNTTJsKTLO5jW3BFTBq//mn0
lJooh7JvX4/i5xTkUptqB9J5T2IypEHv6bsCJUMK9R0Q1BvBwWpk4JHGjMJLYwbV
iBoFpOpzw8CodMewDgg3C8HhOul3ZuY0f3Y3oRowcCyC+TBMqu5IBjm+9lZIrxfu
an6HKYfWws8evp4MBDBK57+gsmOR7Iw8Q5MYXbwiZAfYTbJ3jJGSGrEsfR9p2ELi
c1KMozBwQVjnBPxNZR/n/pp2u1btcXkOws6NNg5hDqla+skFIvb8SV7Csg6BIGlU
j57mKVfB1E+6vzhQd6zWUkOjwAoKz9MVv10SzI/Xfb0MWKuOq5kydflWzaj5nGKt
awT6UJYdge0JBepyPUPJlZMIWYgBplZ7drggZAbJWBw0raWUJj6d2795OmZXpTwv
hgJTl9FFAz0XyMv28YcPtVQ6AdKun3a6aO9CrdCHT9Y/rWJjJw4+oFGGEqK58zFM
QnyMOdZ0yC1gn8wLsmJwvt+lV4FMlZj9/VB/kVDj/I7m3Ak2/uJ9PL+i8fpwHTA6
EmpKd0uy0kNSctw21/KCofXBWyUoEoYKbsnWILPGx9DslrePERxPFJJXhAkZ475s
DfT0wDq3ppuMBu3E5ywOcQmFsq6EwfnBICV8D84e1qgJFs6HCMcnOAX69iwYHRyw
T7J0mJ39MCl5+WuDPq+r5rtisdCavLw+OroPgP8QmVmpEL1sP7qWR5oPlK19eFpx
VBiSGODWo38o5QcDdFkVeY6jhyOxpxdGcnoVgwF95lQKS3ilysQ09hgHPmYu2hX8
2lFD2BReiIWJc0azZYjWARoi+7LgQuCz8pLlp1gpwaIeltIIm+N+/UPoOnmji2ZY
0P4nppdUeykYdGJzJpisZRYzvyj+3V2dQ3q3R2nKk6J8LmrxTchTnA/c8BYsduDG
Q8V8u9oDGGsCuwaDFjfhoXRm80P4o+MFyLfGBXkkP0f4Zab5IUqMQLB0yJHQNmRQ
b11dhYAJenVOGgWP6ZXEFK5EDiHaJgACzTFpGYfwcWHR9nYPvVverwX89v/oi7Kt
dHCdAwieznfUMwO1/Z+viCewabBe/co5axmafDlvvOY/58B9V95IQXDa3RPi7lXw
djAyqeH4Wv8faHxm+XHASp6bGR8KFCE4QlweVVJc6JYbGtB532AXGPxI3x2/xcCd
2PLUniarnWfgMdQOJc1KTCU3Ap9vcJS//or+C5A7Rv4ZpfCS09YZiy0q065pKtzN
txaeUOPSzShOGlwQ7P6xKQsolxyxBzc3Ul3Kj6eP/+xHGlt2Oz/eSuGonkmLybTX
I5YuM3kgv0p7M5GfS0j19jBhGw8xS9pywc5axFRIP2fMm9JF/ifLXgAO+TJOVcWf
NHHlTZvO3rSHrPbiCwibVFj1TXWztzOxz+DRMK0w5O/b05QbGGnLCAS3zUEvuu/l
zYfmVhKYvQ3palcb37Aakl6cUd/mCZt4+9xcRSbcVNGSfS65jjAZnDnY8jr8sNvU
5HBOKBMwGCBUd69R6RefD2YgjC8UZmVaIig2PsDlR8F3RQgYl4khvVEEl+2DWiZd
s15d1ukSBxZ51Z9e+qmW2Ews+GUPdpWZB6us5zGvLkzM8pV6CYdJQ7qyuQwV7PjY
P18aMmQU/EoXzVfgwIJThjYWWzc3K0H/VcjJ2R3N/JjQ20FGRhh2n17MyHWAKjub
pBumGgmGq//cDioAqre09JpZ8NS4xy9Wj49XaLdBOqvH862HCnptP61nSoP6qFVS
NcRKdCg/skfy4Zbwziee57L0EXHFE4+uYmiAhxoWYr+ThGviLlCwFOEuyxe8uwfb
uqB1KjHVLLNSJe1AGp8Xi2AkVPTkPd20kEw8oR25vOVtraHOl6OXqtN7brMtGlAP
uAYzjAhMyZOYR7sY2FeZT03onND4Q4r8Ub5QlCf22ocEAx9ZxaJ05efjIqf51c0I
Eouu/jCpUyzzFEURf//15VmrISSjr8lF7l8Eit2H28LSRMLLxi5nM9nwrLvAhWhG
F11p8R5ER7IwqezvaHe04yu9ig1Gr9OvQ2Vj1s6YYgJATtqYMLVnMMBAf/u5Fbne
BrVNwNRMaxp6NA0qri1/Xy8fKu/SJbqNFsec+qxX/znMC3sLJwdA3aWc5IrXFUMU
mI6d0Yg8Le9tLU6VhxFS5aMG4pNvL9/z2CXKw9AkraLlamxYTaA4ktvUSwKqBxO5
+BVWbukF8ptxAuPi4C9OTjHf2NC6w+H8mqCIo2ByNMI8mqJlKHPoauJT9jUfBLU9
uWo40YcL3yON5L1RejZzVlp2dIfqHLRPDw3WmSvepi61h/qgbBJf2tl0okpM8mx4
+SCTQSoYgeBRyXHpWBJu7df4NhyCULnAIcv/9PxOFYwSpj3WEPQfGAP659CGorva
uawAhJGgW2gsvcsm56qqqg/G/Tzc/EFVEpiij6gugkLXr5Cc+wP6cz2VE53+5Mb6
rmqAQ/CTtSVe9ADu08PmpRkAn0pDo5o+2nThcQPCIZJsdoGTxOd2G4+tNOVIewDR
4u+CBbbABfKay16JlwCrDovXQ9KXQ8UCsonb+7K3YqVHtSx9We6MREE578w0cWjg
3eNN9HZVJVnFBOgl0DCusaOjDEWvJ1UE5zinNx8BXSvzDqS+oBLw8u45mB+94Ktg
tk+dmiqBg9FpmPUGDvHtctMqhJUBFahIBx7QCLcsNdoEo9NsAlADzFTBYpajz+9F
Seb7HbfDG6f5VdG6rATSWb6WYDOTbICbzabpoErqRSuhxMV6M0HdJ92Z3AgYxBeq
9+DQpgh7cmBZirTJEsuVxHlo/Q/PrYLZwSTUsN8e+zJGfuPOSrS3jMbl2/hDEort
dkWmlRKJibvGFA9L62rZ+wCvRf4q98cYByqs49LgK9sMgReSs4F9xz+GR/bl71B2
W5O/joETyTaMeMNPa2POYF13X65zop3FFpGbLRVZ/beSu95CrttoywPFxrlbo+mu
lrQHYII3PgCaNPT4K/hW4jSnRnKmfg+0NG4UtIxi4j55vdcdsmIUvMtctvK1vi8W
JjbnH11SsafcLdPduszB2BYYfbSgqYvEgp8JSUvzM5aGkW8TwLyQIHg9GznN0b4Q
jnBh5Sl22kzgBB52r5e+iOX7TGSgCaB3+i5FvpMawqBrpQb/iplG62lC5dBGonYy
OHCgLnxz9DPVDDzrp62sztQl7kO64+J9qqjPIEpohGN4yqa7/GPCn2HlYKaMWxIX
jlvypOPk+/OFnyy0JM7huFFzFGp+cLR16I4OjJkgLQoffP845MAKikXOqg/SKJIK
T7a23oFubH9GO8iji3a9y1+BA+ZjNL5TqN+7euLYSfI6PCPGG0yheH81UKvj46lj
6YiJ0Qns3sL6KW+25fLi/1GLfFg2h1UDOkZRWY0RUKvw9gm6FCW0I/cxlL0TRa+L
zZ37or8mC31UaQ98rS3NO3XlxxnLs2aglmpHcebz7AnzBiJUb2hIl5UToyEFAK2H
/AisAlldeCn/MvyOdf//cTPSZ2qoghRDVoQc+paa1xiNYT3J+siVBWw7+fnHdYb/
/3Ux4CoPTp/7K0NvZ9STJEFZ09bFde8tz+s+9w3ex35hNyHDhx9NvM3j2E+vSb0U
qLFcb8OvzFM+RG6Rg5HG4Jmx1OertRIPoqpzr8PV5QfW9nGET4JsXTGJnqVI3GYv
x2hRmA/qYLEnVzDm4v75AYE6RHplGoCHyfKn7LWbuWX+Zp7jIX0N3JPMvrmjtdp8
+q3r/qxCJjAhqa65wqoJAm4RsvzBb9pCiE9x57JZKMQTef+d5psvDIb8qLJGr0TC
SWVmGtSC+bJJ61kC8zh12GGK2izuNduTNwVN6l6H/ii7RwzrQMdykcBwdHhnHF7H
pED7ubVdZlETeilvDpAngWw1Sfn6EEprc4h4Le7VDnMIV06CpWdE592Yei339MJy
xs/mRP/yrBFBrDOhVQgKvRHS27/6JVtxL+bbZhFuzQb3WW1g2DVXgcccOdmktKJt
hreYiZ2vcUCjIHmfYw61GKhRr9ZN1SvdMfslLM2akL+GgfJ7ijPfwwnQnuvoC0RS
lbh9PfWO8vw8mo3xMb6zppM0CpGs8vWXov4NH/bgw5SOukGmiluCRapsLsgq4yXt
G8KbMZVFDZhBEEYWvyoMdzkDTJPKpJDFezyYFUkvlLDTqWEbAuwquWFCU/avuQVT
pz4J1wz2cSRTuYEW0uATgYLyGxHU1e+FQLjgUWUlaUW3wZK+Tv3nJOztFOMEI7R7
dOE39BOPtufinm8hbXL/TmicA1LaoX9DcD4OaIN9uBGya7QWLBzIT8cJjW5Q66lx
A4emf3lbc7CTz83ot+awT0lHbKuBtBqR3chaQfSIJlUpJPn0ZuDEEbyHpF10nlEZ
kIKWaU233f6hEJTUi8gXu1N5GRZrDnECzQU6wz7YTzmzAHrDeDS+Z6be5DYC6YfB
lkKLaowSAOT5Q2WaRTZP/nI15IGeZtFWDOFt1pz2mnUIuEXRgP6xt5E4u6pr7lk+
WSB3JlyWja+Mffhk+iihcK7VypiQgCyTILS6vr654E2VUTImO2kTsiSVIQ4jZE2J
h2qMzX5VVUBXO7FQxBUI/0p3+O/vfUjjzGLGlhNe2QClLQBum+MuTtyN7VOYV7Bc
P9CIFG6q1w4GxShEFBI7lS+mW/MAgx227+EBRIxCIyROPMBm1US4J84LB6tvf4fU
2ATHQ+/FT3mVnWrZ9Ooo3KyyZMtnXE/G+kRMjXRGn6QSBt6B1DV6Qtq6uMRX3S0O
ioPVTEuiZocO98kD8U2O2wIPe5GFBGL985gQG1BbWjUZ5+Im0cQIpKdTBaz45TP2
ZO3m0XA1oK6d0r75FH+q5YsFeATG1v+UBQvXnJ+3TWHbuQYrNd2TKQp9Q/Ip3yOY
ZCdFgqq+U4hnnTKBbrgv8MWMfnQCEXOHTkBAQGhegdK/N38KrrPXh3On8X28lgzJ
kYIxaUPDHIbLgaIwq0Ecr/pexPUM93l3LfHON9mVLIZQlH2QWCPCLM4T1+xdRtmI
Y8f6FErTexAlIPUIDuB7oqkTHg00bfw2o/bTHRKavrZygz+npYJY7ZY6dP4bnoT+
J9zH0qUYnEvF/HW5Fv2RQe+XofxskGEud76Zer0hplspxNHglrSegSVozgKHCXHG
8NMNIkGUopcDJJeBwmUGVEdF/N+Vi9AxDdmMRCCJgjXFCKnVdFOhNfgeG1+bSVHd
wU+S5GfxneD6VG59vsVmW2oYzqmfpTxM+CXrBKFYqzBQB1wPDGvLCBUHW2ZZi+MT
5aTDcfLpojVePCgnOa+rxPFAT6+vlqD9XKf1R790HWLxE0gEJtqMQ2UQI+VUxqUB
GGFNxGOAYNR+fB6NY/jnraTRT7+XO1LLh5MZHRAfysw2g+jFVKK9C+PbamLvFSdd
q1N2O2hoU7vAKKUHcjaCWNx+x81Yu4XYIIBCHSHoZqbgUHn/yRP/8Ev9UFZh/oGY
66gDOgAtOMMPBHkqHmAw6cL2VJuyEF3DKNg/4BLmMkaPjllCwOe0niJSbCps2VbT
5WDcev9HCo9ITeWvH6sZDTaCZ9CS+lp8FtCGgIVmRBMYjRfWMFiM1Q7350NS04qB
0K2tBZMoxs+fK7jN+Vk00sn1iFPPCLFhzT3E1JFuQ2uJYlRauYT5dSc2IqDEYWof
yxh6sGm1iiQrJkW9ufEyCS3wa784C4ITbUvbDhXaevS9WcuUZsRkLxCkcTSD5gKp
YOVG4FV8ZOZ6PqrRKEu5T3LiED5spa3cJ+BxqAtVUV74TRTA34tUPkp+hPt4Ifvt
HIZylSYZpICrNTYZVBt5vmXTyEDOXUx8R+hFP3/f1oXzOA0q9kKNsDGoTimHjUqF
QzqOdqGWUoyhEBkxHGR5dAdW2XU6N4gRM5xvRMCTSQ/H965rmRk4g3PZ7X/KjUDo
Xs2Av88l5DJLrzJvu7PP4pK3MJAxYo7Jevlt6NK8u7hjjk3EiUGg6T3/UQgpp9eh
kpdH5mH0rWoaeHTHoz8UUqjBR635oAMIUPiCyBSG+hsmV8QrJxGniOrg0ypmZFvZ
FA3LvpzCyXiIICsAJntebKuIZPMTX0PHlPL/TMMi/5gyl+Y5ujzhmZeZTHXUpsX9
RBG4EcxXcXJ56mI1Tnwtvlivu5a7WM5UQFrgh+2anXusBTLMFgGxnQxL8MSdCGl+
NzyKSHoDX2oXLDwFFb5Q3VxEr9eP5woR6F917rb6+0+8QmaOnc1d4YBDa/A3BHe6
yvMSwcrN8DRz2wi4UshA2ilbJklwsS1wfpMdXRyZ16pgR1kXq4E+Al3c9tf5cNNW
MSICmDqHyQFKescUE32tvTwT8szefH+SMkc0fISUGEg=
`pragma protect end_protected
