// Copyright (C) 2018  Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License 
// Subscription Agreement, the Intel Quartus Prime License Agreement,
// the Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is for
// the sole purpose of programming logic devices manufactured by
// Intel and sold by Intel or its authorized distributors.  Please
// refer to the applicable agreement for further details.

// VENDOR "Altera"
// PROGRAM "Quartus Prime"
// VERSION "Version 18.1.0 Build 625 09/12/2018 SJ Standard Edition"

// DATE "05/21/2019 10:48:37"

// 
// Device: Altera 5AGXMA7G4F31C4 Package FBGA896
// 

// 
// This greybox netlist file is for third party Synthesis Tools
// for timing and resource estimation only.
// 


module cic (
	in_error,
	in_valid,
	in_ready,
	in_data,
	out_data,
	out_error,
	out_valid,
	out_ready,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	[1:0] in_error;
input 	in_valid;
output 	in_ready;
input 	[19:0] in_data;
output 	[27:0] out_data;
output 	[1:0] out_error;
output 	out_valid;
input 	out_ready;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \cic_ii_0|core|input_sink|sink_FIFO|auto_generated|dpfifo|full_dff~q ;
wire \cic_ii_0|core|output_source_0|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[0] ;
wire \cic_ii_0|core|output_source_0|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[1] ;
wire \cic_ii_0|core|output_source_0|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[2] ;
wire \cic_ii_0|core|output_source_0|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[3] ;
wire \cic_ii_0|core|output_source_0|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[4] ;
wire \cic_ii_0|core|output_source_0|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[5] ;
wire \cic_ii_0|core|output_source_0|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[6] ;
wire \cic_ii_0|core|output_source_0|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[7] ;
wire \cic_ii_0|core|output_source_0|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[8] ;
wire \cic_ii_0|core|output_source_0|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[9] ;
wire \cic_ii_0|core|output_source_0|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[10] ;
wire \cic_ii_0|core|output_source_0|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[11] ;
wire \cic_ii_0|core|output_source_0|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[12] ;
wire \cic_ii_0|core|output_source_0|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[13] ;
wire \cic_ii_0|core|output_source_0|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[14] ;
wire \cic_ii_0|core|output_source_0|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[15] ;
wire \cic_ii_0|core|output_source_0|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[16] ;
wire \cic_ii_0|core|output_source_0|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[17] ;
wire \cic_ii_0|core|output_source_0|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[18] ;
wire \cic_ii_0|core|output_source_0|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[19] ;
wire \cic_ii_0|core|output_source_0|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[20] ;
wire \cic_ii_0|core|output_source_0|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[21] ;
wire \cic_ii_0|core|output_source_0|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[22] ;
wire \cic_ii_0|core|output_source_0|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[23] ;
wire \cic_ii_0|core|output_source_0|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[24] ;
wire \cic_ii_0|core|output_source_0|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[25] ;
wire \cic_ii_0|core|output_source_0|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[26] ;
wire \cic_ii_0|core|output_source_0|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[27] ;
wire \cic_ii_0|core|output_source_0|source_valid_s~q ;
wire \clk~input_o ;
wire \in_valid~input_o ;
wire \reset_n~input_o ;
wire \out_ready~input_o ;
wire \in_data[19]~input_o ;
wire \in_data[18]~input_o ;
wire \in_data[17]~input_o ;
wire \in_data[16]~input_o ;
wire \in_data[15]~input_o ;
wire \in_data[14]~input_o ;
wire \in_data[13]~input_o ;
wire \in_data[12]~input_o ;
wire \in_data[11]~input_o ;
wire \in_data[10]~input_o ;
wire \in_data[9]~input_o ;
wire \in_data[8]~input_o ;
wire \in_data[7]~input_o ;
wire \in_data[6]~input_o ;
wire \in_data[5]~input_o ;
wire \in_data[4]~input_o ;
wire \in_data[3]~input_o ;
wire \in_data[2]~input_o ;
wire \in_data[1]~input_o ;
wire \in_data[0]~input_o ;
wire \in_error[0]~input_o ;
wire \in_error[1]~input_o ;


cic_cic_cic_ii_0 cic_ii_0(
	.full_dff(\cic_ii_0|core|input_sink|sink_FIFO|auto_generated|dpfifo|full_dff~q ),
	.q_b_0(\cic_ii_0|core|output_source_0|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[0] ),
	.q_b_1(\cic_ii_0|core|output_source_0|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[1] ),
	.q_b_2(\cic_ii_0|core|output_source_0|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[2] ),
	.q_b_3(\cic_ii_0|core|output_source_0|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[3] ),
	.q_b_4(\cic_ii_0|core|output_source_0|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[4] ),
	.q_b_5(\cic_ii_0|core|output_source_0|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[5] ),
	.q_b_6(\cic_ii_0|core|output_source_0|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[6] ),
	.q_b_7(\cic_ii_0|core|output_source_0|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[7] ),
	.q_b_8(\cic_ii_0|core|output_source_0|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[8] ),
	.q_b_9(\cic_ii_0|core|output_source_0|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[9] ),
	.q_b_10(\cic_ii_0|core|output_source_0|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[10] ),
	.q_b_11(\cic_ii_0|core|output_source_0|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[11] ),
	.q_b_12(\cic_ii_0|core|output_source_0|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[12] ),
	.q_b_13(\cic_ii_0|core|output_source_0|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[13] ),
	.q_b_14(\cic_ii_0|core|output_source_0|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[14] ),
	.q_b_15(\cic_ii_0|core|output_source_0|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[15] ),
	.q_b_16(\cic_ii_0|core|output_source_0|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[16] ),
	.q_b_17(\cic_ii_0|core|output_source_0|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[17] ),
	.q_b_18(\cic_ii_0|core|output_source_0|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[18] ),
	.q_b_19(\cic_ii_0|core|output_source_0|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[19] ),
	.q_b_20(\cic_ii_0|core|output_source_0|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[20] ),
	.q_b_21(\cic_ii_0|core|output_source_0|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[21] ),
	.q_b_22(\cic_ii_0|core|output_source_0|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[22] ),
	.q_b_23(\cic_ii_0|core|output_source_0|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[23] ),
	.q_b_24(\cic_ii_0|core|output_source_0|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[24] ),
	.q_b_25(\cic_ii_0|core|output_source_0|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[25] ),
	.q_b_26(\cic_ii_0|core|output_source_0|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[26] ),
	.q_b_27(\cic_ii_0|core|output_source_0|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[27] ),
	.source_valid_s(\cic_ii_0|core|output_source_0|source_valid_s~q ),
	.clk(\clk~input_o ),
	.in_valid(\in_valid~input_o ),
	.reset_n(\reset_n~input_o ),
	.out_ready(\out_ready~input_o ),
	.in_data_19(\in_data[19]~input_o ),
	.in_data_18(\in_data[18]~input_o ),
	.in_data_17(\in_data[17]~input_o ),
	.in_data_16(\in_data[16]~input_o ),
	.in_data_15(\in_data[15]~input_o ),
	.in_data_14(\in_data[14]~input_o ),
	.in_data_13(\in_data[13]~input_o ),
	.in_data_12(\in_data[12]~input_o ),
	.in_data_11(\in_data[11]~input_o ),
	.in_data_10(\in_data[10]~input_o ),
	.in_data_9(\in_data[9]~input_o ),
	.in_data_8(\in_data[8]~input_o ),
	.in_data_7(\in_data[7]~input_o ),
	.in_data_6(\in_data[6]~input_o ),
	.in_data_5(\in_data[5]~input_o ),
	.in_data_4(\in_data[4]~input_o ),
	.in_data_3(\in_data[3]~input_o ),
	.in_data_2(\in_data[2]~input_o ),
	.in_data_1(\in_data[1]~input_o ),
	.in_data_0(\in_data[0]~input_o ));

assign \clk~input_o  = clk;

assign \in_valid~input_o  = in_valid;

assign \reset_n~input_o  = reset_n;

assign \out_ready~input_o  = out_ready;

assign \in_data[19]~input_o  = in_data[19];

assign \in_data[18]~input_o  = in_data[18];

assign \in_data[17]~input_o  = in_data[17];

assign \in_data[16]~input_o  = in_data[16];

assign \in_data[15]~input_o  = in_data[15];

assign \in_data[14]~input_o  = in_data[14];

assign \in_data[13]~input_o  = in_data[13];

assign \in_data[12]~input_o  = in_data[12];

assign \in_data[11]~input_o  = in_data[11];

assign \in_data[10]~input_o  = in_data[10];

assign \in_data[9]~input_o  = in_data[9];

assign \in_data[8]~input_o  = in_data[8];

assign \in_data[7]~input_o  = in_data[7];

assign \in_data[6]~input_o  = in_data[6];

assign \in_data[5]~input_o  = in_data[5];

assign \in_data[4]~input_o  = in_data[4];

assign \in_data[3]~input_o  = in_data[3];

assign \in_data[2]~input_o  = in_data[2];

assign \in_data[1]~input_o  = in_data[1];

assign \in_data[0]~input_o  = in_data[0];

assign in_ready = ~ \cic_ii_0|core|input_sink|sink_FIFO|auto_generated|dpfifo|full_dff~q ;

assign out_data[0] = \cic_ii_0|core|output_source_0|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[0] ;

assign out_data[1] = \cic_ii_0|core|output_source_0|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[1] ;

assign out_data[2] = \cic_ii_0|core|output_source_0|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[2] ;

assign out_data[3] = \cic_ii_0|core|output_source_0|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[3] ;

assign out_data[4] = \cic_ii_0|core|output_source_0|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[4] ;

assign out_data[5] = \cic_ii_0|core|output_source_0|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[5] ;

assign out_data[6] = \cic_ii_0|core|output_source_0|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[6] ;

assign out_data[7] = \cic_ii_0|core|output_source_0|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[7] ;

assign out_data[8] = \cic_ii_0|core|output_source_0|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[8] ;

assign out_data[9] = \cic_ii_0|core|output_source_0|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[9] ;

assign out_data[10] = \cic_ii_0|core|output_source_0|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[10] ;

assign out_data[11] = \cic_ii_0|core|output_source_0|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[11] ;

assign out_data[12] = \cic_ii_0|core|output_source_0|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[12] ;

assign out_data[13] = \cic_ii_0|core|output_source_0|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[13] ;

assign out_data[14] = \cic_ii_0|core|output_source_0|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[14] ;

assign out_data[15] = \cic_ii_0|core|output_source_0|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[15] ;

assign out_data[16] = \cic_ii_0|core|output_source_0|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[16] ;

assign out_data[17] = \cic_ii_0|core|output_source_0|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[17] ;

assign out_data[18] = \cic_ii_0|core|output_source_0|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[18] ;

assign out_data[19] = \cic_ii_0|core|output_source_0|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[19] ;

assign out_data[20] = \cic_ii_0|core|output_source_0|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[20] ;

assign out_data[21] = \cic_ii_0|core|output_source_0|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[21] ;

assign out_data[22] = \cic_ii_0|core|output_source_0|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[22] ;

assign out_data[23] = \cic_ii_0|core|output_source_0|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[23] ;

assign out_data[24] = \cic_ii_0|core|output_source_0|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[24] ;

assign out_data[25] = \cic_ii_0|core|output_source_0|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[25] ;

assign out_data[26] = \cic_ii_0|core|output_source_0|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[26] ;

assign out_data[27] = \cic_ii_0|core|output_source_0|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[27] ;

assign out_error[0] = \in_error[0]~input_o ;

assign out_error[1] = \in_error[1]~input_o ;

assign out_valid = \cic_ii_0|core|output_source_0|source_valid_s~q ;

assign \in_error[0]~input_o  = in_error[0];

assign \in_error[1]~input_o  = in_error[1];

endmodule

module cic_cic_cic_ii_0 (
	full_dff,
	q_b_0,
	q_b_1,
	q_b_2,
	q_b_3,
	q_b_4,
	q_b_5,
	q_b_6,
	q_b_7,
	q_b_8,
	q_b_9,
	q_b_10,
	q_b_11,
	q_b_12,
	q_b_13,
	q_b_14,
	q_b_15,
	q_b_16,
	q_b_17,
	q_b_18,
	q_b_19,
	q_b_20,
	q_b_21,
	q_b_22,
	q_b_23,
	q_b_24,
	q_b_25,
	q_b_26,
	q_b_27,
	source_valid_s,
	clk,
	in_valid,
	reset_n,
	out_ready,
	in_data_19,
	in_data_18,
	in_data_17,
	in_data_16,
	in_data_15,
	in_data_14,
	in_data_13,
	in_data_12,
	in_data_11,
	in_data_10,
	in_data_9,
	in_data_8,
	in_data_7,
	in_data_6,
	in_data_5,
	in_data_4,
	in_data_3,
	in_data_2,
	in_data_1,
	in_data_0)/* synthesis synthesis_greybox=1 */;
output 	full_dff;
output 	q_b_0;
output 	q_b_1;
output 	q_b_2;
output 	q_b_3;
output 	q_b_4;
output 	q_b_5;
output 	q_b_6;
output 	q_b_7;
output 	q_b_8;
output 	q_b_9;
output 	q_b_10;
output 	q_b_11;
output 	q_b_12;
output 	q_b_13;
output 	q_b_14;
output 	q_b_15;
output 	q_b_16;
output 	q_b_17;
output 	q_b_18;
output 	q_b_19;
output 	q_b_20;
output 	q_b_21;
output 	q_b_22;
output 	q_b_23;
output 	q_b_24;
output 	q_b_25;
output 	q_b_26;
output 	q_b_27;
output 	source_valid_s;
input 	clk;
input 	in_valid;
input 	reset_n;
input 	out_ready;
input 	in_data_19;
input 	in_data_18;
input 	in_data_17;
input 	in_data_16;
input 	in_data_15;
input 	in_data_14;
input 	in_data_13;
input 	in_data_12;
input 	in_data_11;
input 	in_data_10;
input 	in_data_9;
input 	in_data_8;
input 	in_data_7;
input 	in_data_6;
input 	in_data_5;
input 	in_data_4;
input 	in_data_3;
input 	in_data_2;
input 	in_data_1;
input 	in_data_0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cic_alt_cic_core core(
	.full_dff(full_dff),
	.q_b_0(q_b_0),
	.q_b_1(q_b_1),
	.q_b_2(q_b_2),
	.q_b_3(q_b_3),
	.q_b_4(q_b_4),
	.q_b_5(q_b_5),
	.q_b_6(q_b_6),
	.q_b_7(q_b_7),
	.q_b_8(q_b_8),
	.q_b_9(q_b_9),
	.q_b_10(q_b_10),
	.q_b_11(q_b_11),
	.q_b_12(q_b_12),
	.q_b_13(q_b_13),
	.q_b_14(q_b_14),
	.q_b_15(q_b_15),
	.q_b_16(q_b_16),
	.q_b_17(q_b_17),
	.q_b_18(q_b_18),
	.q_b_19(q_b_19),
	.q_b_20(q_b_20),
	.q_b_21(q_b_21),
	.q_b_22(q_b_22),
	.q_b_23(q_b_23),
	.q_b_24(q_b_24),
	.q_b_25(q_b_25),
	.q_b_26(q_b_26),
	.q_b_27(q_b_27),
	.source_valid_s(source_valid_s),
	.clk(clk),
	.in_valid(in_valid),
	.reset_n(reset_n),
	.out_ready(out_ready),
	.in_data_19(in_data_19),
	.in_data_18(in_data_18),
	.in_data_17(in_data_17),
	.in_data_16(in_data_16),
	.in_data_15(in_data_15),
	.in_data_14(in_data_14),
	.in_data_13(in_data_13),
	.in_data_12(in_data_12),
	.in_data_11(in_data_11),
	.in_data_10(in_data_10),
	.in_data_9(in_data_9),
	.in_data_8(in_data_8),
	.in_data_7(in_data_7),
	.in_data_6(in_data_6),
	.in_data_5(in_data_5),
	.in_data_4(in_data_4),
	.in_data_3(in_data_3),
	.in_data_2(in_data_2),
	.in_data_1(in_data_1),
	.in_data_0(in_data_0));

endmodule

module cic_alt_cic_core (
	full_dff,
	q_b_0,
	q_b_1,
	q_b_2,
	q_b_3,
	q_b_4,
	q_b_5,
	q_b_6,
	q_b_7,
	q_b_8,
	q_b_9,
	q_b_10,
	q_b_11,
	q_b_12,
	q_b_13,
	q_b_14,
	q_b_15,
	q_b_16,
	q_b_17,
	q_b_18,
	q_b_19,
	q_b_20,
	q_b_21,
	q_b_22,
	q_b_23,
	q_b_24,
	q_b_25,
	q_b_26,
	q_b_27,
	source_valid_s,
	clk,
	in_valid,
	reset_n,
	out_ready,
	in_data_19,
	in_data_18,
	in_data_17,
	in_data_16,
	in_data_15,
	in_data_14,
	in_data_13,
	in_data_12,
	in_data_11,
	in_data_10,
	in_data_9,
	in_data_8,
	in_data_7,
	in_data_6,
	in_data_5,
	in_data_4,
	in_data_3,
	in_data_2,
	in_data_1,
	in_data_0)/* synthesis synthesis_greybox=1 */;
output 	full_dff;
output 	q_b_0;
output 	q_b_1;
output 	q_b_2;
output 	q_b_3;
output 	q_b_4;
output 	q_b_5;
output 	q_b_6;
output 	q_b_7;
output 	q_b_8;
output 	q_b_9;
output 	q_b_10;
output 	q_b_11;
output 	q_b_12;
output 	q_b_13;
output 	q_b_14;
output 	q_b_15;
output 	q_b_16;
output 	q_b_17;
output 	q_b_18;
output 	q_b_19;
output 	q_b_20;
output 	q_b_21;
output 	q_b_22;
output 	q_b_23;
output 	q_b_24;
output 	q_b_25;
output 	q_b_26;
output 	q_b_27;
output 	source_valid_s;
input 	clk;
input 	in_valid;
input 	reset_n;
input 	out_ready;
input 	in_data_19;
input 	in_data_18;
input 	in_data_17;
input 	in_data_16;
input 	in_data_15;
input 	in_data_14;
input 	in_data_13;
input 	in_data_12;
input 	in_data_11;
input 	in_data_10;
input 	in_data_9;
input 	in_data_8;
input 	in_data_7;
input 	in_data_6;
input 	in_data_5;
input 	in_data_4;
input 	in_data_3;
input 	in_data_2;
input 	in_data_1;
input 	in_data_0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \avalon_controller|ready_FIFO|rd_addr_ptr[2]~q ;
wire \input_sink|sink_FIFO|auto_generated|dffe_nae~q ;
wire \output_source_0|source_FIFO|auto_generated|dffe_af~q ;
wire \dec_one|differentiate_stages[7].auk_dsp_diff|dout_valid~q ;
wire \dec_one|state[0]~q ;
wire \dec_one|differentiate_stages[7].auk_dsp_diff|dout[3]~q ;
wire \dec_one|differentiate_stages[7].auk_dsp_diff|dout[4]~q ;
wire \dec_one|differentiate_stages[7].auk_dsp_diff|dout[5]~q ;
wire \dec_one|differentiate_stages[7].auk_dsp_diff|dout[6]~q ;
wire \dec_one|differentiate_stages[7].auk_dsp_diff|dout[7]~q ;
wire \dec_one|differentiate_stages[7].auk_dsp_diff|dout[8]~q ;
wire \dec_one|differentiate_stages[7].auk_dsp_diff|dout[9]~q ;
wire \dec_one|differentiate_stages[7].auk_dsp_diff|dout[10]~q ;
wire \dec_one|differentiate_stages[7].auk_dsp_diff|dout[11]~q ;
wire \dec_one|differentiate_stages[7].auk_dsp_diff|dout[12]~q ;
wire \dec_one|differentiate_stages[7].auk_dsp_diff|dout[13]~q ;
wire \dec_one|differentiate_stages[7].auk_dsp_diff|dout[14]~q ;
wire \dec_one|differentiate_stages[7].auk_dsp_diff|dout[15]~q ;
wire \dec_one|differentiate_stages[7].auk_dsp_diff|dout[16]~q ;
wire \dec_one|differentiate_stages[7].auk_dsp_diff|dout[17]~q ;
wire \dec_one|differentiate_stages[7].auk_dsp_diff|dout[18]~q ;
wire \dec_one|differentiate_stages[7].auk_dsp_diff|dout[19]~q ;
wire \dec_one|differentiate_stages[7].auk_dsp_diff|dout[20]~q ;
wire \dec_one|differentiate_stages[7].auk_dsp_diff|dout[21]~q ;
wire \dec_one|differentiate_stages[7].auk_dsp_diff|dout[22]~q ;
wire \dec_one|differentiate_stages[7].auk_dsp_diff|dout[23]~q ;
wire \dec_one|differentiate_stages[7].auk_dsp_diff|dout[24]~q ;
wire \dec_one|differentiate_stages[7].auk_dsp_diff|dout[25]~q ;
wire \dec_one|differentiate_stages[7].auk_dsp_diff|dout[26]~q ;
wire \dec_one|differentiate_stages[7].auk_dsp_diff|dout[27]~q ;
wire \dec_one|differentiate_stages[7].auk_dsp_diff|dout[28]~q ;
wire \dec_one|differentiate_stages[7].auk_dsp_diff|dout[29]~q ;
wire \dec_one|differentiate_stages[7].auk_dsp_diff|dout[30]~q ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[19] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[18] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[17] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[16] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[15] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[14] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[13] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[12] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[11] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[10] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[9] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[8] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[7] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[6] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[5] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[4] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[3] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[2] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[1] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[0] ;
wire \avalon_controller|ready_FIFO|Equal2~0_combout ;
wire \avalon_controller|ready_FIFO|Mux0~0_combout ;
wire \avalon_controller|sink_ready_ctrl~0_combout ;
wire \avalon_controller|ready_FIFO|usedw_process~0_combout ;
wire \avalon_controller|stall_reg~q ;
wire \avalon_controller|sink_ready_ctrl~1_combout ;
wire \avalon_controller|sink_ready_ctrl~2_combout ;


cic_auk_dspip_avalon_streaming_source output_source_0(
	.at_source_data({q_b_27,q_b_26,q_b_25,q_b_24,q_b_23,q_b_22,q_b_21,q_b_20,q_b_19,q_b_18,q_b_17,q_b_16,q_b_15,q_b_14,q_b_13,q_b_12,q_b_11,q_b_10,q_b_9,q_b_8,q_b_7,q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.source_valid_s1(source_valid_s),
	.dffe_af(\output_source_0|source_FIFO|auto_generated|dffe_af~q ),
	.dout_valid(\dec_one|differentiate_stages[7].auk_dsp_diff|dout_valid~q ),
	.state_0(\dec_one|state[0]~q ),
	.data({\dec_one|differentiate_stages[7].auk_dsp_diff|dout[30]~q ,\dec_one|differentiate_stages[7].auk_dsp_diff|dout[29]~q ,\dec_one|differentiate_stages[7].auk_dsp_diff|dout[28]~q ,\dec_one|differentiate_stages[7].auk_dsp_diff|dout[27]~q ,
\dec_one|differentiate_stages[7].auk_dsp_diff|dout[26]~q ,\dec_one|differentiate_stages[7].auk_dsp_diff|dout[25]~q ,\dec_one|differentiate_stages[7].auk_dsp_diff|dout[24]~q ,\dec_one|differentiate_stages[7].auk_dsp_diff|dout[23]~q ,
\dec_one|differentiate_stages[7].auk_dsp_diff|dout[22]~q ,\dec_one|differentiate_stages[7].auk_dsp_diff|dout[21]~q ,\dec_one|differentiate_stages[7].auk_dsp_diff|dout[20]~q ,\dec_one|differentiate_stages[7].auk_dsp_diff|dout[19]~q ,
\dec_one|differentiate_stages[7].auk_dsp_diff|dout[18]~q ,\dec_one|differentiate_stages[7].auk_dsp_diff|dout[17]~q ,\dec_one|differentiate_stages[7].auk_dsp_diff|dout[16]~q ,\dec_one|differentiate_stages[7].auk_dsp_diff|dout[15]~q ,
\dec_one|differentiate_stages[7].auk_dsp_diff|dout[14]~q ,\dec_one|differentiate_stages[7].auk_dsp_diff|dout[13]~q ,\dec_one|differentiate_stages[7].auk_dsp_diff|dout[12]~q ,\dec_one|differentiate_stages[7].auk_dsp_diff|dout[11]~q ,
\dec_one|differentiate_stages[7].auk_dsp_diff|dout[10]~q ,\dec_one|differentiate_stages[7].auk_dsp_diff|dout[9]~q ,\dec_one|differentiate_stages[7].auk_dsp_diff|dout[8]~q ,\dec_one|differentiate_stages[7].auk_dsp_diff|dout[7]~q ,
\dec_one|differentiate_stages[7].auk_dsp_diff|dout[6]~q ,\dec_one|differentiate_stages[7].auk_dsp_diff|dout[5]~q ,\dec_one|differentiate_stages[7].auk_dsp_diff|dout[4]~q ,\dec_one|differentiate_stages[7].auk_dsp_diff|dout[3]~q }),
	.stall_reg(\avalon_controller|stall_reg~q ),
	.clk(clk),
	.reset_n(reset_n),
	.out_ready(out_ready));

cic_auk_dspip_avalon_streaming_sink input_sink(
	.full_dff(full_dff),
	.rd_addr_ptr_2(\avalon_controller|ready_FIFO|rd_addr_ptr[2]~q ),
	.dffe_nae(\input_sink|sink_FIFO|auto_generated|dffe_nae~q ),
	.data({\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[19] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[18] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[17] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[16] ,
\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[15] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[14] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[13] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[12] ,
\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[11] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[10] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[9] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[8] ,
\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[7] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[6] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[5] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[4] ,
\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[3] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[2] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[1] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[0] }),
	.Equal2(\avalon_controller|ready_FIFO|Equal2~0_combout ),
	.Mux0(\avalon_controller|ready_FIFO|Mux0~0_combout ),
	.sink_ready_ctrl(\avalon_controller|sink_ready_ctrl~0_combout ),
	.usedw_process(\avalon_controller|ready_FIFO|usedw_process~0_combout ),
	.sink_ready_ctrl1(\avalon_controller|sink_ready_ctrl~1_combout ),
	.sink_ready_ctrl2(\avalon_controller|sink_ready_ctrl~2_combout ),
	.clk(clk),
	.in_valid(in_valid),
	.reset_n(reset_n),
	.at_sink_data({in_data_19,in_data_18,in_data_17,in_data_16,in_data_15,in_data_14,in_data_13,in_data_12,in_data_11,in_data_10,in_data_9,in_data_8,in_data_7,in_data_6,in_data_5,in_data_4,in_data_3,in_data_2,in_data_1,in_data_0}));

cic_alt_cic_dec_siso dec_one(
	.dout_valid(\dec_one|differentiate_stages[7].auk_dsp_diff|dout_valid~q ),
	.state_0(\dec_one|state[0]~q ),
	.dout_3(\dec_one|differentiate_stages[7].auk_dsp_diff|dout[3]~q ),
	.dout_4(\dec_one|differentiate_stages[7].auk_dsp_diff|dout[4]~q ),
	.dout_5(\dec_one|differentiate_stages[7].auk_dsp_diff|dout[5]~q ),
	.dout_6(\dec_one|differentiate_stages[7].auk_dsp_diff|dout[6]~q ),
	.dout_7(\dec_one|differentiate_stages[7].auk_dsp_diff|dout[7]~q ),
	.dout_8(\dec_one|differentiate_stages[7].auk_dsp_diff|dout[8]~q ),
	.dout_9(\dec_one|differentiate_stages[7].auk_dsp_diff|dout[9]~q ),
	.dout_10(\dec_one|differentiate_stages[7].auk_dsp_diff|dout[10]~q ),
	.dout_11(\dec_one|differentiate_stages[7].auk_dsp_diff|dout[11]~q ),
	.dout_12(\dec_one|differentiate_stages[7].auk_dsp_diff|dout[12]~q ),
	.dout_13(\dec_one|differentiate_stages[7].auk_dsp_diff|dout[13]~q ),
	.dout_14(\dec_one|differentiate_stages[7].auk_dsp_diff|dout[14]~q ),
	.dout_15(\dec_one|differentiate_stages[7].auk_dsp_diff|dout[15]~q ),
	.dout_16(\dec_one|differentiate_stages[7].auk_dsp_diff|dout[16]~q ),
	.dout_17(\dec_one|differentiate_stages[7].auk_dsp_diff|dout[17]~q ),
	.dout_18(\dec_one|differentiate_stages[7].auk_dsp_diff|dout[18]~q ),
	.dout_19(\dec_one|differentiate_stages[7].auk_dsp_diff|dout[19]~q ),
	.dout_20(\dec_one|differentiate_stages[7].auk_dsp_diff|dout[20]~q ),
	.dout_21(\dec_one|differentiate_stages[7].auk_dsp_diff|dout[21]~q ),
	.dout_22(\dec_one|differentiate_stages[7].auk_dsp_diff|dout[22]~q ),
	.dout_23(\dec_one|differentiate_stages[7].auk_dsp_diff|dout[23]~q ),
	.dout_24(\dec_one|differentiate_stages[7].auk_dsp_diff|dout[24]~q ),
	.dout_25(\dec_one|differentiate_stages[7].auk_dsp_diff|dout[25]~q ),
	.dout_26(\dec_one|differentiate_stages[7].auk_dsp_diff|dout[26]~q ),
	.dout_27(\dec_one|differentiate_stages[7].auk_dsp_diff|dout[27]~q ),
	.dout_28(\dec_one|differentiate_stages[7].auk_dsp_diff|dout[28]~q ),
	.dout_29(\dec_one|differentiate_stages[7].auk_dsp_diff|dout[29]~q ),
	.dout_30(\dec_one|differentiate_stages[7].auk_dsp_diff|dout[30]~q ),
	.q_b_19(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[19] ),
	.q_b_18(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[18] ),
	.q_b_17(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[17] ),
	.q_b_16(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[16] ),
	.q_b_15(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[15] ),
	.q_b_14(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[14] ),
	.q_b_13(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[13] ),
	.q_b_12(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[12] ),
	.q_b_11(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[11] ),
	.q_b_10(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[10] ),
	.q_b_9(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[9] ),
	.q_b_8(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[8] ),
	.q_b_7(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[7] ),
	.q_b_6(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[6] ),
	.q_b_5(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[5] ),
	.q_b_4(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[4] ),
	.q_b_3(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[3] ),
	.q_b_2(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[2] ),
	.q_b_1(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[1] ),
	.q_b_0(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[0] ),
	.stall_reg(\avalon_controller|stall_reg~q ),
	.clk(clk),
	.reset_n(reset_n));

cic_auk_dspip_avalon_streaming_controller avalon_controller(
	.rd_addr_ptr_2(\avalon_controller|ready_FIFO|rd_addr_ptr[2]~q ),
	.dffe_nae(\input_sink|sink_FIFO|auto_generated|dffe_nae~q ),
	.dffe_af(\output_source_0|source_FIFO|auto_generated|dffe_af~q ),
	.Equal2(\avalon_controller|ready_FIFO|Equal2~0_combout ),
	.Mux0(\avalon_controller|ready_FIFO|Mux0~0_combout ),
	.sink_ready_ctrl(\avalon_controller|sink_ready_ctrl~0_combout ),
	.usedw_process(\avalon_controller|ready_FIFO|usedw_process~0_combout ),
	.stall_reg1(\avalon_controller|stall_reg~q ),
	.sink_ready_ctrl1(\avalon_controller|sink_ready_ctrl~1_combout ),
	.sink_ready_ctrl2(\avalon_controller|sink_ready_ctrl~2_combout ),
	.clk(clk),
	.reset_n(reset_n));

endmodule

module cic_alt_cic_dec_siso (
	dout_valid,
	state_0,
	dout_3,
	dout_4,
	dout_5,
	dout_6,
	dout_7,
	dout_8,
	dout_9,
	dout_10,
	dout_11,
	dout_12,
	dout_13,
	dout_14,
	dout_15,
	dout_16,
	dout_17,
	dout_18,
	dout_19,
	dout_20,
	dout_21,
	dout_22,
	dout_23,
	dout_24,
	dout_25,
	dout_26,
	dout_27,
	dout_28,
	dout_29,
	dout_30,
	q_b_19,
	q_b_18,
	q_b_17,
	q_b_16,
	q_b_15,
	q_b_14,
	q_b_13,
	q_b_12,
	q_b_11,
	q_b_10,
	q_b_9,
	q_b_8,
	q_b_7,
	q_b_6,
	q_b_5,
	q_b_4,
	q_b_3,
	q_b_2,
	q_b_1,
	q_b_0,
	stall_reg,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	dout_valid;
output 	state_0;
output 	dout_3;
output 	dout_4;
output 	dout_5;
output 	dout_6;
output 	dout_7;
output 	dout_8;
output 	dout_9;
output 	dout_10;
output 	dout_11;
output 	dout_12;
output 	dout_13;
output 	dout_14;
output 	dout_15;
output 	dout_16;
output 	dout_17;
output 	dout_18;
output 	dout_19;
output 	dout_20;
output 	dout_21;
output 	dout_22;
output 	dout_23;
output 	dout_24;
output 	dout_25;
output 	dout_26;
output 	dout_27;
output 	dout_28;
output 	dout_29;
output 	dout_30;
input 	q_b_19;
input 	q_b_18;
input 	q_b_17;
input 	q_b_16;
input 	q_b_15;
input 	q_b_14;
input 	q_b_13;
input 	q_b_12;
input 	q_b_11;
input 	q_b_10;
input 	q_b_9;
input 	q_b_8;
input 	q_b_7;
input 	q_b_6;
input 	q_b_5;
input 	q_b_4;
input 	q_b_3;
input 	q_b_2;
input 	q_b_1;
input 	q_b_0;
input 	stall_reg;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \differentiate_stages[6].auk_dsp_diff|dout_valid~q ;
wire \differentiate_stages[5].auk_dsp_diff|dout_valid~q ;
wire \differentiate_stages[6].auk_dsp_diff|dout[4]~q ;
wire \differentiate_stages[6].auk_dsp_diff|dout[5]~q ;
wire \differentiate_stages[6].auk_dsp_diff|dout[6]~q ;
wire \differentiate_stages[6].auk_dsp_diff|dout[7]~q ;
wire \differentiate_stages[6].auk_dsp_diff|dout[8]~q ;
wire \differentiate_stages[6].auk_dsp_diff|dout[9]~q ;
wire \differentiate_stages[6].auk_dsp_diff|dout[10]~q ;
wire \differentiate_stages[6].auk_dsp_diff|dout[11]~q ;
wire \differentiate_stages[6].auk_dsp_diff|dout[12]~q ;
wire \differentiate_stages[6].auk_dsp_diff|dout[13]~q ;
wire \differentiate_stages[6].auk_dsp_diff|dout[14]~q ;
wire \differentiate_stages[6].auk_dsp_diff|dout[15]~q ;
wire \differentiate_stages[6].auk_dsp_diff|dout[16]~q ;
wire \differentiate_stages[6].auk_dsp_diff|dout[17]~q ;
wire \differentiate_stages[6].auk_dsp_diff|dout[18]~q ;
wire \differentiate_stages[6].auk_dsp_diff|dout[19]~q ;
wire \differentiate_stages[6].auk_dsp_diff|dout[20]~q ;
wire \differentiate_stages[6].auk_dsp_diff|dout[21]~q ;
wire \differentiate_stages[6].auk_dsp_diff|dout[22]~q ;
wire \differentiate_stages[6].auk_dsp_diff|dout[23]~q ;
wire \differentiate_stages[6].auk_dsp_diff|dout[24]~q ;
wire \differentiate_stages[6].auk_dsp_diff|dout[25]~q ;
wire \differentiate_stages[6].auk_dsp_diff|dout[26]~q ;
wire \differentiate_stages[6].auk_dsp_diff|dout[27]~q ;
wire \differentiate_stages[6].auk_dsp_diff|dout[28]~q ;
wire \differentiate_stages[6].auk_dsp_diff|dout[29]~q ;
wire \differentiate_stages[6].auk_dsp_diff|dout[30]~q ;
wire \differentiate_stages[6].auk_dsp_diff|dout[31]~q ;
wire \differentiate_stages[4].auk_dsp_diff|dout_valid~q ;
wire \differentiate_stages[6].auk_dsp_diff|dout[3]~q ;
wire \differentiate_stages[3].auk_dsp_diff|dout_valid~q ;
wire \differentiate_stages[5].auk_dsp_diff|dout[5]~q ;
wire \differentiate_stages[6].auk_dsp_diff|dout[2]~q ;
wire \differentiate_stages[5].auk_dsp_diff|dout[6]~q ;
wire \differentiate_stages[5].auk_dsp_diff|dout[7]~q ;
wire \differentiate_stages[5].auk_dsp_diff|dout[8]~q ;
wire \differentiate_stages[5].auk_dsp_diff|dout[9]~q ;
wire \differentiate_stages[5].auk_dsp_diff|dout[10]~q ;
wire \differentiate_stages[5].auk_dsp_diff|dout[11]~q ;
wire \differentiate_stages[5].auk_dsp_diff|dout[12]~q ;
wire \differentiate_stages[5].auk_dsp_diff|dout[13]~q ;
wire \differentiate_stages[5].auk_dsp_diff|dout[14]~q ;
wire \differentiate_stages[5].auk_dsp_diff|dout[15]~q ;
wire \differentiate_stages[5].auk_dsp_diff|dout[16]~q ;
wire \differentiate_stages[5].auk_dsp_diff|dout[17]~q ;
wire \differentiate_stages[5].auk_dsp_diff|dout[18]~q ;
wire \differentiate_stages[5].auk_dsp_diff|dout[19]~q ;
wire \differentiate_stages[5].auk_dsp_diff|dout[20]~q ;
wire \differentiate_stages[5].auk_dsp_diff|dout[21]~q ;
wire \differentiate_stages[5].auk_dsp_diff|dout[22]~q ;
wire \differentiate_stages[5].auk_dsp_diff|dout[23]~q ;
wire \differentiate_stages[5].auk_dsp_diff|dout[24]~q ;
wire \differentiate_stages[5].auk_dsp_diff|dout[25]~q ;
wire \differentiate_stages[5].auk_dsp_diff|dout[26]~q ;
wire \differentiate_stages[5].auk_dsp_diff|dout[27]~q ;
wire \differentiate_stages[5].auk_dsp_diff|dout[28]~q ;
wire \differentiate_stages[5].auk_dsp_diff|dout[29]~q ;
wire \differentiate_stages[5].auk_dsp_diff|dout[30]~q ;
wire \differentiate_stages[5].auk_dsp_diff|dout[31]~q ;
wire \differentiate_stages[5].auk_dsp_diff|dout[32]~q ;
wire \differentiate_stages[2].auk_dsp_diff|dout_valid~q ;
wire \differentiate_stages[5].auk_dsp_diff|dout[4]~q ;
wire \differentiate_stages[6].auk_dsp_diff|dout[1]~q ;
wire \differentiate_stages[1].auk_dsp_diff|dout_valid~q ;
wire \differentiate_stages[4].auk_dsp_diff|dout[6]~q ;
wire \differentiate_stages[5].auk_dsp_diff|dout[3]~q ;
wire \differentiate_stages[4].auk_dsp_diff|dout[7]~q ;
wire \differentiate_stages[4].auk_dsp_diff|dout[8]~q ;
wire \differentiate_stages[4].auk_dsp_diff|dout[9]~q ;
wire \differentiate_stages[4].auk_dsp_diff|dout[10]~q ;
wire \differentiate_stages[4].auk_dsp_diff|dout[11]~q ;
wire \differentiate_stages[4].auk_dsp_diff|dout[12]~q ;
wire \differentiate_stages[4].auk_dsp_diff|dout[13]~q ;
wire \differentiate_stages[4].auk_dsp_diff|dout[14]~q ;
wire \differentiate_stages[4].auk_dsp_diff|dout[15]~q ;
wire \differentiate_stages[4].auk_dsp_diff|dout[16]~q ;
wire \differentiate_stages[4].auk_dsp_diff|dout[17]~q ;
wire \differentiate_stages[4].auk_dsp_diff|dout[18]~q ;
wire \differentiate_stages[4].auk_dsp_diff|dout[19]~q ;
wire \differentiate_stages[4].auk_dsp_diff|dout[20]~q ;
wire \differentiate_stages[4].auk_dsp_diff|dout[21]~q ;
wire \differentiate_stages[4].auk_dsp_diff|dout[22]~q ;
wire \differentiate_stages[4].auk_dsp_diff|dout[23]~q ;
wire \differentiate_stages[4].auk_dsp_diff|dout[24]~q ;
wire \differentiate_stages[4].auk_dsp_diff|dout[25]~q ;
wire \differentiate_stages[4].auk_dsp_diff|dout[26]~q ;
wire \differentiate_stages[4].auk_dsp_diff|dout[27]~q ;
wire \differentiate_stages[4].auk_dsp_diff|dout[28]~q ;
wire \differentiate_stages[4].auk_dsp_diff|dout[29]~q ;
wire \differentiate_stages[4].auk_dsp_diff|dout[30]~q ;
wire \differentiate_stages[4].auk_dsp_diff|dout[31]~q ;
wire \differentiate_stages[4].auk_dsp_diff|dout[32]~q ;
wire \differentiate_stages[4].auk_dsp_diff|dout[33]~q ;
wire \differentiate_stages[0].auk_dsp_diff|dout_valid~q ;
wire \differentiate_stages[4].auk_dsp_diff|dout[5]~q ;
wire \differentiate_stages[5].auk_dsp_diff|dout[2]~q ;
wire \differentiate_stages[3].auk_dsp_diff|dout[6]~q ;
wire \differentiate_stages[4].auk_dsp_diff|dout[4]~q ;
wire \differentiate_stages[5].auk_dsp_diff|dout[1]~q ;
wire \differentiate_stages[3].auk_dsp_diff|dout[7]~q ;
wire \differentiate_stages[3].auk_dsp_diff|dout[8]~q ;
wire \differentiate_stages[3].auk_dsp_diff|dout[9]~q ;
wire \differentiate_stages[3].auk_dsp_diff|dout[10]~q ;
wire \differentiate_stages[3].auk_dsp_diff|dout[11]~q ;
wire \differentiate_stages[3].auk_dsp_diff|dout[12]~q ;
wire \differentiate_stages[3].auk_dsp_diff|dout[13]~q ;
wire \differentiate_stages[3].auk_dsp_diff|dout[14]~q ;
wire \differentiate_stages[3].auk_dsp_diff|dout[15]~q ;
wire \differentiate_stages[3].auk_dsp_diff|dout[16]~q ;
wire \differentiate_stages[3].auk_dsp_diff|dout[17]~q ;
wire \differentiate_stages[3].auk_dsp_diff|dout[18]~q ;
wire \differentiate_stages[3].auk_dsp_diff|dout[19]~q ;
wire \differentiate_stages[3].auk_dsp_diff|dout[20]~q ;
wire \differentiate_stages[3].auk_dsp_diff|dout[21]~q ;
wire \differentiate_stages[3].auk_dsp_diff|dout[22]~q ;
wire \differentiate_stages[3].auk_dsp_diff|dout[23]~q ;
wire \differentiate_stages[3].auk_dsp_diff|dout[24]~q ;
wire \differentiate_stages[3].auk_dsp_diff|dout[25]~q ;
wire \differentiate_stages[3].auk_dsp_diff|dout[26]~q ;
wire \differentiate_stages[3].auk_dsp_diff|dout[27]~q ;
wire \differentiate_stages[3].auk_dsp_diff|dout[28]~q ;
wire \differentiate_stages[3].auk_dsp_diff|dout[29]~q ;
wire \differentiate_stages[3].auk_dsp_diff|dout[30]~q ;
wire \differentiate_stages[3].auk_dsp_diff|dout[31]~q ;
wire \differentiate_stages[3].auk_dsp_diff|dout[32]~q ;
wire \differentiate_stages[3].auk_dsp_diff|dout[33]~q ;
wire \differentiate_stages[3].auk_dsp_diff|dout[5]~q ;
wire \differentiate_stages[4].auk_dsp_diff|dout[3]~q ;
wire \ena_diff_s[0]~q ;
wire \differentiate_stages[2].auk_dsp_diff|dout[7]~q ;
wire \differentiate_stages[3].auk_dsp_diff|dout[4]~q ;
wire \differentiate_stages[4].auk_dsp_diff|dout[2]~q ;
wire \differentiate_stages[2].auk_dsp_diff|dout[8]~q ;
wire \differentiate_stages[2].auk_dsp_diff|dout[9]~q ;
wire \differentiate_stages[2].auk_dsp_diff|dout[10]~q ;
wire \differentiate_stages[2].auk_dsp_diff|dout[11]~q ;
wire \differentiate_stages[2].auk_dsp_diff|dout[12]~q ;
wire \differentiate_stages[2].auk_dsp_diff|dout[13]~q ;
wire \differentiate_stages[2].auk_dsp_diff|dout[14]~q ;
wire \differentiate_stages[2].auk_dsp_diff|dout[15]~q ;
wire \differentiate_stages[2].auk_dsp_diff|dout[16]~q ;
wire \differentiate_stages[2].auk_dsp_diff|dout[17]~q ;
wire \differentiate_stages[2].auk_dsp_diff|dout[18]~q ;
wire \differentiate_stages[2].auk_dsp_diff|dout[19]~q ;
wire \differentiate_stages[2].auk_dsp_diff|dout[20]~q ;
wire \differentiate_stages[2].auk_dsp_diff|dout[21]~q ;
wire \differentiate_stages[2].auk_dsp_diff|dout[22]~q ;
wire \differentiate_stages[2].auk_dsp_diff|dout[23]~q ;
wire \differentiate_stages[2].auk_dsp_diff|dout[24]~q ;
wire \differentiate_stages[2].auk_dsp_diff|dout[25]~q ;
wire \differentiate_stages[2].auk_dsp_diff|dout[26]~q ;
wire \differentiate_stages[2].auk_dsp_diff|dout[27]~q ;
wire \differentiate_stages[2].auk_dsp_diff|dout[28]~q ;
wire \differentiate_stages[2].auk_dsp_diff|dout[29]~q ;
wire \differentiate_stages[2].auk_dsp_diff|dout[30]~q ;
wire \differentiate_stages[2].auk_dsp_diff|dout[31]~q ;
wire \differentiate_stages[2].auk_dsp_diff|dout[32]~q ;
wire \differentiate_stages[2].auk_dsp_diff|dout[33]~q ;
wire \differentiate_stages[2].auk_dsp_diff|dout[34]~q ;
wire \sample_state[0]~q ;
wire \differentiate_stages[2].auk_dsp_diff|dout[6]~q ;
wire \differentiate_stages[3].auk_dsp_diff|dout[3]~q ;
wire \differentiate_stages[4].auk_dsp_diff|dout[1]~q ;
wire \differentiate_stages[1].auk_dsp_diff|dout[8]~q ;
wire \differentiate_stages[2].auk_dsp_diff|dout[5]~q ;
wire \differentiate_stages[3].auk_dsp_diff|dout[2]~q ;
wire \differentiate_stages[1].auk_dsp_diff|dout[9]~q ;
wire \differentiate_stages[1].auk_dsp_diff|dout[10]~q ;
wire \differentiate_stages[1].auk_dsp_diff|dout[11]~q ;
wire \differentiate_stages[1].auk_dsp_diff|dout[12]~q ;
wire \differentiate_stages[1].auk_dsp_diff|dout[13]~q ;
wire \differentiate_stages[1].auk_dsp_diff|dout[14]~q ;
wire \differentiate_stages[1].auk_dsp_diff|dout[15]~q ;
wire \differentiate_stages[1].auk_dsp_diff|dout[16]~q ;
wire \differentiate_stages[1].auk_dsp_diff|dout[17]~q ;
wire \differentiate_stages[1].auk_dsp_diff|dout[18]~q ;
wire \differentiate_stages[1].auk_dsp_diff|dout[19]~q ;
wire \differentiate_stages[1].auk_dsp_diff|dout[20]~q ;
wire \differentiate_stages[1].auk_dsp_diff|dout[21]~q ;
wire \differentiate_stages[1].auk_dsp_diff|dout[22]~q ;
wire \differentiate_stages[1].auk_dsp_diff|dout[23]~q ;
wire \differentiate_stages[1].auk_dsp_diff|dout[24]~q ;
wire \differentiate_stages[1].auk_dsp_diff|dout[25]~q ;
wire \differentiate_stages[1].auk_dsp_diff|dout[26]~q ;
wire \differentiate_stages[1].auk_dsp_diff|dout[27]~q ;
wire \differentiate_stages[1].auk_dsp_diff|dout[28]~q ;
wire \differentiate_stages[1].auk_dsp_diff|dout[29]~q ;
wire \differentiate_stages[1].auk_dsp_diff|dout[30]~q ;
wire \differentiate_stages[1].auk_dsp_diff|dout[31]~q ;
wire \differentiate_stages[1].auk_dsp_diff|dout[32]~q ;
wire \differentiate_stages[1].auk_dsp_diff|dout[33]~q ;
wire \differentiate_stages[1].auk_dsp_diff|dout[34]~q ;
wire \differentiate_stages[1].auk_dsp_diff|dout[35]~q ;
wire \differentiate_stages[1].auk_dsp_diff|dout[7]~q ;
wire \differentiate_stages[2].auk_dsp_diff|dout[4]~q ;
wire \differentiate_stages[3].auk_dsp_diff|dout[1]~q ;
wire \differentiate_stages[0].auk_dsp_diff|dout[9]~q ;
wire \differentiate_stages[1].auk_dsp_diff|dout[6]~q ;
wire \differentiate_stages[2].auk_dsp_diff|dout[3]~q ;
wire \differentiate_stages[3].auk_dsp_diff|dout[0]~q ;
wire \differentiate_stages[0].auk_dsp_diff|dout[10]~q ;
wire \differentiate_stages[0].auk_dsp_diff|dout[11]~q ;
wire \differentiate_stages[0].auk_dsp_diff|dout[12]~q ;
wire \differentiate_stages[0].auk_dsp_diff|dout[13]~q ;
wire \differentiate_stages[0].auk_dsp_diff|dout[14]~q ;
wire \differentiate_stages[0].auk_dsp_diff|dout[15]~q ;
wire \differentiate_stages[0].auk_dsp_diff|dout[16]~q ;
wire \differentiate_stages[0].auk_dsp_diff|dout[17]~q ;
wire \differentiate_stages[0].auk_dsp_diff|dout[18]~q ;
wire \differentiate_stages[0].auk_dsp_diff|dout[19]~q ;
wire \differentiate_stages[0].auk_dsp_diff|dout[20]~q ;
wire \differentiate_stages[0].auk_dsp_diff|dout[21]~q ;
wire \differentiate_stages[0].auk_dsp_diff|dout[22]~q ;
wire \differentiate_stages[0].auk_dsp_diff|dout[23]~q ;
wire \differentiate_stages[0].auk_dsp_diff|dout[24]~q ;
wire \differentiate_stages[0].auk_dsp_diff|dout[25]~q ;
wire \differentiate_stages[0].auk_dsp_diff|dout[26]~q ;
wire \differentiate_stages[0].auk_dsp_diff|dout[27]~q ;
wire \differentiate_stages[0].auk_dsp_diff|dout[28]~q ;
wire \differentiate_stages[0].auk_dsp_diff|dout[29]~q ;
wire \differentiate_stages[0].auk_dsp_diff|dout[30]~q ;
wire \differentiate_stages[0].auk_dsp_diff|dout[31]~q ;
wire \differentiate_stages[0].auk_dsp_diff|dout[32]~q ;
wire \differentiate_stages[0].auk_dsp_diff|dout[33]~q ;
wire \differentiate_stages[0].auk_dsp_diff|dout[34]~q ;
wire \differentiate_stages[0].auk_dsp_diff|dout[35]~q ;
wire \differentiate_stages[0].auk_dsp_diff|dout[36]~q ;
wire \differentiate_stages[0].auk_dsp_diff|dout[8]~q ;
wire \differentiate_stages[1].auk_dsp_diff|dout[5]~q ;
wire \differentiate_stages[2].auk_dsp_diff|dout[2]~q ;
wire \fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[10] ;
wire \differentiate_stages[0].auk_dsp_diff|dout[7]~q ;
wire \differentiate_stages[1].auk_dsp_diff|dout[4]~q ;
wire \differentiate_stages[2].auk_dsp_diff|dout[1]~q ;
wire \fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[11] ;
wire \fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[12] ;
wire \fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[13] ;
wire \fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[14] ;
wire \fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[15] ;
wire \fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[16] ;
wire \fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[17] ;
wire \fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[18] ;
wire \fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[19] ;
wire \fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[20] ;
wire \fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[21] ;
wire \fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[22] ;
wire \fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[23] ;
wire \fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[24] ;
wire \fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[25] ;
wire \fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[26] ;
wire \fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[27] ;
wire \fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[28] ;
wire \fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[29] ;
wire \fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[30] ;
wire \fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[31] ;
wire \fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[32] ;
wire \fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[33] ;
wire \fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[34] ;
wire \fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[35] ;
wire \fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[36] ;
wire \fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[37] ;
wire \fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[9] ;
wire \differentiate_stages[0].auk_dsp_diff|dout[6]~q ;
wire \differentiate_stages[1].auk_dsp_diff|dout[3]~q ;
wire \fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[8] ;
wire \differentiate_stages[0].auk_dsp_diff|dout[5]~q ;
wire \differentiate_stages[1].auk_dsp_diff|dout[2]~q ;
wire \fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[7] ;
wire \differentiate_stages[0].auk_dsp_diff|dout[4]~q ;
wire \differentiate_stages[1].auk_dsp_diff|dout[1]~q ;
wire \fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[6] ;
wire \differentiate_stages[0].auk_dsp_diff|dout[3]~q ;
wire \fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[5] ;
wire \differentiate_stages[0].auk_dsp_diff|dout[2]~q ;
wire \fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[4] ;
wire \differentiate_stages[0].auk_dsp_diff|dout[1]~q ;
wire \fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[3] ;
wire \fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[2] ;
wire \fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[1] ;
wire \differentiate_stages[7].auk_dsp_diff|dout_valid~0_combout ;
wire \latency_cnt_inst|count[0]~q ;
wire \latency_cnt_inst|count[1]~q ;
wire \latency_cnt_inst|count[2]~q ;
wire \latency_cnt_inst|count[3]~q ;
wire \latency_cnt_inst|count[4]~q ;
wire \latency_cnt_inst|Equal0~0_combout ;
wire \sample_state~0_combout ;
wire \ena_diff_s[1]~q ;
wire \fifo_rdreq~q ;
wire \fifo_regulator|buffer_FIFO|auto_generated|dpfifo|valid_rreq~0_combout ;
wire \fifo_rdreq~0_combout ;
wire \vrc_en_0.first_dsample|counter_fs_inst|count[0]~q ;
wire \vrc_en_0.first_dsample|counter_fs_inst|count[3]~q ;
wire \vrc_en_0.first_dsample|counter_fs_inst|count[1]~q ;
wire \vrc_en_0.first_dsample|counter_fs_inst|count[2]~q ;
wire \fifo_regulator|buffer_FIFO|auto_generated|dpfifo|valid_wreq~0_combout ;
wire \ena_diff_s~0_combout ;
wire \sample_state~1_combout ;
wire \integrator[7].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ;
wire \integrator[7].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ;
wire \integrator[7].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ;
wire \integrator[7].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ;
wire \integrator[7].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ;
wire \integrator[7].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ;
wire \integrator[7].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ;
wire \integrator[7].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ;
wire \integrator[7].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ;
wire \integrator[7].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][19]~q ;
wire \integrator[7].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][20]~q ;
wire \integrator[7].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][21]~q ;
wire \integrator[7].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][22]~q ;
wire \integrator[7].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][23]~q ;
wire \integrator[7].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][24]~q ;
wire \integrator[7].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][25]~q ;
wire \integrator[7].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][26]~q ;
wire \integrator[7].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][27]~q ;
wire \integrator[7].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][28]~q ;
wire \integrator[7].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][29]~q ;
wire \integrator[7].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][30]~q ;
wire \integrator[7].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][31]~q ;
wire \integrator[7].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][32]~q ;
wire \integrator[7].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][33]~q ;
wire \integrator[7].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][34]~q ;
wire \integrator[7].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][35]~q ;
wire \integrator[7].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][36]~q ;
wire \integrator[7].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][37]~q ;
wire \integrator[7].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ;
wire \integrator[6].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ;
wire \integrator[7].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ;
wire \integrator[6].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ;
wire \integrator[6].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ;
wire \integrator[6].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ;
wire \integrator[6].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ;
wire \integrator[6].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ;
wire \integrator[6].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ;
wire \integrator[6].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][19]~q ;
wire \integrator[6].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][20]~q ;
wire \integrator[6].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][21]~q ;
wire \integrator[6].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][22]~q ;
wire \integrator[6].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][23]~q ;
wire \integrator[6].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][24]~q ;
wire \integrator[6].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][25]~q ;
wire \integrator[6].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][26]~q ;
wire \integrator[6].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][27]~q ;
wire \integrator[6].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][28]~q ;
wire \integrator[6].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][29]~q ;
wire \integrator[6].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][30]~q ;
wire \integrator[6].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][31]~q ;
wire \integrator[6].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][32]~q ;
wire \integrator[6].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][33]~q ;
wire \integrator[6].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][34]~q ;
wire \integrator[6].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][35]~q ;
wire \integrator[6].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][36]~q ;
wire \integrator[6].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][37]~q ;
wire \integrator[6].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][38]~q ;
wire \integrator[6].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][39]~q ;
wire \integrator[6].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ;
wire \integrator[7].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ;
wire \integrator[5].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ;
wire \integrator[6].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ;
wire \integrator[7].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ;
wire \integrator[5].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ;
wire \integrator[5].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ;
wire \integrator[5].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ;
wire \integrator[5].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ;
wire \integrator[5].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][19]~q ;
wire \integrator[5].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][20]~q ;
wire \integrator[5].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][21]~q ;
wire \integrator[5].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][22]~q ;
wire \integrator[5].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][23]~q ;
wire \integrator[5].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][24]~q ;
wire \integrator[5].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][25]~q ;
wire \integrator[5].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][26]~q ;
wire \integrator[5].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][27]~q ;
wire \integrator[5].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][28]~q ;
wire \integrator[5].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][29]~q ;
wire \integrator[5].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][30]~q ;
wire \integrator[5].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][31]~q ;
wire \integrator[5].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][32]~q ;
wire \integrator[5].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][33]~q ;
wire \integrator[5].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][34]~q ;
wire \integrator[5].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][35]~q ;
wire \integrator[5].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][36]~q ;
wire \integrator[5].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][37]~q ;
wire \integrator[5].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][38]~q ;
wire \integrator[5].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][39]~q ;
wire \integrator[5].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][40]~q ;
wire \integrator[5].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][41]~q ;
wire \integrator[5].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ;
wire \integrator[6].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ;
wire \integrator[7].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ;
wire \integrator[4].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ;
wire \integrator[5].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ;
wire \integrator[6].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ;
wire \integrator[7].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][4]~q ;
wire \integrator[4].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ;
wire \integrator[4].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ;
wire \integrator[4].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][19]~q ;
wire \integrator[4].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][20]~q ;
wire \integrator[4].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][21]~q ;
wire \integrator[4].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][22]~q ;
wire \integrator[4].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][23]~q ;
wire \integrator[4].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][24]~q ;
wire \integrator[4].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][25]~q ;
wire \integrator[4].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][26]~q ;
wire \integrator[4].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][27]~q ;
wire \integrator[4].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][28]~q ;
wire \integrator[4].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][29]~q ;
wire \integrator[4].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][30]~q ;
wire \integrator[4].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][31]~q ;
wire \integrator[4].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][32]~q ;
wire \integrator[4].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][33]~q ;
wire \integrator[4].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][34]~q ;
wire \integrator[4].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][35]~q ;
wire \integrator[4].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][36]~q ;
wire \integrator[4].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][37]~q ;
wire \integrator[4].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][38]~q ;
wire \integrator[4].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][39]~q ;
wire \integrator[4].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][40]~q ;
wire \integrator[4].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][41]~q ;
wire \integrator[4].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][42]~q ;
wire \integrator[4].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][43]~q ;
wire \integrator[4].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ;
wire \integrator[5].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ;
wire \integrator[6].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ;
wire \integrator[7].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][3]~q ;
wire \integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ;
wire \integrator[4].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ;
wire \integrator[5].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ;
wire \integrator[6].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ;
wire \integrator[7].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][2]~q ;
wire \integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][19]~q ;
wire \integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][20]~q ;
wire \integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][21]~q ;
wire \integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][22]~q ;
wire \integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][23]~q ;
wire \integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][24]~q ;
wire \integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][25]~q ;
wire \integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][26]~q ;
wire \integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][27]~q ;
wire \integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][28]~q ;
wire \integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][29]~q ;
wire \integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][30]~q ;
wire \integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][31]~q ;
wire \integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][32]~q ;
wire \integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][33]~q ;
wire \integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][34]~q ;
wire \integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][35]~q ;
wire \integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][36]~q ;
wire \integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][37]~q ;
wire \integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][38]~q ;
wire \integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][39]~q ;
wire \integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][40]~q ;
wire \integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][41]~q ;
wire \integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][42]~q ;
wire \integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][43]~q ;
wire \integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][44]~q ;
wire \integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][45]~q ;
wire \integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ;
wire \integrator[4].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ;
wire \integrator[5].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ;
wire \integrator[6].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ;
wire \integrator[7].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][1]~q ;
wire \integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][19]~q ;
wire \integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ;
wire \integrator[4].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ;
wire \integrator[5].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ;
wire \integrator[6].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][4]~q ;
wire \integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][20]~q ;
wire \integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][21]~q ;
wire \integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][22]~q ;
wire \integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][23]~q ;
wire \integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][24]~q ;
wire \integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][25]~q ;
wire \integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][26]~q ;
wire \integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][27]~q ;
wire \integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][28]~q ;
wire \integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][29]~q ;
wire \integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][30]~q ;
wire \integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][31]~q ;
wire \integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][32]~q ;
wire \integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][33]~q ;
wire \integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][34]~q ;
wire \integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][35]~q ;
wire \integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][36]~q ;
wire \integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][37]~q ;
wire \integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][38]~q ;
wire \integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][39]~q ;
wire \integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][40]~q ;
wire \integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][41]~q ;
wire \integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][42]~q ;
wire \integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][43]~q ;
wire \integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][44]~q ;
wire \integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][45]~q ;
wire \integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][46]~q ;
wire \integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ;
wire \integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ;
wire \integrator[4].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ;
wire \integrator[5].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ;
wire \integrator[6].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][3]~q ;
wire \integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][19]~q ;
wire \integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ;
wire \integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ;
wire \integrator[4].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ;
wire \integrator[5].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ;
wire \integrator[6].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][2]~q ;
wire \integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][20]~q ;
wire \integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][21]~q ;
wire \integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][22]~q ;
wire \integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][23]~q ;
wire \integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][24]~q ;
wire \integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][25]~q ;
wire \integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][26]~q ;
wire \integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][27]~q ;
wire \integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][28]~q ;
wire \integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][29]~q ;
wire \integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][30]~q ;
wire \integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][31]~q ;
wire \integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][32]~q ;
wire \integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][33]~q ;
wire \integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][34]~q ;
wire \integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][35]~q ;
wire \integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][36]~q ;
wire \integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][37]~q ;
wire \integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][38]~q ;
wire \integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][39]~q ;
wire \integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][40]~q ;
wire \integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][41]~q ;
wire \integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][42]~q ;
wire \integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][43]~q ;
wire \integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][44]~q ;
wire \integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][45]~q ;
wire \integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][46]~q ;
wire \integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ;
wire \integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ;
wire \integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ;
wire \integrator[4].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ;
wire \integrator[5].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ;
wire \integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][19]~q ;
wire \integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ;
wire \integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ;
wire \integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ;
wire \integrator[4].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ;
wire \integrator[5].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][4]~q ;
wire \integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][20]~q ;
wire \integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][21]~q ;
wire \integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][22]~q ;
wire \integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][23]~q ;
wire \integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][24]~q ;
wire \integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][25]~q ;
wire \integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][26]~q ;
wire \integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][27]~q ;
wire \integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][28]~q ;
wire \integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][29]~q ;
wire \integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][30]~q ;
wire \integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][31]~q ;
wire \integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][32]~q ;
wire \integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][33]~q ;
wire \integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][34]~q ;
wire \integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][35]~q ;
wire \integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][36]~q ;
wire \integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][37]~q ;
wire \integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][38]~q ;
wire \integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][39]~q ;
wire \integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][40]~q ;
wire \integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][41]~q ;
wire \integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][42]~q ;
wire \integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][43]~q ;
wire \integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][44]~q ;
wire \integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][45]~q ;
wire \integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][46]~q ;
wire \integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ;
wire \integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ;
wire \integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ;
wire \integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ;
wire \integrator[4].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ;
wire \integrator[5].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][3]~q ;
wire \integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ;
wire \integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ;
wire \integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ;
wire \integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ;
wire \integrator[4].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ;
wire \integrator[5].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][2]~q ;
wire \integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ;
wire \integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ;
wire \integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ;
wire \integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ;
wire \integrator[4].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ;
wire \integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ;
wire \integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ;
wire \integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ;
wire \integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ;
wire \integrator[4].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][4]~q ;
wire \integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ;
wire \integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ;
wire \integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ;
wire \integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ;
wire \integrator[4].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][3]~q ;
wire \integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ;
wire \integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ;
wire \integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ;
wire \integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ;
wire \integrator[4].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][2]~q ;
wire \integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ;
wire \integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ;
wire \integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ;
wire \integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ;
wire \integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ;
wire \integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ;
wire \integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ;
wire \integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][4]~q ;
wire \integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ;
wire \integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ;
wire \integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ;
wire \integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][3]~q ;
wire \integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ;
wire \integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ;
wire \integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ;
wire \integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][2]~q ;
wire \integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ;
wire \integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ;
wire \integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][4]~q ;
wire \integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ;
wire \integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ;
wire \integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][3]~q ;
wire \integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ;
wire \integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][4]~q ;
wire \integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][2]~q ;
wire \integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ;
wire \integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][3]~q ;
wire \integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][1]~q ;
wire \integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][4]~q ;
wire \integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][2]~q ;
wire \integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][3]~q ;
wire \integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][1]~q ;
wire \integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][2]~q ;
wire \integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][0]~q ;
wire \integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][1]~q ;
wire \integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][0]~q ;
wire \state~0_combout ;


cic_auk_dspip_integrator \integrator[0].integration (
	.q_b_19(q_b_19),
	.q_b_18(q_b_18),
	.q_b_17(q_b_17),
	.q_b_16(q_b_16),
	.q_b_15(q_b_15),
	.q_b_14(q_b_14),
	.q_b_13(q_b_13),
	.q_b_12(q_b_12),
	.q_b_11(q_b_11),
	.q_b_10(q_b_10),
	.q_b_9(q_b_9),
	.q_b_8(q_b_8),
	.q_b_7(q_b_7),
	.q_b_6(q_b_6),
	.q_b_5(q_b_5),
	.q_b_4(q_b_4),
	.q_b_3(q_b_3),
	.q_b_2(q_b_2),
	.q_b_1(q_b_1),
	.q_b_0(q_b_0),
	.stall_reg(stall_reg),
	.register_fifofifo_data019(\integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][19]~q ),
	.register_fifofifo_data020(\integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][20]~q ),
	.register_fifofifo_data021(\integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][21]~q ),
	.register_fifofifo_data022(\integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][22]~q ),
	.register_fifofifo_data023(\integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][23]~q ),
	.register_fifofifo_data024(\integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][24]~q ),
	.register_fifofifo_data025(\integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][25]~q ),
	.register_fifofifo_data026(\integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][26]~q ),
	.register_fifofifo_data027(\integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][27]~q ),
	.register_fifofifo_data028(\integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][28]~q ),
	.register_fifofifo_data029(\integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][29]~q ),
	.register_fifofifo_data030(\integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][30]~q ),
	.register_fifofifo_data031(\integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][31]~q ),
	.register_fifofifo_data032(\integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][32]~q ),
	.register_fifofifo_data033(\integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][33]~q ),
	.register_fifofifo_data034(\integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][34]~q ),
	.register_fifofifo_data035(\integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][35]~q ),
	.register_fifofifo_data036(\integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][36]~q ),
	.register_fifofifo_data037(\integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][37]~q ),
	.register_fifofifo_data038(\integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][38]~q ),
	.register_fifofifo_data039(\integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][39]~q ),
	.register_fifofifo_data040(\integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][40]~q ),
	.register_fifofifo_data041(\integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][41]~q ),
	.register_fifofifo_data042(\integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][42]~q ),
	.register_fifofifo_data043(\integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][43]~q ),
	.register_fifofifo_data044(\integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][44]~q ),
	.register_fifofifo_data045(\integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][45]~q ),
	.register_fifofifo_data046(\integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][46]~q ),
	.register_fifofifo_data018(\integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ),
	.register_fifofifo_data017(\integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ),
	.register_fifofifo_data016(\integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ),
	.register_fifofifo_data015(\integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ),
	.register_fifofifo_data014(\integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ),
	.register_fifofifo_data013(\integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ),
	.register_fifofifo_data012(\integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ),
	.register_fifofifo_data011(\integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ),
	.register_fifofifo_data010(\integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ),
	.register_fifofifo_data09(\integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ),
	.register_fifofifo_data08(\integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ),
	.register_fifofifo_data07(\integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ),
	.register_fifofifo_data06(\integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ),
	.register_fifofifo_data05(\integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ),
	.register_fifofifo_data04(\integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][4]~q ),
	.register_fifofifo_data03(\integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][3]~q ),
	.register_fifofifo_data02(\integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][2]~q ),
	.register_fifofifo_data01(\integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][1]~q ),
	.register_fifofifo_data00(\integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][0]~q ),
	.clk(clk),
	.reset_n(reset_n));

cic_auk_dspip_integrator_3 \integrator[3].integration (
	.stall_reg(stall_reg),
	.register_fifofifo_data018(\integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ),
	.register_fifofifo_data019(\integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][19]~q ),
	.register_fifofifo_data020(\integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][20]~q ),
	.register_fifofifo_data021(\integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][21]~q ),
	.register_fifofifo_data022(\integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][22]~q ),
	.register_fifofifo_data023(\integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][23]~q ),
	.register_fifofifo_data024(\integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][24]~q ),
	.register_fifofifo_data025(\integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][25]~q ),
	.register_fifofifo_data026(\integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][26]~q ),
	.register_fifofifo_data027(\integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][27]~q ),
	.register_fifofifo_data028(\integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][28]~q ),
	.register_fifofifo_data029(\integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][29]~q ),
	.register_fifofifo_data030(\integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][30]~q ),
	.register_fifofifo_data031(\integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][31]~q ),
	.register_fifofifo_data032(\integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][32]~q ),
	.register_fifofifo_data033(\integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][33]~q ),
	.register_fifofifo_data034(\integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][34]~q ),
	.register_fifofifo_data035(\integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][35]~q ),
	.register_fifofifo_data036(\integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][36]~q ),
	.register_fifofifo_data037(\integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][37]~q ),
	.register_fifofifo_data038(\integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][38]~q ),
	.register_fifofifo_data039(\integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][39]~q ),
	.register_fifofifo_data040(\integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][40]~q ),
	.register_fifofifo_data041(\integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][41]~q ),
	.register_fifofifo_data042(\integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][42]~q ),
	.register_fifofifo_data043(\integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][43]~q ),
	.register_fifofifo_data044(\integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][44]~q ),
	.register_fifofifo_data045(\integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][45]~q ),
	.register_fifofifo_data017(\integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ),
	.register_fifofifo_data0191(\integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][19]~q ),
	.register_fifofifo_data016(\integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ),
	.register_fifofifo_data0201(\integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][20]~q ),
	.register_fifofifo_data0211(\integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][21]~q ),
	.register_fifofifo_data0221(\integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][22]~q ),
	.register_fifofifo_data0231(\integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][23]~q ),
	.register_fifofifo_data0241(\integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][24]~q ),
	.register_fifofifo_data0251(\integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][25]~q ),
	.register_fifofifo_data0261(\integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][26]~q ),
	.register_fifofifo_data0271(\integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][27]~q ),
	.register_fifofifo_data0281(\integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][28]~q ),
	.register_fifofifo_data0291(\integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][29]~q ),
	.register_fifofifo_data0301(\integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][30]~q ),
	.register_fifofifo_data0311(\integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][31]~q ),
	.register_fifofifo_data0321(\integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][32]~q ),
	.register_fifofifo_data0331(\integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][33]~q ),
	.register_fifofifo_data0341(\integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][34]~q ),
	.register_fifofifo_data0351(\integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][35]~q ),
	.register_fifofifo_data0361(\integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][36]~q ),
	.register_fifofifo_data0371(\integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][37]~q ),
	.register_fifofifo_data0381(\integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][38]~q ),
	.register_fifofifo_data0391(\integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][39]~q ),
	.register_fifofifo_data0401(\integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][40]~q ),
	.register_fifofifo_data0411(\integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][41]~q ),
	.register_fifofifo_data0421(\integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][42]~q ),
	.register_fifofifo_data0431(\integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][43]~q ),
	.register_fifofifo_data0441(\integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][44]~q ),
	.register_fifofifo_data0451(\integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][45]~q ),
	.register_fifofifo_data046(\integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][46]~q ),
	.register_fifofifo_data0181(\integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ),
	.register_fifofifo_data015(\integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ),
	.register_fifofifo_data0171(\integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ),
	.register_fifofifo_data014(\integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ),
	.register_fifofifo_data0161(\integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ),
	.register_fifofifo_data013(\integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ),
	.register_fifofifo_data0151(\integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ),
	.register_fifofifo_data012(\integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ),
	.register_fifofifo_data0141(\integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ),
	.register_fifofifo_data011(\integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ),
	.register_fifofifo_data0131(\integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ),
	.register_fifofifo_data010(\integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ),
	.register_fifofifo_data0121(\integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ),
	.register_fifofifo_data09(\integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ),
	.register_fifofifo_data0111(\integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ),
	.register_fifofifo_data08(\integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ),
	.register_fifofifo_data0101(\integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ),
	.register_fifofifo_data07(\integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ),
	.register_fifofifo_data091(\integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ),
	.register_fifofifo_data06(\integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ),
	.register_fifofifo_data081(\integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ),
	.register_fifofifo_data05(\integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ),
	.register_fifofifo_data071(\integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ),
	.register_fifofifo_data04(\integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][4]~q ),
	.register_fifofifo_data061(\integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ),
	.register_fifofifo_data03(\integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][3]~q ),
	.register_fifofifo_data051(\integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ),
	.register_fifofifo_data02(\integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][2]~q ),
	.register_fifofifo_data047(\integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][4]~q ),
	.register_fifofifo_data0310(\integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][3]~q ),
	.register_fifofifo_data0210(\integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][2]~q ),
	.register_fifofifo_data01(\integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][1]~q ),
	.clk(clk),
	.reset_n(reset_n));

cic_auk_dspip_integrator_2 \integrator[2].integration (
	.stall_reg(stall_reg),
	.register_fifofifo_data019(\integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][19]~q ),
	.register_fifofifo_data020(\integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][20]~q ),
	.register_fifofifo_data021(\integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][21]~q ),
	.register_fifofifo_data022(\integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][22]~q ),
	.register_fifofifo_data023(\integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][23]~q ),
	.register_fifofifo_data024(\integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][24]~q ),
	.register_fifofifo_data025(\integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][25]~q ),
	.register_fifofifo_data026(\integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][26]~q ),
	.register_fifofifo_data027(\integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][27]~q ),
	.register_fifofifo_data028(\integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][28]~q ),
	.register_fifofifo_data029(\integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][29]~q ),
	.register_fifofifo_data030(\integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][30]~q ),
	.register_fifofifo_data031(\integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][31]~q ),
	.register_fifofifo_data032(\integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][32]~q ),
	.register_fifofifo_data033(\integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][33]~q ),
	.register_fifofifo_data034(\integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][34]~q ),
	.register_fifofifo_data035(\integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][35]~q ),
	.register_fifofifo_data036(\integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][36]~q ),
	.register_fifofifo_data037(\integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][37]~q ),
	.register_fifofifo_data038(\integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][38]~q ),
	.register_fifofifo_data039(\integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][39]~q ),
	.register_fifofifo_data040(\integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][40]~q ),
	.register_fifofifo_data041(\integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][41]~q ),
	.register_fifofifo_data042(\integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][42]~q ),
	.register_fifofifo_data043(\integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][43]~q ),
	.register_fifofifo_data044(\integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][44]~q ),
	.register_fifofifo_data045(\integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][45]~q ),
	.register_fifofifo_data046(\integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][46]~q ),
	.register_fifofifo_data018(\integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ),
	.register_fifofifo_data0191(\integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][19]~q ),
	.register_fifofifo_data017(\integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ),
	.register_fifofifo_data0201(\integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][20]~q ),
	.register_fifofifo_data0211(\integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][21]~q ),
	.register_fifofifo_data0221(\integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][22]~q ),
	.register_fifofifo_data0231(\integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][23]~q ),
	.register_fifofifo_data0241(\integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][24]~q ),
	.register_fifofifo_data0251(\integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][25]~q ),
	.register_fifofifo_data0261(\integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][26]~q ),
	.register_fifofifo_data0271(\integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][27]~q ),
	.register_fifofifo_data0281(\integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][28]~q ),
	.register_fifofifo_data0291(\integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][29]~q ),
	.register_fifofifo_data0301(\integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][30]~q ),
	.register_fifofifo_data0311(\integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][31]~q ),
	.register_fifofifo_data0321(\integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][32]~q ),
	.register_fifofifo_data0331(\integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][33]~q ),
	.register_fifofifo_data0341(\integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][34]~q ),
	.register_fifofifo_data0351(\integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][35]~q ),
	.register_fifofifo_data0361(\integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][36]~q ),
	.register_fifofifo_data0371(\integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][37]~q ),
	.register_fifofifo_data0381(\integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][38]~q ),
	.register_fifofifo_data0391(\integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][39]~q ),
	.register_fifofifo_data0401(\integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][40]~q ),
	.register_fifofifo_data0411(\integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][41]~q ),
	.register_fifofifo_data0421(\integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][42]~q ),
	.register_fifofifo_data0431(\integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][43]~q ),
	.register_fifofifo_data0441(\integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][44]~q ),
	.register_fifofifo_data0451(\integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][45]~q ),
	.register_fifofifo_data0461(\integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][46]~q ),
	.register_fifofifo_data0181(\integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ),
	.register_fifofifo_data016(\integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ),
	.register_fifofifo_data0171(\integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ),
	.register_fifofifo_data015(\integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ),
	.register_fifofifo_data0161(\integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ),
	.register_fifofifo_data014(\integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ),
	.register_fifofifo_data0151(\integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ),
	.register_fifofifo_data013(\integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ),
	.register_fifofifo_data0141(\integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ),
	.register_fifofifo_data012(\integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ),
	.register_fifofifo_data0131(\integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ),
	.register_fifofifo_data011(\integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ),
	.register_fifofifo_data0121(\integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ),
	.register_fifofifo_data010(\integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ),
	.register_fifofifo_data0111(\integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ),
	.register_fifofifo_data09(\integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ),
	.register_fifofifo_data0101(\integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ),
	.register_fifofifo_data08(\integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ),
	.register_fifofifo_data091(\integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ),
	.register_fifofifo_data07(\integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ),
	.register_fifofifo_data081(\integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ),
	.register_fifofifo_data06(\integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ),
	.register_fifofifo_data071(\integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ),
	.register_fifofifo_data05(\integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ),
	.register_fifofifo_data061(\integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ),
	.register_fifofifo_data04(\integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][4]~q ),
	.register_fifofifo_data051(\integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ),
	.register_fifofifo_data03(\integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][3]~q ),
	.register_fifofifo_data047(\integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][4]~q ),
	.register_fifofifo_data02(\integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][2]~q ),
	.register_fifofifo_data0310(\integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][3]~q ),
	.register_fifofifo_data01(\integrator[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][1]~q ),
	.register_fifofifo_data0210(\integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][2]~q ),
	.register_fifofifo_data0110(\integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][1]~q ),
	.register_fifofifo_data00(\integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][0]~q ),
	.clk(clk),
	.reset_n(reset_n));

cic_auk_dspip_integrator_1 \integrator[1].integration (
	.stall_reg(stall_reg),
	.register_fifofifo_data019(\integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][19]~q ),
	.register_fifofifo_data020(\integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][20]~q ),
	.register_fifofifo_data021(\integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][21]~q ),
	.register_fifofifo_data022(\integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][22]~q ),
	.register_fifofifo_data023(\integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][23]~q ),
	.register_fifofifo_data024(\integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][24]~q ),
	.register_fifofifo_data025(\integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][25]~q ),
	.register_fifofifo_data026(\integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][26]~q ),
	.register_fifofifo_data027(\integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][27]~q ),
	.register_fifofifo_data028(\integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][28]~q ),
	.register_fifofifo_data029(\integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][29]~q ),
	.register_fifofifo_data030(\integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][30]~q ),
	.register_fifofifo_data031(\integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][31]~q ),
	.register_fifofifo_data032(\integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][32]~q ),
	.register_fifofifo_data033(\integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][33]~q ),
	.register_fifofifo_data034(\integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][34]~q ),
	.register_fifofifo_data035(\integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][35]~q ),
	.register_fifofifo_data036(\integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][36]~q ),
	.register_fifofifo_data037(\integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][37]~q ),
	.register_fifofifo_data038(\integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][38]~q ),
	.register_fifofifo_data039(\integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][39]~q ),
	.register_fifofifo_data040(\integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][40]~q ),
	.register_fifofifo_data041(\integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][41]~q ),
	.register_fifofifo_data042(\integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][42]~q ),
	.register_fifofifo_data043(\integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][43]~q ),
	.register_fifofifo_data044(\integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][44]~q ),
	.register_fifofifo_data045(\integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][45]~q ),
	.register_fifofifo_data046(\integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][46]~q ),
	.register_fifofifo_data018(\integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ),
	.register_fifofifo_data0191(\integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][19]~q ),
	.register_fifofifo_data017(\integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ),
	.register_fifofifo_data0201(\integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][20]~q ),
	.register_fifofifo_data0211(\integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][21]~q ),
	.register_fifofifo_data0221(\integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][22]~q ),
	.register_fifofifo_data0231(\integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][23]~q ),
	.register_fifofifo_data0241(\integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][24]~q ),
	.register_fifofifo_data0251(\integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][25]~q ),
	.register_fifofifo_data0261(\integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][26]~q ),
	.register_fifofifo_data0271(\integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][27]~q ),
	.register_fifofifo_data0281(\integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][28]~q ),
	.register_fifofifo_data0291(\integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][29]~q ),
	.register_fifofifo_data0301(\integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][30]~q ),
	.register_fifofifo_data0311(\integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][31]~q ),
	.register_fifofifo_data0321(\integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][32]~q ),
	.register_fifofifo_data0331(\integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][33]~q ),
	.register_fifofifo_data0341(\integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][34]~q ),
	.register_fifofifo_data0351(\integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][35]~q ),
	.register_fifofifo_data0361(\integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][36]~q ),
	.register_fifofifo_data0371(\integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][37]~q ),
	.register_fifofifo_data0381(\integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][38]~q ),
	.register_fifofifo_data0391(\integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][39]~q ),
	.register_fifofifo_data0401(\integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][40]~q ),
	.register_fifofifo_data0411(\integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][41]~q ),
	.register_fifofifo_data0421(\integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][42]~q ),
	.register_fifofifo_data0431(\integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][43]~q ),
	.register_fifofifo_data0441(\integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][44]~q ),
	.register_fifofifo_data0451(\integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][45]~q ),
	.register_fifofifo_data0461(\integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][46]~q ),
	.register_fifofifo_data0181(\integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ),
	.register_fifofifo_data016(\integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ),
	.register_fifofifo_data0171(\integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ),
	.register_fifofifo_data015(\integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ),
	.register_fifofifo_data0161(\integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ),
	.register_fifofifo_data014(\integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ),
	.register_fifofifo_data0151(\integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ),
	.register_fifofifo_data013(\integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ),
	.register_fifofifo_data0141(\integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ),
	.register_fifofifo_data012(\integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ),
	.register_fifofifo_data0131(\integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ),
	.register_fifofifo_data011(\integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ),
	.register_fifofifo_data0121(\integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ),
	.register_fifofifo_data010(\integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ),
	.register_fifofifo_data0111(\integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ),
	.register_fifofifo_data09(\integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ),
	.register_fifofifo_data0101(\integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ),
	.register_fifofifo_data08(\integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ),
	.register_fifofifo_data091(\integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ),
	.register_fifofifo_data07(\integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ),
	.register_fifofifo_data081(\integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ),
	.register_fifofifo_data06(\integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ),
	.register_fifofifo_data071(\integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ),
	.register_fifofifo_data05(\integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ),
	.register_fifofifo_data061(\integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ),
	.register_fifofifo_data04(\integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][4]~q ),
	.register_fifofifo_data051(\integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ),
	.register_fifofifo_data03(\integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][3]~q ),
	.register_fifofifo_data047(\integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][4]~q ),
	.register_fifofifo_data02(\integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][2]~q ),
	.register_fifofifo_data0310(\integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][3]~q ),
	.register_fifofifo_data01(\integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][1]~q ),
	.register_fifofifo_data0210(\integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][2]~q ),
	.register_fifofifo_data00(\integrator[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][0]~q ),
	.register_fifofifo_data0110(\integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][1]~q ),
	.register_fifofifo_data001(\integrator[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][0]~q ),
	.clk(clk),
	.reset_n(reset_n));

cic_auk_dspip_integrator_6 \integrator[6].integration (
	.stall_reg(stall_reg),
	.register_fifofifo_data012(\integrator[6].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ),
	.register_fifofifo_data013(\integrator[6].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ),
	.register_fifofifo_data014(\integrator[6].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ),
	.register_fifofifo_data015(\integrator[6].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ),
	.register_fifofifo_data016(\integrator[6].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ),
	.register_fifofifo_data017(\integrator[6].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ),
	.register_fifofifo_data018(\integrator[6].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ),
	.register_fifofifo_data019(\integrator[6].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][19]~q ),
	.register_fifofifo_data020(\integrator[6].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][20]~q ),
	.register_fifofifo_data021(\integrator[6].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][21]~q ),
	.register_fifofifo_data022(\integrator[6].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][22]~q ),
	.register_fifofifo_data023(\integrator[6].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][23]~q ),
	.register_fifofifo_data024(\integrator[6].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][24]~q ),
	.register_fifofifo_data025(\integrator[6].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][25]~q ),
	.register_fifofifo_data026(\integrator[6].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][26]~q ),
	.register_fifofifo_data027(\integrator[6].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][27]~q ),
	.register_fifofifo_data028(\integrator[6].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][28]~q ),
	.register_fifofifo_data029(\integrator[6].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][29]~q ),
	.register_fifofifo_data030(\integrator[6].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][30]~q ),
	.register_fifofifo_data031(\integrator[6].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][31]~q ),
	.register_fifofifo_data032(\integrator[6].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][32]~q ),
	.register_fifofifo_data033(\integrator[6].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][33]~q ),
	.register_fifofifo_data034(\integrator[6].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][34]~q ),
	.register_fifofifo_data035(\integrator[6].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][35]~q ),
	.register_fifofifo_data036(\integrator[6].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][36]~q ),
	.register_fifofifo_data037(\integrator[6].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][37]~q ),
	.register_fifofifo_data038(\integrator[6].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][38]~q ),
	.register_fifofifo_data039(\integrator[6].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][39]~q ),
	.register_fifofifo_data011(\integrator[6].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ),
	.register_fifofifo_data0141(\integrator[5].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ),
	.register_fifofifo_data010(\integrator[6].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ),
	.register_fifofifo_data0151(\integrator[5].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ),
	.register_fifofifo_data0161(\integrator[5].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ),
	.register_fifofifo_data0171(\integrator[5].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ),
	.register_fifofifo_data0181(\integrator[5].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ),
	.register_fifofifo_data0191(\integrator[5].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][19]~q ),
	.register_fifofifo_data0201(\integrator[5].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][20]~q ),
	.register_fifofifo_data0211(\integrator[5].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][21]~q ),
	.register_fifofifo_data0221(\integrator[5].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][22]~q ),
	.register_fifofifo_data0231(\integrator[5].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][23]~q ),
	.register_fifofifo_data0241(\integrator[5].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][24]~q ),
	.register_fifofifo_data0251(\integrator[5].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][25]~q ),
	.register_fifofifo_data0261(\integrator[5].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][26]~q ),
	.register_fifofifo_data0271(\integrator[5].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][27]~q ),
	.register_fifofifo_data0281(\integrator[5].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][28]~q ),
	.register_fifofifo_data0291(\integrator[5].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][29]~q ),
	.register_fifofifo_data0301(\integrator[5].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][30]~q ),
	.register_fifofifo_data0311(\integrator[5].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][31]~q ),
	.register_fifofifo_data0321(\integrator[5].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][32]~q ),
	.register_fifofifo_data0331(\integrator[5].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][33]~q ),
	.register_fifofifo_data0341(\integrator[5].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][34]~q ),
	.register_fifofifo_data0351(\integrator[5].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][35]~q ),
	.register_fifofifo_data0361(\integrator[5].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][36]~q ),
	.register_fifofifo_data0371(\integrator[5].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][37]~q ),
	.register_fifofifo_data0381(\integrator[5].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][38]~q ),
	.register_fifofifo_data0391(\integrator[5].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][39]~q ),
	.register_fifofifo_data040(\integrator[5].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][40]~q ),
	.register_fifofifo_data041(\integrator[5].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][41]~q ),
	.register_fifofifo_data0131(\integrator[5].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ),
	.register_fifofifo_data09(\integrator[6].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ),
	.register_fifofifo_data0121(\integrator[5].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ),
	.register_fifofifo_data08(\integrator[6].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ),
	.register_fifofifo_data0111(\integrator[5].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ),
	.register_fifofifo_data07(\integrator[6].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ),
	.register_fifofifo_data0101(\integrator[5].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ),
	.register_fifofifo_data06(\integrator[6].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ),
	.register_fifofifo_data091(\integrator[5].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ),
	.register_fifofifo_data05(\integrator[6].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ),
	.register_fifofifo_data081(\integrator[5].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ),
	.register_fifofifo_data04(\integrator[6].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][4]~q ),
	.register_fifofifo_data071(\integrator[5].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ),
	.register_fifofifo_data03(\integrator[6].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][3]~q ),
	.register_fifofifo_data061(\integrator[5].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ),
	.register_fifofifo_data02(\integrator[6].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][2]~q ),
	.register_fifofifo_data051(\integrator[5].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ),
	.register_fifofifo_data042(\integrator[5].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][4]~q ),
	.register_fifofifo_data0310(\integrator[5].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][3]~q ),
	.register_fifofifo_data0210(\integrator[5].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][2]~q ),
	.clk(clk),
	.reset_n(reset_n));

cic_auk_dspip_integrator_5 \integrator[5].integration (
	.stall_reg(stall_reg),
	.register_fifofifo_data014(\integrator[5].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ),
	.register_fifofifo_data015(\integrator[5].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ),
	.register_fifofifo_data016(\integrator[5].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ),
	.register_fifofifo_data017(\integrator[5].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ),
	.register_fifofifo_data018(\integrator[5].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ),
	.register_fifofifo_data019(\integrator[5].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][19]~q ),
	.register_fifofifo_data020(\integrator[5].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][20]~q ),
	.register_fifofifo_data021(\integrator[5].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][21]~q ),
	.register_fifofifo_data022(\integrator[5].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][22]~q ),
	.register_fifofifo_data023(\integrator[5].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][23]~q ),
	.register_fifofifo_data024(\integrator[5].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][24]~q ),
	.register_fifofifo_data025(\integrator[5].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][25]~q ),
	.register_fifofifo_data026(\integrator[5].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][26]~q ),
	.register_fifofifo_data027(\integrator[5].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][27]~q ),
	.register_fifofifo_data028(\integrator[5].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][28]~q ),
	.register_fifofifo_data029(\integrator[5].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][29]~q ),
	.register_fifofifo_data030(\integrator[5].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][30]~q ),
	.register_fifofifo_data031(\integrator[5].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][31]~q ),
	.register_fifofifo_data032(\integrator[5].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][32]~q ),
	.register_fifofifo_data033(\integrator[5].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][33]~q ),
	.register_fifofifo_data034(\integrator[5].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][34]~q ),
	.register_fifofifo_data035(\integrator[5].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][35]~q ),
	.register_fifofifo_data036(\integrator[5].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][36]~q ),
	.register_fifofifo_data037(\integrator[5].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][37]~q ),
	.register_fifofifo_data038(\integrator[5].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][38]~q ),
	.register_fifofifo_data039(\integrator[5].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][39]~q ),
	.register_fifofifo_data040(\integrator[5].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][40]~q ),
	.register_fifofifo_data041(\integrator[5].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][41]~q ),
	.register_fifofifo_data013(\integrator[5].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ),
	.register_fifofifo_data0161(\integrator[4].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ),
	.register_fifofifo_data012(\integrator[5].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ),
	.register_fifofifo_data0171(\integrator[4].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ),
	.register_fifofifo_data0181(\integrator[4].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ),
	.register_fifofifo_data0191(\integrator[4].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][19]~q ),
	.register_fifofifo_data0201(\integrator[4].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][20]~q ),
	.register_fifofifo_data0211(\integrator[4].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][21]~q ),
	.register_fifofifo_data0221(\integrator[4].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][22]~q ),
	.register_fifofifo_data0231(\integrator[4].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][23]~q ),
	.register_fifofifo_data0241(\integrator[4].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][24]~q ),
	.register_fifofifo_data0251(\integrator[4].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][25]~q ),
	.register_fifofifo_data0261(\integrator[4].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][26]~q ),
	.register_fifofifo_data0271(\integrator[4].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][27]~q ),
	.register_fifofifo_data0281(\integrator[4].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][28]~q ),
	.register_fifofifo_data0291(\integrator[4].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][29]~q ),
	.register_fifofifo_data0301(\integrator[4].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][30]~q ),
	.register_fifofifo_data0311(\integrator[4].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][31]~q ),
	.register_fifofifo_data0321(\integrator[4].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][32]~q ),
	.register_fifofifo_data0331(\integrator[4].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][33]~q ),
	.register_fifofifo_data0341(\integrator[4].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][34]~q ),
	.register_fifofifo_data0351(\integrator[4].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][35]~q ),
	.register_fifofifo_data0361(\integrator[4].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][36]~q ),
	.register_fifofifo_data0371(\integrator[4].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][37]~q ),
	.register_fifofifo_data0381(\integrator[4].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][38]~q ),
	.register_fifofifo_data0391(\integrator[4].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][39]~q ),
	.register_fifofifo_data0401(\integrator[4].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][40]~q ),
	.register_fifofifo_data0411(\integrator[4].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][41]~q ),
	.register_fifofifo_data042(\integrator[4].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][42]~q ),
	.register_fifofifo_data043(\integrator[4].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][43]~q ),
	.register_fifofifo_data0151(\integrator[4].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ),
	.register_fifofifo_data011(\integrator[5].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ),
	.register_fifofifo_data0141(\integrator[4].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ),
	.register_fifofifo_data010(\integrator[5].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ),
	.register_fifofifo_data0131(\integrator[4].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ),
	.register_fifofifo_data09(\integrator[5].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ),
	.register_fifofifo_data0121(\integrator[4].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ),
	.register_fifofifo_data08(\integrator[5].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ),
	.register_fifofifo_data0111(\integrator[4].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ),
	.register_fifofifo_data07(\integrator[5].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ),
	.register_fifofifo_data0101(\integrator[4].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ),
	.register_fifofifo_data06(\integrator[5].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ),
	.register_fifofifo_data091(\integrator[4].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ),
	.register_fifofifo_data05(\integrator[5].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ),
	.register_fifofifo_data081(\integrator[4].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ),
	.register_fifofifo_data04(\integrator[5].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][4]~q ),
	.register_fifofifo_data071(\integrator[4].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ),
	.register_fifofifo_data03(\integrator[5].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][3]~q ),
	.register_fifofifo_data061(\integrator[4].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ),
	.register_fifofifo_data02(\integrator[5].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][2]~q ),
	.register_fifofifo_data051(\integrator[4].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ),
	.register_fifofifo_data044(\integrator[4].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][4]~q ),
	.register_fifofifo_data0310(\integrator[4].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][3]~q ),
	.register_fifofifo_data0210(\integrator[4].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][2]~q ),
	.clk(clk),
	.reset_n(reset_n));

cic_auk_dspip_integrator_4 \integrator[4].integration (
	.stall_reg(stall_reg),
	.register_fifofifo_data016(\integrator[4].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ),
	.register_fifofifo_data017(\integrator[4].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ),
	.register_fifofifo_data018(\integrator[4].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ),
	.register_fifofifo_data019(\integrator[4].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][19]~q ),
	.register_fifofifo_data020(\integrator[4].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][20]~q ),
	.register_fifofifo_data021(\integrator[4].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][21]~q ),
	.register_fifofifo_data022(\integrator[4].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][22]~q ),
	.register_fifofifo_data023(\integrator[4].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][23]~q ),
	.register_fifofifo_data024(\integrator[4].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][24]~q ),
	.register_fifofifo_data025(\integrator[4].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][25]~q ),
	.register_fifofifo_data026(\integrator[4].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][26]~q ),
	.register_fifofifo_data027(\integrator[4].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][27]~q ),
	.register_fifofifo_data028(\integrator[4].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][28]~q ),
	.register_fifofifo_data029(\integrator[4].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][29]~q ),
	.register_fifofifo_data030(\integrator[4].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][30]~q ),
	.register_fifofifo_data031(\integrator[4].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][31]~q ),
	.register_fifofifo_data032(\integrator[4].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][32]~q ),
	.register_fifofifo_data033(\integrator[4].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][33]~q ),
	.register_fifofifo_data034(\integrator[4].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][34]~q ),
	.register_fifofifo_data035(\integrator[4].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][35]~q ),
	.register_fifofifo_data036(\integrator[4].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][36]~q ),
	.register_fifofifo_data037(\integrator[4].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][37]~q ),
	.register_fifofifo_data038(\integrator[4].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][38]~q ),
	.register_fifofifo_data039(\integrator[4].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][39]~q ),
	.register_fifofifo_data040(\integrator[4].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][40]~q ),
	.register_fifofifo_data041(\integrator[4].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][41]~q ),
	.register_fifofifo_data042(\integrator[4].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][42]~q ),
	.register_fifofifo_data043(\integrator[4].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][43]~q ),
	.register_fifofifo_data015(\integrator[4].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ),
	.register_fifofifo_data0181(\integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ),
	.register_fifofifo_data014(\integrator[4].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ),
	.register_fifofifo_data0191(\integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][19]~q ),
	.register_fifofifo_data0201(\integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][20]~q ),
	.register_fifofifo_data0211(\integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][21]~q ),
	.register_fifofifo_data0221(\integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][22]~q ),
	.register_fifofifo_data0231(\integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][23]~q ),
	.register_fifofifo_data0241(\integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][24]~q ),
	.register_fifofifo_data0251(\integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][25]~q ),
	.register_fifofifo_data0261(\integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][26]~q ),
	.register_fifofifo_data0271(\integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][27]~q ),
	.register_fifofifo_data0281(\integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][28]~q ),
	.register_fifofifo_data0291(\integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][29]~q ),
	.register_fifofifo_data0301(\integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][30]~q ),
	.register_fifofifo_data0311(\integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][31]~q ),
	.register_fifofifo_data0321(\integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][32]~q ),
	.register_fifofifo_data0331(\integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][33]~q ),
	.register_fifofifo_data0341(\integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][34]~q ),
	.register_fifofifo_data0351(\integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][35]~q ),
	.register_fifofifo_data0361(\integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][36]~q ),
	.register_fifofifo_data0371(\integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][37]~q ),
	.register_fifofifo_data0381(\integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][38]~q ),
	.register_fifofifo_data0391(\integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][39]~q ),
	.register_fifofifo_data0401(\integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][40]~q ),
	.register_fifofifo_data0411(\integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][41]~q ),
	.register_fifofifo_data0421(\integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][42]~q ),
	.register_fifofifo_data0431(\integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][43]~q ),
	.register_fifofifo_data044(\integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][44]~q ),
	.register_fifofifo_data045(\integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][45]~q ),
	.register_fifofifo_data0171(\integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ),
	.register_fifofifo_data013(\integrator[4].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ),
	.register_fifofifo_data0161(\integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ),
	.register_fifofifo_data012(\integrator[4].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ),
	.register_fifofifo_data0151(\integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ),
	.register_fifofifo_data011(\integrator[4].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ),
	.register_fifofifo_data0141(\integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ),
	.register_fifofifo_data010(\integrator[4].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ),
	.register_fifofifo_data0131(\integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ),
	.register_fifofifo_data09(\integrator[4].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ),
	.register_fifofifo_data0121(\integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ),
	.register_fifofifo_data08(\integrator[4].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ),
	.register_fifofifo_data0111(\integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ),
	.register_fifofifo_data07(\integrator[4].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ),
	.register_fifofifo_data0101(\integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ),
	.register_fifofifo_data06(\integrator[4].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ),
	.register_fifofifo_data091(\integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ),
	.register_fifofifo_data05(\integrator[4].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ),
	.register_fifofifo_data081(\integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ),
	.register_fifofifo_data04(\integrator[4].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][4]~q ),
	.register_fifofifo_data071(\integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ),
	.register_fifofifo_data03(\integrator[4].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][3]~q ),
	.register_fifofifo_data061(\integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ),
	.register_fifofifo_data02(\integrator[4].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][2]~q ),
	.register_fifofifo_data051(\integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ),
	.register_fifofifo_data046(\integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][4]~q ),
	.register_fifofifo_data0310(\integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][3]~q ),
	.register_fifofifo_data0210(\integrator[3].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][2]~q ),
	.clk(clk),
	.reset_n(reset_n));

cic_auk_dspip_channel_buffer fifo_regulator(
	.sample_state_0(\sample_state[0]~q ),
	.q({\fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[37] ,\fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[36] ,\fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[35] ,
\fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[34] ,\fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[33] ,\fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[32] ,
\fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[31] ,\fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[30] ,\fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[29] ,
\fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[28] ,\fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[27] ,\fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[26] ,
\fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[25] ,\fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[24] ,\fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[23] ,
\fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[22] ,\fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[21] ,\fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[20] ,
\fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[19] ,\fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[18] ,\fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[17] ,
\fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[16] ,\fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[15] ,\fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[14] ,
\fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[13] ,\fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[12] ,\fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[11] ,
\fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[10] ,\fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[9] ,\fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[8] ,
\fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[7] ,\fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[6] ,\fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[5] ,
\fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[4] ,\fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[3] ,\fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[2] ,
\fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[1] ,q_unconnected_wire_0}),
	.stall_reg(stall_reg),
	.fifo_rdreq(\fifo_rdreq~q ),
	.valid_rreq(\fifo_regulator|buffer_FIFO|auto_generated|dpfifo|valid_rreq~0_combout ),
	.count_0(\vrc_en_0.first_dsample|counter_fs_inst|count[0]~q ),
	.count_3(\vrc_en_0.first_dsample|counter_fs_inst|count[3]~q ),
	.count_1(\vrc_en_0.first_dsample|counter_fs_inst|count[1]~q ),
	.count_2(\vrc_en_0.first_dsample|counter_fs_inst|count[2]~q ),
	.valid_wreq(\fifo_regulator|buffer_FIFO|auto_generated|dpfifo|valid_wreq~0_combout ),
	.data({\integrator[7].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][37]~q ,\integrator[7].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][36]~q ,
\integrator[7].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][35]~q ,\integrator[7].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][34]~q ,
\integrator[7].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][33]~q ,\integrator[7].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][32]~q ,
\integrator[7].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][31]~q ,\integrator[7].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][30]~q ,
\integrator[7].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][29]~q ,\integrator[7].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][28]~q ,
\integrator[7].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][27]~q ,\integrator[7].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][26]~q ,
\integrator[7].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][25]~q ,\integrator[7].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][24]~q ,
\integrator[7].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][23]~q ,\integrator[7].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][22]~q ,
\integrator[7].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][21]~q ,\integrator[7].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][20]~q ,
\integrator[7].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][19]~q ,\integrator[7].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ,
\integrator[7].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ,\integrator[7].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ,
\integrator[7].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ,\integrator[7].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ,
\integrator[7].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ,\integrator[7].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ,
\integrator[7].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ,\integrator[7].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ,
\integrator[7].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ,\integrator[7].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ,
\integrator[7].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ,\integrator[7].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ,
\integrator[7].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ,\integrator[7].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][4]~q ,
\integrator[7].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][3]~q ,\integrator[7].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][2]~q ,
\integrator[7].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][1]~q ,gnd}),
	.clk(clk),
	.clr(reset_n));

cic_auk_dspip_downsample \vrc_en_0.first_dsample (
	.sample_state_0(\sample_state[0]~q ),
	.stall_reg(stall_reg),
	.count_0(\vrc_en_0.first_dsample|counter_fs_inst|count[0]~q ),
	.count_3(\vrc_en_0.first_dsample|counter_fs_inst|count[3]~q ),
	.count_1(\vrc_en_0.first_dsample|counter_fs_inst|count[1]~q ),
	.count_2(\vrc_en_0.first_dsample|counter_fs_inst|count[2]~q ),
	.clk(clk),
	.reset_n(reset_n));

cic_auk_dspip_integrator_7 \integrator[7].integration (
	.stall_reg(stall_reg),
	.register_fifofifo_data010(\integrator[7].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ),
	.register_fifofifo_data011(\integrator[7].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ),
	.register_fifofifo_data012(\integrator[7].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ),
	.register_fifofifo_data013(\integrator[7].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ),
	.register_fifofifo_data014(\integrator[7].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ),
	.register_fifofifo_data015(\integrator[7].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ),
	.register_fifofifo_data016(\integrator[7].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ),
	.register_fifofifo_data017(\integrator[7].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ),
	.register_fifofifo_data018(\integrator[7].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ),
	.register_fifofifo_data019(\integrator[7].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][19]~q ),
	.register_fifofifo_data020(\integrator[7].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][20]~q ),
	.register_fifofifo_data021(\integrator[7].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][21]~q ),
	.register_fifofifo_data022(\integrator[7].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][22]~q ),
	.register_fifofifo_data023(\integrator[7].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][23]~q ),
	.register_fifofifo_data024(\integrator[7].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][24]~q ),
	.register_fifofifo_data025(\integrator[7].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][25]~q ),
	.register_fifofifo_data026(\integrator[7].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][26]~q ),
	.register_fifofifo_data027(\integrator[7].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][27]~q ),
	.register_fifofifo_data028(\integrator[7].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][28]~q ),
	.register_fifofifo_data029(\integrator[7].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][29]~q ),
	.register_fifofifo_data030(\integrator[7].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][30]~q ),
	.register_fifofifo_data031(\integrator[7].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][31]~q ),
	.register_fifofifo_data032(\integrator[7].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][32]~q ),
	.register_fifofifo_data033(\integrator[7].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][33]~q ),
	.register_fifofifo_data034(\integrator[7].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][34]~q ),
	.register_fifofifo_data035(\integrator[7].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][35]~q ),
	.register_fifofifo_data036(\integrator[7].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][36]~q ),
	.register_fifofifo_data037(\integrator[7].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][37]~q ),
	.register_fifofifo_data09(\integrator[7].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ),
	.register_fifofifo_data0121(\integrator[6].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ),
	.register_fifofifo_data08(\integrator[7].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ),
	.register_fifofifo_data0131(\integrator[6].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ),
	.register_fifofifo_data0141(\integrator[6].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ),
	.register_fifofifo_data0151(\integrator[6].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ),
	.register_fifofifo_data0161(\integrator[6].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ),
	.register_fifofifo_data0171(\integrator[6].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ),
	.register_fifofifo_data0181(\integrator[6].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ),
	.register_fifofifo_data0191(\integrator[6].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][19]~q ),
	.register_fifofifo_data0201(\integrator[6].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][20]~q ),
	.register_fifofifo_data0211(\integrator[6].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][21]~q ),
	.register_fifofifo_data0221(\integrator[6].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][22]~q ),
	.register_fifofifo_data0231(\integrator[6].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][23]~q ),
	.register_fifofifo_data0241(\integrator[6].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][24]~q ),
	.register_fifofifo_data0251(\integrator[6].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][25]~q ),
	.register_fifofifo_data0261(\integrator[6].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][26]~q ),
	.register_fifofifo_data0271(\integrator[6].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][27]~q ),
	.register_fifofifo_data0281(\integrator[6].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][28]~q ),
	.register_fifofifo_data0291(\integrator[6].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][29]~q ),
	.register_fifofifo_data0301(\integrator[6].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][30]~q ),
	.register_fifofifo_data0311(\integrator[6].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][31]~q ),
	.register_fifofifo_data0321(\integrator[6].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][32]~q ),
	.register_fifofifo_data0331(\integrator[6].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][33]~q ),
	.register_fifofifo_data0341(\integrator[6].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][34]~q ),
	.register_fifofifo_data0351(\integrator[6].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][35]~q ),
	.register_fifofifo_data0361(\integrator[6].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][36]~q ),
	.register_fifofifo_data0371(\integrator[6].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][37]~q ),
	.register_fifofifo_data038(\integrator[6].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][38]~q ),
	.register_fifofifo_data039(\integrator[6].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][39]~q ),
	.register_fifofifo_data0111(\integrator[6].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ),
	.register_fifofifo_data07(\integrator[7].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ),
	.register_fifofifo_data0101(\integrator[6].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ),
	.register_fifofifo_data06(\integrator[7].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ),
	.register_fifofifo_data091(\integrator[6].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ),
	.register_fifofifo_data05(\integrator[7].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ),
	.register_fifofifo_data081(\integrator[6].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ),
	.register_fifofifo_data04(\integrator[7].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][4]~q ),
	.register_fifofifo_data071(\integrator[6].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ),
	.register_fifofifo_data03(\integrator[7].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][3]~q ),
	.register_fifofifo_data061(\integrator[6].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ),
	.register_fifofifo_data02(\integrator[7].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][2]~q ),
	.register_fifofifo_data051(\integrator[6].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ),
	.register_fifofifo_data01(\integrator[7].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][1]~q ),
	.register_fifofifo_data041(\integrator[6].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][4]~q ),
	.register_fifofifo_data0310(\integrator[6].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][3]~q ),
	.register_fifofifo_data0210(\integrator[6].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][2]~q ),
	.clk(clk),
	.reset_n(reset_n));

cic_auk_dspip_differentiator_1 \differentiate_stages[1].auk_dsp_diff (
	.dout_valid1(\differentiate_stages[1].auk_dsp_diff|dout_valid~q ),
	.dout_valid2(\differentiate_stages[0].auk_dsp_diff|dout_valid~q ),
	.dout_8(\differentiate_stages[1].auk_dsp_diff|dout[8]~q ),
	.dout_9(\differentiate_stages[1].auk_dsp_diff|dout[9]~q ),
	.dout_10(\differentiate_stages[1].auk_dsp_diff|dout[10]~q ),
	.dout_11(\differentiate_stages[1].auk_dsp_diff|dout[11]~q ),
	.dout_12(\differentiate_stages[1].auk_dsp_diff|dout[12]~q ),
	.dout_13(\differentiate_stages[1].auk_dsp_diff|dout[13]~q ),
	.dout_14(\differentiate_stages[1].auk_dsp_diff|dout[14]~q ),
	.dout_15(\differentiate_stages[1].auk_dsp_diff|dout[15]~q ),
	.dout_16(\differentiate_stages[1].auk_dsp_diff|dout[16]~q ),
	.dout_17(\differentiate_stages[1].auk_dsp_diff|dout[17]~q ),
	.dout_18(\differentiate_stages[1].auk_dsp_diff|dout[18]~q ),
	.dout_19(\differentiate_stages[1].auk_dsp_diff|dout[19]~q ),
	.dout_20(\differentiate_stages[1].auk_dsp_diff|dout[20]~q ),
	.dout_21(\differentiate_stages[1].auk_dsp_diff|dout[21]~q ),
	.dout_22(\differentiate_stages[1].auk_dsp_diff|dout[22]~q ),
	.dout_23(\differentiate_stages[1].auk_dsp_diff|dout[23]~q ),
	.dout_24(\differentiate_stages[1].auk_dsp_diff|dout[24]~q ),
	.dout_25(\differentiate_stages[1].auk_dsp_diff|dout[25]~q ),
	.dout_26(\differentiate_stages[1].auk_dsp_diff|dout[26]~q ),
	.dout_27(\differentiate_stages[1].auk_dsp_diff|dout[27]~q ),
	.dout_28(\differentiate_stages[1].auk_dsp_diff|dout[28]~q ),
	.dout_29(\differentiate_stages[1].auk_dsp_diff|dout[29]~q ),
	.dout_30(\differentiate_stages[1].auk_dsp_diff|dout[30]~q ),
	.dout_31(\differentiate_stages[1].auk_dsp_diff|dout[31]~q ),
	.dout_32(\differentiate_stages[1].auk_dsp_diff|dout[32]~q ),
	.dout_33(\differentiate_stages[1].auk_dsp_diff|dout[33]~q ),
	.dout_34(\differentiate_stages[1].auk_dsp_diff|dout[34]~q ),
	.dout_35(\differentiate_stages[1].auk_dsp_diff|dout[35]~q ),
	.dout_7(\differentiate_stages[1].auk_dsp_diff|dout[7]~q ),
	.dout_91(\differentiate_stages[0].auk_dsp_diff|dout[9]~q ),
	.dout_6(\differentiate_stages[1].auk_dsp_diff|dout[6]~q ),
	.dout_101(\differentiate_stages[0].auk_dsp_diff|dout[10]~q ),
	.dout_111(\differentiate_stages[0].auk_dsp_diff|dout[11]~q ),
	.dout_121(\differentiate_stages[0].auk_dsp_diff|dout[12]~q ),
	.dout_131(\differentiate_stages[0].auk_dsp_diff|dout[13]~q ),
	.dout_141(\differentiate_stages[0].auk_dsp_diff|dout[14]~q ),
	.dout_151(\differentiate_stages[0].auk_dsp_diff|dout[15]~q ),
	.dout_161(\differentiate_stages[0].auk_dsp_diff|dout[16]~q ),
	.dout_171(\differentiate_stages[0].auk_dsp_diff|dout[17]~q ),
	.dout_181(\differentiate_stages[0].auk_dsp_diff|dout[18]~q ),
	.dout_191(\differentiate_stages[0].auk_dsp_diff|dout[19]~q ),
	.dout_201(\differentiate_stages[0].auk_dsp_diff|dout[20]~q ),
	.dout_211(\differentiate_stages[0].auk_dsp_diff|dout[21]~q ),
	.dout_221(\differentiate_stages[0].auk_dsp_diff|dout[22]~q ),
	.dout_231(\differentiate_stages[0].auk_dsp_diff|dout[23]~q ),
	.dout_241(\differentiate_stages[0].auk_dsp_diff|dout[24]~q ),
	.dout_251(\differentiate_stages[0].auk_dsp_diff|dout[25]~q ),
	.dout_261(\differentiate_stages[0].auk_dsp_diff|dout[26]~q ),
	.dout_271(\differentiate_stages[0].auk_dsp_diff|dout[27]~q ),
	.dout_281(\differentiate_stages[0].auk_dsp_diff|dout[28]~q ),
	.dout_291(\differentiate_stages[0].auk_dsp_diff|dout[29]~q ),
	.dout_301(\differentiate_stages[0].auk_dsp_diff|dout[30]~q ),
	.dout_311(\differentiate_stages[0].auk_dsp_diff|dout[31]~q ),
	.dout_321(\differentiate_stages[0].auk_dsp_diff|dout[32]~q ),
	.dout_331(\differentiate_stages[0].auk_dsp_diff|dout[33]~q ),
	.dout_341(\differentiate_stages[0].auk_dsp_diff|dout[34]~q ),
	.dout_351(\differentiate_stages[0].auk_dsp_diff|dout[35]~q ),
	.dout_36(\differentiate_stages[0].auk_dsp_diff|dout[36]~q ),
	.dout_81(\differentiate_stages[0].auk_dsp_diff|dout[8]~q ),
	.dout_5(\differentiate_stages[1].auk_dsp_diff|dout[5]~q ),
	.dout_71(\differentiate_stages[0].auk_dsp_diff|dout[7]~q ),
	.dout_4(\differentiate_stages[1].auk_dsp_diff|dout[4]~q ),
	.dout_61(\differentiate_stages[0].auk_dsp_diff|dout[6]~q ),
	.dout_3(\differentiate_stages[1].auk_dsp_diff|dout[3]~q ),
	.dout_51(\differentiate_stages[0].auk_dsp_diff|dout[5]~q ),
	.dout_2(\differentiate_stages[1].auk_dsp_diff|dout[2]~q ),
	.dout_41(\differentiate_stages[0].auk_dsp_diff|dout[4]~q ),
	.dout_1(\differentiate_stages[1].auk_dsp_diff|dout[1]~q ),
	.dout_37(\differentiate_stages[0].auk_dsp_diff|dout[3]~q ),
	.dout_210(\differentiate_stages[0].auk_dsp_diff|dout[2]~q ),
	.dout_110(\differentiate_stages[0].auk_dsp_diff|dout[1]~q ),
	.stall_reg(stall_reg),
	.dout_valid3(\differentiate_stages[7].auk_dsp_diff|dout_valid~0_combout ),
	.clk(clk),
	.reset_n(reset_n));

cic_auk_dspip_differentiator \differentiate_stages[0].auk_dsp_diff (
	.dout_valid1(\differentiate_stages[0].auk_dsp_diff|dout_valid~q ),
	.dout_9(\differentiate_stages[0].auk_dsp_diff|dout[9]~q ),
	.dout_10(\differentiate_stages[0].auk_dsp_diff|dout[10]~q ),
	.dout_11(\differentiate_stages[0].auk_dsp_diff|dout[11]~q ),
	.dout_12(\differentiate_stages[0].auk_dsp_diff|dout[12]~q ),
	.dout_13(\differentiate_stages[0].auk_dsp_diff|dout[13]~q ),
	.dout_14(\differentiate_stages[0].auk_dsp_diff|dout[14]~q ),
	.dout_15(\differentiate_stages[0].auk_dsp_diff|dout[15]~q ),
	.dout_16(\differentiate_stages[0].auk_dsp_diff|dout[16]~q ),
	.dout_17(\differentiate_stages[0].auk_dsp_diff|dout[17]~q ),
	.dout_18(\differentiate_stages[0].auk_dsp_diff|dout[18]~q ),
	.dout_19(\differentiate_stages[0].auk_dsp_diff|dout[19]~q ),
	.dout_20(\differentiate_stages[0].auk_dsp_diff|dout[20]~q ),
	.dout_21(\differentiate_stages[0].auk_dsp_diff|dout[21]~q ),
	.dout_22(\differentiate_stages[0].auk_dsp_diff|dout[22]~q ),
	.dout_23(\differentiate_stages[0].auk_dsp_diff|dout[23]~q ),
	.dout_24(\differentiate_stages[0].auk_dsp_diff|dout[24]~q ),
	.dout_25(\differentiate_stages[0].auk_dsp_diff|dout[25]~q ),
	.dout_26(\differentiate_stages[0].auk_dsp_diff|dout[26]~q ),
	.dout_27(\differentiate_stages[0].auk_dsp_diff|dout[27]~q ),
	.dout_28(\differentiate_stages[0].auk_dsp_diff|dout[28]~q ),
	.dout_29(\differentiate_stages[0].auk_dsp_diff|dout[29]~q ),
	.dout_30(\differentiate_stages[0].auk_dsp_diff|dout[30]~q ),
	.dout_31(\differentiate_stages[0].auk_dsp_diff|dout[31]~q ),
	.dout_32(\differentiate_stages[0].auk_dsp_diff|dout[32]~q ),
	.dout_33(\differentiate_stages[0].auk_dsp_diff|dout[33]~q ),
	.dout_34(\differentiate_stages[0].auk_dsp_diff|dout[34]~q ),
	.dout_35(\differentiate_stages[0].auk_dsp_diff|dout[35]~q ),
	.dout_36(\differentiate_stages[0].auk_dsp_diff|dout[36]~q ),
	.dout_8(\differentiate_stages[0].auk_dsp_diff|dout[8]~q ),
	.q_b_10(\fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[10] ),
	.dout_7(\differentiate_stages[0].auk_dsp_diff|dout[7]~q ),
	.q_b_11(\fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[11] ),
	.q_b_12(\fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[12] ),
	.q_b_13(\fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[13] ),
	.q_b_14(\fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[14] ),
	.q_b_15(\fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[15] ),
	.q_b_16(\fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[16] ),
	.q_b_17(\fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[17] ),
	.q_b_18(\fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[18] ),
	.q_b_19(\fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[19] ),
	.q_b_20(\fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[20] ),
	.q_b_21(\fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[21] ),
	.q_b_22(\fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[22] ),
	.q_b_23(\fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[23] ),
	.q_b_24(\fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[24] ),
	.q_b_25(\fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[25] ),
	.q_b_26(\fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[26] ),
	.q_b_27(\fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[27] ),
	.q_b_28(\fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[28] ),
	.q_b_29(\fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[29] ),
	.q_b_30(\fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[30] ),
	.q_b_31(\fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[31] ),
	.q_b_32(\fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[32] ),
	.q_b_33(\fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[33] ),
	.q_b_34(\fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[34] ),
	.q_b_35(\fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[35] ),
	.q_b_36(\fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[36] ),
	.q_b_37(\fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[37] ),
	.q_b_9(\fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[9] ),
	.dout_6(\differentiate_stages[0].auk_dsp_diff|dout[6]~q ),
	.q_b_8(\fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[8] ),
	.dout_5(\differentiate_stages[0].auk_dsp_diff|dout[5]~q ),
	.q_b_7(\fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[7] ),
	.dout_4(\differentiate_stages[0].auk_dsp_diff|dout[4]~q ),
	.q_b_6(\fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[6] ),
	.dout_3(\differentiate_stages[0].auk_dsp_diff|dout[3]~q ),
	.q_b_5(\fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[5] ),
	.dout_2(\differentiate_stages[0].auk_dsp_diff|dout[2]~q ),
	.q_b_4(\fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[4] ),
	.dout_1(\differentiate_stages[0].auk_dsp_diff|dout[1]~q ),
	.q_b_3(\fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[3] ),
	.q_b_2(\fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[2] ),
	.q_b_1(\fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[1] ),
	.stall_reg(stall_reg),
	.dout_valid2(\differentiate_stages[7].auk_dsp_diff|dout_valid~0_combout ),
	.ena_diff_s_1(\ena_diff_s[1]~q ),
	.clk(clk),
	.reset_n(reset_n));

cic_counter_module_3 latency_cnt_inst(
	.stall_reg(stall_reg),
	.count_0(\latency_cnt_inst|count[0]~q ),
	.count_1(\latency_cnt_inst|count[1]~q ),
	.count_2(\latency_cnt_inst|count[2]~q ),
	.count_3(\latency_cnt_inst|count[3]~q ),
	.count_4(\latency_cnt_inst|count[4]~q ),
	.Equal0(\latency_cnt_inst|Equal0~0_combout ),
	.sample_state(\sample_state~0_combout ),
	.clk(clk),
	.reset_n(reset_n));

cic_auk_dspip_differentiator_5 \differentiate_stages[5].auk_dsp_diff (
	.dout_valid1(\differentiate_stages[5].auk_dsp_diff|dout_valid~q ),
	.dout_valid2(\differentiate_stages[4].auk_dsp_diff|dout_valid~q ),
	.dout_5(\differentiate_stages[5].auk_dsp_diff|dout[5]~q ),
	.dout_6(\differentiate_stages[5].auk_dsp_diff|dout[6]~q ),
	.dout_7(\differentiate_stages[5].auk_dsp_diff|dout[7]~q ),
	.dout_8(\differentiate_stages[5].auk_dsp_diff|dout[8]~q ),
	.dout_9(\differentiate_stages[5].auk_dsp_diff|dout[9]~q ),
	.dout_10(\differentiate_stages[5].auk_dsp_diff|dout[10]~q ),
	.dout_11(\differentiate_stages[5].auk_dsp_diff|dout[11]~q ),
	.dout_12(\differentiate_stages[5].auk_dsp_diff|dout[12]~q ),
	.dout_13(\differentiate_stages[5].auk_dsp_diff|dout[13]~q ),
	.dout_14(\differentiate_stages[5].auk_dsp_diff|dout[14]~q ),
	.dout_15(\differentiate_stages[5].auk_dsp_diff|dout[15]~q ),
	.dout_16(\differentiate_stages[5].auk_dsp_diff|dout[16]~q ),
	.dout_17(\differentiate_stages[5].auk_dsp_diff|dout[17]~q ),
	.dout_18(\differentiate_stages[5].auk_dsp_diff|dout[18]~q ),
	.dout_19(\differentiate_stages[5].auk_dsp_diff|dout[19]~q ),
	.dout_20(\differentiate_stages[5].auk_dsp_diff|dout[20]~q ),
	.dout_21(\differentiate_stages[5].auk_dsp_diff|dout[21]~q ),
	.dout_22(\differentiate_stages[5].auk_dsp_diff|dout[22]~q ),
	.dout_23(\differentiate_stages[5].auk_dsp_diff|dout[23]~q ),
	.dout_24(\differentiate_stages[5].auk_dsp_diff|dout[24]~q ),
	.dout_25(\differentiate_stages[5].auk_dsp_diff|dout[25]~q ),
	.dout_26(\differentiate_stages[5].auk_dsp_diff|dout[26]~q ),
	.dout_27(\differentiate_stages[5].auk_dsp_diff|dout[27]~q ),
	.dout_28(\differentiate_stages[5].auk_dsp_diff|dout[28]~q ),
	.dout_29(\differentiate_stages[5].auk_dsp_diff|dout[29]~q ),
	.dout_30(\differentiate_stages[5].auk_dsp_diff|dout[30]~q ),
	.dout_31(\differentiate_stages[5].auk_dsp_diff|dout[31]~q ),
	.dout_32(\differentiate_stages[5].auk_dsp_diff|dout[32]~q ),
	.dout_4(\differentiate_stages[5].auk_dsp_diff|dout[4]~q ),
	.dout_61(\differentiate_stages[4].auk_dsp_diff|dout[6]~q ),
	.dout_3(\differentiate_stages[5].auk_dsp_diff|dout[3]~q ),
	.dout_71(\differentiate_stages[4].auk_dsp_diff|dout[7]~q ),
	.dout_81(\differentiate_stages[4].auk_dsp_diff|dout[8]~q ),
	.dout_91(\differentiate_stages[4].auk_dsp_diff|dout[9]~q ),
	.dout_101(\differentiate_stages[4].auk_dsp_diff|dout[10]~q ),
	.dout_111(\differentiate_stages[4].auk_dsp_diff|dout[11]~q ),
	.dout_121(\differentiate_stages[4].auk_dsp_diff|dout[12]~q ),
	.dout_131(\differentiate_stages[4].auk_dsp_diff|dout[13]~q ),
	.dout_141(\differentiate_stages[4].auk_dsp_diff|dout[14]~q ),
	.dout_151(\differentiate_stages[4].auk_dsp_diff|dout[15]~q ),
	.dout_161(\differentiate_stages[4].auk_dsp_diff|dout[16]~q ),
	.dout_171(\differentiate_stages[4].auk_dsp_diff|dout[17]~q ),
	.dout_181(\differentiate_stages[4].auk_dsp_diff|dout[18]~q ),
	.dout_191(\differentiate_stages[4].auk_dsp_diff|dout[19]~q ),
	.dout_201(\differentiate_stages[4].auk_dsp_diff|dout[20]~q ),
	.dout_211(\differentiate_stages[4].auk_dsp_diff|dout[21]~q ),
	.dout_221(\differentiate_stages[4].auk_dsp_diff|dout[22]~q ),
	.dout_231(\differentiate_stages[4].auk_dsp_diff|dout[23]~q ),
	.dout_241(\differentiate_stages[4].auk_dsp_diff|dout[24]~q ),
	.dout_251(\differentiate_stages[4].auk_dsp_diff|dout[25]~q ),
	.dout_261(\differentiate_stages[4].auk_dsp_diff|dout[26]~q ),
	.dout_271(\differentiate_stages[4].auk_dsp_diff|dout[27]~q ),
	.dout_281(\differentiate_stages[4].auk_dsp_diff|dout[28]~q ),
	.dout_291(\differentiate_stages[4].auk_dsp_diff|dout[29]~q ),
	.dout_301(\differentiate_stages[4].auk_dsp_diff|dout[30]~q ),
	.dout_311(\differentiate_stages[4].auk_dsp_diff|dout[31]~q ),
	.dout_321(\differentiate_stages[4].auk_dsp_diff|dout[32]~q ),
	.dout_33(\differentiate_stages[4].auk_dsp_diff|dout[33]~q ),
	.dout_51(\differentiate_stages[4].auk_dsp_diff|dout[5]~q ),
	.dout_2(\differentiate_stages[5].auk_dsp_diff|dout[2]~q ),
	.dout_41(\differentiate_stages[4].auk_dsp_diff|dout[4]~q ),
	.dout_1(\differentiate_stages[5].auk_dsp_diff|dout[1]~q ),
	.dout_34(\differentiate_stages[4].auk_dsp_diff|dout[3]~q ),
	.dout_210(\differentiate_stages[4].auk_dsp_diff|dout[2]~q ),
	.dout_110(\differentiate_stages[4].auk_dsp_diff|dout[1]~q ),
	.stall_reg(stall_reg),
	.dout_valid3(\differentiate_stages[7].auk_dsp_diff|dout_valid~0_combout ),
	.clk(clk),
	.reset_n(reset_n));

cic_auk_dspip_differentiator_4 \differentiate_stages[4].auk_dsp_diff (
	.dout_valid1(\differentiate_stages[4].auk_dsp_diff|dout_valid~q ),
	.dout_valid2(\differentiate_stages[3].auk_dsp_diff|dout_valid~q ),
	.dout_6(\differentiate_stages[4].auk_dsp_diff|dout[6]~q ),
	.dout_7(\differentiate_stages[4].auk_dsp_diff|dout[7]~q ),
	.dout_8(\differentiate_stages[4].auk_dsp_diff|dout[8]~q ),
	.dout_9(\differentiate_stages[4].auk_dsp_diff|dout[9]~q ),
	.dout_10(\differentiate_stages[4].auk_dsp_diff|dout[10]~q ),
	.dout_11(\differentiate_stages[4].auk_dsp_diff|dout[11]~q ),
	.dout_12(\differentiate_stages[4].auk_dsp_diff|dout[12]~q ),
	.dout_13(\differentiate_stages[4].auk_dsp_diff|dout[13]~q ),
	.dout_14(\differentiate_stages[4].auk_dsp_diff|dout[14]~q ),
	.dout_15(\differentiate_stages[4].auk_dsp_diff|dout[15]~q ),
	.dout_16(\differentiate_stages[4].auk_dsp_diff|dout[16]~q ),
	.dout_17(\differentiate_stages[4].auk_dsp_diff|dout[17]~q ),
	.dout_18(\differentiate_stages[4].auk_dsp_diff|dout[18]~q ),
	.dout_19(\differentiate_stages[4].auk_dsp_diff|dout[19]~q ),
	.dout_20(\differentiate_stages[4].auk_dsp_diff|dout[20]~q ),
	.dout_21(\differentiate_stages[4].auk_dsp_diff|dout[21]~q ),
	.dout_22(\differentiate_stages[4].auk_dsp_diff|dout[22]~q ),
	.dout_23(\differentiate_stages[4].auk_dsp_diff|dout[23]~q ),
	.dout_24(\differentiate_stages[4].auk_dsp_diff|dout[24]~q ),
	.dout_25(\differentiate_stages[4].auk_dsp_diff|dout[25]~q ),
	.dout_26(\differentiate_stages[4].auk_dsp_diff|dout[26]~q ),
	.dout_27(\differentiate_stages[4].auk_dsp_diff|dout[27]~q ),
	.dout_28(\differentiate_stages[4].auk_dsp_diff|dout[28]~q ),
	.dout_29(\differentiate_stages[4].auk_dsp_diff|dout[29]~q ),
	.dout_30(\differentiate_stages[4].auk_dsp_diff|dout[30]~q ),
	.dout_31(\differentiate_stages[4].auk_dsp_diff|dout[31]~q ),
	.dout_32(\differentiate_stages[4].auk_dsp_diff|dout[32]~q ),
	.dout_33(\differentiate_stages[4].auk_dsp_diff|dout[33]~q ),
	.dout_5(\differentiate_stages[4].auk_dsp_diff|dout[5]~q ),
	.dout_61(\differentiate_stages[3].auk_dsp_diff|dout[6]~q ),
	.dout_4(\differentiate_stages[4].auk_dsp_diff|dout[4]~q ),
	.dout_71(\differentiate_stages[3].auk_dsp_diff|dout[7]~q ),
	.dout_81(\differentiate_stages[3].auk_dsp_diff|dout[8]~q ),
	.dout_91(\differentiate_stages[3].auk_dsp_diff|dout[9]~q ),
	.dout_101(\differentiate_stages[3].auk_dsp_diff|dout[10]~q ),
	.dout_111(\differentiate_stages[3].auk_dsp_diff|dout[11]~q ),
	.dout_121(\differentiate_stages[3].auk_dsp_diff|dout[12]~q ),
	.dout_131(\differentiate_stages[3].auk_dsp_diff|dout[13]~q ),
	.dout_141(\differentiate_stages[3].auk_dsp_diff|dout[14]~q ),
	.dout_151(\differentiate_stages[3].auk_dsp_diff|dout[15]~q ),
	.dout_161(\differentiate_stages[3].auk_dsp_diff|dout[16]~q ),
	.dout_171(\differentiate_stages[3].auk_dsp_diff|dout[17]~q ),
	.dout_181(\differentiate_stages[3].auk_dsp_diff|dout[18]~q ),
	.dout_191(\differentiate_stages[3].auk_dsp_diff|dout[19]~q ),
	.dout_201(\differentiate_stages[3].auk_dsp_diff|dout[20]~q ),
	.dout_211(\differentiate_stages[3].auk_dsp_diff|dout[21]~q ),
	.dout_221(\differentiate_stages[3].auk_dsp_diff|dout[22]~q ),
	.dout_231(\differentiate_stages[3].auk_dsp_diff|dout[23]~q ),
	.dout_241(\differentiate_stages[3].auk_dsp_diff|dout[24]~q ),
	.dout_251(\differentiate_stages[3].auk_dsp_diff|dout[25]~q ),
	.dout_261(\differentiate_stages[3].auk_dsp_diff|dout[26]~q ),
	.dout_271(\differentiate_stages[3].auk_dsp_diff|dout[27]~q ),
	.dout_281(\differentiate_stages[3].auk_dsp_diff|dout[28]~q ),
	.dout_291(\differentiate_stages[3].auk_dsp_diff|dout[29]~q ),
	.dout_301(\differentiate_stages[3].auk_dsp_diff|dout[30]~q ),
	.dout_311(\differentiate_stages[3].auk_dsp_diff|dout[31]~q ),
	.dout_321(\differentiate_stages[3].auk_dsp_diff|dout[32]~q ),
	.dout_331(\differentiate_stages[3].auk_dsp_diff|dout[33]~q ),
	.dout_51(\differentiate_stages[3].auk_dsp_diff|dout[5]~q ),
	.dout_3(\differentiate_stages[4].auk_dsp_diff|dout[3]~q ),
	.dout_41(\differentiate_stages[3].auk_dsp_diff|dout[4]~q ),
	.dout_2(\differentiate_stages[4].auk_dsp_diff|dout[2]~q ),
	.dout_34(\differentiate_stages[3].auk_dsp_diff|dout[3]~q ),
	.dout_1(\differentiate_stages[4].auk_dsp_diff|dout[1]~q ),
	.dout_210(\differentiate_stages[3].auk_dsp_diff|dout[2]~q ),
	.dout_110(\differentiate_stages[3].auk_dsp_diff|dout[1]~q ),
	.dout_0(\differentiate_stages[3].auk_dsp_diff|dout[0]~q ),
	.stall_reg(stall_reg),
	.dout_valid3(\differentiate_stages[7].auk_dsp_diff|dout_valid~0_combout ),
	.clk(clk),
	.reset_n(reset_n));

cic_auk_dspip_differentiator_3 \differentiate_stages[3].auk_dsp_diff (
	.dout_valid1(\differentiate_stages[3].auk_dsp_diff|dout_valid~q ),
	.dout_valid2(\differentiate_stages[2].auk_dsp_diff|dout_valid~q ),
	.dout_6(\differentiate_stages[3].auk_dsp_diff|dout[6]~q ),
	.dout_7(\differentiate_stages[3].auk_dsp_diff|dout[7]~q ),
	.dout_8(\differentiate_stages[3].auk_dsp_diff|dout[8]~q ),
	.dout_9(\differentiate_stages[3].auk_dsp_diff|dout[9]~q ),
	.dout_10(\differentiate_stages[3].auk_dsp_diff|dout[10]~q ),
	.dout_11(\differentiate_stages[3].auk_dsp_diff|dout[11]~q ),
	.dout_12(\differentiate_stages[3].auk_dsp_diff|dout[12]~q ),
	.dout_13(\differentiate_stages[3].auk_dsp_diff|dout[13]~q ),
	.dout_14(\differentiate_stages[3].auk_dsp_diff|dout[14]~q ),
	.dout_15(\differentiate_stages[3].auk_dsp_diff|dout[15]~q ),
	.dout_16(\differentiate_stages[3].auk_dsp_diff|dout[16]~q ),
	.dout_17(\differentiate_stages[3].auk_dsp_diff|dout[17]~q ),
	.dout_18(\differentiate_stages[3].auk_dsp_diff|dout[18]~q ),
	.dout_19(\differentiate_stages[3].auk_dsp_diff|dout[19]~q ),
	.dout_20(\differentiate_stages[3].auk_dsp_diff|dout[20]~q ),
	.dout_21(\differentiate_stages[3].auk_dsp_diff|dout[21]~q ),
	.dout_22(\differentiate_stages[3].auk_dsp_diff|dout[22]~q ),
	.dout_23(\differentiate_stages[3].auk_dsp_diff|dout[23]~q ),
	.dout_24(\differentiate_stages[3].auk_dsp_diff|dout[24]~q ),
	.dout_25(\differentiate_stages[3].auk_dsp_diff|dout[25]~q ),
	.dout_26(\differentiate_stages[3].auk_dsp_diff|dout[26]~q ),
	.dout_27(\differentiate_stages[3].auk_dsp_diff|dout[27]~q ),
	.dout_28(\differentiate_stages[3].auk_dsp_diff|dout[28]~q ),
	.dout_29(\differentiate_stages[3].auk_dsp_diff|dout[29]~q ),
	.dout_30(\differentiate_stages[3].auk_dsp_diff|dout[30]~q ),
	.dout_31(\differentiate_stages[3].auk_dsp_diff|dout[31]~q ),
	.dout_32(\differentiate_stages[3].auk_dsp_diff|dout[32]~q ),
	.dout_33(\differentiate_stages[3].auk_dsp_diff|dout[33]~q ),
	.dout_5(\differentiate_stages[3].auk_dsp_diff|dout[5]~q ),
	.dout_71(\differentiate_stages[2].auk_dsp_diff|dout[7]~q ),
	.dout_4(\differentiate_stages[3].auk_dsp_diff|dout[4]~q ),
	.dout_81(\differentiate_stages[2].auk_dsp_diff|dout[8]~q ),
	.dout_91(\differentiate_stages[2].auk_dsp_diff|dout[9]~q ),
	.dout_101(\differentiate_stages[2].auk_dsp_diff|dout[10]~q ),
	.dout_111(\differentiate_stages[2].auk_dsp_diff|dout[11]~q ),
	.dout_121(\differentiate_stages[2].auk_dsp_diff|dout[12]~q ),
	.dout_131(\differentiate_stages[2].auk_dsp_diff|dout[13]~q ),
	.dout_141(\differentiate_stages[2].auk_dsp_diff|dout[14]~q ),
	.dout_151(\differentiate_stages[2].auk_dsp_diff|dout[15]~q ),
	.dout_161(\differentiate_stages[2].auk_dsp_diff|dout[16]~q ),
	.dout_171(\differentiate_stages[2].auk_dsp_diff|dout[17]~q ),
	.dout_181(\differentiate_stages[2].auk_dsp_diff|dout[18]~q ),
	.dout_191(\differentiate_stages[2].auk_dsp_diff|dout[19]~q ),
	.dout_201(\differentiate_stages[2].auk_dsp_diff|dout[20]~q ),
	.dout_211(\differentiate_stages[2].auk_dsp_diff|dout[21]~q ),
	.dout_221(\differentiate_stages[2].auk_dsp_diff|dout[22]~q ),
	.dout_231(\differentiate_stages[2].auk_dsp_diff|dout[23]~q ),
	.dout_241(\differentiate_stages[2].auk_dsp_diff|dout[24]~q ),
	.dout_251(\differentiate_stages[2].auk_dsp_diff|dout[25]~q ),
	.dout_261(\differentiate_stages[2].auk_dsp_diff|dout[26]~q ),
	.dout_271(\differentiate_stages[2].auk_dsp_diff|dout[27]~q ),
	.dout_281(\differentiate_stages[2].auk_dsp_diff|dout[28]~q ),
	.dout_291(\differentiate_stages[2].auk_dsp_diff|dout[29]~q ),
	.dout_301(\differentiate_stages[2].auk_dsp_diff|dout[30]~q ),
	.dout_311(\differentiate_stages[2].auk_dsp_diff|dout[31]~q ),
	.dout_321(\differentiate_stages[2].auk_dsp_diff|dout[32]~q ),
	.dout_331(\differentiate_stages[2].auk_dsp_diff|dout[33]~q ),
	.dout_34(\differentiate_stages[2].auk_dsp_diff|dout[34]~q ),
	.dout_61(\differentiate_stages[2].auk_dsp_diff|dout[6]~q ),
	.dout_3(\differentiate_stages[3].auk_dsp_diff|dout[3]~q ),
	.dout_51(\differentiate_stages[2].auk_dsp_diff|dout[5]~q ),
	.dout_2(\differentiate_stages[3].auk_dsp_diff|dout[2]~q ),
	.dout_41(\differentiate_stages[2].auk_dsp_diff|dout[4]~q ),
	.dout_1(\differentiate_stages[3].auk_dsp_diff|dout[1]~q ),
	.dout_35(\differentiate_stages[2].auk_dsp_diff|dout[3]~q ),
	.dout_0(\differentiate_stages[3].auk_dsp_diff|dout[0]~q ),
	.dout_210(\differentiate_stages[2].auk_dsp_diff|dout[2]~q ),
	.dout_110(\differentiate_stages[2].auk_dsp_diff|dout[1]~q ),
	.stall_reg(stall_reg),
	.dout_valid3(\differentiate_stages[7].auk_dsp_diff|dout_valid~0_combout ),
	.clk(clk),
	.reset_n(reset_n));

cic_auk_dspip_differentiator_2 \differentiate_stages[2].auk_dsp_diff (
	.dout_valid1(\differentiate_stages[2].auk_dsp_diff|dout_valid~q ),
	.dout_valid2(\differentiate_stages[1].auk_dsp_diff|dout_valid~q ),
	.dout_7(\differentiate_stages[2].auk_dsp_diff|dout[7]~q ),
	.dout_8(\differentiate_stages[2].auk_dsp_diff|dout[8]~q ),
	.dout_9(\differentiate_stages[2].auk_dsp_diff|dout[9]~q ),
	.dout_10(\differentiate_stages[2].auk_dsp_diff|dout[10]~q ),
	.dout_11(\differentiate_stages[2].auk_dsp_diff|dout[11]~q ),
	.dout_12(\differentiate_stages[2].auk_dsp_diff|dout[12]~q ),
	.dout_13(\differentiate_stages[2].auk_dsp_diff|dout[13]~q ),
	.dout_14(\differentiate_stages[2].auk_dsp_diff|dout[14]~q ),
	.dout_15(\differentiate_stages[2].auk_dsp_diff|dout[15]~q ),
	.dout_16(\differentiate_stages[2].auk_dsp_diff|dout[16]~q ),
	.dout_17(\differentiate_stages[2].auk_dsp_diff|dout[17]~q ),
	.dout_18(\differentiate_stages[2].auk_dsp_diff|dout[18]~q ),
	.dout_19(\differentiate_stages[2].auk_dsp_diff|dout[19]~q ),
	.dout_20(\differentiate_stages[2].auk_dsp_diff|dout[20]~q ),
	.dout_21(\differentiate_stages[2].auk_dsp_diff|dout[21]~q ),
	.dout_22(\differentiate_stages[2].auk_dsp_diff|dout[22]~q ),
	.dout_23(\differentiate_stages[2].auk_dsp_diff|dout[23]~q ),
	.dout_24(\differentiate_stages[2].auk_dsp_diff|dout[24]~q ),
	.dout_25(\differentiate_stages[2].auk_dsp_diff|dout[25]~q ),
	.dout_26(\differentiate_stages[2].auk_dsp_diff|dout[26]~q ),
	.dout_27(\differentiate_stages[2].auk_dsp_diff|dout[27]~q ),
	.dout_28(\differentiate_stages[2].auk_dsp_diff|dout[28]~q ),
	.dout_29(\differentiate_stages[2].auk_dsp_diff|dout[29]~q ),
	.dout_30(\differentiate_stages[2].auk_dsp_diff|dout[30]~q ),
	.dout_31(\differentiate_stages[2].auk_dsp_diff|dout[31]~q ),
	.dout_32(\differentiate_stages[2].auk_dsp_diff|dout[32]~q ),
	.dout_33(\differentiate_stages[2].auk_dsp_diff|dout[33]~q ),
	.dout_34(\differentiate_stages[2].auk_dsp_diff|dout[34]~q ),
	.dout_6(\differentiate_stages[2].auk_dsp_diff|dout[6]~q ),
	.dout_81(\differentiate_stages[1].auk_dsp_diff|dout[8]~q ),
	.dout_5(\differentiate_stages[2].auk_dsp_diff|dout[5]~q ),
	.dout_91(\differentiate_stages[1].auk_dsp_diff|dout[9]~q ),
	.dout_101(\differentiate_stages[1].auk_dsp_diff|dout[10]~q ),
	.dout_111(\differentiate_stages[1].auk_dsp_diff|dout[11]~q ),
	.dout_121(\differentiate_stages[1].auk_dsp_diff|dout[12]~q ),
	.dout_131(\differentiate_stages[1].auk_dsp_diff|dout[13]~q ),
	.dout_141(\differentiate_stages[1].auk_dsp_diff|dout[14]~q ),
	.dout_151(\differentiate_stages[1].auk_dsp_diff|dout[15]~q ),
	.dout_161(\differentiate_stages[1].auk_dsp_diff|dout[16]~q ),
	.dout_171(\differentiate_stages[1].auk_dsp_diff|dout[17]~q ),
	.dout_181(\differentiate_stages[1].auk_dsp_diff|dout[18]~q ),
	.dout_191(\differentiate_stages[1].auk_dsp_diff|dout[19]~q ),
	.dout_201(\differentiate_stages[1].auk_dsp_diff|dout[20]~q ),
	.dout_211(\differentiate_stages[1].auk_dsp_diff|dout[21]~q ),
	.dout_221(\differentiate_stages[1].auk_dsp_diff|dout[22]~q ),
	.dout_231(\differentiate_stages[1].auk_dsp_diff|dout[23]~q ),
	.dout_241(\differentiate_stages[1].auk_dsp_diff|dout[24]~q ),
	.dout_251(\differentiate_stages[1].auk_dsp_diff|dout[25]~q ),
	.dout_261(\differentiate_stages[1].auk_dsp_diff|dout[26]~q ),
	.dout_271(\differentiate_stages[1].auk_dsp_diff|dout[27]~q ),
	.dout_281(\differentiate_stages[1].auk_dsp_diff|dout[28]~q ),
	.dout_291(\differentiate_stages[1].auk_dsp_diff|dout[29]~q ),
	.dout_301(\differentiate_stages[1].auk_dsp_diff|dout[30]~q ),
	.dout_311(\differentiate_stages[1].auk_dsp_diff|dout[31]~q ),
	.dout_321(\differentiate_stages[1].auk_dsp_diff|dout[32]~q ),
	.dout_331(\differentiate_stages[1].auk_dsp_diff|dout[33]~q ),
	.dout_341(\differentiate_stages[1].auk_dsp_diff|dout[34]~q ),
	.dout_35(\differentiate_stages[1].auk_dsp_diff|dout[35]~q ),
	.dout_71(\differentiate_stages[1].auk_dsp_diff|dout[7]~q ),
	.dout_4(\differentiate_stages[2].auk_dsp_diff|dout[4]~q ),
	.dout_61(\differentiate_stages[1].auk_dsp_diff|dout[6]~q ),
	.dout_3(\differentiate_stages[2].auk_dsp_diff|dout[3]~q ),
	.dout_51(\differentiate_stages[1].auk_dsp_diff|dout[5]~q ),
	.dout_2(\differentiate_stages[2].auk_dsp_diff|dout[2]~q ),
	.dout_41(\differentiate_stages[1].auk_dsp_diff|dout[4]~q ),
	.dout_1(\differentiate_stages[2].auk_dsp_diff|dout[1]~q ),
	.dout_36(\differentiate_stages[1].auk_dsp_diff|dout[3]~q ),
	.dout_210(\differentiate_stages[1].auk_dsp_diff|dout[2]~q ),
	.dout_110(\differentiate_stages[1].auk_dsp_diff|dout[1]~q ),
	.stall_reg(stall_reg),
	.dout_valid3(\differentiate_stages[7].auk_dsp_diff|dout_valid~0_combout ),
	.clk(clk),
	.reset_n(reset_n));

cic_auk_dspip_differentiator_7 \differentiate_stages[7].auk_dsp_diff (
	.dout_valid1(dout_valid),
	.dout_3(dout_3),
	.dout_4(dout_4),
	.dout_5(dout_5),
	.dout_6(dout_6),
	.dout_7(dout_7),
	.dout_8(dout_8),
	.dout_9(dout_9),
	.dout_10(dout_10),
	.dout_11(dout_11),
	.dout_12(dout_12),
	.dout_13(dout_13),
	.dout_14(dout_14),
	.dout_15(dout_15),
	.dout_16(dout_16),
	.dout_17(dout_17),
	.dout_18(dout_18),
	.dout_19(dout_19),
	.dout_20(dout_20),
	.dout_21(dout_21),
	.dout_22(dout_22),
	.dout_23(dout_23),
	.dout_24(dout_24),
	.dout_25(dout_25),
	.dout_26(dout_26),
	.dout_27(dout_27),
	.dout_28(dout_28),
	.dout_29(dout_29),
	.dout_30(dout_30),
	.dout_valid2(\differentiate_stages[6].auk_dsp_diff|dout_valid~q ),
	.dout_41(\differentiate_stages[6].auk_dsp_diff|dout[4]~q ),
	.dout_51(\differentiate_stages[6].auk_dsp_diff|dout[5]~q ),
	.dout_61(\differentiate_stages[6].auk_dsp_diff|dout[6]~q ),
	.dout_71(\differentiate_stages[6].auk_dsp_diff|dout[7]~q ),
	.dout_81(\differentiate_stages[6].auk_dsp_diff|dout[8]~q ),
	.dout_91(\differentiate_stages[6].auk_dsp_diff|dout[9]~q ),
	.dout_101(\differentiate_stages[6].auk_dsp_diff|dout[10]~q ),
	.dout_111(\differentiate_stages[6].auk_dsp_diff|dout[11]~q ),
	.dout_121(\differentiate_stages[6].auk_dsp_diff|dout[12]~q ),
	.dout_131(\differentiate_stages[6].auk_dsp_diff|dout[13]~q ),
	.dout_141(\differentiate_stages[6].auk_dsp_diff|dout[14]~q ),
	.dout_151(\differentiate_stages[6].auk_dsp_diff|dout[15]~q ),
	.dout_161(\differentiate_stages[6].auk_dsp_diff|dout[16]~q ),
	.dout_171(\differentiate_stages[6].auk_dsp_diff|dout[17]~q ),
	.dout_181(\differentiate_stages[6].auk_dsp_diff|dout[18]~q ),
	.dout_191(\differentiate_stages[6].auk_dsp_diff|dout[19]~q ),
	.dout_201(\differentiate_stages[6].auk_dsp_diff|dout[20]~q ),
	.dout_211(\differentiate_stages[6].auk_dsp_diff|dout[21]~q ),
	.dout_221(\differentiate_stages[6].auk_dsp_diff|dout[22]~q ),
	.dout_231(\differentiate_stages[6].auk_dsp_diff|dout[23]~q ),
	.dout_241(\differentiate_stages[6].auk_dsp_diff|dout[24]~q ),
	.dout_251(\differentiate_stages[6].auk_dsp_diff|dout[25]~q ),
	.dout_261(\differentiate_stages[6].auk_dsp_diff|dout[26]~q ),
	.dout_271(\differentiate_stages[6].auk_dsp_diff|dout[27]~q ),
	.dout_281(\differentiate_stages[6].auk_dsp_diff|dout[28]~q ),
	.dout_291(\differentiate_stages[6].auk_dsp_diff|dout[29]~q ),
	.dout_301(\differentiate_stages[6].auk_dsp_diff|dout[30]~q ),
	.dout_31(\differentiate_stages[6].auk_dsp_diff|dout[31]~q ),
	.dout_32(\differentiate_stages[6].auk_dsp_diff|dout[3]~q ),
	.dout_2(\differentiate_stages[6].auk_dsp_diff|dout[2]~q ),
	.dout_1(\differentiate_stages[6].auk_dsp_diff|dout[1]~q ),
	.stall_reg(stall_reg),
	.dout_valid3(\differentiate_stages[7].auk_dsp_diff|dout_valid~0_combout ),
	.clk(clk),
	.reset_n(reset_n));

cic_auk_dspip_differentiator_6 \differentiate_stages[6].auk_dsp_diff (
	.dout_valid1(\differentiate_stages[6].auk_dsp_diff|dout_valid~q ),
	.dout_valid2(\differentiate_stages[5].auk_dsp_diff|dout_valid~q ),
	.dout_4(\differentiate_stages[6].auk_dsp_diff|dout[4]~q ),
	.dout_5(\differentiate_stages[6].auk_dsp_diff|dout[5]~q ),
	.dout_6(\differentiate_stages[6].auk_dsp_diff|dout[6]~q ),
	.dout_7(\differentiate_stages[6].auk_dsp_diff|dout[7]~q ),
	.dout_8(\differentiate_stages[6].auk_dsp_diff|dout[8]~q ),
	.dout_9(\differentiate_stages[6].auk_dsp_diff|dout[9]~q ),
	.dout_10(\differentiate_stages[6].auk_dsp_diff|dout[10]~q ),
	.dout_11(\differentiate_stages[6].auk_dsp_diff|dout[11]~q ),
	.dout_12(\differentiate_stages[6].auk_dsp_diff|dout[12]~q ),
	.dout_13(\differentiate_stages[6].auk_dsp_diff|dout[13]~q ),
	.dout_14(\differentiate_stages[6].auk_dsp_diff|dout[14]~q ),
	.dout_15(\differentiate_stages[6].auk_dsp_diff|dout[15]~q ),
	.dout_16(\differentiate_stages[6].auk_dsp_diff|dout[16]~q ),
	.dout_17(\differentiate_stages[6].auk_dsp_diff|dout[17]~q ),
	.dout_18(\differentiate_stages[6].auk_dsp_diff|dout[18]~q ),
	.dout_19(\differentiate_stages[6].auk_dsp_diff|dout[19]~q ),
	.dout_20(\differentiate_stages[6].auk_dsp_diff|dout[20]~q ),
	.dout_21(\differentiate_stages[6].auk_dsp_diff|dout[21]~q ),
	.dout_22(\differentiate_stages[6].auk_dsp_diff|dout[22]~q ),
	.dout_23(\differentiate_stages[6].auk_dsp_diff|dout[23]~q ),
	.dout_24(\differentiate_stages[6].auk_dsp_diff|dout[24]~q ),
	.dout_25(\differentiate_stages[6].auk_dsp_diff|dout[25]~q ),
	.dout_26(\differentiate_stages[6].auk_dsp_diff|dout[26]~q ),
	.dout_27(\differentiate_stages[6].auk_dsp_diff|dout[27]~q ),
	.dout_28(\differentiate_stages[6].auk_dsp_diff|dout[28]~q ),
	.dout_29(\differentiate_stages[6].auk_dsp_diff|dout[29]~q ),
	.dout_30(\differentiate_stages[6].auk_dsp_diff|dout[30]~q ),
	.dout_31(\differentiate_stages[6].auk_dsp_diff|dout[31]~q ),
	.dout_3(\differentiate_stages[6].auk_dsp_diff|dout[3]~q ),
	.dout_51(\differentiate_stages[5].auk_dsp_diff|dout[5]~q ),
	.dout_2(\differentiate_stages[6].auk_dsp_diff|dout[2]~q ),
	.dout_61(\differentiate_stages[5].auk_dsp_diff|dout[6]~q ),
	.dout_71(\differentiate_stages[5].auk_dsp_diff|dout[7]~q ),
	.dout_81(\differentiate_stages[5].auk_dsp_diff|dout[8]~q ),
	.dout_91(\differentiate_stages[5].auk_dsp_diff|dout[9]~q ),
	.dout_101(\differentiate_stages[5].auk_dsp_diff|dout[10]~q ),
	.dout_111(\differentiate_stages[5].auk_dsp_diff|dout[11]~q ),
	.dout_121(\differentiate_stages[5].auk_dsp_diff|dout[12]~q ),
	.dout_131(\differentiate_stages[5].auk_dsp_diff|dout[13]~q ),
	.dout_141(\differentiate_stages[5].auk_dsp_diff|dout[14]~q ),
	.dout_151(\differentiate_stages[5].auk_dsp_diff|dout[15]~q ),
	.dout_161(\differentiate_stages[5].auk_dsp_diff|dout[16]~q ),
	.dout_171(\differentiate_stages[5].auk_dsp_diff|dout[17]~q ),
	.dout_181(\differentiate_stages[5].auk_dsp_diff|dout[18]~q ),
	.dout_191(\differentiate_stages[5].auk_dsp_diff|dout[19]~q ),
	.dout_201(\differentiate_stages[5].auk_dsp_diff|dout[20]~q ),
	.dout_211(\differentiate_stages[5].auk_dsp_diff|dout[21]~q ),
	.dout_221(\differentiate_stages[5].auk_dsp_diff|dout[22]~q ),
	.dout_231(\differentiate_stages[5].auk_dsp_diff|dout[23]~q ),
	.dout_241(\differentiate_stages[5].auk_dsp_diff|dout[24]~q ),
	.dout_251(\differentiate_stages[5].auk_dsp_diff|dout[25]~q ),
	.dout_261(\differentiate_stages[5].auk_dsp_diff|dout[26]~q ),
	.dout_271(\differentiate_stages[5].auk_dsp_diff|dout[27]~q ),
	.dout_281(\differentiate_stages[5].auk_dsp_diff|dout[28]~q ),
	.dout_291(\differentiate_stages[5].auk_dsp_diff|dout[29]~q ),
	.dout_301(\differentiate_stages[5].auk_dsp_diff|dout[30]~q ),
	.dout_311(\differentiate_stages[5].auk_dsp_diff|dout[31]~q ),
	.dout_32(\differentiate_stages[5].auk_dsp_diff|dout[32]~q ),
	.dout_41(\differentiate_stages[5].auk_dsp_diff|dout[4]~q ),
	.dout_1(\differentiate_stages[6].auk_dsp_diff|dout[1]~q ),
	.dout_33(\differentiate_stages[5].auk_dsp_diff|dout[3]~q ),
	.dout_210(\differentiate_stages[5].auk_dsp_diff|dout[2]~q ),
	.dout_110(\differentiate_stages[5].auk_dsp_diff|dout[1]~q ),
	.stall_reg(stall_reg),
	.dout_valid3(\differentiate_stages[7].auk_dsp_diff|dout_valid~0_combout ),
	.clk(clk),
	.reset_n(reset_n));

dffeas \ena_diff_s[0] (
	.clk(clk),
	.d(\ena_diff_s~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(vcc),
	.q(\ena_diff_s[0]~q ),
	.prn(vcc));
defparam \ena_diff_s[0] .is_wysiwyg = "true";
defparam \ena_diff_s[0] .power_up = "low";

dffeas \sample_state[0] (
	.clk(clk),
	.d(\sample_state~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(vcc),
	.q(\sample_state[0]~q ),
	.prn(vcc));
defparam \sample_state[0] .is_wysiwyg = "true";
defparam \sample_state[0] .power_up = "low";

arriav_lcell_comb \sample_state~0 (
	.dataa(!\latency_cnt_inst|count[0]~q ),
	.datab(!\latency_cnt_inst|count[1]~q ),
	.datac(!\latency_cnt_inst|count[2]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sample_state~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sample_state~0 .extended_lut = "off";
defparam \sample_state~0 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \sample_state~0 .shared_arith = "off";

dffeas \ena_diff_s[1] (
	.clk(clk),
	.d(\fifo_regulator|buffer_FIFO|auto_generated|dpfifo|valid_rreq~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\differentiate_stages[7].auk_dsp_diff|dout_valid~0_combout ),
	.q(\ena_diff_s[1]~q ),
	.prn(vcc));
defparam \ena_diff_s[1] .is_wysiwyg = "true";
defparam \ena_diff_s[1] .power_up = "low";

dffeas fifo_rdreq(
	.clk(clk),
	.d(\fifo_rdreq~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\differentiate_stages[7].auk_dsp_diff|dout_valid~0_combout ),
	.q(\fifo_rdreq~q ),
	.prn(vcc));
defparam fifo_rdreq.is_wysiwyg = "true";
defparam fifo_rdreq.power_up = "low";

arriav_lcell_comb \fifo_rdreq~0 (
	.dataa(!stall_reg),
	.datab(!\ena_diff_s[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fifo_rdreq~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fifo_rdreq~0 .extended_lut = "off";
defparam \fifo_rdreq~0 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \fifo_rdreq~0 .shared_arith = "off";

arriav_lcell_comb \ena_diff_s~0 (
	.dataa(!stall_reg),
	.datab(!\ena_diff_s[0]~q ),
	.datac(!\sample_state[0]~q ),
	.datad(!\fifo_regulator|buffer_FIFO|auto_generated|dpfifo|valid_wreq~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ena_diff_s~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ena_diff_s~0 .extended_lut = "off";
defparam \ena_diff_s~0 .lut_mask = 64'h7BFF7BFF7BFF7BFF;
defparam \ena_diff_s~0 .shared_arith = "off";

arriav_lcell_comb \sample_state~1 (
	.dataa(!stall_reg),
	.datab(!\latency_cnt_inst|count[3]~q ),
	.datac(!\latency_cnt_inst|count[4]~q ),
	.datad(!\sample_state~0_combout ),
	.datae(!\sample_state[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sample_state~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sample_state~1 .extended_lut = "off";
defparam \sample_state~1 .lut_mask = 64'hBFFFFFFFBFFFFFFF;
defparam \sample_state~1 .shared_arith = "off";

dffeas \state[0] (
	.clk(clk),
	.d(\state~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(vcc),
	.q(state_0),
	.prn(vcc));
defparam \state[0] .is_wysiwyg = "true";
defparam \state[0] .power_up = "low";

arriav_lcell_comb \state~0 (
	.dataa(!stall_reg),
	.datab(!state_0),
	.datac(!\latency_cnt_inst|count[0]~q ),
	.datad(!\latency_cnt_inst|Equal0~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\state~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \state~0 .extended_lut = "off";
defparam \state~0 .lut_mask = 64'hFBFFFBFFFBFFFBFF;
defparam \state~0 .shared_arith = "off";

endmodule

module cic_auk_dspip_channel_buffer (
	sample_state_0,
	q,
	stall_reg,
	fifo_rdreq,
	valid_rreq,
	count_0,
	count_3,
	count_1,
	count_2,
	valid_wreq,
	data,
	clk,
	clr)/* synthesis synthesis_greybox=1 */;
input 	sample_state_0;
output 	[37:0] q;
input 	stall_reg;
input 	fifo_rdreq;
output 	valid_rreq;
input 	count_0;
input 	count_3;
input 	count_1;
input 	count_2;
output 	valid_wreq;
input 	[37:0] data;
input 	clk;
input 	clr;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cic_scfifo_1 buffer_FIFO(
	.sample_state_0(sample_state_0),
	.q({q[37],q[36],q[35],q[34],q[33],q[32],q[31],q[30],q[29],q[28],q[27],q[26],q[25],q[24],q[23],q[22],q[21],q[20],q[19],q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q[4],q[3],q[2],q[1],q_unconnected_wire_0}),
	.stall_reg(stall_reg),
	.fifo_rdreq(fifo_rdreq),
	.valid_rreq(valid_rreq),
	.count_0(count_0),
	.count_3(count_3),
	.count_1(count_1),
	.count_2(count_2),
	.valid_wreq(valid_wreq),
	.data({data[37],data[36],data[35],data[34],data[33],data[32],data[31],data[30],data[29],data[28],data[27],data[26],data[25],data[24],data[23],data[22],data[21],data[20],data[19],data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],data[4],data[3],data[2],data[1],gnd}),
	.clock(clk),
	.sclr(clr));

endmodule

module cic_scfifo_1 (
	sample_state_0,
	q,
	stall_reg,
	fifo_rdreq,
	valid_rreq,
	count_0,
	count_3,
	count_1,
	count_2,
	valid_wreq,
	data,
	clock,
	sclr)/* synthesis synthesis_greybox=1 */;
input 	sample_state_0;
output 	[37:0] q;
input 	stall_reg;
input 	fifo_rdreq;
output 	valid_rreq;
input 	count_0;
input 	count_3;
input 	count_1;
input 	count_2;
output 	valid_wreq;
input 	[37:0] data;
input 	clock;
input 	sclr;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cic_scfifo_9mb1 auto_generated(
	.sample_state_0(sample_state_0),
	.q({q[37],q[36],q[35],q[34],q[33],q[32],q[31],q[30],q[29],q[28],q[27],q[26],q[25],q[24],q[23],q[22],q[21],q[20],q[19],q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q[4],q[3],q[2],q[1],q_unconnected_wire_0}),
	.stall_reg(stall_reg),
	.fifo_rdreq(fifo_rdreq),
	.valid_rreq(valid_rreq),
	.count_0(count_0),
	.count_3(count_3),
	.count_1(count_1),
	.count_2(count_2),
	.valid_wreq(valid_wreq),
	.data({data[37],data[36],data[35],data[34],data[33],data[32],data[31],data[30],data[29],data[28],data[27],data[26],data[25],data[24],data[23],data[22],data[21],data[20],data[19],data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],data[4],data[3],data[2],data[1],gnd}),
	.clock(clock),
	.sclr(sclr));

endmodule

module cic_scfifo_9mb1 (
	sample_state_0,
	q,
	stall_reg,
	fifo_rdreq,
	valid_rreq,
	count_0,
	count_3,
	count_1,
	count_2,
	valid_wreq,
	data,
	clock,
	sclr)/* synthesis synthesis_greybox=1 */;
input 	sample_state_0;
output 	[37:0] q;
input 	stall_reg;
input 	fifo_rdreq;
output 	valid_rreq;
input 	count_0;
input 	count_3;
input 	count_1;
input 	count_2;
output 	valid_wreq;
input 	[37:0] data;
input 	clock;
input 	sclr;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cic_a_dpfifo_kj41 dpfifo(
	.sample_state_0(sample_state_0),
	.q({q[37],q[36],q[35],q[34],q[33],q[32],q[31],q[30],q[29],q[28],q[27],q[26],q[25],q[24],q[23],q[22],q[21],q[20],q[19],q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q[4],q[3],q[2],q[1],q_unconnected_wire_0}),
	.stall_reg(stall_reg),
	.fifo_rdreq(fifo_rdreq),
	.valid_rreq1(valid_rreq),
	.count_0(count_0),
	.count_3(count_3),
	.count_1(count_1),
	.count_2(count_2),
	.valid_wreq(valid_wreq),
	.data({data[37],data[36],data[35],data[34],data[33],data[32],data[31],data[30],data[29],data[28],data[27],data[26],data[25],data[24],data[23],data[22],data[21],data[20],data[19],data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],data[4],data[3],data[2],data[1],gnd}),
	.clock(clock),
	.sclr(sclr));

endmodule

module cic_a_dpfifo_kj41 (
	sample_state_0,
	q,
	stall_reg,
	fifo_rdreq,
	valid_rreq1,
	count_0,
	count_3,
	count_1,
	count_2,
	valid_wreq,
	data,
	clock,
	sclr)/* synthesis synthesis_greybox=1 */;
input 	sample_state_0;
output 	[37:0] q;
input 	stall_reg;
input 	fifo_rdreq;
output 	valid_rreq1;
input 	count_0;
input 	count_3;
input 	count_1;
input 	count_2;
output 	valid_wreq;
input 	[37:0] data;
input 	clock;
input 	sclr;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \full_dff~q ;
wire \wr_ptr|counter_reg_bit[0]~q ;
wire \wr_ptr|counter_reg_bit[1]~q ;
wire \rd_ptr_msb|counter_reg_bit[0]~q ;
wire \usedw_counter|counter_reg_bit[1]~q ;
wire \usedw_counter|counter_reg_bit[0]~q ;
wire \valid_wreq~1_combout ;
wire \empty_dff~q ;
wire \valid_rreq~combout ;
wire \low_addressa[0]~q ;
wire \rd_ptr_lsb~q ;
wire \ram_read_address[0]~0_combout ;
wire \low_addressa[1]~q ;
wire \ram_read_address[1]~1_combout ;
wire \valid_wreq~2_combout ;
wire \_~0_combout ;
wire \_~1_combout ;
wire \usedw_is_1_dff~q ;
wire \usedw_is_0_dff~q ;
wire \empty_dff~0_combout ;
wire \low_addressa[0]~0_combout ;
wire \rd_ptr_lsb~0_combout ;
wire \rd_ptr_lsb~1_combout ;
wire \low_addressa[1]~1_combout ;
wire \usedw_will_be_1~0_combout ;
wire \empty_dff~1_combout ;


cic_cntr_rr6 usedw_counter(
	.sample_state_0(sample_state_0),
	.full_dff(\full_dff~q ),
	.counter_reg_bit_1(\usedw_counter|counter_reg_bit[1]~q ),
	.counter_reg_bit_0(\usedw_counter|counter_reg_bit[0]~q ),
	.stall_reg(stall_reg),
	.valid_wreq(valid_wreq),
	.valid_wreq1(\valid_wreq~1_combout ),
	.valid_rreq(\valid_rreq~combout ),
	.clock(clock),
	.sclr(sclr));

cic_cntr_era rd_ptr_msb(
	.counter_reg_bit_0(\rd_ptr_msb|counter_reg_bit[0]~q ),
	.stall_reg(stall_reg),
	.fifo_rdreq(fifo_rdreq),
	.empty_dff(\empty_dff~q ),
	.rd_ptr_lsb(\rd_ptr_lsb~q ),
	.clock(clock),
	.sclr(sclr));

cic_altsyncram_17n1 FIFOram(
	.q_b({q[37],q[36],q[35],q[34],q[33],q[32],q[31],q[30],q[29],q[28],q[27],q[26],q[25],q[24],q[23],q[22],q[21],q[20],q[19],q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q[4],q[3],q[2],q[1],q_b_unconnected_wire_0}),
	.address_a({\wr_ptr|counter_reg_bit[1]~q ,\wr_ptr|counter_reg_bit[0]~q }),
	.wren_a(\valid_wreq~1_combout ),
	.clocken1(\valid_rreq~combout ),
	.data_a({data[37],data[36],data[35],data[34],data[33],data[32],data[31],data[30],data[29],data[28],data[27],data[26],data[25],data[24],data[23],data[22],data[21],data[20],data[19],data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],data[4],data[3],data[2],data[1],gnd}),
	.address_b({\ram_read_address[1]~1_combout ,\ram_read_address[0]~0_combout }),
	.clock1(clock),
	.clock0(clock));

cic_cntr_fra wr_ptr(
	.sample_state_0(sample_state_0),
	.full_dff(\full_dff~q ),
	.counter_reg_bit_0(\wr_ptr|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\wr_ptr|counter_reg_bit[1]~q ),
	.stall_reg(stall_reg),
	.valid_wreq(valid_wreq),
	.clock(clock),
	.sclr(sclr));

dffeas full_dff(
	.clk(clock),
	.d(\_~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!sclr),
	.sload(gnd),
	.ena(vcc),
	.q(\full_dff~q ),
	.prn(vcc));
defparam full_dff.is_wysiwyg = "true";
defparam full_dff.power_up = "low";

arriav_lcell_comb \valid_wreq~1 (
	.dataa(!stall_reg),
	.datab(!sample_state_0),
	.datac(!valid_wreq),
	.datad(!\full_dff~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\valid_wreq~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \valid_wreq~1 .extended_lut = "off";
defparam \valid_wreq~1 .lut_mask = 64'hFFBFFFBFFFBFFFBF;
defparam \valid_wreq~1 .shared_arith = "off";

dffeas empty_dff(
	.clk(clock),
	.d(\empty_dff~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\empty_dff~q ),
	.prn(vcc));
defparam empty_dff.is_wysiwyg = "true";
defparam empty_dff.power_up = "low";

arriav_lcell_comb valid_rreq(
	.dataa(!stall_reg),
	.datab(!fifo_rdreq),
	.datac(!\empty_dff~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\valid_rreq~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam valid_rreq.extended_lut = "off";
defparam valid_rreq.lut_mask = 64'hBFBFBFBFBFBFBFBF;
defparam valid_rreq.shared_arith = "off";

dffeas \low_addressa[0] (
	.clk(clock),
	.d(\low_addressa[0]~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[0]~q ),
	.prn(vcc));
defparam \low_addressa[0] .is_wysiwyg = "true";
defparam \low_addressa[0] .power_up = "low";

dffeas rd_ptr_lsb(
	.clk(clock),
	.d(\rd_ptr_lsb~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\rd_ptr_lsb~1_combout ),
	.q(\rd_ptr_lsb~q ),
	.prn(vcc));
defparam rd_ptr_lsb.is_wysiwyg = "true";
defparam rd_ptr_lsb.power_up = "low";

arriav_lcell_comb \ram_read_address[0]~0 (
	.dataa(!stall_reg),
	.datab(!fifo_rdreq),
	.datac(!\empty_dff~q ),
	.datad(!\low_addressa[0]~q ),
	.datae(!\rd_ptr_lsb~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ram_read_address[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ram_read_address[0]~0 .extended_lut = "off";
defparam \ram_read_address[0]~0 .lut_mask = 64'hFFFF96FFFFFF96FF;
defparam \ram_read_address[0]~0 .shared_arith = "off";

dffeas \low_addressa[1] (
	.clk(clock),
	.d(\low_addressa[1]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[1]~q ),
	.prn(vcc));
defparam \low_addressa[1] .is_wysiwyg = "true";
defparam \low_addressa[1] .power_up = "low";

arriav_lcell_comb \ram_read_address[1]~1 (
	.dataa(!stall_reg),
	.datab(!fifo_rdreq),
	.datac(!\empty_dff~q ),
	.datad(!\rd_ptr_msb|counter_reg_bit[0]~q ),
	.datae(!\low_addressa[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ram_read_address[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ram_read_address[1]~1 .extended_lut = "off";
defparam \ram_read_address[1]~1 .lut_mask = 64'h96FFFFFF96FFFFFF;
defparam \ram_read_address[1]~1 .shared_arith = "off";

arriav_lcell_comb \valid_wreq~2 (
	.dataa(!stall_reg),
	.datab(!sample_state_0),
	.datac(!count_0),
	.datad(!count_3),
	.datae(!count_1),
	.dataf(!count_2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\valid_wreq~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \valid_wreq~2 .extended_lut = "off";
defparam \valid_wreq~2 .lut_mask = 64'hFFFFFFFFFFFFFFFB;
defparam \valid_wreq~2 .shared_arith = "off";

arriav_lcell_comb \_~0 (
	.dataa(!\usedw_counter|counter_reg_bit[1]~q ),
	.datab(!\usedw_counter|counter_reg_bit[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\_~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \_~0 .extended_lut = "off";
defparam \_~0 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \_~0 .shared_arith = "off";

arriav_lcell_comb \_~1 (
	.dataa(!\valid_wreq~2_combout ),
	.datab(!\full_dff~q ),
	.datac(!\valid_rreq~combout ),
	.datad(!\_~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\_~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \_~1 .extended_lut = "off";
defparam \_~1 .lut_mask = 64'hF7FFF7FFF7FFF7FF;
defparam \_~1 .shared_arith = "off";

dffeas usedw_is_1_dff(
	.clk(clock),
	.d(\usedw_will_be_1~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\usedw_is_1_dff~q ),
	.prn(vcc));
defparam usedw_is_1_dff.is_wysiwyg = "true";
defparam usedw_is_1_dff.power_up = "low";

dffeas usedw_is_0_dff(
	.clk(clock),
	.d(\empty_dff~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\usedw_is_0_dff~q ),
	.prn(vcc));
defparam usedw_is_0_dff.is_wysiwyg = "true";
defparam usedw_is_0_dff.power_up = "low";

arriav_lcell_comb \empty_dff~0 (
	.dataa(!sclr),
	.datab(!\valid_wreq~1_combout ),
	.datac(!\valid_rreq~combout ),
	.datad(gnd),
	.datae(!\usedw_is_1_dff~q ),
	.dataf(!\usedw_is_0_dff~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\empty_dff~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \empty_dff~0 .extended_lut = "off";
defparam \empty_dff~0 .lut_mask = 64'hDFDFD5D5FFFFFFFF;
defparam \empty_dff~0 .shared_arith = "off";

arriav_lcell_comb \low_addressa[0]~0 (
	.dataa(!sclr),
	.datab(!stall_reg),
	.datac(!fifo_rdreq),
	.datad(!\empty_dff~q ),
	.datae(!\low_addressa[0]~q ),
	.dataf(!\rd_ptr_lsb~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\low_addressa[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \low_addressa[0]~0 .extended_lut = "off";
defparam \low_addressa[0]~0 .lut_mask = 64'hFFFFFFFFD77DFFFF;
defparam \low_addressa[0]~0 .shared_arith = "off";

arriav_lcell_comb \rd_ptr_lsb~0 (
	.dataa(!sclr),
	.datab(!\rd_ptr_lsb~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rd_ptr_lsb~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rd_ptr_lsb~0 .extended_lut = "off";
defparam \rd_ptr_lsb~0 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \rd_ptr_lsb~0 .shared_arith = "off";

arriav_lcell_comb \rd_ptr_lsb~1 (
	.dataa(!sclr),
	.datab(!stall_reg),
	.datac(!fifo_rdreq),
	.datad(!\empty_dff~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rd_ptr_lsb~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rd_ptr_lsb~1 .extended_lut = "off";
defparam \rd_ptr_lsb~1 .lut_mask = 64'hEFFFEFFFEFFFEFFF;
defparam \rd_ptr_lsb~1 .shared_arith = "off";

arriav_lcell_comb \low_addressa[1]~1 (
	.dataa(!sclr),
	.datab(!stall_reg),
	.datac(!fifo_rdreq),
	.datad(!\empty_dff~q ),
	.datae(!\rd_ptr_msb|counter_reg_bit[0]~q ),
	.dataf(!\low_addressa[1]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\low_addressa[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \low_addressa[1]~1 .extended_lut = "off";
defparam \low_addressa[1]~1 .lut_mask = 64'hD77DFFFFFFFFFFFF;
defparam \low_addressa[1]~1 .shared_arith = "off";

arriav_lcell_comb \usedw_will_be_1~0 (
	.dataa(!sclr),
	.datab(!\valid_wreq~1_combout ),
	.datac(!\valid_rreq~combout ),
	.datad(!\_~0_combout ),
	.datae(!\usedw_is_1_dff~q ),
	.dataf(!\usedw_is_0_dff~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\usedw_will_be_1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \usedw_will_be_1~0 .extended_lut = "off";
defparam \usedw_will_be_1~0 .lut_mask = 64'hFFFFFFFF7DFFFFFF;
defparam \usedw_will_be_1~0 .shared_arith = "off";

arriav_lcell_comb \empty_dff~1 (
	.dataa(!sclr),
	.datab(!\valid_wreq~2_combout ),
	.datac(!\full_dff~q ),
	.datad(!\valid_rreq~combout ),
	.datae(!\usedw_is_1_dff~q ),
	.dataf(!\usedw_is_0_dff~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\empty_dff~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \empty_dff~1 .extended_lut = "off";
defparam \empty_dff~1 .lut_mask = 64'hFFFFD77DFFFFFFFF;
defparam \empty_dff~1 .shared_arith = "off";

arriav_lcell_comb \valid_rreq~0 (
	.dataa(!stall_reg),
	.datab(!fifo_rdreq),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(valid_rreq1),
	.sumout(),
	.cout(),
	.shareout());
defparam \valid_rreq~0 .extended_lut = "off";
defparam \valid_rreq~0 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \valid_rreq~0 .shared_arith = "off";

arriav_lcell_comb \valid_wreq~0 (
	.dataa(!count_0),
	.datab(!count_3),
	.datac(!count_1),
	.datad(!count_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(valid_wreq),
	.sumout(),
	.cout(),
	.shareout());
defparam \valid_wreq~0 .extended_lut = "off";
defparam \valid_wreq~0 .lut_mask = 64'hFFFEFFFEFFFEFFFE;
defparam \valid_wreq~0 .shared_arith = "off";

endmodule

module cic_altsyncram_17n1 (
	q_b,
	address_a,
	wren_a,
	clocken1,
	data_a,
	address_b,
	clock1,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[37:0] q_b;
input 	[1:0] address_a;
input 	wren_a;
input 	clocken1;
input 	[37:0] data_a;
input 	[1:0] address_b;
input 	clock1;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a10_PORTBDATAOUT_bus;
wire [143:0] ram_block1a11_PORTBDATAOUT_bus;
wire [143:0] ram_block1a12_PORTBDATAOUT_bus;
wire [143:0] ram_block1a13_PORTBDATAOUT_bus;
wire [143:0] ram_block1a14_PORTBDATAOUT_bus;
wire [143:0] ram_block1a15_PORTBDATAOUT_bus;
wire [143:0] ram_block1a16_PORTBDATAOUT_bus;
wire [143:0] ram_block1a17_PORTBDATAOUT_bus;
wire [143:0] ram_block1a18_PORTBDATAOUT_bus;
wire [143:0] ram_block1a19_PORTBDATAOUT_bus;
wire [143:0] ram_block1a20_PORTBDATAOUT_bus;
wire [143:0] ram_block1a21_PORTBDATAOUT_bus;
wire [143:0] ram_block1a22_PORTBDATAOUT_bus;
wire [143:0] ram_block1a23_PORTBDATAOUT_bus;
wire [143:0] ram_block1a24_PORTBDATAOUT_bus;
wire [143:0] ram_block1a25_PORTBDATAOUT_bus;
wire [143:0] ram_block1a26_PORTBDATAOUT_bus;
wire [143:0] ram_block1a27_PORTBDATAOUT_bus;
wire [143:0] ram_block1a28_PORTBDATAOUT_bus;
wire [143:0] ram_block1a29_PORTBDATAOUT_bus;
wire [143:0] ram_block1a30_PORTBDATAOUT_bus;
wire [143:0] ram_block1a31_PORTBDATAOUT_bus;
wire [143:0] ram_block1a32_PORTBDATAOUT_bus;
wire [143:0] ram_block1a33_PORTBDATAOUT_bus;
wire [143:0] ram_block1a34_PORTBDATAOUT_bus;
wire [143:0] ram_block1a35_PORTBDATAOUT_bus;
wire [143:0] ram_block1a36_PORTBDATAOUT_bus;
wire [143:0] ram_block1a37_PORTBDATAOUT_bus;
wire [143:0] ram_block1a9_PORTBDATAOUT_bus;
wire [143:0] ram_block1a8_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a1_PORTBDATAOUT_bus;

assign q_b[10] = ram_block1a10_PORTBDATAOUT_bus[0];

assign q_b[11] = ram_block1a11_PORTBDATAOUT_bus[0];

assign q_b[12] = ram_block1a12_PORTBDATAOUT_bus[0];

assign q_b[13] = ram_block1a13_PORTBDATAOUT_bus[0];

assign q_b[14] = ram_block1a14_PORTBDATAOUT_bus[0];

assign q_b[15] = ram_block1a15_PORTBDATAOUT_bus[0];

assign q_b[16] = ram_block1a16_PORTBDATAOUT_bus[0];

assign q_b[17] = ram_block1a17_PORTBDATAOUT_bus[0];

assign q_b[18] = ram_block1a18_PORTBDATAOUT_bus[0];

assign q_b[19] = ram_block1a19_PORTBDATAOUT_bus[0];

assign q_b[20] = ram_block1a20_PORTBDATAOUT_bus[0];

assign q_b[21] = ram_block1a21_PORTBDATAOUT_bus[0];

assign q_b[22] = ram_block1a22_PORTBDATAOUT_bus[0];

assign q_b[23] = ram_block1a23_PORTBDATAOUT_bus[0];

assign q_b[24] = ram_block1a24_PORTBDATAOUT_bus[0];

assign q_b[25] = ram_block1a25_PORTBDATAOUT_bus[0];

assign q_b[26] = ram_block1a26_PORTBDATAOUT_bus[0];

assign q_b[27] = ram_block1a27_PORTBDATAOUT_bus[0];

assign q_b[28] = ram_block1a28_PORTBDATAOUT_bus[0];

assign q_b[29] = ram_block1a29_PORTBDATAOUT_bus[0];

assign q_b[30] = ram_block1a30_PORTBDATAOUT_bus[0];

assign q_b[31] = ram_block1a31_PORTBDATAOUT_bus[0];

assign q_b[32] = ram_block1a32_PORTBDATAOUT_bus[0];

assign q_b[33] = ram_block1a33_PORTBDATAOUT_bus[0];

assign q_b[34] = ram_block1a34_PORTBDATAOUT_bus[0];

assign q_b[35] = ram_block1a35_PORTBDATAOUT_bus[0];

assign q_b[36] = ram_block1a36_PORTBDATAOUT_bus[0];

assign q_b[37] = ram_block1a37_PORTBDATAOUT_bus[0];

assign q_b[9] = ram_block1a9_PORTBDATAOUT_bus[0];

assign q_b[8] = ram_block1a8_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

arriav_ram_block ram_block1a10(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a10_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a10.clk1_output_clock_enable = "ena1";
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_siso:dec_one|auk_dspip_channel_buffer:fifo_regulator|scfifo:buffer_FIFO|scfifo_9mb1:auto_generated|a_dpfifo_kj41:dpfifo|altsyncram_17n1:FIFOram|ALTSYNCRAM";
defparam ram_block1a10.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a10.operation_mode = "dual_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 2;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 3;
defparam ram_block1a10.port_a_logical_ram_depth = 4;
defparam ram_block1a10.port_a_logical_ram_width = 38;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a10.port_b_address_clear = "none";
defparam ram_block1a10.port_b_address_clock = "clock1";
defparam ram_block1a10.port_b_address_width = 2;
defparam ram_block1a10.port_b_data_out_clear = "none";
defparam ram_block1a10.port_b_data_out_clock = "clock1";
defparam ram_block1a10.port_b_data_width = 1;
defparam ram_block1a10.port_b_first_address = 0;
defparam ram_block1a10.port_b_first_bit_number = 10;
defparam ram_block1a10.port_b_last_address = 3;
defparam ram_block1a10.port_b_logical_ram_depth = 4;
defparam ram_block1a10.port_b_logical_ram_width = 38;
defparam ram_block1a10.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a10.port_b_read_enable_clock = "clock1";
defparam ram_block1a10.ram_block_type = "auto";

arriav_ram_block ram_block1a11(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a11_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a11.clk1_output_clock_enable = "ena1";
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_siso:dec_one|auk_dspip_channel_buffer:fifo_regulator|scfifo:buffer_FIFO|scfifo_9mb1:auto_generated|a_dpfifo_kj41:dpfifo|altsyncram_17n1:FIFOram|ALTSYNCRAM";
defparam ram_block1a11.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a11.operation_mode = "dual_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 2;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 3;
defparam ram_block1a11.port_a_logical_ram_depth = 4;
defparam ram_block1a11.port_a_logical_ram_width = 38;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a11.port_b_address_clear = "none";
defparam ram_block1a11.port_b_address_clock = "clock1";
defparam ram_block1a11.port_b_address_width = 2;
defparam ram_block1a11.port_b_data_out_clear = "none";
defparam ram_block1a11.port_b_data_out_clock = "clock1";
defparam ram_block1a11.port_b_data_width = 1;
defparam ram_block1a11.port_b_first_address = 0;
defparam ram_block1a11.port_b_first_bit_number = 11;
defparam ram_block1a11.port_b_last_address = 3;
defparam ram_block1a11.port_b_logical_ram_depth = 4;
defparam ram_block1a11.port_b_logical_ram_width = 38;
defparam ram_block1a11.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a11.port_b_read_enable_clock = "clock1";
defparam ram_block1a11.ram_block_type = "auto";

arriav_ram_block ram_block1a12(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a12_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a12.clk1_output_clock_enable = "ena1";
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_siso:dec_one|auk_dspip_channel_buffer:fifo_regulator|scfifo:buffer_FIFO|scfifo_9mb1:auto_generated|a_dpfifo_kj41:dpfifo|altsyncram_17n1:FIFOram|ALTSYNCRAM";
defparam ram_block1a12.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a12.operation_mode = "dual_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 2;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 3;
defparam ram_block1a12.port_a_logical_ram_depth = 4;
defparam ram_block1a12.port_a_logical_ram_width = 38;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a12.port_b_address_clear = "none";
defparam ram_block1a12.port_b_address_clock = "clock1";
defparam ram_block1a12.port_b_address_width = 2;
defparam ram_block1a12.port_b_data_out_clear = "none";
defparam ram_block1a12.port_b_data_out_clock = "clock1";
defparam ram_block1a12.port_b_data_width = 1;
defparam ram_block1a12.port_b_first_address = 0;
defparam ram_block1a12.port_b_first_bit_number = 12;
defparam ram_block1a12.port_b_last_address = 3;
defparam ram_block1a12.port_b_logical_ram_depth = 4;
defparam ram_block1a12.port_b_logical_ram_width = 38;
defparam ram_block1a12.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a12.port_b_read_enable_clock = "clock1";
defparam ram_block1a12.ram_block_type = "auto";

arriav_ram_block ram_block1a13(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a13_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a13.clk1_output_clock_enable = "ena1";
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_siso:dec_one|auk_dspip_channel_buffer:fifo_regulator|scfifo:buffer_FIFO|scfifo_9mb1:auto_generated|a_dpfifo_kj41:dpfifo|altsyncram_17n1:FIFOram|ALTSYNCRAM";
defparam ram_block1a13.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a13.operation_mode = "dual_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 2;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 3;
defparam ram_block1a13.port_a_logical_ram_depth = 4;
defparam ram_block1a13.port_a_logical_ram_width = 38;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a13.port_b_address_clear = "none";
defparam ram_block1a13.port_b_address_clock = "clock1";
defparam ram_block1a13.port_b_address_width = 2;
defparam ram_block1a13.port_b_data_out_clear = "none";
defparam ram_block1a13.port_b_data_out_clock = "clock1";
defparam ram_block1a13.port_b_data_width = 1;
defparam ram_block1a13.port_b_first_address = 0;
defparam ram_block1a13.port_b_first_bit_number = 13;
defparam ram_block1a13.port_b_last_address = 3;
defparam ram_block1a13.port_b_logical_ram_depth = 4;
defparam ram_block1a13.port_b_logical_ram_width = 38;
defparam ram_block1a13.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a13.port_b_read_enable_clock = "clock1";
defparam ram_block1a13.ram_block_type = "auto";

arriav_ram_block ram_block1a14(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a14_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a14.clk1_output_clock_enable = "ena1";
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_siso:dec_one|auk_dspip_channel_buffer:fifo_regulator|scfifo:buffer_FIFO|scfifo_9mb1:auto_generated|a_dpfifo_kj41:dpfifo|altsyncram_17n1:FIFOram|ALTSYNCRAM";
defparam ram_block1a14.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a14.operation_mode = "dual_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 2;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 3;
defparam ram_block1a14.port_a_logical_ram_depth = 4;
defparam ram_block1a14.port_a_logical_ram_width = 38;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a14.port_b_address_clear = "none";
defparam ram_block1a14.port_b_address_clock = "clock1";
defparam ram_block1a14.port_b_address_width = 2;
defparam ram_block1a14.port_b_data_out_clear = "none";
defparam ram_block1a14.port_b_data_out_clock = "clock1";
defparam ram_block1a14.port_b_data_width = 1;
defparam ram_block1a14.port_b_first_address = 0;
defparam ram_block1a14.port_b_first_bit_number = 14;
defparam ram_block1a14.port_b_last_address = 3;
defparam ram_block1a14.port_b_logical_ram_depth = 4;
defparam ram_block1a14.port_b_logical_ram_width = 38;
defparam ram_block1a14.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a14.port_b_read_enable_clock = "clock1";
defparam ram_block1a14.ram_block_type = "auto";

arriav_ram_block ram_block1a15(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a15_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a15.clk1_output_clock_enable = "ena1";
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_siso:dec_one|auk_dspip_channel_buffer:fifo_regulator|scfifo:buffer_FIFO|scfifo_9mb1:auto_generated|a_dpfifo_kj41:dpfifo|altsyncram_17n1:FIFOram|ALTSYNCRAM";
defparam ram_block1a15.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a15.operation_mode = "dual_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 2;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 3;
defparam ram_block1a15.port_a_logical_ram_depth = 4;
defparam ram_block1a15.port_a_logical_ram_width = 38;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a15.port_b_address_clear = "none";
defparam ram_block1a15.port_b_address_clock = "clock1";
defparam ram_block1a15.port_b_address_width = 2;
defparam ram_block1a15.port_b_data_out_clear = "none";
defparam ram_block1a15.port_b_data_out_clock = "clock1";
defparam ram_block1a15.port_b_data_width = 1;
defparam ram_block1a15.port_b_first_address = 0;
defparam ram_block1a15.port_b_first_bit_number = 15;
defparam ram_block1a15.port_b_last_address = 3;
defparam ram_block1a15.port_b_logical_ram_depth = 4;
defparam ram_block1a15.port_b_logical_ram_width = 38;
defparam ram_block1a15.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a15.port_b_read_enable_clock = "clock1";
defparam ram_block1a15.ram_block_type = "auto";

arriav_ram_block ram_block1a16(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a16_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a16.clk1_output_clock_enable = "ena1";
defparam ram_block1a16.data_interleave_offset_in_bits = 1;
defparam ram_block1a16.data_interleave_width_in_bits = 1;
defparam ram_block1a16.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_siso:dec_one|auk_dspip_channel_buffer:fifo_regulator|scfifo:buffer_FIFO|scfifo_9mb1:auto_generated|a_dpfifo_kj41:dpfifo|altsyncram_17n1:FIFOram|ALTSYNCRAM";
defparam ram_block1a16.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a16.operation_mode = "dual_port";
defparam ram_block1a16.port_a_address_clear = "none";
defparam ram_block1a16.port_a_address_width = 2;
defparam ram_block1a16.port_a_data_out_clear = "none";
defparam ram_block1a16.port_a_data_out_clock = "none";
defparam ram_block1a16.port_a_data_width = 1;
defparam ram_block1a16.port_a_first_address = 0;
defparam ram_block1a16.port_a_first_bit_number = 16;
defparam ram_block1a16.port_a_last_address = 3;
defparam ram_block1a16.port_a_logical_ram_depth = 4;
defparam ram_block1a16.port_a_logical_ram_width = 38;
defparam ram_block1a16.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a16.port_b_address_clear = "none";
defparam ram_block1a16.port_b_address_clock = "clock1";
defparam ram_block1a16.port_b_address_width = 2;
defparam ram_block1a16.port_b_data_out_clear = "none";
defparam ram_block1a16.port_b_data_out_clock = "clock1";
defparam ram_block1a16.port_b_data_width = 1;
defparam ram_block1a16.port_b_first_address = 0;
defparam ram_block1a16.port_b_first_bit_number = 16;
defparam ram_block1a16.port_b_last_address = 3;
defparam ram_block1a16.port_b_logical_ram_depth = 4;
defparam ram_block1a16.port_b_logical_ram_width = 38;
defparam ram_block1a16.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a16.port_b_read_enable_clock = "clock1";
defparam ram_block1a16.ram_block_type = "auto";

arriav_ram_block ram_block1a17(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[17]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a17_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a17.clk1_output_clock_enable = "ena1";
defparam ram_block1a17.data_interleave_offset_in_bits = 1;
defparam ram_block1a17.data_interleave_width_in_bits = 1;
defparam ram_block1a17.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_siso:dec_one|auk_dspip_channel_buffer:fifo_regulator|scfifo:buffer_FIFO|scfifo_9mb1:auto_generated|a_dpfifo_kj41:dpfifo|altsyncram_17n1:FIFOram|ALTSYNCRAM";
defparam ram_block1a17.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a17.operation_mode = "dual_port";
defparam ram_block1a17.port_a_address_clear = "none";
defparam ram_block1a17.port_a_address_width = 2;
defparam ram_block1a17.port_a_data_out_clear = "none";
defparam ram_block1a17.port_a_data_out_clock = "none";
defparam ram_block1a17.port_a_data_width = 1;
defparam ram_block1a17.port_a_first_address = 0;
defparam ram_block1a17.port_a_first_bit_number = 17;
defparam ram_block1a17.port_a_last_address = 3;
defparam ram_block1a17.port_a_logical_ram_depth = 4;
defparam ram_block1a17.port_a_logical_ram_width = 38;
defparam ram_block1a17.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a17.port_b_address_clear = "none";
defparam ram_block1a17.port_b_address_clock = "clock1";
defparam ram_block1a17.port_b_address_width = 2;
defparam ram_block1a17.port_b_data_out_clear = "none";
defparam ram_block1a17.port_b_data_out_clock = "clock1";
defparam ram_block1a17.port_b_data_width = 1;
defparam ram_block1a17.port_b_first_address = 0;
defparam ram_block1a17.port_b_first_bit_number = 17;
defparam ram_block1a17.port_b_last_address = 3;
defparam ram_block1a17.port_b_logical_ram_depth = 4;
defparam ram_block1a17.port_b_logical_ram_width = 38;
defparam ram_block1a17.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a17.port_b_read_enable_clock = "clock1";
defparam ram_block1a17.ram_block_type = "auto";

arriav_ram_block ram_block1a18(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[18]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a18_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a18.clk1_output_clock_enable = "ena1";
defparam ram_block1a18.data_interleave_offset_in_bits = 1;
defparam ram_block1a18.data_interleave_width_in_bits = 1;
defparam ram_block1a18.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_siso:dec_one|auk_dspip_channel_buffer:fifo_regulator|scfifo:buffer_FIFO|scfifo_9mb1:auto_generated|a_dpfifo_kj41:dpfifo|altsyncram_17n1:FIFOram|ALTSYNCRAM";
defparam ram_block1a18.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a18.operation_mode = "dual_port";
defparam ram_block1a18.port_a_address_clear = "none";
defparam ram_block1a18.port_a_address_width = 2;
defparam ram_block1a18.port_a_data_out_clear = "none";
defparam ram_block1a18.port_a_data_out_clock = "none";
defparam ram_block1a18.port_a_data_width = 1;
defparam ram_block1a18.port_a_first_address = 0;
defparam ram_block1a18.port_a_first_bit_number = 18;
defparam ram_block1a18.port_a_last_address = 3;
defparam ram_block1a18.port_a_logical_ram_depth = 4;
defparam ram_block1a18.port_a_logical_ram_width = 38;
defparam ram_block1a18.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a18.port_b_address_clear = "none";
defparam ram_block1a18.port_b_address_clock = "clock1";
defparam ram_block1a18.port_b_address_width = 2;
defparam ram_block1a18.port_b_data_out_clear = "none";
defparam ram_block1a18.port_b_data_out_clock = "clock1";
defparam ram_block1a18.port_b_data_width = 1;
defparam ram_block1a18.port_b_first_address = 0;
defparam ram_block1a18.port_b_first_bit_number = 18;
defparam ram_block1a18.port_b_last_address = 3;
defparam ram_block1a18.port_b_logical_ram_depth = 4;
defparam ram_block1a18.port_b_logical_ram_width = 38;
defparam ram_block1a18.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a18.port_b_read_enable_clock = "clock1";
defparam ram_block1a18.ram_block_type = "auto";

arriav_ram_block ram_block1a19(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[19]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a19_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a19.clk1_output_clock_enable = "ena1";
defparam ram_block1a19.data_interleave_offset_in_bits = 1;
defparam ram_block1a19.data_interleave_width_in_bits = 1;
defparam ram_block1a19.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_siso:dec_one|auk_dspip_channel_buffer:fifo_regulator|scfifo:buffer_FIFO|scfifo_9mb1:auto_generated|a_dpfifo_kj41:dpfifo|altsyncram_17n1:FIFOram|ALTSYNCRAM";
defparam ram_block1a19.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a19.operation_mode = "dual_port";
defparam ram_block1a19.port_a_address_clear = "none";
defparam ram_block1a19.port_a_address_width = 2;
defparam ram_block1a19.port_a_data_out_clear = "none";
defparam ram_block1a19.port_a_data_out_clock = "none";
defparam ram_block1a19.port_a_data_width = 1;
defparam ram_block1a19.port_a_first_address = 0;
defparam ram_block1a19.port_a_first_bit_number = 19;
defparam ram_block1a19.port_a_last_address = 3;
defparam ram_block1a19.port_a_logical_ram_depth = 4;
defparam ram_block1a19.port_a_logical_ram_width = 38;
defparam ram_block1a19.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a19.port_b_address_clear = "none";
defparam ram_block1a19.port_b_address_clock = "clock1";
defparam ram_block1a19.port_b_address_width = 2;
defparam ram_block1a19.port_b_data_out_clear = "none";
defparam ram_block1a19.port_b_data_out_clock = "clock1";
defparam ram_block1a19.port_b_data_width = 1;
defparam ram_block1a19.port_b_first_address = 0;
defparam ram_block1a19.port_b_first_bit_number = 19;
defparam ram_block1a19.port_b_last_address = 3;
defparam ram_block1a19.port_b_logical_ram_depth = 4;
defparam ram_block1a19.port_b_logical_ram_width = 38;
defparam ram_block1a19.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a19.port_b_read_enable_clock = "clock1";
defparam ram_block1a19.ram_block_type = "auto";

arriav_ram_block ram_block1a20(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[20]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a20_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a20.clk1_output_clock_enable = "ena1";
defparam ram_block1a20.data_interleave_offset_in_bits = 1;
defparam ram_block1a20.data_interleave_width_in_bits = 1;
defparam ram_block1a20.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_siso:dec_one|auk_dspip_channel_buffer:fifo_regulator|scfifo:buffer_FIFO|scfifo_9mb1:auto_generated|a_dpfifo_kj41:dpfifo|altsyncram_17n1:FIFOram|ALTSYNCRAM";
defparam ram_block1a20.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a20.operation_mode = "dual_port";
defparam ram_block1a20.port_a_address_clear = "none";
defparam ram_block1a20.port_a_address_width = 2;
defparam ram_block1a20.port_a_data_out_clear = "none";
defparam ram_block1a20.port_a_data_out_clock = "none";
defparam ram_block1a20.port_a_data_width = 1;
defparam ram_block1a20.port_a_first_address = 0;
defparam ram_block1a20.port_a_first_bit_number = 20;
defparam ram_block1a20.port_a_last_address = 3;
defparam ram_block1a20.port_a_logical_ram_depth = 4;
defparam ram_block1a20.port_a_logical_ram_width = 38;
defparam ram_block1a20.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a20.port_b_address_clear = "none";
defparam ram_block1a20.port_b_address_clock = "clock1";
defparam ram_block1a20.port_b_address_width = 2;
defparam ram_block1a20.port_b_data_out_clear = "none";
defparam ram_block1a20.port_b_data_out_clock = "clock1";
defparam ram_block1a20.port_b_data_width = 1;
defparam ram_block1a20.port_b_first_address = 0;
defparam ram_block1a20.port_b_first_bit_number = 20;
defparam ram_block1a20.port_b_last_address = 3;
defparam ram_block1a20.port_b_logical_ram_depth = 4;
defparam ram_block1a20.port_b_logical_ram_width = 38;
defparam ram_block1a20.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a20.port_b_read_enable_clock = "clock1";
defparam ram_block1a20.ram_block_type = "auto";

arriav_ram_block ram_block1a21(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[21]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a21_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a21.clk1_output_clock_enable = "ena1";
defparam ram_block1a21.data_interleave_offset_in_bits = 1;
defparam ram_block1a21.data_interleave_width_in_bits = 1;
defparam ram_block1a21.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_siso:dec_one|auk_dspip_channel_buffer:fifo_regulator|scfifo:buffer_FIFO|scfifo_9mb1:auto_generated|a_dpfifo_kj41:dpfifo|altsyncram_17n1:FIFOram|ALTSYNCRAM";
defparam ram_block1a21.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a21.operation_mode = "dual_port";
defparam ram_block1a21.port_a_address_clear = "none";
defparam ram_block1a21.port_a_address_width = 2;
defparam ram_block1a21.port_a_data_out_clear = "none";
defparam ram_block1a21.port_a_data_out_clock = "none";
defparam ram_block1a21.port_a_data_width = 1;
defparam ram_block1a21.port_a_first_address = 0;
defparam ram_block1a21.port_a_first_bit_number = 21;
defparam ram_block1a21.port_a_last_address = 3;
defparam ram_block1a21.port_a_logical_ram_depth = 4;
defparam ram_block1a21.port_a_logical_ram_width = 38;
defparam ram_block1a21.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a21.port_b_address_clear = "none";
defparam ram_block1a21.port_b_address_clock = "clock1";
defparam ram_block1a21.port_b_address_width = 2;
defparam ram_block1a21.port_b_data_out_clear = "none";
defparam ram_block1a21.port_b_data_out_clock = "clock1";
defparam ram_block1a21.port_b_data_width = 1;
defparam ram_block1a21.port_b_first_address = 0;
defparam ram_block1a21.port_b_first_bit_number = 21;
defparam ram_block1a21.port_b_last_address = 3;
defparam ram_block1a21.port_b_logical_ram_depth = 4;
defparam ram_block1a21.port_b_logical_ram_width = 38;
defparam ram_block1a21.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a21.port_b_read_enable_clock = "clock1";
defparam ram_block1a21.ram_block_type = "auto";

arriav_ram_block ram_block1a22(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[22]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a22_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a22.clk1_output_clock_enable = "ena1";
defparam ram_block1a22.data_interleave_offset_in_bits = 1;
defparam ram_block1a22.data_interleave_width_in_bits = 1;
defparam ram_block1a22.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_siso:dec_one|auk_dspip_channel_buffer:fifo_regulator|scfifo:buffer_FIFO|scfifo_9mb1:auto_generated|a_dpfifo_kj41:dpfifo|altsyncram_17n1:FIFOram|ALTSYNCRAM";
defparam ram_block1a22.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a22.operation_mode = "dual_port";
defparam ram_block1a22.port_a_address_clear = "none";
defparam ram_block1a22.port_a_address_width = 2;
defparam ram_block1a22.port_a_data_out_clear = "none";
defparam ram_block1a22.port_a_data_out_clock = "none";
defparam ram_block1a22.port_a_data_width = 1;
defparam ram_block1a22.port_a_first_address = 0;
defparam ram_block1a22.port_a_first_bit_number = 22;
defparam ram_block1a22.port_a_last_address = 3;
defparam ram_block1a22.port_a_logical_ram_depth = 4;
defparam ram_block1a22.port_a_logical_ram_width = 38;
defparam ram_block1a22.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a22.port_b_address_clear = "none";
defparam ram_block1a22.port_b_address_clock = "clock1";
defparam ram_block1a22.port_b_address_width = 2;
defparam ram_block1a22.port_b_data_out_clear = "none";
defparam ram_block1a22.port_b_data_out_clock = "clock1";
defparam ram_block1a22.port_b_data_width = 1;
defparam ram_block1a22.port_b_first_address = 0;
defparam ram_block1a22.port_b_first_bit_number = 22;
defparam ram_block1a22.port_b_last_address = 3;
defparam ram_block1a22.port_b_logical_ram_depth = 4;
defparam ram_block1a22.port_b_logical_ram_width = 38;
defparam ram_block1a22.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a22.port_b_read_enable_clock = "clock1";
defparam ram_block1a22.ram_block_type = "auto";

arriav_ram_block ram_block1a23(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[23]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a23_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a23.clk1_output_clock_enable = "ena1";
defparam ram_block1a23.data_interleave_offset_in_bits = 1;
defparam ram_block1a23.data_interleave_width_in_bits = 1;
defparam ram_block1a23.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_siso:dec_one|auk_dspip_channel_buffer:fifo_regulator|scfifo:buffer_FIFO|scfifo_9mb1:auto_generated|a_dpfifo_kj41:dpfifo|altsyncram_17n1:FIFOram|ALTSYNCRAM";
defparam ram_block1a23.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a23.operation_mode = "dual_port";
defparam ram_block1a23.port_a_address_clear = "none";
defparam ram_block1a23.port_a_address_width = 2;
defparam ram_block1a23.port_a_data_out_clear = "none";
defparam ram_block1a23.port_a_data_out_clock = "none";
defparam ram_block1a23.port_a_data_width = 1;
defparam ram_block1a23.port_a_first_address = 0;
defparam ram_block1a23.port_a_first_bit_number = 23;
defparam ram_block1a23.port_a_last_address = 3;
defparam ram_block1a23.port_a_logical_ram_depth = 4;
defparam ram_block1a23.port_a_logical_ram_width = 38;
defparam ram_block1a23.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a23.port_b_address_clear = "none";
defparam ram_block1a23.port_b_address_clock = "clock1";
defparam ram_block1a23.port_b_address_width = 2;
defparam ram_block1a23.port_b_data_out_clear = "none";
defparam ram_block1a23.port_b_data_out_clock = "clock1";
defparam ram_block1a23.port_b_data_width = 1;
defparam ram_block1a23.port_b_first_address = 0;
defparam ram_block1a23.port_b_first_bit_number = 23;
defparam ram_block1a23.port_b_last_address = 3;
defparam ram_block1a23.port_b_logical_ram_depth = 4;
defparam ram_block1a23.port_b_logical_ram_width = 38;
defparam ram_block1a23.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a23.port_b_read_enable_clock = "clock1";
defparam ram_block1a23.ram_block_type = "auto";

arriav_ram_block ram_block1a24(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[24]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a24_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a24.clk1_output_clock_enable = "ena1";
defparam ram_block1a24.data_interleave_offset_in_bits = 1;
defparam ram_block1a24.data_interleave_width_in_bits = 1;
defparam ram_block1a24.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_siso:dec_one|auk_dspip_channel_buffer:fifo_regulator|scfifo:buffer_FIFO|scfifo_9mb1:auto_generated|a_dpfifo_kj41:dpfifo|altsyncram_17n1:FIFOram|ALTSYNCRAM";
defparam ram_block1a24.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a24.operation_mode = "dual_port";
defparam ram_block1a24.port_a_address_clear = "none";
defparam ram_block1a24.port_a_address_width = 2;
defparam ram_block1a24.port_a_data_out_clear = "none";
defparam ram_block1a24.port_a_data_out_clock = "none";
defparam ram_block1a24.port_a_data_width = 1;
defparam ram_block1a24.port_a_first_address = 0;
defparam ram_block1a24.port_a_first_bit_number = 24;
defparam ram_block1a24.port_a_last_address = 3;
defparam ram_block1a24.port_a_logical_ram_depth = 4;
defparam ram_block1a24.port_a_logical_ram_width = 38;
defparam ram_block1a24.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a24.port_b_address_clear = "none";
defparam ram_block1a24.port_b_address_clock = "clock1";
defparam ram_block1a24.port_b_address_width = 2;
defparam ram_block1a24.port_b_data_out_clear = "none";
defparam ram_block1a24.port_b_data_out_clock = "clock1";
defparam ram_block1a24.port_b_data_width = 1;
defparam ram_block1a24.port_b_first_address = 0;
defparam ram_block1a24.port_b_first_bit_number = 24;
defparam ram_block1a24.port_b_last_address = 3;
defparam ram_block1a24.port_b_logical_ram_depth = 4;
defparam ram_block1a24.port_b_logical_ram_width = 38;
defparam ram_block1a24.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a24.port_b_read_enable_clock = "clock1";
defparam ram_block1a24.ram_block_type = "auto";

arriav_ram_block ram_block1a25(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[25]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a25_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a25.clk1_output_clock_enable = "ena1";
defparam ram_block1a25.data_interleave_offset_in_bits = 1;
defparam ram_block1a25.data_interleave_width_in_bits = 1;
defparam ram_block1a25.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_siso:dec_one|auk_dspip_channel_buffer:fifo_regulator|scfifo:buffer_FIFO|scfifo_9mb1:auto_generated|a_dpfifo_kj41:dpfifo|altsyncram_17n1:FIFOram|ALTSYNCRAM";
defparam ram_block1a25.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a25.operation_mode = "dual_port";
defparam ram_block1a25.port_a_address_clear = "none";
defparam ram_block1a25.port_a_address_width = 2;
defparam ram_block1a25.port_a_data_out_clear = "none";
defparam ram_block1a25.port_a_data_out_clock = "none";
defparam ram_block1a25.port_a_data_width = 1;
defparam ram_block1a25.port_a_first_address = 0;
defparam ram_block1a25.port_a_first_bit_number = 25;
defparam ram_block1a25.port_a_last_address = 3;
defparam ram_block1a25.port_a_logical_ram_depth = 4;
defparam ram_block1a25.port_a_logical_ram_width = 38;
defparam ram_block1a25.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a25.port_b_address_clear = "none";
defparam ram_block1a25.port_b_address_clock = "clock1";
defparam ram_block1a25.port_b_address_width = 2;
defparam ram_block1a25.port_b_data_out_clear = "none";
defparam ram_block1a25.port_b_data_out_clock = "clock1";
defparam ram_block1a25.port_b_data_width = 1;
defparam ram_block1a25.port_b_first_address = 0;
defparam ram_block1a25.port_b_first_bit_number = 25;
defparam ram_block1a25.port_b_last_address = 3;
defparam ram_block1a25.port_b_logical_ram_depth = 4;
defparam ram_block1a25.port_b_logical_ram_width = 38;
defparam ram_block1a25.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a25.port_b_read_enable_clock = "clock1";
defparam ram_block1a25.ram_block_type = "auto";

arriav_ram_block ram_block1a26(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[26]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a26_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a26.clk1_output_clock_enable = "ena1";
defparam ram_block1a26.data_interleave_offset_in_bits = 1;
defparam ram_block1a26.data_interleave_width_in_bits = 1;
defparam ram_block1a26.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_siso:dec_one|auk_dspip_channel_buffer:fifo_regulator|scfifo:buffer_FIFO|scfifo_9mb1:auto_generated|a_dpfifo_kj41:dpfifo|altsyncram_17n1:FIFOram|ALTSYNCRAM";
defparam ram_block1a26.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a26.operation_mode = "dual_port";
defparam ram_block1a26.port_a_address_clear = "none";
defparam ram_block1a26.port_a_address_width = 2;
defparam ram_block1a26.port_a_data_out_clear = "none";
defparam ram_block1a26.port_a_data_out_clock = "none";
defparam ram_block1a26.port_a_data_width = 1;
defparam ram_block1a26.port_a_first_address = 0;
defparam ram_block1a26.port_a_first_bit_number = 26;
defparam ram_block1a26.port_a_last_address = 3;
defparam ram_block1a26.port_a_logical_ram_depth = 4;
defparam ram_block1a26.port_a_logical_ram_width = 38;
defparam ram_block1a26.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a26.port_b_address_clear = "none";
defparam ram_block1a26.port_b_address_clock = "clock1";
defparam ram_block1a26.port_b_address_width = 2;
defparam ram_block1a26.port_b_data_out_clear = "none";
defparam ram_block1a26.port_b_data_out_clock = "clock1";
defparam ram_block1a26.port_b_data_width = 1;
defparam ram_block1a26.port_b_first_address = 0;
defparam ram_block1a26.port_b_first_bit_number = 26;
defparam ram_block1a26.port_b_last_address = 3;
defparam ram_block1a26.port_b_logical_ram_depth = 4;
defparam ram_block1a26.port_b_logical_ram_width = 38;
defparam ram_block1a26.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a26.port_b_read_enable_clock = "clock1";
defparam ram_block1a26.ram_block_type = "auto";

arriav_ram_block ram_block1a27(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[27]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a27_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a27.clk1_output_clock_enable = "ena1";
defparam ram_block1a27.data_interleave_offset_in_bits = 1;
defparam ram_block1a27.data_interleave_width_in_bits = 1;
defparam ram_block1a27.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_siso:dec_one|auk_dspip_channel_buffer:fifo_regulator|scfifo:buffer_FIFO|scfifo_9mb1:auto_generated|a_dpfifo_kj41:dpfifo|altsyncram_17n1:FIFOram|ALTSYNCRAM";
defparam ram_block1a27.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a27.operation_mode = "dual_port";
defparam ram_block1a27.port_a_address_clear = "none";
defparam ram_block1a27.port_a_address_width = 2;
defparam ram_block1a27.port_a_data_out_clear = "none";
defparam ram_block1a27.port_a_data_out_clock = "none";
defparam ram_block1a27.port_a_data_width = 1;
defparam ram_block1a27.port_a_first_address = 0;
defparam ram_block1a27.port_a_first_bit_number = 27;
defparam ram_block1a27.port_a_last_address = 3;
defparam ram_block1a27.port_a_logical_ram_depth = 4;
defparam ram_block1a27.port_a_logical_ram_width = 38;
defparam ram_block1a27.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a27.port_b_address_clear = "none";
defparam ram_block1a27.port_b_address_clock = "clock1";
defparam ram_block1a27.port_b_address_width = 2;
defparam ram_block1a27.port_b_data_out_clear = "none";
defparam ram_block1a27.port_b_data_out_clock = "clock1";
defparam ram_block1a27.port_b_data_width = 1;
defparam ram_block1a27.port_b_first_address = 0;
defparam ram_block1a27.port_b_first_bit_number = 27;
defparam ram_block1a27.port_b_last_address = 3;
defparam ram_block1a27.port_b_logical_ram_depth = 4;
defparam ram_block1a27.port_b_logical_ram_width = 38;
defparam ram_block1a27.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a27.port_b_read_enable_clock = "clock1";
defparam ram_block1a27.ram_block_type = "auto";

arriav_ram_block ram_block1a28(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[28]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a28_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a28.clk1_output_clock_enable = "ena1";
defparam ram_block1a28.data_interleave_offset_in_bits = 1;
defparam ram_block1a28.data_interleave_width_in_bits = 1;
defparam ram_block1a28.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_siso:dec_one|auk_dspip_channel_buffer:fifo_regulator|scfifo:buffer_FIFO|scfifo_9mb1:auto_generated|a_dpfifo_kj41:dpfifo|altsyncram_17n1:FIFOram|ALTSYNCRAM";
defparam ram_block1a28.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a28.operation_mode = "dual_port";
defparam ram_block1a28.port_a_address_clear = "none";
defparam ram_block1a28.port_a_address_width = 2;
defparam ram_block1a28.port_a_data_out_clear = "none";
defparam ram_block1a28.port_a_data_out_clock = "none";
defparam ram_block1a28.port_a_data_width = 1;
defparam ram_block1a28.port_a_first_address = 0;
defparam ram_block1a28.port_a_first_bit_number = 28;
defparam ram_block1a28.port_a_last_address = 3;
defparam ram_block1a28.port_a_logical_ram_depth = 4;
defparam ram_block1a28.port_a_logical_ram_width = 38;
defparam ram_block1a28.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a28.port_b_address_clear = "none";
defparam ram_block1a28.port_b_address_clock = "clock1";
defparam ram_block1a28.port_b_address_width = 2;
defparam ram_block1a28.port_b_data_out_clear = "none";
defparam ram_block1a28.port_b_data_out_clock = "clock1";
defparam ram_block1a28.port_b_data_width = 1;
defparam ram_block1a28.port_b_first_address = 0;
defparam ram_block1a28.port_b_first_bit_number = 28;
defparam ram_block1a28.port_b_last_address = 3;
defparam ram_block1a28.port_b_logical_ram_depth = 4;
defparam ram_block1a28.port_b_logical_ram_width = 38;
defparam ram_block1a28.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a28.port_b_read_enable_clock = "clock1";
defparam ram_block1a28.ram_block_type = "auto";

arriav_ram_block ram_block1a29(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[29]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a29_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a29.clk1_output_clock_enable = "ena1";
defparam ram_block1a29.data_interleave_offset_in_bits = 1;
defparam ram_block1a29.data_interleave_width_in_bits = 1;
defparam ram_block1a29.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_siso:dec_one|auk_dspip_channel_buffer:fifo_regulator|scfifo:buffer_FIFO|scfifo_9mb1:auto_generated|a_dpfifo_kj41:dpfifo|altsyncram_17n1:FIFOram|ALTSYNCRAM";
defparam ram_block1a29.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a29.operation_mode = "dual_port";
defparam ram_block1a29.port_a_address_clear = "none";
defparam ram_block1a29.port_a_address_width = 2;
defparam ram_block1a29.port_a_data_out_clear = "none";
defparam ram_block1a29.port_a_data_out_clock = "none";
defparam ram_block1a29.port_a_data_width = 1;
defparam ram_block1a29.port_a_first_address = 0;
defparam ram_block1a29.port_a_first_bit_number = 29;
defparam ram_block1a29.port_a_last_address = 3;
defparam ram_block1a29.port_a_logical_ram_depth = 4;
defparam ram_block1a29.port_a_logical_ram_width = 38;
defparam ram_block1a29.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a29.port_b_address_clear = "none";
defparam ram_block1a29.port_b_address_clock = "clock1";
defparam ram_block1a29.port_b_address_width = 2;
defparam ram_block1a29.port_b_data_out_clear = "none";
defparam ram_block1a29.port_b_data_out_clock = "clock1";
defparam ram_block1a29.port_b_data_width = 1;
defparam ram_block1a29.port_b_first_address = 0;
defparam ram_block1a29.port_b_first_bit_number = 29;
defparam ram_block1a29.port_b_last_address = 3;
defparam ram_block1a29.port_b_logical_ram_depth = 4;
defparam ram_block1a29.port_b_logical_ram_width = 38;
defparam ram_block1a29.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a29.port_b_read_enable_clock = "clock1";
defparam ram_block1a29.ram_block_type = "auto";

arriav_ram_block ram_block1a30(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[30]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a30_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a30.clk1_output_clock_enable = "ena1";
defparam ram_block1a30.data_interleave_offset_in_bits = 1;
defparam ram_block1a30.data_interleave_width_in_bits = 1;
defparam ram_block1a30.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_siso:dec_one|auk_dspip_channel_buffer:fifo_regulator|scfifo:buffer_FIFO|scfifo_9mb1:auto_generated|a_dpfifo_kj41:dpfifo|altsyncram_17n1:FIFOram|ALTSYNCRAM";
defparam ram_block1a30.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a30.operation_mode = "dual_port";
defparam ram_block1a30.port_a_address_clear = "none";
defparam ram_block1a30.port_a_address_width = 2;
defparam ram_block1a30.port_a_data_out_clear = "none";
defparam ram_block1a30.port_a_data_out_clock = "none";
defparam ram_block1a30.port_a_data_width = 1;
defparam ram_block1a30.port_a_first_address = 0;
defparam ram_block1a30.port_a_first_bit_number = 30;
defparam ram_block1a30.port_a_last_address = 3;
defparam ram_block1a30.port_a_logical_ram_depth = 4;
defparam ram_block1a30.port_a_logical_ram_width = 38;
defparam ram_block1a30.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a30.port_b_address_clear = "none";
defparam ram_block1a30.port_b_address_clock = "clock1";
defparam ram_block1a30.port_b_address_width = 2;
defparam ram_block1a30.port_b_data_out_clear = "none";
defparam ram_block1a30.port_b_data_out_clock = "clock1";
defparam ram_block1a30.port_b_data_width = 1;
defparam ram_block1a30.port_b_first_address = 0;
defparam ram_block1a30.port_b_first_bit_number = 30;
defparam ram_block1a30.port_b_last_address = 3;
defparam ram_block1a30.port_b_logical_ram_depth = 4;
defparam ram_block1a30.port_b_logical_ram_width = 38;
defparam ram_block1a30.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a30.port_b_read_enable_clock = "clock1";
defparam ram_block1a30.ram_block_type = "auto";

arriav_ram_block ram_block1a31(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[31]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a31_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a31.clk1_output_clock_enable = "ena1";
defparam ram_block1a31.data_interleave_offset_in_bits = 1;
defparam ram_block1a31.data_interleave_width_in_bits = 1;
defparam ram_block1a31.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_siso:dec_one|auk_dspip_channel_buffer:fifo_regulator|scfifo:buffer_FIFO|scfifo_9mb1:auto_generated|a_dpfifo_kj41:dpfifo|altsyncram_17n1:FIFOram|ALTSYNCRAM";
defparam ram_block1a31.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a31.operation_mode = "dual_port";
defparam ram_block1a31.port_a_address_clear = "none";
defparam ram_block1a31.port_a_address_width = 2;
defparam ram_block1a31.port_a_data_out_clear = "none";
defparam ram_block1a31.port_a_data_out_clock = "none";
defparam ram_block1a31.port_a_data_width = 1;
defparam ram_block1a31.port_a_first_address = 0;
defparam ram_block1a31.port_a_first_bit_number = 31;
defparam ram_block1a31.port_a_last_address = 3;
defparam ram_block1a31.port_a_logical_ram_depth = 4;
defparam ram_block1a31.port_a_logical_ram_width = 38;
defparam ram_block1a31.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a31.port_b_address_clear = "none";
defparam ram_block1a31.port_b_address_clock = "clock1";
defparam ram_block1a31.port_b_address_width = 2;
defparam ram_block1a31.port_b_data_out_clear = "none";
defparam ram_block1a31.port_b_data_out_clock = "clock1";
defparam ram_block1a31.port_b_data_width = 1;
defparam ram_block1a31.port_b_first_address = 0;
defparam ram_block1a31.port_b_first_bit_number = 31;
defparam ram_block1a31.port_b_last_address = 3;
defparam ram_block1a31.port_b_logical_ram_depth = 4;
defparam ram_block1a31.port_b_logical_ram_width = 38;
defparam ram_block1a31.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a31.port_b_read_enable_clock = "clock1";
defparam ram_block1a31.ram_block_type = "auto";

arriav_ram_block ram_block1a32(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[32]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a32_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a32.clk1_output_clock_enable = "ena1";
defparam ram_block1a32.data_interleave_offset_in_bits = 1;
defparam ram_block1a32.data_interleave_width_in_bits = 1;
defparam ram_block1a32.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_siso:dec_one|auk_dspip_channel_buffer:fifo_regulator|scfifo:buffer_FIFO|scfifo_9mb1:auto_generated|a_dpfifo_kj41:dpfifo|altsyncram_17n1:FIFOram|ALTSYNCRAM";
defparam ram_block1a32.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a32.operation_mode = "dual_port";
defparam ram_block1a32.port_a_address_clear = "none";
defparam ram_block1a32.port_a_address_width = 2;
defparam ram_block1a32.port_a_data_out_clear = "none";
defparam ram_block1a32.port_a_data_out_clock = "none";
defparam ram_block1a32.port_a_data_width = 1;
defparam ram_block1a32.port_a_first_address = 0;
defparam ram_block1a32.port_a_first_bit_number = 32;
defparam ram_block1a32.port_a_last_address = 3;
defparam ram_block1a32.port_a_logical_ram_depth = 4;
defparam ram_block1a32.port_a_logical_ram_width = 38;
defparam ram_block1a32.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a32.port_b_address_clear = "none";
defparam ram_block1a32.port_b_address_clock = "clock1";
defparam ram_block1a32.port_b_address_width = 2;
defparam ram_block1a32.port_b_data_out_clear = "none";
defparam ram_block1a32.port_b_data_out_clock = "clock1";
defparam ram_block1a32.port_b_data_width = 1;
defparam ram_block1a32.port_b_first_address = 0;
defparam ram_block1a32.port_b_first_bit_number = 32;
defparam ram_block1a32.port_b_last_address = 3;
defparam ram_block1a32.port_b_logical_ram_depth = 4;
defparam ram_block1a32.port_b_logical_ram_width = 38;
defparam ram_block1a32.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a32.port_b_read_enable_clock = "clock1";
defparam ram_block1a32.ram_block_type = "auto";

arriav_ram_block ram_block1a33(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[33]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a33_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a33.clk1_output_clock_enable = "ena1";
defparam ram_block1a33.data_interleave_offset_in_bits = 1;
defparam ram_block1a33.data_interleave_width_in_bits = 1;
defparam ram_block1a33.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_siso:dec_one|auk_dspip_channel_buffer:fifo_regulator|scfifo:buffer_FIFO|scfifo_9mb1:auto_generated|a_dpfifo_kj41:dpfifo|altsyncram_17n1:FIFOram|ALTSYNCRAM";
defparam ram_block1a33.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a33.operation_mode = "dual_port";
defparam ram_block1a33.port_a_address_clear = "none";
defparam ram_block1a33.port_a_address_width = 2;
defparam ram_block1a33.port_a_data_out_clear = "none";
defparam ram_block1a33.port_a_data_out_clock = "none";
defparam ram_block1a33.port_a_data_width = 1;
defparam ram_block1a33.port_a_first_address = 0;
defparam ram_block1a33.port_a_first_bit_number = 33;
defparam ram_block1a33.port_a_last_address = 3;
defparam ram_block1a33.port_a_logical_ram_depth = 4;
defparam ram_block1a33.port_a_logical_ram_width = 38;
defparam ram_block1a33.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a33.port_b_address_clear = "none";
defparam ram_block1a33.port_b_address_clock = "clock1";
defparam ram_block1a33.port_b_address_width = 2;
defparam ram_block1a33.port_b_data_out_clear = "none";
defparam ram_block1a33.port_b_data_out_clock = "clock1";
defparam ram_block1a33.port_b_data_width = 1;
defparam ram_block1a33.port_b_first_address = 0;
defparam ram_block1a33.port_b_first_bit_number = 33;
defparam ram_block1a33.port_b_last_address = 3;
defparam ram_block1a33.port_b_logical_ram_depth = 4;
defparam ram_block1a33.port_b_logical_ram_width = 38;
defparam ram_block1a33.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a33.port_b_read_enable_clock = "clock1";
defparam ram_block1a33.ram_block_type = "auto";

arriav_ram_block ram_block1a34(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[34]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a34_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a34.clk1_output_clock_enable = "ena1";
defparam ram_block1a34.data_interleave_offset_in_bits = 1;
defparam ram_block1a34.data_interleave_width_in_bits = 1;
defparam ram_block1a34.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_siso:dec_one|auk_dspip_channel_buffer:fifo_regulator|scfifo:buffer_FIFO|scfifo_9mb1:auto_generated|a_dpfifo_kj41:dpfifo|altsyncram_17n1:FIFOram|ALTSYNCRAM";
defparam ram_block1a34.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a34.operation_mode = "dual_port";
defparam ram_block1a34.port_a_address_clear = "none";
defparam ram_block1a34.port_a_address_width = 2;
defparam ram_block1a34.port_a_data_out_clear = "none";
defparam ram_block1a34.port_a_data_out_clock = "none";
defparam ram_block1a34.port_a_data_width = 1;
defparam ram_block1a34.port_a_first_address = 0;
defparam ram_block1a34.port_a_first_bit_number = 34;
defparam ram_block1a34.port_a_last_address = 3;
defparam ram_block1a34.port_a_logical_ram_depth = 4;
defparam ram_block1a34.port_a_logical_ram_width = 38;
defparam ram_block1a34.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a34.port_b_address_clear = "none";
defparam ram_block1a34.port_b_address_clock = "clock1";
defparam ram_block1a34.port_b_address_width = 2;
defparam ram_block1a34.port_b_data_out_clear = "none";
defparam ram_block1a34.port_b_data_out_clock = "clock1";
defparam ram_block1a34.port_b_data_width = 1;
defparam ram_block1a34.port_b_first_address = 0;
defparam ram_block1a34.port_b_first_bit_number = 34;
defparam ram_block1a34.port_b_last_address = 3;
defparam ram_block1a34.port_b_logical_ram_depth = 4;
defparam ram_block1a34.port_b_logical_ram_width = 38;
defparam ram_block1a34.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a34.port_b_read_enable_clock = "clock1";
defparam ram_block1a34.ram_block_type = "auto";

arriav_ram_block ram_block1a35(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[35]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a35_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a35.clk1_output_clock_enable = "ena1";
defparam ram_block1a35.data_interleave_offset_in_bits = 1;
defparam ram_block1a35.data_interleave_width_in_bits = 1;
defparam ram_block1a35.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_siso:dec_one|auk_dspip_channel_buffer:fifo_regulator|scfifo:buffer_FIFO|scfifo_9mb1:auto_generated|a_dpfifo_kj41:dpfifo|altsyncram_17n1:FIFOram|ALTSYNCRAM";
defparam ram_block1a35.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a35.operation_mode = "dual_port";
defparam ram_block1a35.port_a_address_clear = "none";
defparam ram_block1a35.port_a_address_width = 2;
defparam ram_block1a35.port_a_data_out_clear = "none";
defparam ram_block1a35.port_a_data_out_clock = "none";
defparam ram_block1a35.port_a_data_width = 1;
defparam ram_block1a35.port_a_first_address = 0;
defparam ram_block1a35.port_a_first_bit_number = 35;
defparam ram_block1a35.port_a_last_address = 3;
defparam ram_block1a35.port_a_logical_ram_depth = 4;
defparam ram_block1a35.port_a_logical_ram_width = 38;
defparam ram_block1a35.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a35.port_b_address_clear = "none";
defparam ram_block1a35.port_b_address_clock = "clock1";
defparam ram_block1a35.port_b_address_width = 2;
defparam ram_block1a35.port_b_data_out_clear = "none";
defparam ram_block1a35.port_b_data_out_clock = "clock1";
defparam ram_block1a35.port_b_data_width = 1;
defparam ram_block1a35.port_b_first_address = 0;
defparam ram_block1a35.port_b_first_bit_number = 35;
defparam ram_block1a35.port_b_last_address = 3;
defparam ram_block1a35.port_b_logical_ram_depth = 4;
defparam ram_block1a35.port_b_logical_ram_width = 38;
defparam ram_block1a35.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a35.port_b_read_enable_clock = "clock1";
defparam ram_block1a35.ram_block_type = "auto";

arriav_ram_block ram_block1a36(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[36]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a36_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a36.clk1_output_clock_enable = "ena1";
defparam ram_block1a36.data_interleave_offset_in_bits = 1;
defparam ram_block1a36.data_interleave_width_in_bits = 1;
defparam ram_block1a36.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_siso:dec_one|auk_dspip_channel_buffer:fifo_regulator|scfifo:buffer_FIFO|scfifo_9mb1:auto_generated|a_dpfifo_kj41:dpfifo|altsyncram_17n1:FIFOram|ALTSYNCRAM";
defparam ram_block1a36.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a36.operation_mode = "dual_port";
defparam ram_block1a36.port_a_address_clear = "none";
defparam ram_block1a36.port_a_address_width = 2;
defparam ram_block1a36.port_a_data_out_clear = "none";
defparam ram_block1a36.port_a_data_out_clock = "none";
defparam ram_block1a36.port_a_data_width = 1;
defparam ram_block1a36.port_a_first_address = 0;
defparam ram_block1a36.port_a_first_bit_number = 36;
defparam ram_block1a36.port_a_last_address = 3;
defparam ram_block1a36.port_a_logical_ram_depth = 4;
defparam ram_block1a36.port_a_logical_ram_width = 38;
defparam ram_block1a36.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a36.port_b_address_clear = "none";
defparam ram_block1a36.port_b_address_clock = "clock1";
defparam ram_block1a36.port_b_address_width = 2;
defparam ram_block1a36.port_b_data_out_clear = "none";
defparam ram_block1a36.port_b_data_out_clock = "clock1";
defparam ram_block1a36.port_b_data_width = 1;
defparam ram_block1a36.port_b_first_address = 0;
defparam ram_block1a36.port_b_first_bit_number = 36;
defparam ram_block1a36.port_b_last_address = 3;
defparam ram_block1a36.port_b_logical_ram_depth = 4;
defparam ram_block1a36.port_b_logical_ram_width = 38;
defparam ram_block1a36.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a36.port_b_read_enable_clock = "clock1";
defparam ram_block1a36.ram_block_type = "auto";

arriav_ram_block ram_block1a37(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[37]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a37_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a37.clk1_output_clock_enable = "ena1";
defparam ram_block1a37.data_interleave_offset_in_bits = 1;
defparam ram_block1a37.data_interleave_width_in_bits = 1;
defparam ram_block1a37.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_siso:dec_one|auk_dspip_channel_buffer:fifo_regulator|scfifo:buffer_FIFO|scfifo_9mb1:auto_generated|a_dpfifo_kj41:dpfifo|altsyncram_17n1:FIFOram|ALTSYNCRAM";
defparam ram_block1a37.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a37.operation_mode = "dual_port";
defparam ram_block1a37.port_a_address_clear = "none";
defparam ram_block1a37.port_a_address_width = 2;
defparam ram_block1a37.port_a_data_out_clear = "none";
defparam ram_block1a37.port_a_data_out_clock = "none";
defparam ram_block1a37.port_a_data_width = 1;
defparam ram_block1a37.port_a_first_address = 0;
defparam ram_block1a37.port_a_first_bit_number = 37;
defparam ram_block1a37.port_a_last_address = 3;
defparam ram_block1a37.port_a_logical_ram_depth = 4;
defparam ram_block1a37.port_a_logical_ram_width = 38;
defparam ram_block1a37.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a37.port_b_address_clear = "none";
defparam ram_block1a37.port_b_address_clock = "clock1";
defparam ram_block1a37.port_b_address_width = 2;
defparam ram_block1a37.port_b_data_out_clear = "none";
defparam ram_block1a37.port_b_data_out_clock = "clock1";
defparam ram_block1a37.port_b_data_width = 1;
defparam ram_block1a37.port_b_first_address = 0;
defparam ram_block1a37.port_b_first_bit_number = 37;
defparam ram_block1a37.port_b_last_address = 3;
defparam ram_block1a37.port_b_logical_ram_depth = 4;
defparam ram_block1a37.port_b_logical_ram_width = 38;
defparam ram_block1a37.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a37.port_b_read_enable_clock = "clock1";
defparam ram_block1a37.ram_block_type = "auto";

arriav_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a9.clk1_output_clock_enable = "ena1";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_siso:dec_one|auk_dspip_channel_buffer:fifo_regulator|scfifo:buffer_FIFO|scfifo_9mb1:auto_generated|a_dpfifo_kj41:dpfifo|altsyncram_17n1:FIFOram|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a9.operation_mode = "dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 2;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 3;
defparam ram_block1a9.port_a_logical_ram_depth = 4;
defparam ram_block1a9.port_a_logical_ram_width = 38;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a9.port_b_address_clear = "none";
defparam ram_block1a9.port_b_address_clock = "clock1";
defparam ram_block1a9.port_b_address_width = 2;
defparam ram_block1a9.port_b_data_out_clear = "none";
defparam ram_block1a9.port_b_data_out_clock = "clock1";
defparam ram_block1a9.port_b_data_width = 1;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 3;
defparam ram_block1a9.port_b_logical_ram_depth = 4;
defparam ram_block1a9.port_b_logical_ram_width = 38;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock1";
defparam ram_block1a9.ram_block_type = "auto";

arriav_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a8.clk1_output_clock_enable = "ena1";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_siso:dec_one|auk_dspip_channel_buffer:fifo_regulator|scfifo:buffer_FIFO|scfifo_9mb1:auto_generated|a_dpfifo_kj41:dpfifo|altsyncram_17n1:FIFOram|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a8.operation_mode = "dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 2;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 3;
defparam ram_block1a8.port_a_logical_ram_depth = 4;
defparam ram_block1a8.port_a_logical_ram_width = 38;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a8.port_b_address_clear = "none";
defparam ram_block1a8.port_b_address_clock = "clock1";
defparam ram_block1a8.port_b_address_width = 2;
defparam ram_block1a8.port_b_data_out_clear = "none";
defparam ram_block1a8.port_b_data_out_clock = "clock1";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 3;
defparam ram_block1a8.port_b_logical_ram_depth = 4;
defparam ram_block1a8.port_b_logical_ram_width = 38;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock1";
defparam ram_block1a8.ram_block_type = "auto";

arriav_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a7.clk1_output_clock_enable = "ena1";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_siso:dec_one|auk_dspip_channel_buffer:fifo_regulator|scfifo:buffer_FIFO|scfifo_9mb1:auto_generated|a_dpfifo_kj41:dpfifo|altsyncram_17n1:FIFOram|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 2;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 3;
defparam ram_block1a7.port_a_logical_ram_depth = 4;
defparam ram_block1a7.port_a_logical_ram_width = 38;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock1";
defparam ram_block1a7.port_b_address_width = 2;
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "clock1";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 3;
defparam ram_block1a7.port_b_logical_ram_depth = 4;
defparam ram_block1a7.port_b_logical_ram_width = 38;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock1";
defparam ram_block1a7.ram_block_type = "auto";

arriav_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a6.clk1_output_clock_enable = "ena1";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_siso:dec_one|auk_dspip_channel_buffer:fifo_regulator|scfifo:buffer_FIFO|scfifo_9mb1:auto_generated|a_dpfifo_kj41:dpfifo|altsyncram_17n1:FIFOram|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 2;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 3;
defparam ram_block1a6.port_a_logical_ram_depth = 4;
defparam ram_block1a6.port_a_logical_ram_width = 38;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock1";
defparam ram_block1a6.port_b_address_width = 2;
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "clock1";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 3;
defparam ram_block1a6.port_b_logical_ram_depth = 4;
defparam ram_block1a6.port_b_logical_ram_width = 38;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock1";
defparam ram_block1a6.ram_block_type = "auto";

arriav_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a5.clk1_output_clock_enable = "ena1";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_siso:dec_one|auk_dspip_channel_buffer:fifo_regulator|scfifo:buffer_FIFO|scfifo_9mb1:auto_generated|a_dpfifo_kj41:dpfifo|altsyncram_17n1:FIFOram|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 2;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 3;
defparam ram_block1a5.port_a_logical_ram_depth = 4;
defparam ram_block1a5.port_a_logical_ram_width = 38;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock1";
defparam ram_block1a5.port_b_address_width = 2;
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "clock1";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 3;
defparam ram_block1a5.port_b_logical_ram_depth = 4;
defparam ram_block1a5.port_b_logical_ram_width = 38;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock1";
defparam ram_block1a5.ram_block_type = "auto";

arriav_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a4.clk1_output_clock_enable = "ena1";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_siso:dec_one|auk_dspip_channel_buffer:fifo_regulator|scfifo:buffer_FIFO|scfifo_9mb1:auto_generated|a_dpfifo_kj41:dpfifo|altsyncram_17n1:FIFOram|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a4.operation_mode = "dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 2;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 3;
defparam ram_block1a4.port_a_logical_ram_depth = 4;
defparam ram_block1a4.port_a_logical_ram_width = 38;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_address_clear = "none";
defparam ram_block1a4.port_b_address_clock = "clock1";
defparam ram_block1a4.port_b_address_width = 2;
defparam ram_block1a4.port_b_data_out_clear = "none";
defparam ram_block1a4.port_b_data_out_clock = "clock1";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 3;
defparam ram_block1a4.port_b_logical_ram_depth = 4;
defparam ram_block1a4.port_b_logical_ram_width = 38;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock1";
defparam ram_block1a4.ram_block_type = "auto";

arriav_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a3.clk1_output_clock_enable = "ena1";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_siso:dec_one|auk_dspip_channel_buffer:fifo_regulator|scfifo:buffer_FIFO|scfifo_9mb1:auto_generated|a_dpfifo_kj41:dpfifo|altsyncram_17n1:FIFOram|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a3.operation_mode = "dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 2;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 3;
defparam ram_block1a3.port_a_logical_ram_depth = 4;
defparam ram_block1a3.port_a_logical_ram_width = 38;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_address_clear = "none";
defparam ram_block1a3.port_b_address_clock = "clock1";
defparam ram_block1a3.port_b_address_width = 2;
defparam ram_block1a3.port_b_data_out_clear = "none";
defparam ram_block1a3.port_b_data_out_clock = "clock1";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 3;
defparam ram_block1a3.port_b_logical_ram_depth = 4;
defparam ram_block1a3.port_b_logical_ram_width = 38;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock1";
defparam ram_block1a3.ram_block_type = "auto";

arriav_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a2.clk1_output_clock_enable = "ena1";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_siso:dec_one|auk_dspip_channel_buffer:fifo_regulator|scfifo:buffer_FIFO|scfifo_9mb1:auto_generated|a_dpfifo_kj41:dpfifo|altsyncram_17n1:FIFOram|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a2.operation_mode = "dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 2;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 3;
defparam ram_block1a2.port_a_logical_ram_depth = 4;
defparam ram_block1a2.port_a_logical_ram_width = 38;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_address_clear = "none";
defparam ram_block1a2.port_b_address_clock = "clock1";
defparam ram_block1a2.port_b_address_width = 2;
defparam ram_block1a2.port_b_data_out_clear = "none";
defparam ram_block1a2.port_b_data_out_clock = "clock1";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 3;
defparam ram_block1a2.port_b_logical_ram_depth = 4;
defparam ram_block1a2.port_b_logical_ram_width = 38;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock1";
defparam ram_block1a2.ram_block_type = "auto";

arriav_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a1.clk1_output_clock_enable = "ena1";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_siso:dec_one|auk_dspip_channel_buffer:fifo_regulator|scfifo:buffer_FIFO|scfifo_9mb1:auto_generated|a_dpfifo_kj41:dpfifo|altsyncram_17n1:FIFOram|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 2;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 3;
defparam ram_block1a1.port_a_logical_ram_depth = 4;
defparam ram_block1a1.port_a_logical_ram_width = 38;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_address_clear = "none";
defparam ram_block1a1.port_b_address_clock = "clock1";
defparam ram_block1a1.port_b_address_width = 2;
defparam ram_block1a1.port_b_data_out_clear = "none";
defparam ram_block1a1.port_b_data_out_clock = "clock1";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 3;
defparam ram_block1a1.port_b_logical_ram_depth = 4;
defparam ram_block1a1.port_b_logical_ram_width = 38;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock1";
defparam ram_block1a1.ram_block_type = "auto";

endmodule

module cic_cntr_era (
	counter_reg_bit_0,
	stall_reg,
	fifo_rdreq,
	empty_dff,
	rd_ptr_lsb,
	clock,
	sclr)/* synthesis synthesis_greybox=1 */;
output 	counter_reg_bit_0;
input 	stall_reg;
input 	fifo_rdreq;
input 	empty_dff;
input 	rd_ptr_lsb;
input 	clock;
input 	sclr;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~COMBOUT ;
wire \_~0_combout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~COMBOUT ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!sclr),
	.sload(gnd),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

arriav_lcell_comb counter_comb_bita0(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\counter_comb_bita0~COMBOUT ),
	.sumout(),
	.cout(),
	.shareout());
defparam counter_comb_bita0.extended_lut = "off";
defparam counter_comb_bita0.lut_mask = 64'hFF00FF00FF00FF00;
defparam counter_comb_bita0.shared_arith = "off";

arriav_lcell_comb \_~0 (
	.dataa(!sclr),
	.datab(!stall_reg),
	.datac(!fifo_rdreq),
	.datad(!empty_dff),
	.datae(!rd_ptr_lsb),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\_~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \_~0 .extended_lut = "off";
defparam \_~0 .lut_mask = 64'hFFFFEFFFFFFFEFFF;
defparam \_~0 .shared_arith = "off";

endmodule

module cic_cntr_fra (
	sample_state_0,
	full_dff,
	counter_reg_bit_0,
	counter_reg_bit_1,
	stall_reg,
	valid_wreq,
	clock,
	sclr)/* synthesis synthesis_greybox=1 */;
input 	sample_state_0;
input 	full_dff;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
input 	stall_reg;
input 	valid_wreq;
input 	clock;
input 	sclr;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~sumout ;
wire \_~0_combout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~sumout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!sclr),
	.sload(gnd),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!sclr),
	.sload(gnd),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

arriav_lcell_comb counter_comb_bita0(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita0~sumout ),
	.cout(\counter_comb_bita0~COUT ),
	.shareout());
defparam counter_comb_bita0.extended_lut = "off";
defparam counter_comb_bita0.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita0.shared_arith = "off";

arriav_lcell_comb \_~0 (
	.dataa(!sclr),
	.datab(!stall_reg),
	.datac(!sample_state_0),
	.datad(!valid_wreq),
	.datae(!full_dff),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\_~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \_~0 .extended_lut = "off";
defparam \_~0 .lut_mask = 64'hFFFFEFFFFFFFEFFF;
defparam \_~0 .shared_arith = "off";

arriav_lcell_comb counter_comb_bita1(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita0~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita1~sumout ),
	.cout(),
	.shareout());
defparam counter_comb_bita1.extended_lut = "off";
defparam counter_comb_bita1.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita1.shared_arith = "off";

endmodule

module cic_cntr_rr6 (
	sample_state_0,
	full_dff,
	counter_reg_bit_1,
	counter_reg_bit_0,
	stall_reg,
	valid_wreq,
	valid_wreq1,
	valid_rreq,
	clock,
	sclr)/* synthesis synthesis_greybox=1 */;
input 	sample_state_0;
input 	full_dff;
output 	counter_reg_bit_1;
output 	counter_reg_bit_0;
input 	stall_reg;
input 	valid_wreq;
input 	valid_wreq1;
input 	valid_rreq;
input 	clock;
input 	sclr;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~sumout ;
wire \_~0_combout ;
wire \counter_comb_bita0~sumout ;


dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!sclr),
	.sload(gnd),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!sclr),
	.sload(gnd),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

arriav_lcell_comb counter_comb_bita0(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita0~sumout ),
	.cout(\counter_comb_bita0~COUT ),
	.shareout());
defparam counter_comb_bita0.extended_lut = "off";
defparam counter_comb_bita0.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita0.shared_arith = "off";

arriav_lcell_comb counter_comb_bita1(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_1),
	.datae(gnd),
	.dataf(!valid_wreq1),
	.datag(gnd),
	.cin(\counter_comb_bita0~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita1~sumout ),
	.cout(),
	.shareout());
defparam counter_comb_bita1.extended_lut = "off";
defparam counter_comb_bita1.lut_mask = 64'h000000FF000000FF;
defparam counter_comb_bita1.shared_arith = "off";

arriav_lcell_comb \_~0 (
	.dataa(!sclr),
	.datab(!stall_reg),
	.datac(!sample_state_0),
	.datad(!valid_wreq),
	.datae(!full_dff),
	.dataf(!valid_rreq),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\_~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \_~0 .extended_lut = "off";
defparam \_~0 .lut_mask = 64'hEBBEBEEBBEEBEBBE;
defparam \_~0 .shared_arith = "off";

endmodule

module cic_auk_dspip_differentiator (
	dout_valid1,
	dout_9,
	dout_10,
	dout_11,
	dout_12,
	dout_13,
	dout_14,
	dout_15,
	dout_16,
	dout_17,
	dout_18,
	dout_19,
	dout_20,
	dout_21,
	dout_22,
	dout_23,
	dout_24,
	dout_25,
	dout_26,
	dout_27,
	dout_28,
	dout_29,
	dout_30,
	dout_31,
	dout_32,
	dout_33,
	dout_34,
	dout_35,
	dout_36,
	dout_8,
	q_b_10,
	dout_7,
	q_b_11,
	q_b_12,
	q_b_13,
	q_b_14,
	q_b_15,
	q_b_16,
	q_b_17,
	q_b_18,
	q_b_19,
	q_b_20,
	q_b_21,
	q_b_22,
	q_b_23,
	q_b_24,
	q_b_25,
	q_b_26,
	q_b_27,
	q_b_28,
	q_b_29,
	q_b_30,
	q_b_31,
	q_b_32,
	q_b_33,
	q_b_34,
	q_b_35,
	q_b_36,
	q_b_37,
	q_b_9,
	dout_6,
	q_b_8,
	dout_5,
	q_b_7,
	dout_4,
	q_b_6,
	dout_3,
	q_b_5,
	dout_2,
	q_b_4,
	dout_1,
	q_b_3,
	q_b_2,
	q_b_1,
	stall_reg,
	dout_valid2,
	ena_diff_s_1,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	dout_valid1;
output 	dout_9;
output 	dout_10;
output 	dout_11;
output 	dout_12;
output 	dout_13;
output 	dout_14;
output 	dout_15;
output 	dout_16;
output 	dout_17;
output 	dout_18;
output 	dout_19;
output 	dout_20;
output 	dout_21;
output 	dout_22;
output 	dout_23;
output 	dout_24;
output 	dout_25;
output 	dout_26;
output 	dout_27;
output 	dout_28;
output 	dout_29;
output 	dout_30;
output 	dout_31;
output 	dout_32;
output 	dout_33;
output 	dout_34;
output 	dout_35;
output 	dout_36;
output 	dout_8;
input 	q_b_10;
output 	dout_7;
input 	q_b_11;
input 	q_b_12;
input 	q_b_13;
input 	q_b_14;
input 	q_b_15;
input 	q_b_16;
input 	q_b_17;
input 	q_b_18;
input 	q_b_19;
input 	q_b_20;
input 	q_b_21;
input 	q_b_22;
input 	q_b_23;
input 	q_b_24;
input 	q_b_25;
input 	q_b_26;
input 	q_b_27;
input 	q_b_28;
input 	q_b_29;
input 	q_b_30;
input 	q_b_31;
input 	q_b_32;
input 	q_b_33;
input 	q_b_34;
input 	q_b_35;
input 	q_b_36;
input 	q_b_37;
input 	q_b_9;
output 	dout_6;
input 	q_b_8;
output 	dout_5;
input 	q_b_7;
output 	dout_4;
input 	q_b_6;
output 	dout_3;
input 	q_b_5;
output 	dout_2;
input 	q_b_4;
output 	dout_1;
input 	q_b_3;
input 	q_b_2;
input 	q_b_1;
input 	stall_reg;
input 	dout_valid2;
input 	ena_diff_s_1;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \glogic:u0|register_fifo:fifo_data[0][9]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][10]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][11]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][12]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][13]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][14]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][15]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][16]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][17]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][18]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][19]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][20]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][21]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][22]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][23]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][24]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][25]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][26]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][27]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][28]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][29]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][30]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][31]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][32]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][33]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][34]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][35]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][36]~q ;
wire \dout~1_combout ;
wire \glogic:u0|register_fifo:fifo_data[0][8]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][7]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][6]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][5]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][4]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][3]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][2]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][1]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][0]~q ;
wire \resq[0]~146_cout ;
wire \resq[0]~147 ;
wire \resq[1]~142 ;
wire \resq[1]~143 ;
wire \resq[2]~138 ;
wire \resq[2]~139 ;
wire \resq[3]~134 ;
wire \resq[3]~135 ;
wire \resq[4]~130 ;
wire \resq[4]~131 ;
wire \resq[5]~126 ;
wire \resq[5]~127 ;
wire \resq[6]~122 ;
wire \resq[6]~123 ;
wire \resq[7]~118 ;
wire \resq[7]~119 ;
wire \resq[8]~114 ;
wire \resq[8]~115 ;
wire \resq[9]~1_sumout ;
wire \dout[36]~0_combout ;
wire \resq[9]~2 ;
wire \resq[9]~3 ;
wire \resq[10]~5_sumout ;
wire \resq[10]~6 ;
wire \resq[10]~7 ;
wire \resq[11]~9_sumout ;
wire \resq[11]~10 ;
wire \resq[11]~11 ;
wire \resq[12]~13_sumout ;
wire \resq[12]~14 ;
wire \resq[12]~15 ;
wire \resq[13]~17_sumout ;
wire \resq[13]~18 ;
wire \resq[13]~19 ;
wire \resq[14]~21_sumout ;
wire \resq[14]~22 ;
wire \resq[14]~23 ;
wire \resq[15]~25_sumout ;
wire \resq[15]~26 ;
wire \resq[15]~27 ;
wire \resq[16]~29_sumout ;
wire \resq[16]~30 ;
wire \resq[16]~31 ;
wire \resq[17]~33_sumout ;
wire \resq[17]~34 ;
wire \resq[17]~35 ;
wire \resq[18]~37_sumout ;
wire \resq[18]~38 ;
wire \resq[18]~39 ;
wire \resq[19]~41_sumout ;
wire \resq[19]~42 ;
wire \resq[19]~43 ;
wire \resq[20]~45_sumout ;
wire \resq[20]~46 ;
wire \resq[20]~47 ;
wire \resq[21]~49_sumout ;
wire \resq[21]~50 ;
wire \resq[21]~51 ;
wire \resq[22]~53_sumout ;
wire \resq[22]~54 ;
wire \resq[22]~55 ;
wire \resq[23]~57_sumout ;
wire \resq[23]~58 ;
wire \resq[23]~59 ;
wire \resq[24]~61_sumout ;
wire \resq[24]~62 ;
wire \resq[24]~63 ;
wire \resq[25]~65_sumout ;
wire \resq[25]~66 ;
wire \resq[25]~67 ;
wire \resq[26]~69_sumout ;
wire \resq[26]~70 ;
wire \resq[26]~71 ;
wire \resq[27]~73_sumout ;
wire \resq[27]~74 ;
wire \resq[27]~75 ;
wire \resq[28]~77_sumout ;
wire \resq[28]~78 ;
wire \resq[28]~79 ;
wire \resq[29]~81_sumout ;
wire \resq[29]~82 ;
wire \resq[29]~83 ;
wire \resq[30]~85_sumout ;
wire \resq[30]~86 ;
wire \resq[30]~87 ;
wire \resq[31]~89_sumout ;
wire \resq[31]~90 ;
wire \resq[31]~91 ;
wire \resq[32]~93_sumout ;
wire \resq[32]~94 ;
wire \resq[32]~95 ;
wire \resq[33]~97_sumout ;
wire \resq[33]~98 ;
wire \resq[33]~99 ;
wire \resq[34]~101_sumout ;
wire \resq[34]~102 ;
wire \resq[34]~103 ;
wire \resq[35]~105_sumout ;
wire \resq[35]~106 ;
wire \resq[35]~107 ;
wire \resq[36]~109_sumout ;
wire \resq[8]~113_sumout ;
wire \resq[7]~117_sumout ;
wire \resq[6]~121_sumout ;
wire \resq[5]~125_sumout ;
wire \resq[4]~129_sumout ;
wire \resq[3]~133_sumout ;
wire \resq[2]~137_sumout ;
wire \resq[1]~141_sumout ;


cic_auk_dspip_delay \glogic:u0 (
	.datain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,q_b_37,q_b_36,q_b_35,q_b_34,q_b_33,q_b_32,q_b_31,q_b_30,q_b_29,q_b_28,q_b_27,q_b_26,q_b_25,q_b_24,q_b_23,q_b_22,q_b_21,q_b_20,q_b_19,q_b_18,q_b_17,q_b_16,q_b_15,q_b_14,q_b_13,q_b_12,q_b_11,q_b_10,q_b_9,q_b_8,q_b_7,q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,q_b_1}),
	.register_fifofifo_data09(\glogic:u0|register_fifo:fifo_data[0][9]~q ),
	.register_fifofifo_data010(\glogic:u0|register_fifo:fifo_data[0][10]~q ),
	.register_fifofifo_data011(\glogic:u0|register_fifo:fifo_data[0][11]~q ),
	.register_fifofifo_data012(\glogic:u0|register_fifo:fifo_data[0][12]~q ),
	.register_fifofifo_data013(\glogic:u0|register_fifo:fifo_data[0][13]~q ),
	.register_fifofifo_data014(\glogic:u0|register_fifo:fifo_data[0][14]~q ),
	.register_fifofifo_data015(\glogic:u0|register_fifo:fifo_data[0][15]~q ),
	.register_fifofifo_data016(\glogic:u0|register_fifo:fifo_data[0][16]~q ),
	.register_fifofifo_data017(\glogic:u0|register_fifo:fifo_data[0][17]~q ),
	.register_fifofifo_data018(\glogic:u0|register_fifo:fifo_data[0][18]~q ),
	.register_fifofifo_data019(\glogic:u0|register_fifo:fifo_data[0][19]~q ),
	.register_fifofifo_data020(\glogic:u0|register_fifo:fifo_data[0][20]~q ),
	.register_fifofifo_data021(\glogic:u0|register_fifo:fifo_data[0][21]~q ),
	.register_fifofifo_data022(\glogic:u0|register_fifo:fifo_data[0][22]~q ),
	.register_fifofifo_data023(\glogic:u0|register_fifo:fifo_data[0][23]~q ),
	.register_fifofifo_data024(\glogic:u0|register_fifo:fifo_data[0][24]~q ),
	.register_fifofifo_data025(\glogic:u0|register_fifo:fifo_data[0][25]~q ),
	.register_fifofifo_data026(\glogic:u0|register_fifo:fifo_data[0][26]~q ),
	.register_fifofifo_data027(\glogic:u0|register_fifo:fifo_data[0][27]~q ),
	.register_fifofifo_data028(\glogic:u0|register_fifo:fifo_data[0][28]~q ),
	.register_fifofifo_data029(\glogic:u0|register_fifo:fifo_data[0][29]~q ),
	.register_fifofifo_data030(\glogic:u0|register_fifo:fifo_data[0][30]~q ),
	.register_fifofifo_data031(\glogic:u0|register_fifo:fifo_data[0][31]~q ),
	.register_fifofifo_data032(\glogic:u0|register_fifo:fifo_data[0][32]~q ),
	.register_fifofifo_data033(\glogic:u0|register_fifo:fifo_data[0][33]~q ),
	.register_fifofifo_data034(\glogic:u0|register_fifo:fifo_data[0][34]~q ),
	.register_fifofifo_data035(\glogic:u0|register_fifo:fifo_data[0][35]~q ),
	.register_fifofifo_data036(\glogic:u0|register_fifo:fifo_data[0][36]~q ),
	.enable(\dout~1_combout ),
	.register_fifofifo_data08(\glogic:u0|register_fifo:fifo_data[0][8]~q ),
	.register_fifofifo_data07(\glogic:u0|register_fifo:fifo_data[0][7]~q ),
	.register_fifofifo_data06(\glogic:u0|register_fifo:fifo_data[0][6]~q ),
	.register_fifofifo_data05(\glogic:u0|register_fifo:fifo_data[0][5]~q ),
	.register_fifofifo_data04(\glogic:u0|register_fifo:fifo_data[0][4]~q ),
	.register_fifofifo_data03(\glogic:u0|register_fifo:fifo_data[0][3]~q ),
	.register_fifofifo_data02(\glogic:u0|register_fifo:fifo_data[0][2]~q ),
	.register_fifofifo_data01(\glogic:u0|register_fifo:fifo_data[0][1]~q ),
	.register_fifofifo_data00(\glogic:u0|register_fifo:fifo_data[0][0]~q ),
	.clk(clk),
	.reset(reset_n));

arriav_lcell_comb \dout~1 (
	.dataa(!stall_reg),
	.datab(!ena_diff_s_1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dout~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dout~1 .extended_lut = "off";
defparam \dout~1 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \dout~1 .shared_arith = "off";

dffeas dout_valid(
	.clk(clk),
	.d(ena_diff_s_1),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(dout_valid2),
	.q(dout_valid1),
	.prn(vcc));
defparam dout_valid.is_wysiwyg = "true";
defparam dout_valid.power_up = "low";

dffeas \dout[9] (
	.clk(clk),
	.d(\resq[9]~1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[36]~0_combout ),
	.q(dout_9),
	.prn(vcc));
defparam \dout[9] .is_wysiwyg = "true";
defparam \dout[9] .power_up = "low";

dffeas \dout[10] (
	.clk(clk),
	.d(\resq[10]~5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[36]~0_combout ),
	.q(dout_10),
	.prn(vcc));
defparam \dout[10] .is_wysiwyg = "true";
defparam \dout[10] .power_up = "low";

dffeas \dout[11] (
	.clk(clk),
	.d(\resq[11]~9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[36]~0_combout ),
	.q(dout_11),
	.prn(vcc));
defparam \dout[11] .is_wysiwyg = "true";
defparam \dout[11] .power_up = "low";

dffeas \dout[12] (
	.clk(clk),
	.d(\resq[12]~13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[36]~0_combout ),
	.q(dout_12),
	.prn(vcc));
defparam \dout[12] .is_wysiwyg = "true";
defparam \dout[12] .power_up = "low";

dffeas \dout[13] (
	.clk(clk),
	.d(\resq[13]~17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[36]~0_combout ),
	.q(dout_13),
	.prn(vcc));
defparam \dout[13] .is_wysiwyg = "true";
defparam \dout[13] .power_up = "low";

dffeas \dout[14] (
	.clk(clk),
	.d(\resq[14]~21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[36]~0_combout ),
	.q(dout_14),
	.prn(vcc));
defparam \dout[14] .is_wysiwyg = "true";
defparam \dout[14] .power_up = "low";

dffeas \dout[15] (
	.clk(clk),
	.d(\resq[15]~25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[36]~0_combout ),
	.q(dout_15),
	.prn(vcc));
defparam \dout[15] .is_wysiwyg = "true";
defparam \dout[15] .power_up = "low";

dffeas \dout[16] (
	.clk(clk),
	.d(\resq[16]~29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[36]~0_combout ),
	.q(dout_16),
	.prn(vcc));
defparam \dout[16] .is_wysiwyg = "true";
defparam \dout[16] .power_up = "low";

dffeas \dout[17] (
	.clk(clk),
	.d(\resq[17]~33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[36]~0_combout ),
	.q(dout_17),
	.prn(vcc));
defparam \dout[17] .is_wysiwyg = "true";
defparam \dout[17] .power_up = "low";

dffeas \dout[18] (
	.clk(clk),
	.d(\resq[18]~37_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[36]~0_combout ),
	.q(dout_18),
	.prn(vcc));
defparam \dout[18] .is_wysiwyg = "true";
defparam \dout[18] .power_up = "low";

dffeas \dout[19] (
	.clk(clk),
	.d(\resq[19]~41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[36]~0_combout ),
	.q(dout_19),
	.prn(vcc));
defparam \dout[19] .is_wysiwyg = "true";
defparam \dout[19] .power_up = "low";

dffeas \dout[20] (
	.clk(clk),
	.d(\resq[20]~45_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[36]~0_combout ),
	.q(dout_20),
	.prn(vcc));
defparam \dout[20] .is_wysiwyg = "true";
defparam \dout[20] .power_up = "low";

dffeas \dout[21] (
	.clk(clk),
	.d(\resq[21]~49_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[36]~0_combout ),
	.q(dout_21),
	.prn(vcc));
defparam \dout[21] .is_wysiwyg = "true";
defparam \dout[21] .power_up = "low";

dffeas \dout[22] (
	.clk(clk),
	.d(\resq[22]~53_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[36]~0_combout ),
	.q(dout_22),
	.prn(vcc));
defparam \dout[22] .is_wysiwyg = "true";
defparam \dout[22] .power_up = "low";

dffeas \dout[23] (
	.clk(clk),
	.d(\resq[23]~57_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[36]~0_combout ),
	.q(dout_23),
	.prn(vcc));
defparam \dout[23] .is_wysiwyg = "true";
defparam \dout[23] .power_up = "low";

dffeas \dout[24] (
	.clk(clk),
	.d(\resq[24]~61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[36]~0_combout ),
	.q(dout_24),
	.prn(vcc));
defparam \dout[24] .is_wysiwyg = "true";
defparam \dout[24] .power_up = "low";

dffeas \dout[25] (
	.clk(clk),
	.d(\resq[25]~65_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[36]~0_combout ),
	.q(dout_25),
	.prn(vcc));
defparam \dout[25] .is_wysiwyg = "true";
defparam \dout[25] .power_up = "low";

dffeas \dout[26] (
	.clk(clk),
	.d(\resq[26]~69_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[36]~0_combout ),
	.q(dout_26),
	.prn(vcc));
defparam \dout[26] .is_wysiwyg = "true";
defparam \dout[26] .power_up = "low";

dffeas \dout[27] (
	.clk(clk),
	.d(\resq[27]~73_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[36]~0_combout ),
	.q(dout_27),
	.prn(vcc));
defparam \dout[27] .is_wysiwyg = "true";
defparam \dout[27] .power_up = "low";

dffeas \dout[28] (
	.clk(clk),
	.d(\resq[28]~77_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[36]~0_combout ),
	.q(dout_28),
	.prn(vcc));
defparam \dout[28] .is_wysiwyg = "true";
defparam \dout[28] .power_up = "low";

dffeas \dout[29] (
	.clk(clk),
	.d(\resq[29]~81_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[36]~0_combout ),
	.q(dout_29),
	.prn(vcc));
defparam \dout[29] .is_wysiwyg = "true";
defparam \dout[29] .power_up = "low";

dffeas \dout[30] (
	.clk(clk),
	.d(\resq[30]~85_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[36]~0_combout ),
	.q(dout_30),
	.prn(vcc));
defparam \dout[30] .is_wysiwyg = "true";
defparam \dout[30] .power_up = "low";

dffeas \dout[31] (
	.clk(clk),
	.d(\resq[31]~89_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[36]~0_combout ),
	.q(dout_31),
	.prn(vcc));
defparam \dout[31] .is_wysiwyg = "true";
defparam \dout[31] .power_up = "low";

dffeas \dout[32] (
	.clk(clk),
	.d(\resq[32]~93_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[36]~0_combout ),
	.q(dout_32),
	.prn(vcc));
defparam \dout[32] .is_wysiwyg = "true";
defparam \dout[32] .power_up = "low";

dffeas \dout[33] (
	.clk(clk),
	.d(\resq[33]~97_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[36]~0_combout ),
	.q(dout_33),
	.prn(vcc));
defparam \dout[33] .is_wysiwyg = "true";
defparam \dout[33] .power_up = "low";

dffeas \dout[34] (
	.clk(clk),
	.d(\resq[34]~101_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[36]~0_combout ),
	.q(dout_34),
	.prn(vcc));
defparam \dout[34] .is_wysiwyg = "true";
defparam \dout[34] .power_up = "low";

dffeas \dout[35] (
	.clk(clk),
	.d(\resq[35]~105_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[36]~0_combout ),
	.q(dout_35),
	.prn(vcc));
defparam \dout[35] .is_wysiwyg = "true";
defparam \dout[35] .power_up = "low";

dffeas \dout[36] (
	.clk(clk),
	.d(\resq[36]~109_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[36]~0_combout ),
	.q(dout_36),
	.prn(vcc));
defparam \dout[36] .is_wysiwyg = "true";
defparam \dout[36] .power_up = "low";

dffeas \dout[8] (
	.clk(clk),
	.d(\resq[8]~113_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[36]~0_combout ),
	.q(dout_8),
	.prn(vcc));
defparam \dout[8] .is_wysiwyg = "true";
defparam \dout[8] .power_up = "low";

dffeas \dout[7] (
	.clk(clk),
	.d(\resq[7]~117_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[36]~0_combout ),
	.q(dout_7),
	.prn(vcc));
defparam \dout[7] .is_wysiwyg = "true";
defparam \dout[7] .power_up = "low";

dffeas \dout[6] (
	.clk(clk),
	.d(\resq[6]~121_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[36]~0_combout ),
	.q(dout_6),
	.prn(vcc));
defparam \dout[6] .is_wysiwyg = "true";
defparam \dout[6] .power_up = "low";

dffeas \dout[5] (
	.clk(clk),
	.d(\resq[5]~125_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[36]~0_combout ),
	.q(dout_5),
	.prn(vcc));
defparam \dout[5] .is_wysiwyg = "true";
defparam \dout[5] .power_up = "low";

dffeas \dout[4] (
	.clk(clk),
	.d(\resq[4]~129_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[36]~0_combout ),
	.q(dout_4),
	.prn(vcc));
defparam \dout[4] .is_wysiwyg = "true";
defparam \dout[4] .power_up = "low";

dffeas \dout[3] (
	.clk(clk),
	.d(\resq[3]~133_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[36]~0_combout ),
	.q(dout_3),
	.prn(vcc));
defparam \dout[3] .is_wysiwyg = "true";
defparam \dout[3] .power_up = "low";

dffeas \dout[2] (
	.clk(clk),
	.d(\resq[2]~137_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[36]~0_combout ),
	.q(dout_2),
	.prn(vcc));
defparam \dout[2] .is_wysiwyg = "true";
defparam \dout[2] .power_up = "low";

dffeas \dout[1] (
	.clk(clk),
	.d(\resq[1]~141_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[36]~0_combout ),
	.q(dout_1),
	.prn(vcc));
defparam \dout[1] .is_wysiwyg = "true";
defparam \dout[1] .power_up = "low";

arriav_lcell_comb \resq[0]~146 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!q_b_1),
	.datad(!\glogic:u0|register_fifo:fifo_data[0][0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\resq[0]~146_cout ),
	.shareout(\resq[0]~147 ));
defparam \resq[0]~146 .extended_lut = "off";
defparam \resq[0]~146 .lut_mask = 64'h0000FF0F00000FF0;
defparam \resq[0]~146 .shared_arith = "on";

arriav_lcell_comb \resq[1]~141 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!q_b_2),
	.datad(!\glogic:u0|register_fifo:fifo_data[0][1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[0]~146_cout ),
	.sharein(\resq[0]~147 ),
	.combout(),
	.sumout(\resq[1]~141_sumout ),
	.cout(\resq[1]~142 ),
	.shareout(\resq[1]~143 ));
defparam \resq[1]~141 .extended_lut = "off";
defparam \resq[1]~141 .lut_mask = 64'h0000FF0F00000FF0;
defparam \resq[1]~141 .shared_arith = "on";

arriav_lcell_comb \resq[2]~137 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!q_b_3),
	.datad(!\glogic:u0|register_fifo:fifo_data[0][2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[1]~142 ),
	.sharein(\resq[1]~143 ),
	.combout(),
	.sumout(\resq[2]~137_sumout ),
	.cout(\resq[2]~138 ),
	.shareout(\resq[2]~139 ));
defparam \resq[2]~137 .extended_lut = "off";
defparam \resq[2]~137 .lut_mask = 64'h0000FF0F00000FF0;
defparam \resq[2]~137 .shared_arith = "on";

arriav_lcell_comb \resq[3]~133 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!q_b_4),
	.datad(!\glogic:u0|register_fifo:fifo_data[0][3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[2]~138 ),
	.sharein(\resq[2]~139 ),
	.combout(),
	.sumout(\resq[3]~133_sumout ),
	.cout(\resq[3]~134 ),
	.shareout(\resq[3]~135 ));
defparam \resq[3]~133 .extended_lut = "off";
defparam \resq[3]~133 .lut_mask = 64'h0000FF0F00000FF0;
defparam \resq[3]~133 .shared_arith = "on";

arriav_lcell_comb \resq[4]~129 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!q_b_5),
	.datad(!\glogic:u0|register_fifo:fifo_data[0][4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[3]~134 ),
	.sharein(\resq[3]~135 ),
	.combout(),
	.sumout(\resq[4]~129_sumout ),
	.cout(\resq[4]~130 ),
	.shareout(\resq[4]~131 ));
defparam \resq[4]~129 .extended_lut = "off";
defparam \resq[4]~129 .lut_mask = 64'h0000FF0F00000FF0;
defparam \resq[4]~129 .shared_arith = "on";

arriav_lcell_comb \resq[5]~125 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!q_b_6),
	.datad(!\glogic:u0|register_fifo:fifo_data[0][5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[4]~130 ),
	.sharein(\resq[4]~131 ),
	.combout(),
	.sumout(\resq[5]~125_sumout ),
	.cout(\resq[5]~126 ),
	.shareout(\resq[5]~127 ));
defparam \resq[5]~125 .extended_lut = "off";
defparam \resq[5]~125 .lut_mask = 64'h0000FF0F00000FF0;
defparam \resq[5]~125 .shared_arith = "on";

arriav_lcell_comb \resq[6]~121 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!q_b_7),
	.datad(!\glogic:u0|register_fifo:fifo_data[0][6]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[5]~126 ),
	.sharein(\resq[5]~127 ),
	.combout(),
	.sumout(\resq[6]~121_sumout ),
	.cout(\resq[6]~122 ),
	.shareout(\resq[6]~123 ));
defparam \resq[6]~121 .extended_lut = "off";
defparam \resq[6]~121 .lut_mask = 64'h0000FF0F00000FF0;
defparam \resq[6]~121 .shared_arith = "on";

arriav_lcell_comb \resq[7]~117 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!q_b_8),
	.datad(!\glogic:u0|register_fifo:fifo_data[0][7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[6]~122 ),
	.sharein(\resq[6]~123 ),
	.combout(),
	.sumout(\resq[7]~117_sumout ),
	.cout(\resq[7]~118 ),
	.shareout(\resq[7]~119 ));
defparam \resq[7]~117 .extended_lut = "off";
defparam \resq[7]~117 .lut_mask = 64'h0000FF0F00000FF0;
defparam \resq[7]~117 .shared_arith = "on";

arriav_lcell_comb \resq[8]~113 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!q_b_9),
	.datad(!\glogic:u0|register_fifo:fifo_data[0][8]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[7]~118 ),
	.sharein(\resq[7]~119 ),
	.combout(),
	.sumout(\resq[8]~113_sumout ),
	.cout(\resq[8]~114 ),
	.shareout(\resq[8]~115 ));
defparam \resq[8]~113 .extended_lut = "off";
defparam \resq[8]~113 .lut_mask = 64'h0000FF0F00000FF0;
defparam \resq[8]~113 .shared_arith = "on";

arriav_lcell_comb \resq[9]~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!q_b_10),
	.datad(!\glogic:u0|register_fifo:fifo_data[0][9]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[8]~114 ),
	.sharein(\resq[8]~115 ),
	.combout(),
	.sumout(\resq[9]~1_sumout ),
	.cout(\resq[9]~2 ),
	.shareout(\resq[9]~3 ));
defparam \resq[9]~1 .extended_lut = "off";
defparam \resq[9]~1 .lut_mask = 64'h0000FF0F00000FF0;
defparam \resq[9]~1 .shared_arith = "on";

arriav_lcell_comb \dout[36]~0 (
	.dataa(!reset_n),
	.datab(!stall_reg),
	.datac(!ena_diff_s_1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dout[36]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dout[36]~0 .extended_lut = "off";
defparam \dout[36]~0 .lut_mask = 64'hEFEFEFEFEFEFEFEF;
defparam \dout[36]~0 .shared_arith = "off";

arriav_lcell_comb \resq[10]~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!q_b_11),
	.datad(!\glogic:u0|register_fifo:fifo_data[0][10]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[9]~2 ),
	.sharein(\resq[9]~3 ),
	.combout(),
	.sumout(\resq[10]~5_sumout ),
	.cout(\resq[10]~6 ),
	.shareout(\resq[10]~7 ));
defparam \resq[10]~5 .extended_lut = "off";
defparam \resq[10]~5 .lut_mask = 64'h0000FF0F00000FF0;
defparam \resq[10]~5 .shared_arith = "on";

arriav_lcell_comb \resq[11]~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!q_b_12),
	.datad(!\glogic:u0|register_fifo:fifo_data[0][11]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[10]~6 ),
	.sharein(\resq[10]~7 ),
	.combout(),
	.sumout(\resq[11]~9_sumout ),
	.cout(\resq[11]~10 ),
	.shareout(\resq[11]~11 ));
defparam \resq[11]~9 .extended_lut = "off";
defparam \resq[11]~9 .lut_mask = 64'h0000FF0F00000FF0;
defparam \resq[11]~9 .shared_arith = "on";

arriav_lcell_comb \resq[12]~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!q_b_13),
	.datad(!\glogic:u0|register_fifo:fifo_data[0][12]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[11]~10 ),
	.sharein(\resq[11]~11 ),
	.combout(),
	.sumout(\resq[12]~13_sumout ),
	.cout(\resq[12]~14 ),
	.shareout(\resq[12]~15 ));
defparam \resq[12]~13 .extended_lut = "off";
defparam \resq[12]~13 .lut_mask = 64'h0000FF0F00000FF0;
defparam \resq[12]~13 .shared_arith = "on";

arriav_lcell_comb \resq[13]~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!q_b_14),
	.datad(!\glogic:u0|register_fifo:fifo_data[0][13]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[12]~14 ),
	.sharein(\resq[12]~15 ),
	.combout(),
	.sumout(\resq[13]~17_sumout ),
	.cout(\resq[13]~18 ),
	.shareout(\resq[13]~19 ));
defparam \resq[13]~17 .extended_lut = "off";
defparam \resq[13]~17 .lut_mask = 64'h0000FF0F00000FF0;
defparam \resq[13]~17 .shared_arith = "on";

arriav_lcell_comb \resq[14]~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!q_b_15),
	.datad(!\glogic:u0|register_fifo:fifo_data[0][14]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[13]~18 ),
	.sharein(\resq[13]~19 ),
	.combout(),
	.sumout(\resq[14]~21_sumout ),
	.cout(\resq[14]~22 ),
	.shareout(\resq[14]~23 ));
defparam \resq[14]~21 .extended_lut = "off";
defparam \resq[14]~21 .lut_mask = 64'h0000FF0F00000FF0;
defparam \resq[14]~21 .shared_arith = "on";

arriav_lcell_comb \resq[15]~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!q_b_16),
	.datad(!\glogic:u0|register_fifo:fifo_data[0][15]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[14]~22 ),
	.sharein(\resq[14]~23 ),
	.combout(),
	.sumout(\resq[15]~25_sumout ),
	.cout(\resq[15]~26 ),
	.shareout(\resq[15]~27 ));
defparam \resq[15]~25 .extended_lut = "off";
defparam \resq[15]~25 .lut_mask = 64'h0000FF0F00000FF0;
defparam \resq[15]~25 .shared_arith = "on";

arriav_lcell_comb \resq[16]~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!q_b_17),
	.datad(!\glogic:u0|register_fifo:fifo_data[0][16]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[15]~26 ),
	.sharein(\resq[15]~27 ),
	.combout(),
	.sumout(\resq[16]~29_sumout ),
	.cout(\resq[16]~30 ),
	.shareout(\resq[16]~31 ));
defparam \resq[16]~29 .extended_lut = "off";
defparam \resq[16]~29 .lut_mask = 64'h0000FF0F00000FF0;
defparam \resq[16]~29 .shared_arith = "on";

arriav_lcell_comb \resq[17]~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!q_b_18),
	.datad(!\glogic:u0|register_fifo:fifo_data[0][17]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[16]~30 ),
	.sharein(\resq[16]~31 ),
	.combout(),
	.sumout(\resq[17]~33_sumout ),
	.cout(\resq[17]~34 ),
	.shareout(\resq[17]~35 ));
defparam \resq[17]~33 .extended_lut = "off";
defparam \resq[17]~33 .lut_mask = 64'h0000FF0F00000FF0;
defparam \resq[17]~33 .shared_arith = "on";

arriav_lcell_comb \resq[18]~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!q_b_19),
	.datad(!\glogic:u0|register_fifo:fifo_data[0][18]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[17]~34 ),
	.sharein(\resq[17]~35 ),
	.combout(),
	.sumout(\resq[18]~37_sumout ),
	.cout(\resq[18]~38 ),
	.shareout(\resq[18]~39 ));
defparam \resq[18]~37 .extended_lut = "off";
defparam \resq[18]~37 .lut_mask = 64'h0000FF0F00000FF0;
defparam \resq[18]~37 .shared_arith = "on";

arriav_lcell_comb \resq[19]~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!q_b_20),
	.datad(!\glogic:u0|register_fifo:fifo_data[0][19]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[18]~38 ),
	.sharein(\resq[18]~39 ),
	.combout(),
	.sumout(\resq[19]~41_sumout ),
	.cout(\resq[19]~42 ),
	.shareout(\resq[19]~43 ));
defparam \resq[19]~41 .extended_lut = "off";
defparam \resq[19]~41 .lut_mask = 64'h0000FF0F00000FF0;
defparam \resq[19]~41 .shared_arith = "on";

arriav_lcell_comb \resq[20]~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!q_b_21),
	.datad(!\glogic:u0|register_fifo:fifo_data[0][20]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[19]~42 ),
	.sharein(\resq[19]~43 ),
	.combout(),
	.sumout(\resq[20]~45_sumout ),
	.cout(\resq[20]~46 ),
	.shareout(\resq[20]~47 ));
defparam \resq[20]~45 .extended_lut = "off";
defparam \resq[20]~45 .lut_mask = 64'h0000FF0F00000FF0;
defparam \resq[20]~45 .shared_arith = "on";

arriav_lcell_comb \resq[21]~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!q_b_22),
	.datad(!\glogic:u0|register_fifo:fifo_data[0][21]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[20]~46 ),
	.sharein(\resq[20]~47 ),
	.combout(),
	.sumout(\resq[21]~49_sumout ),
	.cout(\resq[21]~50 ),
	.shareout(\resq[21]~51 ));
defparam \resq[21]~49 .extended_lut = "off";
defparam \resq[21]~49 .lut_mask = 64'h0000FF0F00000FF0;
defparam \resq[21]~49 .shared_arith = "on";

arriav_lcell_comb \resq[22]~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!q_b_23),
	.datad(!\glogic:u0|register_fifo:fifo_data[0][22]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[21]~50 ),
	.sharein(\resq[21]~51 ),
	.combout(),
	.sumout(\resq[22]~53_sumout ),
	.cout(\resq[22]~54 ),
	.shareout(\resq[22]~55 ));
defparam \resq[22]~53 .extended_lut = "off";
defparam \resq[22]~53 .lut_mask = 64'h0000FF0F00000FF0;
defparam \resq[22]~53 .shared_arith = "on";

arriav_lcell_comb \resq[23]~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!q_b_24),
	.datad(!\glogic:u0|register_fifo:fifo_data[0][23]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[22]~54 ),
	.sharein(\resq[22]~55 ),
	.combout(),
	.sumout(\resq[23]~57_sumout ),
	.cout(\resq[23]~58 ),
	.shareout(\resq[23]~59 ));
defparam \resq[23]~57 .extended_lut = "off";
defparam \resq[23]~57 .lut_mask = 64'h0000FF0F00000FF0;
defparam \resq[23]~57 .shared_arith = "on";

arriav_lcell_comb \resq[24]~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!q_b_25),
	.datad(!\glogic:u0|register_fifo:fifo_data[0][24]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[23]~58 ),
	.sharein(\resq[23]~59 ),
	.combout(),
	.sumout(\resq[24]~61_sumout ),
	.cout(\resq[24]~62 ),
	.shareout(\resq[24]~63 ));
defparam \resq[24]~61 .extended_lut = "off";
defparam \resq[24]~61 .lut_mask = 64'h0000FF0F00000FF0;
defparam \resq[24]~61 .shared_arith = "on";

arriav_lcell_comb \resq[25]~65 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!q_b_26),
	.datad(!\glogic:u0|register_fifo:fifo_data[0][25]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[24]~62 ),
	.sharein(\resq[24]~63 ),
	.combout(),
	.sumout(\resq[25]~65_sumout ),
	.cout(\resq[25]~66 ),
	.shareout(\resq[25]~67 ));
defparam \resq[25]~65 .extended_lut = "off";
defparam \resq[25]~65 .lut_mask = 64'h0000FF0F00000FF0;
defparam \resq[25]~65 .shared_arith = "on";

arriav_lcell_comb \resq[26]~69 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!q_b_27),
	.datad(!\glogic:u0|register_fifo:fifo_data[0][26]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[25]~66 ),
	.sharein(\resq[25]~67 ),
	.combout(),
	.sumout(\resq[26]~69_sumout ),
	.cout(\resq[26]~70 ),
	.shareout(\resq[26]~71 ));
defparam \resq[26]~69 .extended_lut = "off";
defparam \resq[26]~69 .lut_mask = 64'h0000FF0F00000FF0;
defparam \resq[26]~69 .shared_arith = "on";

arriav_lcell_comb \resq[27]~73 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!q_b_28),
	.datad(!\glogic:u0|register_fifo:fifo_data[0][27]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[26]~70 ),
	.sharein(\resq[26]~71 ),
	.combout(),
	.sumout(\resq[27]~73_sumout ),
	.cout(\resq[27]~74 ),
	.shareout(\resq[27]~75 ));
defparam \resq[27]~73 .extended_lut = "off";
defparam \resq[27]~73 .lut_mask = 64'h0000FF0F00000FF0;
defparam \resq[27]~73 .shared_arith = "on";

arriav_lcell_comb \resq[28]~77 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!q_b_29),
	.datad(!\glogic:u0|register_fifo:fifo_data[0][28]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[27]~74 ),
	.sharein(\resq[27]~75 ),
	.combout(),
	.sumout(\resq[28]~77_sumout ),
	.cout(\resq[28]~78 ),
	.shareout(\resq[28]~79 ));
defparam \resq[28]~77 .extended_lut = "off";
defparam \resq[28]~77 .lut_mask = 64'h0000FF0F00000FF0;
defparam \resq[28]~77 .shared_arith = "on";

arriav_lcell_comb \resq[29]~81 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!q_b_30),
	.datad(!\glogic:u0|register_fifo:fifo_data[0][29]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[28]~78 ),
	.sharein(\resq[28]~79 ),
	.combout(),
	.sumout(\resq[29]~81_sumout ),
	.cout(\resq[29]~82 ),
	.shareout(\resq[29]~83 ));
defparam \resq[29]~81 .extended_lut = "off";
defparam \resq[29]~81 .lut_mask = 64'h0000FF0F00000FF0;
defparam \resq[29]~81 .shared_arith = "on";

arriav_lcell_comb \resq[30]~85 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!q_b_31),
	.datad(!\glogic:u0|register_fifo:fifo_data[0][30]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[29]~82 ),
	.sharein(\resq[29]~83 ),
	.combout(),
	.sumout(\resq[30]~85_sumout ),
	.cout(\resq[30]~86 ),
	.shareout(\resq[30]~87 ));
defparam \resq[30]~85 .extended_lut = "off";
defparam \resq[30]~85 .lut_mask = 64'h0000FF0F00000FF0;
defparam \resq[30]~85 .shared_arith = "on";

arriav_lcell_comb \resq[31]~89 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!q_b_32),
	.datad(!\glogic:u0|register_fifo:fifo_data[0][31]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[30]~86 ),
	.sharein(\resq[30]~87 ),
	.combout(),
	.sumout(\resq[31]~89_sumout ),
	.cout(\resq[31]~90 ),
	.shareout(\resq[31]~91 ));
defparam \resq[31]~89 .extended_lut = "off";
defparam \resq[31]~89 .lut_mask = 64'h0000FF0F00000FF0;
defparam \resq[31]~89 .shared_arith = "on";

arriav_lcell_comb \resq[32]~93 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!q_b_33),
	.datad(!\glogic:u0|register_fifo:fifo_data[0][32]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[31]~90 ),
	.sharein(\resq[31]~91 ),
	.combout(),
	.sumout(\resq[32]~93_sumout ),
	.cout(\resq[32]~94 ),
	.shareout(\resq[32]~95 ));
defparam \resq[32]~93 .extended_lut = "off";
defparam \resq[32]~93 .lut_mask = 64'h0000FF0F00000FF0;
defparam \resq[32]~93 .shared_arith = "on";

arriav_lcell_comb \resq[33]~97 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!q_b_34),
	.datad(!\glogic:u0|register_fifo:fifo_data[0][33]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[32]~94 ),
	.sharein(\resq[32]~95 ),
	.combout(),
	.sumout(\resq[33]~97_sumout ),
	.cout(\resq[33]~98 ),
	.shareout(\resq[33]~99 ));
defparam \resq[33]~97 .extended_lut = "off";
defparam \resq[33]~97 .lut_mask = 64'h0000FF0F00000FF0;
defparam \resq[33]~97 .shared_arith = "on";

arriav_lcell_comb \resq[34]~101 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!q_b_35),
	.datad(!\glogic:u0|register_fifo:fifo_data[0][34]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[33]~98 ),
	.sharein(\resq[33]~99 ),
	.combout(),
	.sumout(\resq[34]~101_sumout ),
	.cout(\resq[34]~102 ),
	.shareout(\resq[34]~103 ));
defparam \resq[34]~101 .extended_lut = "off";
defparam \resq[34]~101 .lut_mask = 64'h0000FF0F00000FF0;
defparam \resq[34]~101 .shared_arith = "on";

arriav_lcell_comb \resq[35]~105 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!q_b_36),
	.datad(!\glogic:u0|register_fifo:fifo_data[0][35]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[34]~102 ),
	.sharein(\resq[34]~103 ),
	.combout(),
	.sumout(\resq[35]~105_sumout ),
	.cout(\resq[35]~106 ),
	.shareout(\resq[35]~107 ));
defparam \resq[35]~105 .extended_lut = "off";
defparam \resq[35]~105 .lut_mask = 64'h0000FF0F00000FF0;
defparam \resq[35]~105 .shared_arith = "on";

arriav_lcell_comb \resq[36]~109 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!q_b_37),
	.datad(!\glogic:u0|register_fifo:fifo_data[0][36]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[35]~106 ),
	.sharein(\resq[35]~107 ),
	.combout(),
	.sumout(\resq[36]~109_sumout ),
	.cout(),
	.shareout());
defparam \resq[36]~109 .extended_lut = "off";
defparam \resq[36]~109 .lut_mask = 64'h0000000000000FF0;
defparam \resq[36]~109 .shared_arith = "on";

endmodule

module cic_auk_dspip_delay (
	datain,
	register_fifofifo_data09,
	register_fifofifo_data010,
	register_fifofifo_data011,
	register_fifofifo_data012,
	register_fifofifo_data013,
	register_fifofifo_data014,
	register_fifofifo_data015,
	register_fifofifo_data016,
	register_fifofifo_data017,
	register_fifofifo_data018,
	register_fifofifo_data019,
	register_fifofifo_data020,
	register_fifofifo_data021,
	register_fifofifo_data022,
	register_fifofifo_data023,
	register_fifofifo_data024,
	register_fifofifo_data025,
	register_fifofifo_data026,
	register_fifofifo_data027,
	register_fifofifo_data028,
	register_fifofifo_data029,
	register_fifofifo_data030,
	register_fifofifo_data031,
	register_fifofifo_data032,
	register_fifofifo_data033,
	register_fifofifo_data034,
	register_fifofifo_data035,
	register_fifofifo_data036,
	enable,
	register_fifofifo_data08,
	register_fifofifo_data07,
	register_fifofifo_data06,
	register_fifofifo_data05,
	register_fifofifo_data04,
	register_fifofifo_data03,
	register_fifofifo_data02,
	register_fifofifo_data01,
	register_fifofifo_data00,
	clk,
	reset)/* synthesis synthesis_greybox=1 */;
input 	[46:0] datain;
output 	register_fifofifo_data09;
output 	register_fifofifo_data010;
output 	register_fifofifo_data011;
output 	register_fifofifo_data012;
output 	register_fifofifo_data013;
output 	register_fifofifo_data014;
output 	register_fifofifo_data015;
output 	register_fifofifo_data016;
output 	register_fifofifo_data017;
output 	register_fifofifo_data018;
output 	register_fifofifo_data019;
output 	register_fifofifo_data020;
output 	register_fifofifo_data021;
output 	register_fifofifo_data022;
output 	register_fifofifo_data023;
output 	register_fifofifo_data024;
output 	register_fifofifo_data025;
output 	register_fifofifo_data026;
output 	register_fifofifo_data027;
output 	register_fifofifo_data028;
output 	register_fifofifo_data029;
output 	register_fifofifo_data030;
output 	register_fifofifo_data031;
output 	register_fifofifo_data032;
output 	register_fifofifo_data033;
output 	register_fifofifo_data034;
output 	register_fifofifo_data035;
output 	register_fifofifo_data036;
input 	enable;
output 	register_fifofifo_data08;
output 	register_fifofifo_data07;
output 	register_fifofifo_data06;
output 	register_fifofifo_data05;
output 	register_fifofifo_data04;
output 	register_fifofifo_data03;
output 	register_fifofifo_data02;
output 	register_fifofifo_data01;
output 	register_fifofifo_data00;
input 	clk;
input 	reset;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \register_fifo:fifo_data[0][9] (
	.clk(clk),
	.d(datain[9]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data09),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][9] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][9] .power_up = "low";

dffeas \register_fifo:fifo_data[0][10] (
	.clk(clk),
	.d(datain[10]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data010),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][10] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][10] .power_up = "low";

dffeas \register_fifo:fifo_data[0][11] (
	.clk(clk),
	.d(datain[11]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data011),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][11] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][11] .power_up = "low";

dffeas \register_fifo:fifo_data[0][12] (
	.clk(clk),
	.d(datain[12]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data012),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][12] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][12] .power_up = "low";

dffeas \register_fifo:fifo_data[0][13] (
	.clk(clk),
	.d(datain[13]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data013),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][13] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][13] .power_up = "low";

dffeas \register_fifo:fifo_data[0][14] (
	.clk(clk),
	.d(datain[14]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data014),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][14] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][14] .power_up = "low";

dffeas \register_fifo:fifo_data[0][15] (
	.clk(clk),
	.d(datain[15]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data015),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][15] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][15] .power_up = "low";

dffeas \register_fifo:fifo_data[0][16] (
	.clk(clk),
	.d(datain[16]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data016),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][16] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][16] .power_up = "low";

dffeas \register_fifo:fifo_data[0][17] (
	.clk(clk),
	.d(datain[17]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data017),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][17] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][17] .power_up = "low";

dffeas \register_fifo:fifo_data[0][18] (
	.clk(clk),
	.d(datain[18]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data018),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][18] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][18] .power_up = "low";

dffeas \register_fifo:fifo_data[0][19] (
	.clk(clk),
	.d(datain[19]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data019),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][19] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][19] .power_up = "low";

dffeas \register_fifo:fifo_data[0][20] (
	.clk(clk),
	.d(datain[20]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data020),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][20] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][20] .power_up = "low";

dffeas \register_fifo:fifo_data[0][21] (
	.clk(clk),
	.d(datain[21]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data021),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][21] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][21] .power_up = "low";

dffeas \register_fifo:fifo_data[0][22] (
	.clk(clk),
	.d(datain[22]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data022),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][22] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][22] .power_up = "low";

dffeas \register_fifo:fifo_data[0][23] (
	.clk(clk),
	.d(datain[23]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data023),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][23] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][23] .power_up = "low";

dffeas \register_fifo:fifo_data[0][24] (
	.clk(clk),
	.d(datain[24]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data024),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][24] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][24] .power_up = "low";

dffeas \register_fifo:fifo_data[0][25] (
	.clk(clk),
	.d(datain[25]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data025),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][25] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][25] .power_up = "low";

dffeas \register_fifo:fifo_data[0][26] (
	.clk(clk),
	.d(datain[26]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data026),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][26] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][26] .power_up = "low";

dffeas \register_fifo:fifo_data[0][27] (
	.clk(clk),
	.d(datain[27]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data027),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][27] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][27] .power_up = "low";

dffeas \register_fifo:fifo_data[0][28] (
	.clk(clk),
	.d(datain[28]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data028),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][28] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][28] .power_up = "low";

dffeas \register_fifo:fifo_data[0][29] (
	.clk(clk),
	.d(datain[29]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data029),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][29] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][29] .power_up = "low";

dffeas \register_fifo:fifo_data[0][30] (
	.clk(clk),
	.d(datain[30]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data030),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][30] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][30] .power_up = "low";

dffeas \register_fifo:fifo_data[0][31] (
	.clk(clk),
	.d(datain[31]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data031),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][31] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][31] .power_up = "low";

dffeas \register_fifo:fifo_data[0][32] (
	.clk(clk),
	.d(datain[32]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data032),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][32] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][32] .power_up = "low";

dffeas \register_fifo:fifo_data[0][33] (
	.clk(clk),
	.d(datain[33]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data033),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][33] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][33] .power_up = "low";

dffeas \register_fifo:fifo_data[0][34] (
	.clk(clk),
	.d(datain[34]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data034),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][34] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][34] .power_up = "low";

dffeas \register_fifo:fifo_data[0][35] (
	.clk(clk),
	.d(datain[35]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data035),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][35] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][35] .power_up = "low";

dffeas \register_fifo:fifo_data[0][36] (
	.clk(clk),
	.d(datain[36]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data036),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][36] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][36] .power_up = "low";

dffeas \register_fifo:fifo_data[0][8] (
	.clk(clk),
	.d(datain[8]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data08),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][8] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][8] .power_up = "low";

dffeas \register_fifo:fifo_data[0][7] (
	.clk(clk),
	.d(datain[7]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data07),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][7] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][7] .power_up = "low";

dffeas \register_fifo:fifo_data[0][6] (
	.clk(clk),
	.d(datain[6]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data06),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][6] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][6] .power_up = "low";

dffeas \register_fifo:fifo_data[0][5] (
	.clk(clk),
	.d(datain[5]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data05),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][5] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][5] .power_up = "low";

dffeas \register_fifo:fifo_data[0][4] (
	.clk(clk),
	.d(datain[4]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data04),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][4] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][4] .power_up = "low";

dffeas \register_fifo:fifo_data[0][3] (
	.clk(clk),
	.d(datain[3]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data03),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][3] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][3] .power_up = "low";

dffeas \register_fifo:fifo_data[0][2] (
	.clk(clk),
	.d(datain[2]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data02),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][2] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][2] .power_up = "low";

dffeas \register_fifo:fifo_data[0][1] (
	.clk(clk),
	.d(datain[1]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data01),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][1] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][1] .power_up = "low";

dffeas \register_fifo:fifo_data[0][0] (
	.clk(clk),
	.d(datain[0]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data00),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][0] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][0] .power_up = "low";

endmodule

module cic_auk_dspip_differentiator_1 (
	dout_valid1,
	dout_valid2,
	dout_8,
	dout_9,
	dout_10,
	dout_11,
	dout_12,
	dout_13,
	dout_14,
	dout_15,
	dout_16,
	dout_17,
	dout_18,
	dout_19,
	dout_20,
	dout_21,
	dout_22,
	dout_23,
	dout_24,
	dout_25,
	dout_26,
	dout_27,
	dout_28,
	dout_29,
	dout_30,
	dout_31,
	dout_32,
	dout_33,
	dout_34,
	dout_35,
	dout_7,
	dout_91,
	dout_6,
	dout_101,
	dout_111,
	dout_121,
	dout_131,
	dout_141,
	dout_151,
	dout_161,
	dout_171,
	dout_181,
	dout_191,
	dout_201,
	dout_211,
	dout_221,
	dout_231,
	dout_241,
	dout_251,
	dout_261,
	dout_271,
	dout_281,
	dout_291,
	dout_301,
	dout_311,
	dout_321,
	dout_331,
	dout_341,
	dout_351,
	dout_36,
	dout_81,
	dout_5,
	dout_71,
	dout_4,
	dout_61,
	dout_3,
	dout_51,
	dout_2,
	dout_41,
	dout_1,
	dout_37,
	dout_210,
	dout_110,
	stall_reg,
	dout_valid3,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	dout_valid1;
input 	dout_valid2;
output 	dout_8;
output 	dout_9;
output 	dout_10;
output 	dout_11;
output 	dout_12;
output 	dout_13;
output 	dout_14;
output 	dout_15;
output 	dout_16;
output 	dout_17;
output 	dout_18;
output 	dout_19;
output 	dout_20;
output 	dout_21;
output 	dout_22;
output 	dout_23;
output 	dout_24;
output 	dout_25;
output 	dout_26;
output 	dout_27;
output 	dout_28;
output 	dout_29;
output 	dout_30;
output 	dout_31;
output 	dout_32;
output 	dout_33;
output 	dout_34;
output 	dout_35;
output 	dout_7;
input 	dout_91;
output 	dout_6;
input 	dout_101;
input 	dout_111;
input 	dout_121;
input 	dout_131;
input 	dout_141;
input 	dout_151;
input 	dout_161;
input 	dout_171;
input 	dout_181;
input 	dout_191;
input 	dout_201;
input 	dout_211;
input 	dout_221;
input 	dout_231;
input 	dout_241;
input 	dout_251;
input 	dout_261;
input 	dout_271;
input 	dout_281;
input 	dout_291;
input 	dout_301;
input 	dout_311;
input 	dout_321;
input 	dout_331;
input 	dout_341;
input 	dout_351;
input 	dout_36;
input 	dout_81;
output 	dout_5;
input 	dout_71;
output 	dout_4;
input 	dout_61;
output 	dout_3;
input 	dout_51;
output 	dout_2;
input 	dout_41;
output 	dout_1;
input 	dout_37;
input 	dout_210;
input 	dout_110;
input 	stall_reg;
input 	dout_valid3;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \glogic:u0|register_fifo:fifo_data[0][8]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][9]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][10]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][11]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][12]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][13]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][14]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][15]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][16]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][17]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][18]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][19]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][20]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][21]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][22]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][23]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][24]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][25]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][26]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][27]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][28]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][29]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][30]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][31]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][32]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][33]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][34]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][35]~q ;
wire \dout~1_combout ;
wire \glogic:u0|register_fifo:fifo_data[0][7]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][6]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][5]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][4]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][3]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][2]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][1]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][0]~q ;
wire \resq[0]~142_cout ;
wire \resq[0]~143 ;
wire \resq[1]~138 ;
wire \resq[1]~139 ;
wire \resq[2]~134 ;
wire \resq[2]~135 ;
wire \resq[3]~130 ;
wire \resq[3]~131 ;
wire \resq[4]~126 ;
wire \resq[4]~127 ;
wire \resq[5]~122 ;
wire \resq[5]~123 ;
wire \resq[6]~118 ;
wire \resq[6]~119 ;
wire \resq[7]~114 ;
wire \resq[7]~115 ;
wire \resq[8]~1_sumout ;
wire \dout[32]~0_combout ;
wire \resq[8]~2 ;
wire \resq[8]~3 ;
wire \resq[9]~5_sumout ;
wire \resq[9]~6 ;
wire \resq[9]~7 ;
wire \resq[10]~9_sumout ;
wire \resq[10]~10 ;
wire \resq[10]~11 ;
wire \resq[11]~13_sumout ;
wire \resq[11]~14 ;
wire \resq[11]~15 ;
wire \resq[12]~17_sumout ;
wire \resq[12]~18 ;
wire \resq[12]~19 ;
wire \resq[13]~21_sumout ;
wire \resq[13]~22 ;
wire \resq[13]~23 ;
wire \resq[14]~25_sumout ;
wire \resq[14]~26 ;
wire \resq[14]~27 ;
wire \resq[15]~29_sumout ;
wire \resq[15]~30 ;
wire \resq[15]~31 ;
wire \resq[16]~33_sumout ;
wire \resq[16]~34 ;
wire \resq[16]~35 ;
wire \resq[17]~37_sumout ;
wire \resq[17]~38 ;
wire \resq[17]~39 ;
wire \resq[18]~41_sumout ;
wire \resq[18]~42 ;
wire \resq[18]~43 ;
wire \resq[19]~45_sumout ;
wire \resq[19]~46 ;
wire \resq[19]~47 ;
wire \resq[20]~49_sumout ;
wire \resq[20]~50 ;
wire \resq[20]~51 ;
wire \resq[21]~53_sumout ;
wire \resq[21]~54 ;
wire \resq[21]~55 ;
wire \resq[22]~57_sumout ;
wire \resq[22]~58 ;
wire \resq[22]~59 ;
wire \resq[23]~61_sumout ;
wire \resq[23]~62 ;
wire \resq[23]~63 ;
wire \resq[24]~65_sumout ;
wire \resq[24]~66 ;
wire \resq[24]~67 ;
wire \resq[25]~69_sumout ;
wire \resq[25]~70 ;
wire \resq[25]~71 ;
wire \resq[26]~73_sumout ;
wire \resq[26]~74 ;
wire \resq[26]~75 ;
wire \resq[27]~77_sumout ;
wire \resq[27]~78 ;
wire \resq[27]~79 ;
wire \resq[28]~81_sumout ;
wire \resq[28]~82 ;
wire \resq[28]~83 ;
wire \resq[29]~85_sumout ;
wire \resq[29]~86 ;
wire \resq[29]~87 ;
wire \resq[30]~89_sumout ;
wire \resq[30]~90 ;
wire \resq[30]~91 ;
wire \resq[31]~93_sumout ;
wire \resq[31]~94 ;
wire \resq[31]~95 ;
wire \resq[32]~97_sumout ;
wire \resq[32]~98 ;
wire \resq[32]~99 ;
wire \resq[33]~101_sumout ;
wire \resq[33]~102 ;
wire \resq[33]~103 ;
wire \resq[34]~105_sumout ;
wire \resq[34]~106 ;
wire \resq[34]~107 ;
wire \resq[35]~109_sumout ;
wire \resq[7]~113_sumout ;
wire \resq[6]~117_sumout ;
wire \resq[5]~121_sumout ;
wire \resq[4]~125_sumout ;
wire \resq[3]~129_sumout ;
wire \resq[2]~133_sumout ;
wire \resq[1]~137_sumout ;


cic_auk_dspip_delay_1 \glogic:u0 (
	.datain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,dout_36,dout_351,dout_341,dout_331,dout_321,dout_311,dout_301,dout_291,dout_281,dout_271,dout_261,dout_251,dout_241,dout_231,dout_221,dout_211,dout_201,dout_191,dout_181,dout_171,dout_161,dout_151,dout_141,dout_131,dout_121,dout_111,dout_101,dout_91,
dout_81,dout_71,dout_61,dout_51,dout_41,dout_37,dout_210,dout_110}),
	.register_fifofifo_data08(\glogic:u0|register_fifo:fifo_data[0][8]~q ),
	.register_fifofifo_data09(\glogic:u0|register_fifo:fifo_data[0][9]~q ),
	.register_fifofifo_data010(\glogic:u0|register_fifo:fifo_data[0][10]~q ),
	.register_fifofifo_data011(\glogic:u0|register_fifo:fifo_data[0][11]~q ),
	.register_fifofifo_data012(\glogic:u0|register_fifo:fifo_data[0][12]~q ),
	.register_fifofifo_data013(\glogic:u0|register_fifo:fifo_data[0][13]~q ),
	.register_fifofifo_data014(\glogic:u0|register_fifo:fifo_data[0][14]~q ),
	.register_fifofifo_data015(\glogic:u0|register_fifo:fifo_data[0][15]~q ),
	.register_fifofifo_data016(\glogic:u0|register_fifo:fifo_data[0][16]~q ),
	.register_fifofifo_data017(\glogic:u0|register_fifo:fifo_data[0][17]~q ),
	.register_fifofifo_data018(\glogic:u0|register_fifo:fifo_data[0][18]~q ),
	.register_fifofifo_data019(\glogic:u0|register_fifo:fifo_data[0][19]~q ),
	.register_fifofifo_data020(\glogic:u0|register_fifo:fifo_data[0][20]~q ),
	.register_fifofifo_data021(\glogic:u0|register_fifo:fifo_data[0][21]~q ),
	.register_fifofifo_data022(\glogic:u0|register_fifo:fifo_data[0][22]~q ),
	.register_fifofifo_data023(\glogic:u0|register_fifo:fifo_data[0][23]~q ),
	.register_fifofifo_data024(\glogic:u0|register_fifo:fifo_data[0][24]~q ),
	.register_fifofifo_data025(\glogic:u0|register_fifo:fifo_data[0][25]~q ),
	.register_fifofifo_data026(\glogic:u0|register_fifo:fifo_data[0][26]~q ),
	.register_fifofifo_data027(\glogic:u0|register_fifo:fifo_data[0][27]~q ),
	.register_fifofifo_data028(\glogic:u0|register_fifo:fifo_data[0][28]~q ),
	.register_fifofifo_data029(\glogic:u0|register_fifo:fifo_data[0][29]~q ),
	.register_fifofifo_data030(\glogic:u0|register_fifo:fifo_data[0][30]~q ),
	.register_fifofifo_data031(\glogic:u0|register_fifo:fifo_data[0][31]~q ),
	.register_fifofifo_data032(\glogic:u0|register_fifo:fifo_data[0][32]~q ),
	.register_fifofifo_data033(\glogic:u0|register_fifo:fifo_data[0][33]~q ),
	.register_fifofifo_data034(\glogic:u0|register_fifo:fifo_data[0][34]~q ),
	.register_fifofifo_data035(\glogic:u0|register_fifo:fifo_data[0][35]~q ),
	.enable(\dout~1_combout ),
	.register_fifofifo_data07(\glogic:u0|register_fifo:fifo_data[0][7]~q ),
	.register_fifofifo_data06(\glogic:u0|register_fifo:fifo_data[0][6]~q ),
	.register_fifofifo_data05(\glogic:u0|register_fifo:fifo_data[0][5]~q ),
	.register_fifofifo_data04(\glogic:u0|register_fifo:fifo_data[0][4]~q ),
	.register_fifofifo_data03(\glogic:u0|register_fifo:fifo_data[0][3]~q ),
	.register_fifofifo_data02(\glogic:u0|register_fifo:fifo_data[0][2]~q ),
	.register_fifofifo_data01(\glogic:u0|register_fifo:fifo_data[0][1]~q ),
	.register_fifofifo_data00(\glogic:u0|register_fifo:fifo_data[0][0]~q ),
	.clk(clk),
	.reset(reset_n));

arriav_lcell_comb \dout~1 (
	.dataa(!stall_reg),
	.datab(!dout_valid2),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dout~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dout~1 .extended_lut = "off";
defparam \dout~1 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \dout~1 .shared_arith = "off";

dffeas dout_valid(
	.clk(clk),
	.d(dout_valid2),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(dout_valid3),
	.q(dout_valid1),
	.prn(vcc));
defparam dout_valid.is_wysiwyg = "true";
defparam dout_valid.power_up = "low";

dffeas \dout[8] (
	.clk(clk),
	.d(\resq[8]~1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[32]~0_combout ),
	.q(dout_8),
	.prn(vcc));
defparam \dout[8] .is_wysiwyg = "true";
defparam \dout[8] .power_up = "low";

dffeas \dout[9] (
	.clk(clk),
	.d(\resq[9]~5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[32]~0_combout ),
	.q(dout_9),
	.prn(vcc));
defparam \dout[9] .is_wysiwyg = "true";
defparam \dout[9] .power_up = "low";

dffeas \dout[10] (
	.clk(clk),
	.d(\resq[10]~9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[32]~0_combout ),
	.q(dout_10),
	.prn(vcc));
defparam \dout[10] .is_wysiwyg = "true";
defparam \dout[10] .power_up = "low";

dffeas \dout[11] (
	.clk(clk),
	.d(\resq[11]~13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[32]~0_combout ),
	.q(dout_11),
	.prn(vcc));
defparam \dout[11] .is_wysiwyg = "true";
defparam \dout[11] .power_up = "low";

dffeas \dout[12] (
	.clk(clk),
	.d(\resq[12]~17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[32]~0_combout ),
	.q(dout_12),
	.prn(vcc));
defparam \dout[12] .is_wysiwyg = "true";
defparam \dout[12] .power_up = "low";

dffeas \dout[13] (
	.clk(clk),
	.d(\resq[13]~21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[32]~0_combout ),
	.q(dout_13),
	.prn(vcc));
defparam \dout[13] .is_wysiwyg = "true";
defparam \dout[13] .power_up = "low";

dffeas \dout[14] (
	.clk(clk),
	.d(\resq[14]~25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[32]~0_combout ),
	.q(dout_14),
	.prn(vcc));
defparam \dout[14] .is_wysiwyg = "true";
defparam \dout[14] .power_up = "low";

dffeas \dout[15] (
	.clk(clk),
	.d(\resq[15]~29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[32]~0_combout ),
	.q(dout_15),
	.prn(vcc));
defparam \dout[15] .is_wysiwyg = "true";
defparam \dout[15] .power_up = "low";

dffeas \dout[16] (
	.clk(clk),
	.d(\resq[16]~33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[32]~0_combout ),
	.q(dout_16),
	.prn(vcc));
defparam \dout[16] .is_wysiwyg = "true";
defparam \dout[16] .power_up = "low";

dffeas \dout[17] (
	.clk(clk),
	.d(\resq[17]~37_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[32]~0_combout ),
	.q(dout_17),
	.prn(vcc));
defparam \dout[17] .is_wysiwyg = "true";
defparam \dout[17] .power_up = "low";

dffeas \dout[18] (
	.clk(clk),
	.d(\resq[18]~41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[32]~0_combout ),
	.q(dout_18),
	.prn(vcc));
defparam \dout[18] .is_wysiwyg = "true";
defparam \dout[18] .power_up = "low";

dffeas \dout[19] (
	.clk(clk),
	.d(\resq[19]~45_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[32]~0_combout ),
	.q(dout_19),
	.prn(vcc));
defparam \dout[19] .is_wysiwyg = "true";
defparam \dout[19] .power_up = "low";

dffeas \dout[20] (
	.clk(clk),
	.d(\resq[20]~49_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[32]~0_combout ),
	.q(dout_20),
	.prn(vcc));
defparam \dout[20] .is_wysiwyg = "true";
defparam \dout[20] .power_up = "low";

dffeas \dout[21] (
	.clk(clk),
	.d(\resq[21]~53_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[32]~0_combout ),
	.q(dout_21),
	.prn(vcc));
defparam \dout[21] .is_wysiwyg = "true";
defparam \dout[21] .power_up = "low";

dffeas \dout[22] (
	.clk(clk),
	.d(\resq[22]~57_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[32]~0_combout ),
	.q(dout_22),
	.prn(vcc));
defparam \dout[22] .is_wysiwyg = "true";
defparam \dout[22] .power_up = "low";

dffeas \dout[23] (
	.clk(clk),
	.d(\resq[23]~61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[32]~0_combout ),
	.q(dout_23),
	.prn(vcc));
defparam \dout[23] .is_wysiwyg = "true";
defparam \dout[23] .power_up = "low";

dffeas \dout[24] (
	.clk(clk),
	.d(\resq[24]~65_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[32]~0_combout ),
	.q(dout_24),
	.prn(vcc));
defparam \dout[24] .is_wysiwyg = "true";
defparam \dout[24] .power_up = "low";

dffeas \dout[25] (
	.clk(clk),
	.d(\resq[25]~69_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[32]~0_combout ),
	.q(dout_25),
	.prn(vcc));
defparam \dout[25] .is_wysiwyg = "true";
defparam \dout[25] .power_up = "low";

dffeas \dout[26] (
	.clk(clk),
	.d(\resq[26]~73_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[32]~0_combout ),
	.q(dout_26),
	.prn(vcc));
defparam \dout[26] .is_wysiwyg = "true";
defparam \dout[26] .power_up = "low";

dffeas \dout[27] (
	.clk(clk),
	.d(\resq[27]~77_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[32]~0_combout ),
	.q(dout_27),
	.prn(vcc));
defparam \dout[27] .is_wysiwyg = "true";
defparam \dout[27] .power_up = "low";

dffeas \dout[28] (
	.clk(clk),
	.d(\resq[28]~81_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[32]~0_combout ),
	.q(dout_28),
	.prn(vcc));
defparam \dout[28] .is_wysiwyg = "true";
defparam \dout[28] .power_up = "low";

dffeas \dout[29] (
	.clk(clk),
	.d(\resq[29]~85_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[32]~0_combout ),
	.q(dout_29),
	.prn(vcc));
defparam \dout[29] .is_wysiwyg = "true";
defparam \dout[29] .power_up = "low";

dffeas \dout[30] (
	.clk(clk),
	.d(\resq[30]~89_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[32]~0_combout ),
	.q(dout_30),
	.prn(vcc));
defparam \dout[30] .is_wysiwyg = "true";
defparam \dout[30] .power_up = "low";

dffeas \dout[31] (
	.clk(clk),
	.d(\resq[31]~93_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[32]~0_combout ),
	.q(dout_31),
	.prn(vcc));
defparam \dout[31] .is_wysiwyg = "true";
defparam \dout[31] .power_up = "low";

dffeas \dout[32] (
	.clk(clk),
	.d(\resq[32]~97_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[32]~0_combout ),
	.q(dout_32),
	.prn(vcc));
defparam \dout[32] .is_wysiwyg = "true";
defparam \dout[32] .power_up = "low";

dffeas \dout[33] (
	.clk(clk),
	.d(\resq[33]~101_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[32]~0_combout ),
	.q(dout_33),
	.prn(vcc));
defparam \dout[33] .is_wysiwyg = "true";
defparam \dout[33] .power_up = "low";

dffeas \dout[34] (
	.clk(clk),
	.d(\resq[34]~105_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[32]~0_combout ),
	.q(dout_34),
	.prn(vcc));
defparam \dout[34] .is_wysiwyg = "true";
defparam \dout[34] .power_up = "low";

dffeas \dout[35] (
	.clk(clk),
	.d(\resq[35]~109_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[32]~0_combout ),
	.q(dout_35),
	.prn(vcc));
defparam \dout[35] .is_wysiwyg = "true";
defparam \dout[35] .power_up = "low";

dffeas \dout[7] (
	.clk(clk),
	.d(\resq[7]~113_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[32]~0_combout ),
	.q(dout_7),
	.prn(vcc));
defparam \dout[7] .is_wysiwyg = "true";
defparam \dout[7] .power_up = "low";

dffeas \dout[6] (
	.clk(clk),
	.d(\resq[6]~117_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[32]~0_combout ),
	.q(dout_6),
	.prn(vcc));
defparam \dout[6] .is_wysiwyg = "true";
defparam \dout[6] .power_up = "low";

dffeas \dout[5] (
	.clk(clk),
	.d(\resq[5]~121_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[32]~0_combout ),
	.q(dout_5),
	.prn(vcc));
defparam \dout[5] .is_wysiwyg = "true";
defparam \dout[5] .power_up = "low";

dffeas \dout[4] (
	.clk(clk),
	.d(\resq[4]~125_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[32]~0_combout ),
	.q(dout_4),
	.prn(vcc));
defparam \dout[4] .is_wysiwyg = "true";
defparam \dout[4] .power_up = "low";

dffeas \dout[3] (
	.clk(clk),
	.d(\resq[3]~129_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[32]~0_combout ),
	.q(dout_3),
	.prn(vcc));
defparam \dout[3] .is_wysiwyg = "true";
defparam \dout[3] .power_up = "low";

dffeas \dout[2] (
	.clk(clk),
	.d(\resq[2]~133_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[32]~0_combout ),
	.q(dout_2),
	.prn(vcc));
defparam \dout[2] .is_wysiwyg = "true";
defparam \dout[2] .power_up = "low";

dffeas \dout[1] (
	.clk(clk),
	.d(\resq[1]~137_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[32]~0_combout ),
	.q(dout_1),
	.prn(vcc));
defparam \dout[1] .is_wysiwyg = "true";
defparam \dout[1] .power_up = "low";

arriav_lcell_comb \resq[0]~142 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][0]~q ),
	.datad(!dout_110),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\resq[0]~142_cout ),
	.shareout(\resq[0]~143 ));
defparam \resq[0]~142 .extended_lut = "off";
defparam \resq[0]~142 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[0]~142 .shared_arith = "on";

arriav_lcell_comb \resq[1]~137 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][1]~q ),
	.datad(!dout_210),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[0]~142_cout ),
	.sharein(\resq[0]~143 ),
	.combout(),
	.sumout(\resq[1]~137_sumout ),
	.cout(\resq[1]~138 ),
	.shareout(\resq[1]~139 ));
defparam \resq[1]~137 .extended_lut = "off";
defparam \resq[1]~137 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[1]~137 .shared_arith = "on";

arriav_lcell_comb \resq[2]~133 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][2]~q ),
	.datad(!dout_37),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[1]~138 ),
	.sharein(\resq[1]~139 ),
	.combout(),
	.sumout(\resq[2]~133_sumout ),
	.cout(\resq[2]~134 ),
	.shareout(\resq[2]~135 ));
defparam \resq[2]~133 .extended_lut = "off";
defparam \resq[2]~133 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[2]~133 .shared_arith = "on";

arriav_lcell_comb \resq[3]~129 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][3]~q ),
	.datad(!dout_41),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[2]~134 ),
	.sharein(\resq[2]~135 ),
	.combout(),
	.sumout(\resq[3]~129_sumout ),
	.cout(\resq[3]~130 ),
	.shareout(\resq[3]~131 ));
defparam \resq[3]~129 .extended_lut = "off";
defparam \resq[3]~129 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[3]~129 .shared_arith = "on";

arriav_lcell_comb \resq[4]~125 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][4]~q ),
	.datad(!dout_51),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[3]~130 ),
	.sharein(\resq[3]~131 ),
	.combout(),
	.sumout(\resq[4]~125_sumout ),
	.cout(\resq[4]~126 ),
	.shareout(\resq[4]~127 ));
defparam \resq[4]~125 .extended_lut = "off";
defparam \resq[4]~125 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[4]~125 .shared_arith = "on";

arriav_lcell_comb \resq[5]~121 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][5]~q ),
	.datad(!dout_61),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[4]~126 ),
	.sharein(\resq[4]~127 ),
	.combout(),
	.sumout(\resq[5]~121_sumout ),
	.cout(\resq[5]~122 ),
	.shareout(\resq[5]~123 ));
defparam \resq[5]~121 .extended_lut = "off";
defparam \resq[5]~121 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[5]~121 .shared_arith = "on";

arriav_lcell_comb \resq[6]~117 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][6]~q ),
	.datad(!dout_71),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[5]~122 ),
	.sharein(\resq[5]~123 ),
	.combout(),
	.sumout(\resq[6]~117_sumout ),
	.cout(\resq[6]~118 ),
	.shareout(\resq[6]~119 ));
defparam \resq[6]~117 .extended_lut = "off";
defparam \resq[6]~117 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[6]~117 .shared_arith = "on";

arriav_lcell_comb \resq[7]~113 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][7]~q ),
	.datad(!dout_81),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[6]~118 ),
	.sharein(\resq[6]~119 ),
	.combout(),
	.sumout(\resq[7]~113_sumout ),
	.cout(\resq[7]~114 ),
	.shareout(\resq[7]~115 ));
defparam \resq[7]~113 .extended_lut = "off";
defparam \resq[7]~113 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[7]~113 .shared_arith = "on";

arriav_lcell_comb \resq[8]~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][8]~q ),
	.datad(!dout_91),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[7]~114 ),
	.sharein(\resq[7]~115 ),
	.combout(),
	.sumout(\resq[8]~1_sumout ),
	.cout(\resq[8]~2 ),
	.shareout(\resq[8]~3 ));
defparam \resq[8]~1 .extended_lut = "off";
defparam \resq[8]~1 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[8]~1 .shared_arith = "on";

arriav_lcell_comb \dout[32]~0 (
	.dataa(!reset_n),
	.datab(!stall_reg),
	.datac(!dout_valid2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dout[32]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dout[32]~0 .extended_lut = "off";
defparam \dout[32]~0 .lut_mask = 64'hEFEFEFEFEFEFEFEF;
defparam \dout[32]~0 .shared_arith = "off";

arriav_lcell_comb \resq[9]~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][9]~q ),
	.datad(!dout_101),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[8]~2 ),
	.sharein(\resq[8]~3 ),
	.combout(),
	.sumout(\resq[9]~5_sumout ),
	.cout(\resq[9]~6 ),
	.shareout(\resq[9]~7 ));
defparam \resq[9]~5 .extended_lut = "off";
defparam \resq[9]~5 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[9]~5 .shared_arith = "on";

arriav_lcell_comb \resq[10]~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][10]~q ),
	.datad(!dout_111),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[9]~6 ),
	.sharein(\resq[9]~7 ),
	.combout(),
	.sumout(\resq[10]~9_sumout ),
	.cout(\resq[10]~10 ),
	.shareout(\resq[10]~11 ));
defparam \resq[10]~9 .extended_lut = "off";
defparam \resq[10]~9 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[10]~9 .shared_arith = "on";

arriav_lcell_comb \resq[11]~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][11]~q ),
	.datad(!dout_121),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[10]~10 ),
	.sharein(\resq[10]~11 ),
	.combout(),
	.sumout(\resq[11]~13_sumout ),
	.cout(\resq[11]~14 ),
	.shareout(\resq[11]~15 ));
defparam \resq[11]~13 .extended_lut = "off";
defparam \resq[11]~13 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[11]~13 .shared_arith = "on";

arriav_lcell_comb \resq[12]~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][12]~q ),
	.datad(!dout_131),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[11]~14 ),
	.sharein(\resq[11]~15 ),
	.combout(),
	.sumout(\resq[12]~17_sumout ),
	.cout(\resq[12]~18 ),
	.shareout(\resq[12]~19 ));
defparam \resq[12]~17 .extended_lut = "off";
defparam \resq[12]~17 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[12]~17 .shared_arith = "on";

arriav_lcell_comb \resq[13]~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][13]~q ),
	.datad(!dout_141),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[12]~18 ),
	.sharein(\resq[12]~19 ),
	.combout(),
	.sumout(\resq[13]~21_sumout ),
	.cout(\resq[13]~22 ),
	.shareout(\resq[13]~23 ));
defparam \resq[13]~21 .extended_lut = "off";
defparam \resq[13]~21 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[13]~21 .shared_arith = "on";

arriav_lcell_comb \resq[14]~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][14]~q ),
	.datad(!dout_151),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[13]~22 ),
	.sharein(\resq[13]~23 ),
	.combout(),
	.sumout(\resq[14]~25_sumout ),
	.cout(\resq[14]~26 ),
	.shareout(\resq[14]~27 ));
defparam \resq[14]~25 .extended_lut = "off";
defparam \resq[14]~25 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[14]~25 .shared_arith = "on";

arriav_lcell_comb \resq[15]~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][15]~q ),
	.datad(!dout_161),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[14]~26 ),
	.sharein(\resq[14]~27 ),
	.combout(),
	.sumout(\resq[15]~29_sumout ),
	.cout(\resq[15]~30 ),
	.shareout(\resq[15]~31 ));
defparam \resq[15]~29 .extended_lut = "off";
defparam \resq[15]~29 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[15]~29 .shared_arith = "on";

arriav_lcell_comb \resq[16]~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][16]~q ),
	.datad(!dout_171),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[15]~30 ),
	.sharein(\resq[15]~31 ),
	.combout(),
	.sumout(\resq[16]~33_sumout ),
	.cout(\resq[16]~34 ),
	.shareout(\resq[16]~35 ));
defparam \resq[16]~33 .extended_lut = "off";
defparam \resq[16]~33 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[16]~33 .shared_arith = "on";

arriav_lcell_comb \resq[17]~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][17]~q ),
	.datad(!dout_181),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[16]~34 ),
	.sharein(\resq[16]~35 ),
	.combout(),
	.sumout(\resq[17]~37_sumout ),
	.cout(\resq[17]~38 ),
	.shareout(\resq[17]~39 ));
defparam \resq[17]~37 .extended_lut = "off";
defparam \resq[17]~37 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[17]~37 .shared_arith = "on";

arriav_lcell_comb \resq[18]~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][18]~q ),
	.datad(!dout_191),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[17]~38 ),
	.sharein(\resq[17]~39 ),
	.combout(),
	.sumout(\resq[18]~41_sumout ),
	.cout(\resq[18]~42 ),
	.shareout(\resq[18]~43 ));
defparam \resq[18]~41 .extended_lut = "off";
defparam \resq[18]~41 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[18]~41 .shared_arith = "on";

arriav_lcell_comb \resq[19]~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][19]~q ),
	.datad(!dout_201),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[18]~42 ),
	.sharein(\resq[18]~43 ),
	.combout(),
	.sumout(\resq[19]~45_sumout ),
	.cout(\resq[19]~46 ),
	.shareout(\resq[19]~47 ));
defparam \resq[19]~45 .extended_lut = "off";
defparam \resq[19]~45 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[19]~45 .shared_arith = "on";

arriav_lcell_comb \resq[20]~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][20]~q ),
	.datad(!dout_211),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[19]~46 ),
	.sharein(\resq[19]~47 ),
	.combout(),
	.sumout(\resq[20]~49_sumout ),
	.cout(\resq[20]~50 ),
	.shareout(\resq[20]~51 ));
defparam \resq[20]~49 .extended_lut = "off";
defparam \resq[20]~49 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[20]~49 .shared_arith = "on";

arriav_lcell_comb \resq[21]~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][21]~q ),
	.datad(!dout_221),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[20]~50 ),
	.sharein(\resq[20]~51 ),
	.combout(),
	.sumout(\resq[21]~53_sumout ),
	.cout(\resq[21]~54 ),
	.shareout(\resq[21]~55 ));
defparam \resq[21]~53 .extended_lut = "off";
defparam \resq[21]~53 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[21]~53 .shared_arith = "on";

arriav_lcell_comb \resq[22]~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][22]~q ),
	.datad(!dout_231),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[21]~54 ),
	.sharein(\resq[21]~55 ),
	.combout(),
	.sumout(\resq[22]~57_sumout ),
	.cout(\resq[22]~58 ),
	.shareout(\resq[22]~59 ));
defparam \resq[22]~57 .extended_lut = "off";
defparam \resq[22]~57 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[22]~57 .shared_arith = "on";

arriav_lcell_comb \resq[23]~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][23]~q ),
	.datad(!dout_241),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[22]~58 ),
	.sharein(\resq[22]~59 ),
	.combout(),
	.sumout(\resq[23]~61_sumout ),
	.cout(\resq[23]~62 ),
	.shareout(\resq[23]~63 ));
defparam \resq[23]~61 .extended_lut = "off";
defparam \resq[23]~61 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[23]~61 .shared_arith = "on";

arriav_lcell_comb \resq[24]~65 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][24]~q ),
	.datad(!dout_251),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[23]~62 ),
	.sharein(\resq[23]~63 ),
	.combout(),
	.sumout(\resq[24]~65_sumout ),
	.cout(\resq[24]~66 ),
	.shareout(\resq[24]~67 ));
defparam \resq[24]~65 .extended_lut = "off";
defparam \resq[24]~65 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[24]~65 .shared_arith = "on";

arriav_lcell_comb \resq[25]~69 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][25]~q ),
	.datad(!dout_261),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[24]~66 ),
	.sharein(\resq[24]~67 ),
	.combout(),
	.sumout(\resq[25]~69_sumout ),
	.cout(\resq[25]~70 ),
	.shareout(\resq[25]~71 ));
defparam \resq[25]~69 .extended_lut = "off";
defparam \resq[25]~69 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[25]~69 .shared_arith = "on";

arriav_lcell_comb \resq[26]~73 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][26]~q ),
	.datad(!dout_271),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[25]~70 ),
	.sharein(\resq[25]~71 ),
	.combout(),
	.sumout(\resq[26]~73_sumout ),
	.cout(\resq[26]~74 ),
	.shareout(\resq[26]~75 ));
defparam \resq[26]~73 .extended_lut = "off";
defparam \resq[26]~73 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[26]~73 .shared_arith = "on";

arriav_lcell_comb \resq[27]~77 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][27]~q ),
	.datad(!dout_281),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[26]~74 ),
	.sharein(\resq[26]~75 ),
	.combout(),
	.sumout(\resq[27]~77_sumout ),
	.cout(\resq[27]~78 ),
	.shareout(\resq[27]~79 ));
defparam \resq[27]~77 .extended_lut = "off";
defparam \resq[27]~77 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[27]~77 .shared_arith = "on";

arriav_lcell_comb \resq[28]~81 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][28]~q ),
	.datad(!dout_291),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[27]~78 ),
	.sharein(\resq[27]~79 ),
	.combout(),
	.sumout(\resq[28]~81_sumout ),
	.cout(\resq[28]~82 ),
	.shareout(\resq[28]~83 ));
defparam \resq[28]~81 .extended_lut = "off";
defparam \resq[28]~81 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[28]~81 .shared_arith = "on";

arriav_lcell_comb \resq[29]~85 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][29]~q ),
	.datad(!dout_301),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[28]~82 ),
	.sharein(\resq[28]~83 ),
	.combout(),
	.sumout(\resq[29]~85_sumout ),
	.cout(\resq[29]~86 ),
	.shareout(\resq[29]~87 ));
defparam \resq[29]~85 .extended_lut = "off";
defparam \resq[29]~85 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[29]~85 .shared_arith = "on";

arriav_lcell_comb \resq[30]~89 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][30]~q ),
	.datad(!dout_311),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[29]~86 ),
	.sharein(\resq[29]~87 ),
	.combout(),
	.sumout(\resq[30]~89_sumout ),
	.cout(\resq[30]~90 ),
	.shareout(\resq[30]~91 ));
defparam \resq[30]~89 .extended_lut = "off";
defparam \resq[30]~89 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[30]~89 .shared_arith = "on";

arriav_lcell_comb \resq[31]~93 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][31]~q ),
	.datad(!dout_321),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[30]~90 ),
	.sharein(\resq[30]~91 ),
	.combout(),
	.sumout(\resq[31]~93_sumout ),
	.cout(\resq[31]~94 ),
	.shareout(\resq[31]~95 ));
defparam \resq[31]~93 .extended_lut = "off";
defparam \resq[31]~93 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[31]~93 .shared_arith = "on";

arriav_lcell_comb \resq[32]~97 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][32]~q ),
	.datad(!dout_331),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[31]~94 ),
	.sharein(\resq[31]~95 ),
	.combout(),
	.sumout(\resq[32]~97_sumout ),
	.cout(\resq[32]~98 ),
	.shareout(\resq[32]~99 ));
defparam \resq[32]~97 .extended_lut = "off";
defparam \resq[32]~97 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[32]~97 .shared_arith = "on";

arriav_lcell_comb \resq[33]~101 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][33]~q ),
	.datad(!dout_341),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[32]~98 ),
	.sharein(\resq[32]~99 ),
	.combout(),
	.sumout(\resq[33]~101_sumout ),
	.cout(\resq[33]~102 ),
	.shareout(\resq[33]~103 ));
defparam \resq[33]~101 .extended_lut = "off";
defparam \resq[33]~101 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[33]~101 .shared_arith = "on";

arriav_lcell_comb \resq[34]~105 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][34]~q ),
	.datad(!dout_351),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[33]~102 ),
	.sharein(\resq[33]~103 ),
	.combout(),
	.sumout(\resq[34]~105_sumout ),
	.cout(\resq[34]~106 ),
	.shareout(\resq[34]~107 ));
defparam \resq[34]~105 .extended_lut = "off";
defparam \resq[34]~105 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[34]~105 .shared_arith = "on";

arriav_lcell_comb \resq[35]~109 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][35]~q ),
	.datad(!dout_36),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[34]~106 ),
	.sharein(\resq[34]~107 ),
	.combout(),
	.sumout(\resq[35]~109_sumout ),
	.cout(),
	.shareout());
defparam \resq[35]~109 .extended_lut = "off";
defparam \resq[35]~109 .lut_mask = 64'h0000000000000FF0;
defparam \resq[35]~109 .shared_arith = "on";

endmodule

module cic_auk_dspip_delay_1 (
	datain,
	register_fifofifo_data08,
	register_fifofifo_data09,
	register_fifofifo_data010,
	register_fifofifo_data011,
	register_fifofifo_data012,
	register_fifofifo_data013,
	register_fifofifo_data014,
	register_fifofifo_data015,
	register_fifofifo_data016,
	register_fifofifo_data017,
	register_fifofifo_data018,
	register_fifofifo_data019,
	register_fifofifo_data020,
	register_fifofifo_data021,
	register_fifofifo_data022,
	register_fifofifo_data023,
	register_fifofifo_data024,
	register_fifofifo_data025,
	register_fifofifo_data026,
	register_fifofifo_data027,
	register_fifofifo_data028,
	register_fifofifo_data029,
	register_fifofifo_data030,
	register_fifofifo_data031,
	register_fifofifo_data032,
	register_fifofifo_data033,
	register_fifofifo_data034,
	register_fifofifo_data035,
	enable,
	register_fifofifo_data07,
	register_fifofifo_data06,
	register_fifofifo_data05,
	register_fifofifo_data04,
	register_fifofifo_data03,
	register_fifofifo_data02,
	register_fifofifo_data01,
	register_fifofifo_data00,
	clk,
	reset)/* synthesis synthesis_greybox=1 */;
input 	[46:0] datain;
output 	register_fifofifo_data08;
output 	register_fifofifo_data09;
output 	register_fifofifo_data010;
output 	register_fifofifo_data011;
output 	register_fifofifo_data012;
output 	register_fifofifo_data013;
output 	register_fifofifo_data014;
output 	register_fifofifo_data015;
output 	register_fifofifo_data016;
output 	register_fifofifo_data017;
output 	register_fifofifo_data018;
output 	register_fifofifo_data019;
output 	register_fifofifo_data020;
output 	register_fifofifo_data021;
output 	register_fifofifo_data022;
output 	register_fifofifo_data023;
output 	register_fifofifo_data024;
output 	register_fifofifo_data025;
output 	register_fifofifo_data026;
output 	register_fifofifo_data027;
output 	register_fifofifo_data028;
output 	register_fifofifo_data029;
output 	register_fifofifo_data030;
output 	register_fifofifo_data031;
output 	register_fifofifo_data032;
output 	register_fifofifo_data033;
output 	register_fifofifo_data034;
output 	register_fifofifo_data035;
input 	enable;
output 	register_fifofifo_data07;
output 	register_fifofifo_data06;
output 	register_fifofifo_data05;
output 	register_fifofifo_data04;
output 	register_fifofifo_data03;
output 	register_fifofifo_data02;
output 	register_fifofifo_data01;
output 	register_fifofifo_data00;
input 	clk;
input 	reset;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \register_fifo:fifo_data[0][8] (
	.clk(clk),
	.d(datain[8]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data08),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][8] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][8] .power_up = "low";

dffeas \register_fifo:fifo_data[0][9] (
	.clk(clk),
	.d(datain[9]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data09),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][9] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][9] .power_up = "low";

dffeas \register_fifo:fifo_data[0][10] (
	.clk(clk),
	.d(datain[10]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data010),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][10] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][10] .power_up = "low";

dffeas \register_fifo:fifo_data[0][11] (
	.clk(clk),
	.d(datain[11]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data011),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][11] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][11] .power_up = "low";

dffeas \register_fifo:fifo_data[0][12] (
	.clk(clk),
	.d(datain[12]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data012),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][12] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][12] .power_up = "low";

dffeas \register_fifo:fifo_data[0][13] (
	.clk(clk),
	.d(datain[13]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data013),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][13] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][13] .power_up = "low";

dffeas \register_fifo:fifo_data[0][14] (
	.clk(clk),
	.d(datain[14]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data014),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][14] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][14] .power_up = "low";

dffeas \register_fifo:fifo_data[0][15] (
	.clk(clk),
	.d(datain[15]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data015),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][15] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][15] .power_up = "low";

dffeas \register_fifo:fifo_data[0][16] (
	.clk(clk),
	.d(datain[16]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data016),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][16] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][16] .power_up = "low";

dffeas \register_fifo:fifo_data[0][17] (
	.clk(clk),
	.d(datain[17]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data017),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][17] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][17] .power_up = "low";

dffeas \register_fifo:fifo_data[0][18] (
	.clk(clk),
	.d(datain[18]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data018),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][18] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][18] .power_up = "low";

dffeas \register_fifo:fifo_data[0][19] (
	.clk(clk),
	.d(datain[19]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data019),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][19] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][19] .power_up = "low";

dffeas \register_fifo:fifo_data[0][20] (
	.clk(clk),
	.d(datain[20]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data020),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][20] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][20] .power_up = "low";

dffeas \register_fifo:fifo_data[0][21] (
	.clk(clk),
	.d(datain[21]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data021),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][21] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][21] .power_up = "low";

dffeas \register_fifo:fifo_data[0][22] (
	.clk(clk),
	.d(datain[22]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data022),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][22] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][22] .power_up = "low";

dffeas \register_fifo:fifo_data[0][23] (
	.clk(clk),
	.d(datain[23]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data023),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][23] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][23] .power_up = "low";

dffeas \register_fifo:fifo_data[0][24] (
	.clk(clk),
	.d(datain[24]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data024),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][24] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][24] .power_up = "low";

dffeas \register_fifo:fifo_data[0][25] (
	.clk(clk),
	.d(datain[25]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data025),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][25] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][25] .power_up = "low";

dffeas \register_fifo:fifo_data[0][26] (
	.clk(clk),
	.d(datain[26]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data026),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][26] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][26] .power_up = "low";

dffeas \register_fifo:fifo_data[0][27] (
	.clk(clk),
	.d(datain[27]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data027),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][27] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][27] .power_up = "low";

dffeas \register_fifo:fifo_data[0][28] (
	.clk(clk),
	.d(datain[28]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data028),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][28] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][28] .power_up = "low";

dffeas \register_fifo:fifo_data[0][29] (
	.clk(clk),
	.d(datain[29]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data029),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][29] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][29] .power_up = "low";

dffeas \register_fifo:fifo_data[0][30] (
	.clk(clk),
	.d(datain[30]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data030),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][30] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][30] .power_up = "low";

dffeas \register_fifo:fifo_data[0][31] (
	.clk(clk),
	.d(datain[31]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data031),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][31] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][31] .power_up = "low";

dffeas \register_fifo:fifo_data[0][32] (
	.clk(clk),
	.d(datain[32]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data032),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][32] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][32] .power_up = "low";

dffeas \register_fifo:fifo_data[0][33] (
	.clk(clk),
	.d(datain[33]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data033),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][33] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][33] .power_up = "low";

dffeas \register_fifo:fifo_data[0][34] (
	.clk(clk),
	.d(datain[34]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data034),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][34] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][34] .power_up = "low";

dffeas \register_fifo:fifo_data[0][35] (
	.clk(clk),
	.d(datain[35]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data035),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][35] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][35] .power_up = "low";

dffeas \register_fifo:fifo_data[0][7] (
	.clk(clk),
	.d(datain[7]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data07),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][7] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][7] .power_up = "low";

dffeas \register_fifo:fifo_data[0][6] (
	.clk(clk),
	.d(datain[6]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data06),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][6] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][6] .power_up = "low";

dffeas \register_fifo:fifo_data[0][5] (
	.clk(clk),
	.d(datain[5]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data05),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][5] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][5] .power_up = "low";

dffeas \register_fifo:fifo_data[0][4] (
	.clk(clk),
	.d(datain[4]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data04),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][4] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][4] .power_up = "low";

dffeas \register_fifo:fifo_data[0][3] (
	.clk(clk),
	.d(datain[3]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data03),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][3] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][3] .power_up = "low";

dffeas \register_fifo:fifo_data[0][2] (
	.clk(clk),
	.d(datain[2]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data02),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][2] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][2] .power_up = "low";

dffeas \register_fifo:fifo_data[0][1] (
	.clk(clk),
	.d(datain[1]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data01),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][1] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][1] .power_up = "low";

dffeas \register_fifo:fifo_data[0][0] (
	.clk(clk),
	.d(datain[0]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data00),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][0] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][0] .power_up = "low";

endmodule

module cic_auk_dspip_differentiator_2 (
	dout_valid1,
	dout_valid2,
	dout_7,
	dout_8,
	dout_9,
	dout_10,
	dout_11,
	dout_12,
	dout_13,
	dout_14,
	dout_15,
	dout_16,
	dout_17,
	dout_18,
	dout_19,
	dout_20,
	dout_21,
	dout_22,
	dout_23,
	dout_24,
	dout_25,
	dout_26,
	dout_27,
	dout_28,
	dout_29,
	dout_30,
	dout_31,
	dout_32,
	dout_33,
	dout_34,
	dout_6,
	dout_81,
	dout_5,
	dout_91,
	dout_101,
	dout_111,
	dout_121,
	dout_131,
	dout_141,
	dout_151,
	dout_161,
	dout_171,
	dout_181,
	dout_191,
	dout_201,
	dout_211,
	dout_221,
	dout_231,
	dout_241,
	dout_251,
	dout_261,
	dout_271,
	dout_281,
	dout_291,
	dout_301,
	dout_311,
	dout_321,
	dout_331,
	dout_341,
	dout_35,
	dout_71,
	dout_4,
	dout_61,
	dout_3,
	dout_51,
	dout_2,
	dout_41,
	dout_1,
	dout_36,
	dout_210,
	dout_110,
	stall_reg,
	dout_valid3,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	dout_valid1;
input 	dout_valid2;
output 	dout_7;
output 	dout_8;
output 	dout_9;
output 	dout_10;
output 	dout_11;
output 	dout_12;
output 	dout_13;
output 	dout_14;
output 	dout_15;
output 	dout_16;
output 	dout_17;
output 	dout_18;
output 	dout_19;
output 	dout_20;
output 	dout_21;
output 	dout_22;
output 	dout_23;
output 	dout_24;
output 	dout_25;
output 	dout_26;
output 	dout_27;
output 	dout_28;
output 	dout_29;
output 	dout_30;
output 	dout_31;
output 	dout_32;
output 	dout_33;
output 	dout_34;
output 	dout_6;
input 	dout_81;
output 	dout_5;
input 	dout_91;
input 	dout_101;
input 	dout_111;
input 	dout_121;
input 	dout_131;
input 	dout_141;
input 	dout_151;
input 	dout_161;
input 	dout_171;
input 	dout_181;
input 	dout_191;
input 	dout_201;
input 	dout_211;
input 	dout_221;
input 	dout_231;
input 	dout_241;
input 	dout_251;
input 	dout_261;
input 	dout_271;
input 	dout_281;
input 	dout_291;
input 	dout_301;
input 	dout_311;
input 	dout_321;
input 	dout_331;
input 	dout_341;
input 	dout_35;
input 	dout_71;
output 	dout_4;
input 	dout_61;
output 	dout_3;
input 	dout_51;
output 	dout_2;
input 	dout_41;
output 	dout_1;
input 	dout_36;
input 	dout_210;
input 	dout_110;
input 	stall_reg;
input 	dout_valid3;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \glogic:u0|register_fifo:fifo_data[0][7]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][8]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][9]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][10]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][11]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][12]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][13]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][14]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][15]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][16]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][17]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][18]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][19]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][20]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][21]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][22]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][23]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][24]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][25]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][26]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][27]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][28]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][29]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][30]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][31]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][32]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][33]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][34]~q ;
wire \dout~1_combout ;
wire \glogic:u0|register_fifo:fifo_data[0][6]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][5]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][4]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][3]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][2]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][1]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][0]~q ;
wire \resq[0]~138_cout ;
wire \resq[0]~139 ;
wire \resq[1]~134 ;
wire \resq[1]~135 ;
wire \resq[2]~130 ;
wire \resq[2]~131 ;
wire \resq[3]~126 ;
wire \resq[3]~127 ;
wire \resq[4]~122 ;
wire \resq[4]~123 ;
wire \resq[5]~118 ;
wire \resq[5]~119 ;
wire \resq[6]~114 ;
wire \resq[6]~115 ;
wire \resq[7]~1_sumout ;
wire \dout[31]~0_combout ;
wire \resq[7]~2 ;
wire \resq[7]~3 ;
wire \resq[8]~5_sumout ;
wire \resq[8]~6 ;
wire \resq[8]~7 ;
wire \resq[9]~9_sumout ;
wire \resq[9]~10 ;
wire \resq[9]~11 ;
wire \resq[10]~13_sumout ;
wire \resq[10]~14 ;
wire \resq[10]~15 ;
wire \resq[11]~17_sumout ;
wire \resq[11]~18 ;
wire \resq[11]~19 ;
wire \resq[12]~21_sumout ;
wire \resq[12]~22 ;
wire \resq[12]~23 ;
wire \resq[13]~25_sumout ;
wire \resq[13]~26 ;
wire \resq[13]~27 ;
wire \resq[14]~29_sumout ;
wire \resq[14]~30 ;
wire \resq[14]~31 ;
wire \resq[15]~33_sumout ;
wire \resq[15]~34 ;
wire \resq[15]~35 ;
wire \resq[16]~37_sumout ;
wire \resq[16]~38 ;
wire \resq[16]~39 ;
wire \resq[17]~41_sumout ;
wire \resq[17]~42 ;
wire \resq[17]~43 ;
wire \resq[18]~45_sumout ;
wire \resq[18]~46 ;
wire \resq[18]~47 ;
wire \resq[19]~49_sumout ;
wire \resq[19]~50 ;
wire \resq[19]~51 ;
wire \resq[20]~53_sumout ;
wire \resq[20]~54 ;
wire \resq[20]~55 ;
wire \resq[21]~57_sumout ;
wire \resq[21]~58 ;
wire \resq[21]~59 ;
wire \resq[22]~61_sumout ;
wire \resq[22]~62 ;
wire \resq[22]~63 ;
wire \resq[23]~65_sumout ;
wire \resq[23]~66 ;
wire \resq[23]~67 ;
wire \resq[24]~69_sumout ;
wire \resq[24]~70 ;
wire \resq[24]~71 ;
wire \resq[25]~73_sumout ;
wire \resq[25]~74 ;
wire \resq[25]~75 ;
wire \resq[26]~77_sumout ;
wire \resq[26]~78 ;
wire \resq[26]~79 ;
wire \resq[27]~81_sumout ;
wire \resq[27]~82 ;
wire \resq[27]~83 ;
wire \resq[28]~85_sumout ;
wire \resq[28]~86 ;
wire \resq[28]~87 ;
wire \resq[29]~89_sumout ;
wire \resq[29]~90 ;
wire \resq[29]~91 ;
wire \resq[30]~93_sumout ;
wire \resq[30]~94 ;
wire \resq[30]~95 ;
wire \resq[31]~97_sumout ;
wire \resq[31]~98 ;
wire \resq[31]~99 ;
wire \resq[32]~101_sumout ;
wire \resq[32]~102 ;
wire \resq[32]~103 ;
wire \resq[33]~105_sumout ;
wire \resq[33]~106 ;
wire \resq[33]~107 ;
wire \resq[34]~109_sumout ;
wire \resq[6]~113_sumout ;
wire \resq[5]~117_sumout ;
wire \resq[4]~121_sumout ;
wire \resq[3]~125_sumout ;
wire \resq[2]~129_sumout ;
wire \resq[1]~133_sumout ;


cic_auk_dspip_delay_2 \glogic:u0 (
	.datain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,dout_35,dout_341,dout_331,dout_321,dout_311,dout_301,dout_291,dout_281,dout_271,dout_261,dout_251,dout_241,dout_231,dout_221,dout_211,dout_201,dout_191,dout_181,dout_171,dout_161,dout_151,dout_141,dout_131,dout_121,dout_111,dout_101,dout_91,
dout_81,dout_71,dout_61,dout_51,dout_41,dout_36,dout_210,dout_110}),
	.register_fifofifo_data07(\glogic:u0|register_fifo:fifo_data[0][7]~q ),
	.register_fifofifo_data08(\glogic:u0|register_fifo:fifo_data[0][8]~q ),
	.register_fifofifo_data09(\glogic:u0|register_fifo:fifo_data[0][9]~q ),
	.register_fifofifo_data010(\glogic:u0|register_fifo:fifo_data[0][10]~q ),
	.register_fifofifo_data011(\glogic:u0|register_fifo:fifo_data[0][11]~q ),
	.register_fifofifo_data012(\glogic:u0|register_fifo:fifo_data[0][12]~q ),
	.register_fifofifo_data013(\glogic:u0|register_fifo:fifo_data[0][13]~q ),
	.register_fifofifo_data014(\glogic:u0|register_fifo:fifo_data[0][14]~q ),
	.register_fifofifo_data015(\glogic:u0|register_fifo:fifo_data[0][15]~q ),
	.register_fifofifo_data016(\glogic:u0|register_fifo:fifo_data[0][16]~q ),
	.register_fifofifo_data017(\glogic:u0|register_fifo:fifo_data[0][17]~q ),
	.register_fifofifo_data018(\glogic:u0|register_fifo:fifo_data[0][18]~q ),
	.register_fifofifo_data019(\glogic:u0|register_fifo:fifo_data[0][19]~q ),
	.register_fifofifo_data020(\glogic:u0|register_fifo:fifo_data[0][20]~q ),
	.register_fifofifo_data021(\glogic:u0|register_fifo:fifo_data[0][21]~q ),
	.register_fifofifo_data022(\glogic:u0|register_fifo:fifo_data[0][22]~q ),
	.register_fifofifo_data023(\glogic:u0|register_fifo:fifo_data[0][23]~q ),
	.register_fifofifo_data024(\glogic:u0|register_fifo:fifo_data[0][24]~q ),
	.register_fifofifo_data025(\glogic:u0|register_fifo:fifo_data[0][25]~q ),
	.register_fifofifo_data026(\glogic:u0|register_fifo:fifo_data[0][26]~q ),
	.register_fifofifo_data027(\glogic:u0|register_fifo:fifo_data[0][27]~q ),
	.register_fifofifo_data028(\glogic:u0|register_fifo:fifo_data[0][28]~q ),
	.register_fifofifo_data029(\glogic:u0|register_fifo:fifo_data[0][29]~q ),
	.register_fifofifo_data030(\glogic:u0|register_fifo:fifo_data[0][30]~q ),
	.register_fifofifo_data031(\glogic:u0|register_fifo:fifo_data[0][31]~q ),
	.register_fifofifo_data032(\glogic:u0|register_fifo:fifo_data[0][32]~q ),
	.register_fifofifo_data033(\glogic:u0|register_fifo:fifo_data[0][33]~q ),
	.register_fifofifo_data034(\glogic:u0|register_fifo:fifo_data[0][34]~q ),
	.enable(\dout~1_combout ),
	.register_fifofifo_data06(\glogic:u0|register_fifo:fifo_data[0][6]~q ),
	.register_fifofifo_data05(\glogic:u0|register_fifo:fifo_data[0][5]~q ),
	.register_fifofifo_data04(\glogic:u0|register_fifo:fifo_data[0][4]~q ),
	.register_fifofifo_data03(\glogic:u0|register_fifo:fifo_data[0][3]~q ),
	.register_fifofifo_data02(\glogic:u0|register_fifo:fifo_data[0][2]~q ),
	.register_fifofifo_data01(\glogic:u0|register_fifo:fifo_data[0][1]~q ),
	.register_fifofifo_data00(\glogic:u0|register_fifo:fifo_data[0][0]~q ),
	.clk(clk),
	.reset(reset_n));

arriav_lcell_comb \dout~1 (
	.dataa(!stall_reg),
	.datab(!dout_valid2),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dout~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dout~1 .extended_lut = "off";
defparam \dout~1 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \dout~1 .shared_arith = "off";

dffeas dout_valid(
	.clk(clk),
	.d(dout_valid2),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(dout_valid3),
	.q(dout_valid1),
	.prn(vcc));
defparam dout_valid.is_wysiwyg = "true";
defparam dout_valid.power_up = "low";

dffeas \dout[7] (
	.clk(clk),
	.d(\resq[7]~1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[31]~0_combout ),
	.q(dout_7),
	.prn(vcc));
defparam \dout[7] .is_wysiwyg = "true";
defparam \dout[7] .power_up = "low";

dffeas \dout[8] (
	.clk(clk),
	.d(\resq[8]~5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[31]~0_combout ),
	.q(dout_8),
	.prn(vcc));
defparam \dout[8] .is_wysiwyg = "true";
defparam \dout[8] .power_up = "low";

dffeas \dout[9] (
	.clk(clk),
	.d(\resq[9]~9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[31]~0_combout ),
	.q(dout_9),
	.prn(vcc));
defparam \dout[9] .is_wysiwyg = "true";
defparam \dout[9] .power_up = "low";

dffeas \dout[10] (
	.clk(clk),
	.d(\resq[10]~13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[31]~0_combout ),
	.q(dout_10),
	.prn(vcc));
defparam \dout[10] .is_wysiwyg = "true";
defparam \dout[10] .power_up = "low";

dffeas \dout[11] (
	.clk(clk),
	.d(\resq[11]~17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[31]~0_combout ),
	.q(dout_11),
	.prn(vcc));
defparam \dout[11] .is_wysiwyg = "true";
defparam \dout[11] .power_up = "low";

dffeas \dout[12] (
	.clk(clk),
	.d(\resq[12]~21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[31]~0_combout ),
	.q(dout_12),
	.prn(vcc));
defparam \dout[12] .is_wysiwyg = "true";
defparam \dout[12] .power_up = "low";

dffeas \dout[13] (
	.clk(clk),
	.d(\resq[13]~25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[31]~0_combout ),
	.q(dout_13),
	.prn(vcc));
defparam \dout[13] .is_wysiwyg = "true";
defparam \dout[13] .power_up = "low";

dffeas \dout[14] (
	.clk(clk),
	.d(\resq[14]~29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[31]~0_combout ),
	.q(dout_14),
	.prn(vcc));
defparam \dout[14] .is_wysiwyg = "true";
defparam \dout[14] .power_up = "low";

dffeas \dout[15] (
	.clk(clk),
	.d(\resq[15]~33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[31]~0_combout ),
	.q(dout_15),
	.prn(vcc));
defparam \dout[15] .is_wysiwyg = "true";
defparam \dout[15] .power_up = "low";

dffeas \dout[16] (
	.clk(clk),
	.d(\resq[16]~37_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[31]~0_combout ),
	.q(dout_16),
	.prn(vcc));
defparam \dout[16] .is_wysiwyg = "true";
defparam \dout[16] .power_up = "low";

dffeas \dout[17] (
	.clk(clk),
	.d(\resq[17]~41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[31]~0_combout ),
	.q(dout_17),
	.prn(vcc));
defparam \dout[17] .is_wysiwyg = "true";
defparam \dout[17] .power_up = "low";

dffeas \dout[18] (
	.clk(clk),
	.d(\resq[18]~45_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[31]~0_combout ),
	.q(dout_18),
	.prn(vcc));
defparam \dout[18] .is_wysiwyg = "true";
defparam \dout[18] .power_up = "low";

dffeas \dout[19] (
	.clk(clk),
	.d(\resq[19]~49_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[31]~0_combout ),
	.q(dout_19),
	.prn(vcc));
defparam \dout[19] .is_wysiwyg = "true";
defparam \dout[19] .power_up = "low";

dffeas \dout[20] (
	.clk(clk),
	.d(\resq[20]~53_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[31]~0_combout ),
	.q(dout_20),
	.prn(vcc));
defparam \dout[20] .is_wysiwyg = "true";
defparam \dout[20] .power_up = "low";

dffeas \dout[21] (
	.clk(clk),
	.d(\resq[21]~57_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[31]~0_combout ),
	.q(dout_21),
	.prn(vcc));
defparam \dout[21] .is_wysiwyg = "true";
defparam \dout[21] .power_up = "low";

dffeas \dout[22] (
	.clk(clk),
	.d(\resq[22]~61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[31]~0_combout ),
	.q(dout_22),
	.prn(vcc));
defparam \dout[22] .is_wysiwyg = "true";
defparam \dout[22] .power_up = "low";

dffeas \dout[23] (
	.clk(clk),
	.d(\resq[23]~65_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[31]~0_combout ),
	.q(dout_23),
	.prn(vcc));
defparam \dout[23] .is_wysiwyg = "true";
defparam \dout[23] .power_up = "low";

dffeas \dout[24] (
	.clk(clk),
	.d(\resq[24]~69_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[31]~0_combout ),
	.q(dout_24),
	.prn(vcc));
defparam \dout[24] .is_wysiwyg = "true";
defparam \dout[24] .power_up = "low";

dffeas \dout[25] (
	.clk(clk),
	.d(\resq[25]~73_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[31]~0_combout ),
	.q(dout_25),
	.prn(vcc));
defparam \dout[25] .is_wysiwyg = "true";
defparam \dout[25] .power_up = "low";

dffeas \dout[26] (
	.clk(clk),
	.d(\resq[26]~77_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[31]~0_combout ),
	.q(dout_26),
	.prn(vcc));
defparam \dout[26] .is_wysiwyg = "true";
defparam \dout[26] .power_up = "low";

dffeas \dout[27] (
	.clk(clk),
	.d(\resq[27]~81_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[31]~0_combout ),
	.q(dout_27),
	.prn(vcc));
defparam \dout[27] .is_wysiwyg = "true";
defparam \dout[27] .power_up = "low";

dffeas \dout[28] (
	.clk(clk),
	.d(\resq[28]~85_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[31]~0_combout ),
	.q(dout_28),
	.prn(vcc));
defparam \dout[28] .is_wysiwyg = "true";
defparam \dout[28] .power_up = "low";

dffeas \dout[29] (
	.clk(clk),
	.d(\resq[29]~89_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[31]~0_combout ),
	.q(dout_29),
	.prn(vcc));
defparam \dout[29] .is_wysiwyg = "true";
defparam \dout[29] .power_up = "low";

dffeas \dout[30] (
	.clk(clk),
	.d(\resq[30]~93_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[31]~0_combout ),
	.q(dout_30),
	.prn(vcc));
defparam \dout[30] .is_wysiwyg = "true";
defparam \dout[30] .power_up = "low";

dffeas \dout[31] (
	.clk(clk),
	.d(\resq[31]~97_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[31]~0_combout ),
	.q(dout_31),
	.prn(vcc));
defparam \dout[31] .is_wysiwyg = "true";
defparam \dout[31] .power_up = "low";

dffeas \dout[32] (
	.clk(clk),
	.d(\resq[32]~101_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[31]~0_combout ),
	.q(dout_32),
	.prn(vcc));
defparam \dout[32] .is_wysiwyg = "true";
defparam \dout[32] .power_up = "low";

dffeas \dout[33] (
	.clk(clk),
	.d(\resq[33]~105_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[31]~0_combout ),
	.q(dout_33),
	.prn(vcc));
defparam \dout[33] .is_wysiwyg = "true";
defparam \dout[33] .power_up = "low";

dffeas \dout[34] (
	.clk(clk),
	.d(\resq[34]~109_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[31]~0_combout ),
	.q(dout_34),
	.prn(vcc));
defparam \dout[34] .is_wysiwyg = "true";
defparam \dout[34] .power_up = "low";

dffeas \dout[6] (
	.clk(clk),
	.d(\resq[6]~113_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[31]~0_combout ),
	.q(dout_6),
	.prn(vcc));
defparam \dout[6] .is_wysiwyg = "true";
defparam \dout[6] .power_up = "low";

dffeas \dout[5] (
	.clk(clk),
	.d(\resq[5]~117_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[31]~0_combout ),
	.q(dout_5),
	.prn(vcc));
defparam \dout[5] .is_wysiwyg = "true";
defparam \dout[5] .power_up = "low";

dffeas \dout[4] (
	.clk(clk),
	.d(\resq[4]~121_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[31]~0_combout ),
	.q(dout_4),
	.prn(vcc));
defparam \dout[4] .is_wysiwyg = "true";
defparam \dout[4] .power_up = "low";

dffeas \dout[3] (
	.clk(clk),
	.d(\resq[3]~125_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[31]~0_combout ),
	.q(dout_3),
	.prn(vcc));
defparam \dout[3] .is_wysiwyg = "true";
defparam \dout[3] .power_up = "low";

dffeas \dout[2] (
	.clk(clk),
	.d(\resq[2]~129_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[31]~0_combout ),
	.q(dout_2),
	.prn(vcc));
defparam \dout[2] .is_wysiwyg = "true";
defparam \dout[2] .power_up = "low";

dffeas \dout[1] (
	.clk(clk),
	.d(\resq[1]~133_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[31]~0_combout ),
	.q(dout_1),
	.prn(vcc));
defparam \dout[1] .is_wysiwyg = "true";
defparam \dout[1] .power_up = "low";

arriav_lcell_comb \resq[0]~138 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][0]~q ),
	.datad(!dout_110),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\resq[0]~138_cout ),
	.shareout(\resq[0]~139 ));
defparam \resq[0]~138 .extended_lut = "off";
defparam \resq[0]~138 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[0]~138 .shared_arith = "on";

arriav_lcell_comb \resq[1]~133 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][1]~q ),
	.datad(!dout_210),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[0]~138_cout ),
	.sharein(\resq[0]~139 ),
	.combout(),
	.sumout(\resq[1]~133_sumout ),
	.cout(\resq[1]~134 ),
	.shareout(\resq[1]~135 ));
defparam \resq[1]~133 .extended_lut = "off";
defparam \resq[1]~133 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[1]~133 .shared_arith = "on";

arriav_lcell_comb \resq[2]~129 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][2]~q ),
	.datad(!dout_36),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[1]~134 ),
	.sharein(\resq[1]~135 ),
	.combout(),
	.sumout(\resq[2]~129_sumout ),
	.cout(\resq[2]~130 ),
	.shareout(\resq[2]~131 ));
defparam \resq[2]~129 .extended_lut = "off";
defparam \resq[2]~129 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[2]~129 .shared_arith = "on";

arriav_lcell_comb \resq[3]~125 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][3]~q ),
	.datad(!dout_41),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[2]~130 ),
	.sharein(\resq[2]~131 ),
	.combout(),
	.sumout(\resq[3]~125_sumout ),
	.cout(\resq[3]~126 ),
	.shareout(\resq[3]~127 ));
defparam \resq[3]~125 .extended_lut = "off";
defparam \resq[3]~125 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[3]~125 .shared_arith = "on";

arriav_lcell_comb \resq[4]~121 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][4]~q ),
	.datad(!dout_51),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[3]~126 ),
	.sharein(\resq[3]~127 ),
	.combout(),
	.sumout(\resq[4]~121_sumout ),
	.cout(\resq[4]~122 ),
	.shareout(\resq[4]~123 ));
defparam \resq[4]~121 .extended_lut = "off";
defparam \resq[4]~121 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[4]~121 .shared_arith = "on";

arriav_lcell_comb \resq[5]~117 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][5]~q ),
	.datad(!dout_61),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[4]~122 ),
	.sharein(\resq[4]~123 ),
	.combout(),
	.sumout(\resq[5]~117_sumout ),
	.cout(\resq[5]~118 ),
	.shareout(\resq[5]~119 ));
defparam \resq[5]~117 .extended_lut = "off";
defparam \resq[5]~117 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[5]~117 .shared_arith = "on";

arriav_lcell_comb \resq[6]~113 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][6]~q ),
	.datad(!dout_71),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[5]~118 ),
	.sharein(\resq[5]~119 ),
	.combout(),
	.sumout(\resq[6]~113_sumout ),
	.cout(\resq[6]~114 ),
	.shareout(\resq[6]~115 ));
defparam \resq[6]~113 .extended_lut = "off";
defparam \resq[6]~113 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[6]~113 .shared_arith = "on";

arriav_lcell_comb \resq[7]~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][7]~q ),
	.datad(!dout_81),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[6]~114 ),
	.sharein(\resq[6]~115 ),
	.combout(),
	.sumout(\resq[7]~1_sumout ),
	.cout(\resq[7]~2 ),
	.shareout(\resq[7]~3 ));
defparam \resq[7]~1 .extended_lut = "off";
defparam \resq[7]~1 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[7]~1 .shared_arith = "on";

arriav_lcell_comb \dout[31]~0 (
	.dataa(!reset_n),
	.datab(!stall_reg),
	.datac(!dout_valid2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dout[31]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dout[31]~0 .extended_lut = "off";
defparam \dout[31]~0 .lut_mask = 64'hEFEFEFEFEFEFEFEF;
defparam \dout[31]~0 .shared_arith = "off";

arriav_lcell_comb \resq[8]~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][8]~q ),
	.datad(!dout_91),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[7]~2 ),
	.sharein(\resq[7]~3 ),
	.combout(),
	.sumout(\resq[8]~5_sumout ),
	.cout(\resq[8]~6 ),
	.shareout(\resq[8]~7 ));
defparam \resq[8]~5 .extended_lut = "off";
defparam \resq[8]~5 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[8]~5 .shared_arith = "on";

arriav_lcell_comb \resq[9]~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][9]~q ),
	.datad(!dout_101),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[8]~6 ),
	.sharein(\resq[8]~7 ),
	.combout(),
	.sumout(\resq[9]~9_sumout ),
	.cout(\resq[9]~10 ),
	.shareout(\resq[9]~11 ));
defparam \resq[9]~9 .extended_lut = "off";
defparam \resq[9]~9 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[9]~9 .shared_arith = "on";

arriav_lcell_comb \resq[10]~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][10]~q ),
	.datad(!dout_111),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[9]~10 ),
	.sharein(\resq[9]~11 ),
	.combout(),
	.sumout(\resq[10]~13_sumout ),
	.cout(\resq[10]~14 ),
	.shareout(\resq[10]~15 ));
defparam \resq[10]~13 .extended_lut = "off";
defparam \resq[10]~13 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[10]~13 .shared_arith = "on";

arriav_lcell_comb \resq[11]~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][11]~q ),
	.datad(!dout_121),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[10]~14 ),
	.sharein(\resq[10]~15 ),
	.combout(),
	.sumout(\resq[11]~17_sumout ),
	.cout(\resq[11]~18 ),
	.shareout(\resq[11]~19 ));
defparam \resq[11]~17 .extended_lut = "off";
defparam \resq[11]~17 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[11]~17 .shared_arith = "on";

arriav_lcell_comb \resq[12]~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][12]~q ),
	.datad(!dout_131),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[11]~18 ),
	.sharein(\resq[11]~19 ),
	.combout(),
	.sumout(\resq[12]~21_sumout ),
	.cout(\resq[12]~22 ),
	.shareout(\resq[12]~23 ));
defparam \resq[12]~21 .extended_lut = "off";
defparam \resq[12]~21 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[12]~21 .shared_arith = "on";

arriav_lcell_comb \resq[13]~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][13]~q ),
	.datad(!dout_141),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[12]~22 ),
	.sharein(\resq[12]~23 ),
	.combout(),
	.sumout(\resq[13]~25_sumout ),
	.cout(\resq[13]~26 ),
	.shareout(\resq[13]~27 ));
defparam \resq[13]~25 .extended_lut = "off";
defparam \resq[13]~25 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[13]~25 .shared_arith = "on";

arriav_lcell_comb \resq[14]~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][14]~q ),
	.datad(!dout_151),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[13]~26 ),
	.sharein(\resq[13]~27 ),
	.combout(),
	.sumout(\resq[14]~29_sumout ),
	.cout(\resq[14]~30 ),
	.shareout(\resq[14]~31 ));
defparam \resq[14]~29 .extended_lut = "off";
defparam \resq[14]~29 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[14]~29 .shared_arith = "on";

arriav_lcell_comb \resq[15]~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][15]~q ),
	.datad(!dout_161),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[14]~30 ),
	.sharein(\resq[14]~31 ),
	.combout(),
	.sumout(\resq[15]~33_sumout ),
	.cout(\resq[15]~34 ),
	.shareout(\resq[15]~35 ));
defparam \resq[15]~33 .extended_lut = "off";
defparam \resq[15]~33 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[15]~33 .shared_arith = "on";

arriav_lcell_comb \resq[16]~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][16]~q ),
	.datad(!dout_171),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[15]~34 ),
	.sharein(\resq[15]~35 ),
	.combout(),
	.sumout(\resq[16]~37_sumout ),
	.cout(\resq[16]~38 ),
	.shareout(\resq[16]~39 ));
defparam \resq[16]~37 .extended_lut = "off";
defparam \resq[16]~37 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[16]~37 .shared_arith = "on";

arriav_lcell_comb \resq[17]~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][17]~q ),
	.datad(!dout_181),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[16]~38 ),
	.sharein(\resq[16]~39 ),
	.combout(),
	.sumout(\resq[17]~41_sumout ),
	.cout(\resq[17]~42 ),
	.shareout(\resq[17]~43 ));
defparam \resq[17]~41 .extended_lut = "off";
defparam \resq[17]~41 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[17]~41 .shared_arith = "on";

arriav_lcell_comb \resq[18]~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][18]~q ),
	.datad(!dout_191),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[17]~42 ),
	.sharein(\resq[17]~43 ),
	.combout(),
	.sumout(\resq[18]~45_sumout ),
	.cout(\resq[18]~46 ),
	.shareout(\resq[18]~47 ));
defparam \resq[18]~45 .extended_lut = "off";
defparam \resq[18]~45 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[18]~45 .shared_arith = "on";

arriav_lcell_comb \resq[19]~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][19]~q ),
	.datad(!dout_201),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[18]~46 ),
	.sharein(\resq[18]~47 ),
	.combout(),
	.sumout(\resq[19]~49_sumout ),
	.cout(\resq[19]~50 ),
	.shareout(\resq[19]~51 ));
defparam \resq[19]~49 .extended_lut = "off";
defparam \resq[19]~49 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[19]~49 .shared_arith = "on";

arriav_lcell_comb \resq[20]~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][20]~q ),
	.datad(!dout_211),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[19]~50 ),
	.sharein(\resq[19]~51 ),
	.combout(),
	.sumout(\resq[20]~53_sumout ),
	.cout(\resq[20]~54 ),
	.shareout(\resq[20]~55 ));
defparam \resq[20]~53 .extended_lut = "off";
defparam \resq[20]~53 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[20]~53 .shared_arith = "on";

arriav_lcell_comb \resq[21]~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][21]~q ),
	.datad(!dout_221),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[20]~54 ),
	.sharein(\resq[20]~55 ),
	.combout(),
	.sumout(\resq[21]~57_sumout ),
	.cout(\resq[21]~58 ),
	.shareout(\resq[21]~59 ));
defparam \resq[21]~57 .extended_lut = "off";
defparam \resq[21]~57 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[21]~57 .shared_arith = "on";

arriav_lcell_comb \resq[22]~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][22]~q ),
	.datad(!dout_231),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[21]~58 ),
	.sharein(\resq[21]~59 ),
	.combout(),
	.sumout(\resq[22]~61_sumout ),
	.cout(\resq[22]~62 ),
	.shareout(\resq[22]~63 ));
defparam \resq[22]~61 .extended_lut = "off";
defparam \resq[22]~61 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[22]~61 .shared_arith = "on";

arriav_lcell_comb \resq[23]~65 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][23]~q ),
	.datad(!dout_241),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[22]~62 ),
	.sharein(\resq[22]~63 ),
	.combout(),
	.sumout(\resq[23]~65_sumout ),
	.cout(\resq[23]~66 ),
	.shareout(\resq[23]~67 ));
defparam \resq[23]~65 .extended_lut = "off";
defparam \resq[23]~65 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[23]~65 .shared_arith = "on";

arriav_lcell_comb \resq[24]~69 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][24]~q ),
	.datad(!dout_251),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[23]~66 ),
	.sharein(\resq[23]~67 ),
	.combout(),
	.sumout(\resq[24]~69_sumout ),
	.cout(\resq[24]~70 ),
	.shareout(\resq[24]~71 ));
defparam \resq[24]~69 .extended_lut = "off";
defparam \resq[24]~69 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[24]~69 .shared_arith = "on";

arriav_lcell_comb \resq[25]~73 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][25]~q ),
	.datad(!dout_261),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[24]~70 ),
	.sharein(\resq[24]~71 ),
	.combout(),
	.sumout(\resq[25]~73_sumout ),
	.cout(\resq[25]~74 ),
	.shareout(\resq[25]~75 ));
defparam \resq[25]~73 .extended_lut = "off";
defparam \resq[25]~73 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[25]~73 .shared_arith = "on";

arriav_lcell_comb \resq[26]~77 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][26]~q ),
	.datad(!dout_271),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[25]~74 ),
	.sharein(\resq[25]~75 ),
	.combout(),
	.sumout(\resq[26]~77_sumout ),
	.cout(\resq[26]~78 ),
	.shareout(\resq[26]~79 ));
defparam \resq[26]~77 .extended_lut = "off";
defparam \resq[26]~77 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[26]~77 .shared_arith = "on";

arriav_lcell_comb \resq[27]~81 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][27]~q ),
	.datad(!dout_281),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[26]~78 ),
	.sharein(\resq[26]~79 ),
	.combout(),
	.sumout(\resq[27]~81_sumout ),
	.cout(\resq[27]~82 ),
	.shareout(\resq[27]~83 ));
defparam \resq[27]~81 .extended_lut = "off";
defparam \resq[27]~81 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[27]~81 .shared_arith = "on";

arriav_lcell_comb \resq[28]~85 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][28]~q ),
	.datad(!dout_291),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[27]~82 ),
	.sharein(\resq[27]~83 ),
	.combout(),
	.sumout(\resq[28]~85_sumout ),
	.cout(\resq[28]~86 ),
	.shareout(\resq[28]~87 ));
defparam \resq[28]~85 .extended_lut = "off";
defparam \resq[28]~85 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[28]~85 .shared_arith = "on";

arriav_lcell_comb \resq[29]~89 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][29]~q ),
	.datad(!dout_301),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[28]~86 ),
	.sharein(\resq[28]~87 ),
	.combout(),
	.sumout(\resq[29]~89_sumout ),
	.cout(\resq[29]~90 ),
	.shareout(\resq[29]~91 ));
defparam \resq[29]~89 .extended_lut = "off";
defparam \resq[29]~89 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[29]~89 .shared_arith = "on";

arriav_lcell_comb \resq[30]~93 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][30]~q ),
	.datad(!dout_311),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[29]~90 ),
	.sharein(\resq[29]~91 ),
	.combout(),
	.sumout(\resq[30]~93_sumout ),
	.cout(\resq[30]~94 ),
	.shareout(\resq[30]~95 ));
defparam \resq[30]~93 .extended_lut = "off";
defparam \resq[30]~93 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[30]~93 .shared_arith = "on";

arriav_lcell_comb \resq[31]~97 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][31]~q ),
	.datad(!dout_321),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[30]~94 ),
	.sharein(\resq[30]~95 ),
	.combout(),
	.sumout(\resq[31]~97_sumout ),
	.cout(\resq[31]~98 ),
	.shareout(\resq[31]~99 ));
defparam \resq[31]~97 .extended_lut = "off";
defparam \resq[31]~97 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[31]~97 .shared_arith = "on";

arriav_lcell_comb \resq[32]~101 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][32]~q ),
	.datad(!dout_331),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[31]~98 ),
	.sharein(\resq[31]~99 ),
	.combout(),
	.sumout(\resq[32]~101_sumout ),
	.cout(\resq[32]~102 ),
	.shareout(\resq[32]~103 ));
defparam \resq[32]~101 .extended_lut = "off";
defparam \resq[32]~101 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[32]~101 .shared_arith = "on";

arriav_lcell_comb \resq[33]~105 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][33]~q ),
	.datad(!dout_341),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[32]~102 ),
	.sharein(\resq[32]~103 ),
	.combout(),
	.sumout(\resq[33]~105_sumout ),
	.cout(\resq[33]~106 ),
	.shareout(\resq[33]~107 ));
defparam \resq[33]~105 .extended_lut = "off";
defparam \resq[33]~105 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[33]~105 .shared_arith = "on";

arriav_lcell_comb \resq[34]~109 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][34]~q ),
	.datad(!dout_35),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[33]~106 ),
	.sharein(\resq[33]~107 ),
	.combout(),
	.sumout(\resq[34]~109_sumout ),
	.cout(),
	.shareout());
defparam \resq[34]~109 .extended_lut = "off";
defparam \resq[34]~109 .lut_mask = 64'h0000000000000FF0;
defparam \resq[34]~109 .shared_arith = "on";

endmodule

module cic_auk_dspip_delay_2 (
	datain,
	register_fifofifo_data07,
	register_fifofifo_data08,
	register_fifofifo_data09,
	register_fifofifo_data010,
	register_fifofifo_data011,
	register_fifofifo_data012,
	register_fifofifo_data013,
	register_fifofifo_data014,
	register_fifofifo_data015,
	register_fifofifo_data016,
	register_fifofifo_data017,
	register_fifofifo_data018,
	register_fifofifo_data019,
	register_fifofifo_data020,
	register_fifofifo_data021,
	register_fifofifo_data022,
	register_fifofifo_data023,
	register_fifofifo_data024,
	register_fifofifo_data025,
	register_fifofifo_data026,
	register_fifofifo_data027,
	register_fifofifo_data028,
	register_fifofifo_data029,
	register_fifofifo_data030,
	register_fifofifo_data031,
	register_fifofifo_data032,
	register_fifofifo_data033,
	register_fifofifo_data034,
	enable,
	register_fifofifo_data06,
	register_fifofifo_data05,
	register_fifofifo_data04,
	register_fifofifo_data03,
	register_fifofifo_data02,
	register_fifofifo_data01,
	register_fifofifo_data00,
	clk,
	reset)/* synthesis synthesis_greybox=1 */;
input 	[46:0] datain;
output 	register_fifofifo_data07;
output 	register_fifofifo_data08;
output 	register_fifofifo_data09;
output 	register_fifofifo_data010;
output 	register_fifofifo_data011;
output 	register_fifofifo_data012;
output 	register_fifofifo_data013;
output 	register_fifofifo_data014;
output 	register_fifofifo_data015;
output 	register_fifofifo_data016;
output 	register_fifofifo_data017;
output 	register_fifofifo_data018;
output 	register_fifofifo_data019;
output 	register_fifofifo_data020;
output 	register_fifofifo_data021;
output 	register_fifofifo_data022;
output 	register_fifofifo_data023;
output 	register_fifofifo_data024;
output 	register_fifofifo_data025;
output 	register_fifofifo_data026;
output 	register_fifofifo_data027;
output 	register_fifofifo_data028;
output 	register_fifofifo_data029;
output 	register_fifofifo_data030;
output 	register_fifofifo_data031;
output 	register_fifofifo_data032;
output 	register_fifofifo_data033;
output 	register_fifofifo_data034;
input 	enable;
output 	register_fifofifo_data06;
output 	register_fifofifo_data05;
output 	register_fifofifo_data04;
output 	register_fifofifo_data03;
output 	register_fifofifo_data02;
output 	register_fifofifo_data01;
output 	register_fifofifo_data00;
input 	clk;
input 	reset;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \register_fifo:fifo_data[0][7] (
	.clk(clk),
	.d(datain[7]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data07),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][7] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][7] .power_up = "low";

dffeas \register_fifo:fifo_data[0][8] (
	.clk(clk),
	.d(datain[8]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data08),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][8] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][8] .power_up = "low";

dffeas \register_fifo:fifo_data[0][9] (
	.clk(clk),
	.d(datain[9]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data09),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][9] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][9] .power_up = "low";

dffeas \register_fifo:fifo_data[0][10] (
	.clk(clk),
	.d(datain[10]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data010),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][10] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][10] .power_up = "low";

dffeas \register_fifo:fifo_data[0][11] (
	.clk(clk),
	.d(datain[11]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data011),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][11] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][11] .power_up = "low";

dffeas \register_fifo:fifo_data[0][12] (
	.clk(clk),
	.d(datain[12]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data012),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][12] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][12] .power_up = "low";

dffeas \register_fifo:fifo_data[0][13] (
	.clk(clk),
	.d(datain[13]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data013),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][13] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][13] .power_up = "low";

dffeas \register_fifo:fifo_data[0][14] (
	.clk(clk),
	.d(datain[14]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data014),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][14] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][14] .power_up = "low";

dffeas \register_fifo:fifo_data[0][15] (
	.clk(clk),
	.d(datain[15]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data015),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][15] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][15] .power_up = "low";

dffeas \register_fifo:fifo_data[0][16] (
	.clk(clk),
	.d(datain[16]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data016),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][16] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][16] .power_up = "low";

dffeas \register_fifo:fifo_data[0][17] (
	.clk(clk),
	.d(datain[17]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data017),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][17] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][17] .power_up = "low";

dffeas \register_fifo:fifo_data[0][18] (
	.clk(clk),
	.d(datain[18]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data018),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][18] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][18] .power_up = "low";

dffeas \register_fifo:fifo_data[0][19] (
	.clk(clk),
	.d(datain[19]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data019),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][19] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][19] .power_up = "low";

dffeas \register_fifo:fifo_data[0][20] (
	.clk(clk),
	.d(datain[20]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data020),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][20] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][20] .power_up = "low";

dffeas \register_fifo:fifo_data[0][21] (
	.clk(clk),
	.d(datain[21]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data021),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][21] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][21] .power_up = "low";

dffeas \register_fifo:fifo_data[0][22] (
	.clk(clk),
	.d(datain[22]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data022),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][22] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][22] .power_up = "low";

dffeas \register_fifo:fifo_data[0][23] (
	.clk(clk),
	.d(datain[23]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data023),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][23] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][23] .power_up = "low";

dffeas \register_fifo:fifo_data[0][24] (
	.clk(clk),
	.d(datain[24]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data024),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][24] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][24] .power_up = "low";

dffeas \register_fifo:fifo_data[0][25] (
	.clk(clk),
	.d(datain[25]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data025),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][25] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][25] .power_up = "low";

dffeas \register_fifo:fifo_data[0][26] (
	.clk(clk),
	.d(datain[26]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data026),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][26] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][26] .power_up = "low";

dffeas \register_fifo:fifo_data[0][27] (
	.clk(clk),
	.d(datain[27]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data027),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][27] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][27] .power_up = "low";

dffeas \register_fifo:fifo_data[0][28] (
	.clk(clk),
	.d(datain[28]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data028),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][28] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][28] .power_up = "low";

dffeas \register_fifo:fifo_data[0][29] (
	.clk(clk),
	.d(datain[29]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data029),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][29] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][29] .power_up = "low";

dffeas \register_fifo:fifo_data[0][30] (
	.clk(clk),
	.d(datain[30]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data030),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][30] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][30] .power_up = "low";

dffeas \register_fifo:fifo_data[0][31] (
	.clk(clk),
	.d(datain[31]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data031),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][31] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][31] .power_up = "low";

dffeas \register_fifo:fifo_data[0][32] (
	.clk(clk),
	.d(datain[32]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data032),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][32] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][32] .power_up = "low";

dffeas \register_fifo:fifo_data[0][33] (
	.clk(clk),
	.d(datain[33]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data033),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][33] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][33] .power_up = "low";

dffeas \register_fifo:fifo_data[0][34] (
	.clk(clk),
	.d(datain[34]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data034),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][34] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][34] .power_up = "low";

dffeas \register_fifo:fifo_data[0][6] (
	.clk(clk),
	.d(datain[6]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data06),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][6] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][6] .power_up = "low";

dffeas \register_fifo:fifo_data[0][5] (
	.clk(clk),
	.d(datain[5]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data05),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][5] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][5] .power_up = "low";

dffeas \register_fifo:fifo_data[0][4] (
	.clk(clk),
	.d(datain[4]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data04),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][4] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][4] .power_up = "low";

dffeas \register_fifo:fifo_data[0][3] (
	.clk(clk),
	.d(datain[3]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data03),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][3] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][3] .power_up = "low";

dffeas \register_fifo:fifo_data[0][2] (
	.clk(clk),
	.d(datain[2]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data02),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][2] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][2] .power_up = "low";

dffeas \register_fifo:fifo_data[0][1] (
	.clk(clk),
	.d(datain[1]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data01),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][1] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][1] .power_up = "low";

dffeas \register_fifo:fifo_data[0][0] (
	.clk(clk),
	.d(datain[0]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data00),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][0] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][0] .power_up = "low";

endmodule

module cic_auk_dspip_differentiator_3 (
	dout_valid1,
	dout_valid2,
	dout_6,
	dout_7,
	dout_8,
	dout_9,
	dout_10,
	dout_11,
	dout_12,
	dout_13,
	dout_14,
	dout_15,
	dout_16,
	dout_17,
	dout_18,
	dout_19,
	dout_20,
	dout_21,
	dout_22,
	dout_23,
	dout_24,
	dout_25,
	dout_26,
	dout_27,
	dout_28,
	dout_29,
	dout_30,
	dout_31,
	dout_32,
	dout_33,
	dout_5,
	dout_71,
	dout_4,
	dout_81,
	dout_91,
	dout_101,
	dout_111,
	dout_121,
	dout_131,
	dout_141,
	dout_151,
	dout_161,
	dout_171,
	dout_181,
	dout_191,
	dout_201,
	dout_211,
	dout_221,
	dout_231,
	dout_241,
	dout_251,
	dout_261,
	dout_271,
	dout_281,
	dout_291,
	dout_301,
	dout_311,
	dout_321,
	dout_331,
	dout_34,
	dout_61,
	dout_3,
	dout_51,
	dout_2,
	dout_41,
	dout_1,
	dout_35,
	dout_0,
	dout_210,
	dout_110,
	stall_reg,
	dout_valid3,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	dout_valid1;
input 	dout_valid2;
output 	dout_6;
output 	dout_7;
output 	dout_8;
output 	dout_9;
output 	dout_10;
output 	dout_11;
output 	dout_12;
output 	dout_13;
output 	dout_14;
output 	dout_15;
output 	dout_16;
output 	dout_17;
output 	dout_18;
output 	dout_19;
output 	dout_20;
output 	dout_21;
output 	dout_22;
output 	dout_23;
output 	dout_24;
output 	dout_25;
output 	dout_26;
output 	dout_27;
output 	dout_28;
output 	dout_29;
output 	dout_30;
output 	dout_31;
output 	dout_32;
output 	dout_33;
output 	dout_5;
input 	dout_71;
output 	dout_4;
input 	dout_81;
input 	dout_91;
input 	dout_101;
input 	dout_111;
input 	dout_121;
input 	dout_131;
input 	dout_141;
input 	dout_151;
input 	dout_161;
input 	dout_171;
input 	dout_181;
input 	dout_191;
input 	dout_201;
input 	dout_211;
input 	dout_221;
input 	dout_231;
input 	dout_241;
input 	dout_251;
input 	dout_261;
input 	dout_271;
input 	dout_281;
input 	dout_291;
input 	dout_301;
input 	dout_311;
input 	dout_321;
input 	dout_331;
input 	dout_34;
input 	dout_61;
output 	dout_3;
input 	dout_51;
output 	dout_2;
input 	dout_41;
output 	dout_1;
input 	dout_35;
output 	dout_0;
input 	dout_210;
input 	dout_110;
input 	stall_reg;
input 	dout_valid3;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \glogic:u0|register_fifo:fifo_data[0][6]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][7]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][8]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][9]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][10]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][11]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][12]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][13]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][14]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][15]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][16]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][17]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][18]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][19]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][20]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][21]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][22]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][23]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][24]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][25]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][26]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][27]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][28]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][29]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][30]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][31]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][32]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][33]~q ;
wire \dout~1_combout ;
wire \glogic:u0|register_fifo:fifo_data[0][5]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][4]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][3]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][2]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][1]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][0]~q ;
wire \resq[0]~134 ;
wire \resq[0]~135 ;
wire \resq[1]~130 ;
wire \resq[1]~131 ;
wire \resq[2]~126 ;
wire \resq[2]~127 ;
wire \resq[3]~122 ;
wire \resq[3]~123 ;
wire \resq[4]~118 ;
wire \resq[4]~119 ;
wire \resq[5]~114 ;
wire \resq[5]~115 ;
wire \resq[6]~1_sumout ;
wire \dout[13]~0_combout ;
wire \resq[6]~2 ;
wire \resq[6]~3 ;
wire \resq[7]~5_sumout ;
wire \resq[7]~6 ;
wire \resq[7]~7 ;
wire \resq[8]~9_sumout ;
wire \resq[8]~10 ;
wire \resq[8]~11 ;
wire \resq[9]~13_sumout ;
wire \resq[9]~14 ;
wire \resq[9]~15 ;
wire \resq[10]~17_sumout ;
wire \resq[10]~18 ;
wire \resq[10]~19 ;
wire \resq[11]~21_sumout ;
wire \resq[11]~22 ;
wire \resq[11]~23 ;
wire \resq[12]~25_sumout ;
wire \resq[12]~26 ;
wire \resq[12]~27 ;
wire \resq[13]~29_sumout ;
wire \resq[13]~30 ;
wire \resq[13]~31 ;
wire \resq[14]~33_sumout ;
wire \resq[14]~34 ;
wire \resq[14]~35 ;
wire \resq[15]~37_sumout ;
wire \resq[15]~38 ;
wire \resq[15]~39 ;
wire \resq[16]~41_sumout ;
wire \resq[16]~42 ;
wire \resq[16]~43 ;
wire \resq[17]~45_sumout ;
wire \resq[17]~46 ;
wire \resq[17]~47 ;
wire \resq[18]~49_sumout ;
wire \resq[18]~50 ;
wire \resq[18]~51 ;
wire \resq[19]~53_sumout ;
wire \resq[19]~54 ;
wire \resq[19]~55 ;
wire \resq[20]~57_sumout ;
wire \resq[20]~58 ;
wire \resq[20]~59 ;
wire \resq[21]~61_sumout ;
wire \resq[21]~62 ;
wire \resq[21]~63 ;
wire \resq[22]~65_sumout ;
wire \resq[22]~66 ;
wire \resq[22]~67 ;
wire \resq[23]~69_sumout ;
wire \resq[23]~70 ;
wire \resq[23]~71 ;
wire \resq[24]~73_sumout ;
wire \resq[24]~74 ;
wire \resq[24]~75 ;
wire \resq[25]~77_sumout ;
wire \resq[25]~78 ;
wire \resq[25]~79 ;
wire \resq[26]~81_sumout ;
wire \resq[26]~82 ;
wire \resq[26]~83 ;
wire \resq[27]~85_sumout ;
wire \resq[27]~86 ;
wire \resq[27]~87 ;
wire \resq[28]~89_sumout ;
wire \resq[28]~90 ;
wire \resq[28]~91 ;
wire \resq[29]~93_sumout ;
wire \resq[29]~94 ;
wire \resq[29]~95 ;
wire \resq[30]~97_sumout ;
wire \resq[30]~98 ;
wire \resq[30]~99 ;
wire \resq[31]~101_sumout ;
wire \resq[31]~102 ;
wire \resq[31]~103 ;
wire \resq[32]~105_sumout ;
wire \resq[32]~106 ;
wire \resq[32]~107 ;
wire \resq[33]~109_sumout ;
wire \resq[5]~113_sumout ;
wire \resq[4]~117_sumout ;
wire \resq[3]~121_sumout ;
wire \resq[2]~125_sumout ;
wire \resq[1]~129_sumout ;
wire \resq[0]~133_sumout ;


cic_auk_dspip_delay_3 \glogic:u0 (
	.datain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,dout_34,dout_331,dout_321,dout_311,dout_301,dout_291,dout_281,dout_271,dout_261,dout_251,dout_241,dout_231,dout_221,dout_211,dout_201,dout_191,dout_181,dout_171,dout_161,dout_151,dout_141,dout_131,dout_121,dout_111,dout_101,dout_91,dout_81,
dout_71,dout_61,dout_51,dout_41,dout_35,dout_210,dout_110}),
	.register_fifofifo_data06(\glogic:u0|register_fifo:fifo_data[0][6]~q ),
	.register_fifofifo_data07(\glogic:u0|register_fifo:fifo_data[0][7]~q ),
	.register_fifofifo_data08(\glogic:u0|register_fifo:fifo_data[0][8]~q ),
	.register_fifofifo_data09(\glogic:u0|register_fifo:fifo_data[0][9]~q ),
	.register_fifofifo_data010(\glogic:u0|register_fifo:fifo_data[0][10]~q ),
	.register_fifofifo_data011(\glogic:u0|register_fifo:fifo_data[0][11]~q ),
	.register_fifofifo_data012(\glogic:u0|register_fifo:fifo_data[0][12]~q ),
	.register_fifofifo_data013(\glogic:u0|register_fifo:fifo_data[0][13]~q ),
	.register_fifofifo_data014(\glogic:u0|register_fifo:fifo_data[0][14]~q ),
	.register_fifofifo_data015(\glogic:u0|register_fifo:fifo_data[0][15]~q ),
	.register_fifofifo_data016(\glogic:u0|register_fifo:fifo_data[0][16]~q ),
	.register_fifofifo_data017(\glogic:u0|register_fifo:fifo_data[0][17]~q ),
	.register_fifofifo_data018(\glogic:u0|register_fifo:fifo_data[0][18]~q ),
	.register_fifofifo_data019(\glogic:u0|register_fifo:fifo_data[0][19]~q ),
	.register_fifofifo_data020(\glogic:u0|register_fifo:fifo_data[0][20]~q ),
	.register_fifofifo_data021(\glogic:u0|register_fifo:fifo_data[0][21]~q ),
	.register_fifofifo_data022(\glogic:u0|register_fifo:fifo_data[0][22]~q ),
	.register_fifofifo_data023(\glogic:u0|register_fifo:fifo_data[0][23]~q ),
	.register_fifofifo_data024(\glogic:u0|register_fifo:fifo_data[0][24]~q ),
	.register_fifofifo_data025(\glogic:u0|register_fifo:fifo_data[0][25]~q ),
	.register_fifofifo_data026(\glogic:u0|register_fifo:fifo_data[0][26]~q ),
	.register_fifofifo_data027(\glogic:u0|register_fifo:fifo_data[0][27]~q ),
	.register_fifofifo_data028(\glogic:u0|register_fifo:fifo_data[0][28]~q ),
	.register_fifofifo_data029(\glogic:u0|register_fifo:fifo_data[0][29]~q ),
	.register_fifofifo_data030(\glogic:u0|register_fifo:fifo_data[0][30]~q ),
	.register_fifofifo_data031(\glogic:u0|register_fifo:fifo_data[0][31]~q ),
	.register_fifofifo_data032(\glogic:u0|register_fifo:fifo_data[0][32]~q ),
	.register_fifofifo_data033(\glogic:u0|register_fifo:fifo_data[0][33]~q ),
	.enable(\dout~1_combout ),
	.register_fifofifo_data05(\glogic:u0|register_fifo:fifo_data[0][5]~q ),
	.register_fifofifo_data04(\glogic:u0|register_fifo:fifo_data[0][4]~q ),
	.register_fifofifo_data03(\glogic:u0|register_fifo:fifo_data[0][3]~q ),
	.register_fifofifo_data02(\glogic:u0|register_fifo:fifo_data[0][2]~q ),
	.register_fifofifo_data01(\glogic:u0|register_fifo:fifo_data[0][1]~q ),
	.register_fifofifo_data00(\glogic:u0|register_fifo:fifo_data[0][0]~q ),
	.clk(clk),
	.reset(reset_n));

arriav_lcell_comb \dout~1 (
	.dataa(!stall_reg),
	.datab(!dout_valid2),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dout~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dout~1 .extended_lut = "off";
defparam \dout~1 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \dout~1 .shared_arith = "off";

dffeas dout_valid(
	.clk(clk),
	.d(dout_valid2),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(dout_valid3),
	.q(dout_valid1),
	.prn(vcc));
defparam dout_valid.is_wysiwyg = "true";
defparam dout_valid.power_up = "low";

dffeas \dout[6] (
	.clk(clk),
	.d(\resq[6]~1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[13]~0_combout ),
	.q(dout_6),
	.prn(vcc));
defparam \dout[6] .is_wysiwyg = "true";
defparam \dout[6] .power_up = "low";

dffeas \dout[7] (
	.clk(clk),
	.d(\resq[7]~5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[13]~0_combout ),
	.q(dout_7),
	.prn(vcc));
defparam \dout[7] .is_wysiwyg = "true";
defparam \dout[7] .power_up = "low";

dffeas \dout[8] (
	.clk(clk),
	.d(\resq[8]~9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[13]~0_combout ),
	.q(dout_8),
	.prn(vcc));
defparam \dout[8] .is_wysiwyg = "true";
defparam \dout[8] .power_up = "low";

dffeas \dout[9] (
	.clk(clk),
	.d(\resq[9]~13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[13]~0_combout ),
	.q(dout_9),
	.prn(vcc));
defparam \dout[9] .is_wysiwyg = "true";
defparam \dout[9] .power_up = "low";

dffeas \dout[10] (
	.clk(clk),
	.d(\resq[10]~17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[13]~0_combout ),
	.q(dout_10),
	.prn(vcc));
defparam \dout[10] .is_wysiwyg = "true";
defparam \dout[10] .power_up = "low";

dffeas \dout[11] (
	.clk(clk),
	.d(\resq[11]~21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[13]~0_combout ),
	.q(dout_11),
	.prn(vcc));
defparam \dout[11] .is_wysiwyg = "true";
defparam \dout[11] .power_up = "low";

dffeas \dout[12] (
	.clk(clk),
	.d(\resq[12]~25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[13]~0_combout ),
	.q(dout_12),
	.prn(vcc));
defparam \dout[12] .is_wysiwyg = "true";
defparam \dout[12] .power_up = "low";

dffeas \dout[13] (
	.clk(clk),
	.d(\resq[13]~29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[13]~0_combout ),
	.q(dout_13),
	.prn(vcc));
defparam \dout[13] .is_wysiwyg = "true";
defparam \dout[13] .power_up = "low";

dffeas \dout[14] (
	.clk(clk),
	.d(\resq[14]~33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[13]~0_combout ),
	.q(dout_14),
	.prn(vcc));
defparam \dout[14] .is_wysiwyg = "true";
defparam \dout[14] .power_up = "low";

dffeas \dout[15] (
	.clk(clk),
	.d(\resq[15]~37_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[13]~0_combout ),
	.q(dout_15),
	.prn(vcc));
defparam \dout[15] .is_wysiwyg = "true";
defparam \dout[15] .power_up = "low";

dffeas \dout[16] (
	.clk(clk),
	.d(\resq[16]~41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[13]~0_combout ),
	.q(dout_16),
	.prn(vcc));
defparam \dout[16] .is_wysiwyg = "true";
defparam \dout[16] .power_up = "low";

dffeas \dout[17] (
	.clk(clk),
	.d(\resq[17]~45_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[13]~0_combout ),
	.q(dout_17),
	.prn(vcc));
defparam \dout[17] .is_wysiwyg = "true";
defparam \dout[17] .power_up = "low";

dffeas \dout[18] (
	.clk(clk),
	.d(\resq[18]~49_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[13]~0_combout ),
	.q(dout_18),
	.prn(vcc));
defparam \dout[18] .is_wysiwyg = "true";
defparam \dout[18] .power_up = "low";

dffeas \dout[19] (
	.clk(clk),
	.d(\resq[19]~53_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[13]~0_combout ),
	.q(dout_19),
	.prn(vcc));
defparam \dout[19] .is_wysiwyg = "true";
defparam \dout[19] .power_up = "low";

dffeas \dout[20] (
	.clk(clk),
	.d(\resq[20]~57_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[13]~0_combout ),
	.q(dout_20),
	.prn(vcc));
defparam \dout[20] .is_wysiwyg = "true";
defparam \dout[20] .power_up = "low";

dffeas \dout[21] (
	.clk(clk),
	.d(\resq[21]~61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[13]~0_combout ),
	.q(dout_21),
	.prn(vcc));
defparam \dout[21] .is_wysiwyg = "true";
defparam \dout[21] .power_up = "low";

dffeas \dout[22] (
	.clk(clk),
	.d(\resq[22]~65_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[13]~0_combout ),
	.q(dout_22),
	.prn(vcc));
defparam \dout[22] .is_wysiwyg = "true";
defparam \dout[22] .power_up = "low";

dffeas \dout[23] (
	.clk(clk),
	.d(\resq[23]~69_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[13]~0_combout ),
	.q(dout_23),
	.prn(vcc));
defparam \dout[23] .is_wysiwyg = "true";
defparam \dout[23] .power_up = "low";

dffeas \dout[24] (
	.clk(clk),
	.d(\resq[24]~73_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[13]~0_combout ),
	.q(dout_24),
	.prn(vcc));
defparam \dout[24] .is_wysiwyg = "true";
defparam \dout[24] .power_up = "low";

dffeas \dout[25] (
	.clk(clk),
	.d(\resq[25]~77_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[13]~0_combout ),
	.q(dout_25),
	.prn(vcc));
defparam \dout[25] .is_wysiwyg = "true";
defparam \dout[25] .power_up = "low";

dffeas \dout[26] (
	.clk(clk),
	.d(\resq[26]~81_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[13]~0_combout ),
	.q(dout_26),
	.prn(vcc));
defparam \dout[26] .is_wysiwyg = "true";
defparam \dout[26] .power_up = "low";

dffeas \dout[27] (
	.clk(clk),
	.d(\resq[27]~85_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[13]~0_combout ),
	.q(dout_27),
	.prn(vcc));
defparam \dout[27] .is_wysiwyg = "true";
defparam \dout[27] .power_up = "low";

dffeas \dout[28] (
	.clk(clk),
	.d(\resq[28]~89_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[13]~0_combout ),
	.q(dout_28),
	.prn(vcc));
defparam \dout[28] .is_wysiwyg = "true";
defparam \dout[28] .power_up = "low";

dffeas \dout[29] (
	.clk(clk),
	.d(\resq[29]~93_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[13]~0_combout ),
	.q(dout_29),
	.prn(vcc));
defparam \dout[29] .is_wysiwyg = "true";
defparam \dout[29] .power_up = "low";

dffeas \dout[30] (
	.clk(clk),
	.d(\resq[30]~97_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[13]~0_combout ),
	.q(dout_30),
	.prn(vcc));
defparam \dout[30] .is_wysiwyg = "true";
defparam \dout[30] .power_up = "low";

dffeas \dout[31] (
	.clk(clk),
	.d(\resq[31]~101_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[13]~0_combout ),
	.q(dout_31),
	.prn(vcc));
defparam \dout[31] .is_wysiwyg = "true";
defparam \dout[31] .power_up = "low";

dffeas \dout[32] (
	.clk(clk),
	.d(\resq[32]~105_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[13]~0_combout ),
	.q(dout_32),
	.prn(vcc));
defparam \dout[32] .is_wysiwyg = "true";
defparam \dout[32] .power_up = "low";

dffeas \dout[33] (
	.clk(clk),
	.d(\resq[33]~109_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[13]~0_combout ),
	.q(dout_33),
	.prn(vcc));
defparam \dout[33] .is_wysiwyg = "true";
defparam \dout[33] .power_up = "low";

dffeas \dout[5] (
	.clk(clk),
	.d(\resq[5]~113_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[13]~0_combout ),
	.q(dout_5),
	.prn(vcc));
defparam \dout[5] .is_wysiwyg = "true";
defparam \dout[5] .power_up = "low";

dffeas \dout[4] (
	.clk(clk),
	.d(\resq[4]~117_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[13]~0_combout ),
	.q(dout_4),
	.prn(vcc));
defparam \dout[4] .is_wysiwyg = "true";
defparam \dout[4] .power_up = "low";

dffeas \dout[3] (
	.clk(clk),
	.d(\resq[3]~121_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[13]~0_combout ),
	.q(dout_3),
	.prn(vcc));
defparam \dout[3] .is_wysiwyg = "true";
defparam \dout[3] .power_up = "low";

dffeas \dout[2] (
	.clk(clk),
	.d(\resq[2]~125_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[13]~0_combout ),
	.q(dout_2),
	.prn(vcc));
defparam \dout[2] .is_wysiwyg = "true";
defparam \dout[2] .power_up = "low";

dffeas \dout[1] (
	.clk(clk),
	.d(\resq[1]~129_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[13]~0_combout ),
	.q(dout_1),
	.prn(vcc));
defparam \dout[1] .is_wysiwyg = "true";
defparam \dout[1] .power_up = "low";

dffeas \dout[0] (
	.clk(clk),
	.d(\resq[0]~133_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[13]~0_combout ),
	.q(dout_0),
	.prn(vcc));
defparam \dout[0] .is_wysiwyg = "true";
defparam \dout[0] .power_up = "low";

arriav_lcell_comb \resq[0]~133 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][0]~q ),
	.datad(!dout_110),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\resq[0]~133_sumout ),
	.cout(\resq[0]~134 ),
	.shareout(\resq[0]~135 ));
defparam \resq[0]~133 .extended_lut = "off";
defparam \resq[0]~133 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[0]~133 .shared_arith = "on";

arriav_lcell_comb \resq[1]~129 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][1]~q ),
	.datad(!dout_210),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[0]~134 ),
	.sharein(\resq[0]~135 ),
	.combout(),
	.sumout(\resq[1]~129_sumout ),
	.cout(\resq[1]~130 ),
	.shareout(\resq[1]~131 ));
defparam \resq[1]~129 .extended_lut = "off";
defparam \resq[1]~129 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[1]~129 .shared_arith = "on";

arriav_lcell_comb \resq[2]~125 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][2]~q ),
	.datad(!dout_35),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[1]~130 ),
	.sharein(\resq[1]~131 ),
	.combout(),
	.sumout(\resq[2]~125_sumout ),
	.cout(\resq[2]~126 ),
	.shareout(\resq[2]~127 ));
defparam \resq[2]~125 .extended_lut = "off";
defparam \resq[2]~125 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[2]~125 .shared_arith = "on";

arriav_lcell_comb \resq[3]~121 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][3]~q ),
	.datad(!dout_41),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[2]~126 ),
	.sharein(\resq[2]~127 ),
	.combout(),
	.sumout(\resq[3]~121_sumout ),
	.cout(\resq[3]~122 ),
	.shareout(\resq[3]~123 ));
defparam \resq[3]~121 .extended_lut = "off";
defparam \resq[3]~121 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[3]~121 .shared_arith = "on";

arriav_lcell_comb \resq[4]~117 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][4]~q ),
	.datad(!dout_51),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[3]~122 ),
	.sharein(\resq[3]~123 ),
	.combout(),
	.sumout(\resq[4]~117_sumout ),
	.cout(\resq[4]~118 ),
	.shareout(\resq[4]~119 ));
defparam \resq[4]~117 .extended_lut = "off";
defparam \resq[4]~117 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[4]~117 .shared_arith = "on";

arriav_lcell_comb \resq[5]~113 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][5]~q ),
	.datad(!dout_61),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[4]~118 ),
	.sharein(\resq[4]~119 ),
	.combout(),
	.sumout(\resq[5]~113_sumout ),
	.cout(\resq[5]~114 ),
	.shareout(\resq[5]~115 ));
defparam \resq[5]~113 .extended_lut = "off";
defparam \resq[5]~113 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[5]~113 .shared_arith = "on";

arriav_lcell_comb \resq[6]~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][6]~q ),
	.datad(!dout_71),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[5]~114 ),
	.sharein(\resq[5]~115 ),
	.combout(),
	.sumout(\resq[6]~1_sumout ),
	.cout(\resq[6]~2 ),
	.shareout(\resq[6]~3 ));
defparam \resq[6]~1 .extended_lut = "off";
defparam \resq[6]~1 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[6]~1 .shared_arith = "on";

arriav_lcell_comb \dout[13]~0 (
	.dataa(!reset_n),
	.datab(!stall_reg),
	.datac(!dout_valid2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dout[13]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dout[13]~0 .extended_lut = "off";
defparam \dout[13]~0 .lut_mask = 64'hEFEFEFEFEFEFEFEF;
defparam \dout[13]~0 .shared_arith = "off";

arriav_lcell_comb \resq[7]~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][7]~q ),
	.datad(!dout_81),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[6]~2 ),
	.sharein(\resq[6]~3 ),
	.combout(),
	.sumout(\resq[7]~5_sumout ),
	.cout(\resq[7]~6 ),
	.shareout(\resq[7]~7 ));
defparam \resq[7]~5 .extended_lut = "off";
defparam \resq[7]~5 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[7]~5 .shared_arith = "on";

arriav_lcell_comb \resq[8]~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][8]~q ),
	.datad(!dout_91),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[7]~6 ),
	.sharein(\resq[7]~7 ),
	.combout(),
	.sumout(\resq[8]~9_sumout ),
	.cout(\resq[8]~10 ),
	.shareout(\resq[8]~11 ));
defparam \resq[8]~9 .extended_lut = "off";
defparam \resq[8]~9 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[8]~9 .shared_arith = "on";

arriav_lcell_comb \resq[9]~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][9]~q ),
	.datad(!dout_101),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[8]~10 ),
	.sharein(\resq[8]~11 ),
	.combout(),
	.sumout(\resq[9]~13_sumout ),
	.cout(\resq[9]~14 ),
	.shareout(\resq[9]~15 ));
defparam \resq[9]~13 .extended_lut = "off";
defparam \resq[9]~13 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[9]~13 .shared_arith = "on";

arriav_lcell_comb \resq[10]~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][10]~q ),
	.datad(!dout_111),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[9]~14 ),
	.sharein(\resq[9]~15 ),
	.combout(),
	.sumout(\resq[10]~17_sumout ),
	.cout(\resq[10]~18 ),
	.shareout(\resq[10]~19 ));
defparam \resq[10]~17 .extended_lut = "off";
defparam \resq[10]~17 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[10]~17 .shared_arith = "on";

arriav_lcell_comb \resq[11]~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][11]~q ),
	.datad(!dout_121),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[10]~18 ),
	.sharein(\resq[10]~19 ),
	.combout(),
	.sumout(\resq[11]~21_sumout ),
	.cout(\resq[11]~22 ),
	.shareout(\resq[11]~23 ));
defparam \resq[11]~21 .extended_lut = "off";
defparam \resq[11]~21 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[11]~21 .shared_arith = "on";

arriav_lcell_comb \resq[12]~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][12]~q ),
	.datad(!dout_131),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[11]~22 ),
	.sharein(\resq[11]~23 ),
	.combout(),
	.sumout(\resq[12]~25_sumout ),
	.cout(\resq[12]~26 ),
	.shareout(\resq[12]~27 ));
defparam \resq[12]~25 .extended_lut = "off";
defparam \resq[12]~25 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[12]~25 .shared_arith = "on";

arriav_lcell_comb \resq[13]~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][13]~q ),
	.datad(!dout_141),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[12]~26 ),
	.sharein(\resq[12]~27 ),
	.combout(),
	.sumout(\resq[13]~29_sumout ),
	.cout(\resq[13]~30 ),
	.shareout(\resq[13]~31 ));
defparam \resq[13]~29 .extended_lut = "off";
defparam \resq[13]~29 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[13]~29 .shared_arith = "on";

arriav_lcell_comb \resq[14]~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][14]~q ),
	.datad(!dout_151),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[13]~30 ),
	.sharein(\resq[13]~31 ),
	.combout(),
	.sumout(\resq[14]~33_sumout ),
	.cout(\resq[14]~34 ),
	.shareout(\resq[14]~35 ));
defparam \resq[14]~33 .extended_lut = "off";
defparam \resq[14]~33 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[14]~33 .shared_arith = "on";

arriav_lcell_comb \resq[15]~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][15]~q ),
	.datad(!dout_161),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[14]~34 ),
	.sharein(\resq[14]~35 ),
	.combout(),
	.sumout(\resq[15]~37_sumout ),
	.cout(\resq[15]~38 ),
	.shareout(\resq[15]~39 ));
defparam \resq[15]~37 .extended_lut = "off";
defparam \resq[15]~37 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[15]~37 .shared_arith = "on";

arriav_lcell_comb \resq[16]~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][16]~q ),
	.datad(!dout_171),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[15]~38 ),
	.sharein(\resq[15]~39 ),
	.combout(),
	.sumout(\resq[16]~41_sumout ),
	.cout(\resq[16]~42 ),
	.shareout(\resq[16]~43 ));
defparam \resq[16]~41 .extended_lut = "off";
defparam \resq[16]~41 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[16]~41 .shared_arith = "on";

arriav_lcell_comb \resq[17]~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][17]~q ),
	.datad(!dout_181),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[16]~42 ),
	.sharein(\resq[16]~43 ),
	.combout(),
	.sumout(\resq[17]~45_sumout ),
	.cout(\resq[17]~46 ),
	.shareout(\resq[17]~47 ));
defparam \resq[17]~45 .extended_lut = "off";
defparam \resq[17]~45 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[17]~45 .shared_arith = "on";

arriav_lcell_comb \resq[18]~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][18]~q ),
	.datad(!dout_191),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[17]~46 ),
	.sharein(\resq[17]~47 ),
	.combout(),
	.sumout(\resq[18]~49_sumout ),
	.cout(\resq[18]~50 ),
	.shareout(\resq[18]~51 ));
defparam \resq[18]~49 .extended_lut = "off";
defparam \resq[18]~49 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[18]~49 .shared_arith = "on";

arriav_lcell_comb \resq[19]~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][19]~q ),
	.datad(!dout_201),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[18]~50 ),
	.sharein(\resq[18]~51 ),
	.combout(),
	.sumout(\resq[19]~53_sumout ),
	.cout(\resq[19]~54 ),
	.shareout(\resq[19]~55 ));
defparam \resq[19]~53 .extended_lut = "off";
defparam \resq[19]~53 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[19]~53 .shared_arith = "on";

arriav_lcell_comb \resq[20]~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][20]~q ),
	.datad(!dout_211),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[19]~54 ),
	.sharein(\resq[19]~55 ),
	.combout(),
	.sumout(\resq[20]~57_sumout ),
	.cout(\resq[20]~58 ),
	.shareout(\resq[20]~59 ));
defparam \resq[20]~57 .extended_lut = "off";
defparam \resq[20]~57 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[20]~57 .shared_arith = "on";

arriav_lcell_comb \resq[21]~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][21]~q ),
	.datad(!dout_221),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[20]~58 ),
	.sharein(\resq[20]~59 ),
	.combout(),
	.sumout(\resq[21]~61_sumout ),
	.cout(\resq[21]~62 ),
	.shareout(\resq[21]~63 ));
defparam \resq[21]~61 .extended_lut = "off";
defparam \resq[21]~61 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[21]~61 .shared_arith = "on";

arriav_lcell_comb \resq[22]~65 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][22]~q ),
	.datad(!dout_231),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[21]~62 ),
	.sharein(\resq[21]~63 ),
	.combout(),
	.sumout(\resq[22]~65_sumout ),
	.cout(\resq[22]~66 ),
	.shareout(\resq[22]~67 ));
defparam \resq[22]~65 .extended_lut = "off";
defparam \resq[22]~65 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[22]~65 .shared_arith = "on";

arriav_lcell_comb \resq[23]~69 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][23]~q ),
	.datad(!dout_241),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[22]~66 ),
	.sharein(\resq[22]~67 ),
	.combout(),
	.sumout(\resq[23]~69_sumout ),
	.cout(\resq[23]~70 ),
	.shareout(\resq[23]~71 ));
defparam \resq[23]~69 .extended_lut = "off";
defparam \resq[23]~69 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[23]~69 .shared_arith = "on";

arriav_lcell_comb \resq[24]~73 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][24]~q ),
	.datad(!dout_251),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[23]~70 ),
	.sharein(\resq[23]~71 ),
	.combout(),
	.sumout(\resq[24]~73_sumout ),
	.cout(\resq[24]~74 ),
	.shareout(\resq[24]~75 ));
defparam \resq[24]~73 .extended_lut = "off";
defparam \resq[24]~73 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[24]~73 .shared_arith = "on";

arriav_lcell_comb \resq[25]~77 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][25]~q ),
	.datad(!dout_261),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[24]~74 ),
	.sharein(\resq[24]~75 ),
	.combout(),
	.sumout(\resq[25]~77_sumout ),
	.cout(\resq[25]~78 ),
	.shareout(\resq[25]~79 ));
defparam \resq[25]~77 .extended_lut = "off";
defparam \resq[25]~77 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[25]~77 .shared_arith = "on";

arriav_lcell_comb \resq[26]~81 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][26]~q ),
	.datad(!dout_271),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[25]~78 ),
	.sharein(\resq[25]~79 ),
	.combout(),
	.sumout(\resq[26]~81_sumout ),
	.cout(\resq[26]~82 ),
	.shareout(\resq[26]~83 ));
defparam \resq[26]~81 .extended_lut = "off";
defparam \resq[26]~81 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[26]~81 .shared_arith = "on";

arriav_lcell_comb \resq[27]~85 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][27]~q ),
	.datad(!dout_281),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[26]~82 ),
	.sharein(\resq[26]~83 ),
	.combout(),
	.sumout(\resq[27]~85_sumout ),
	.cout(\resq[27]~86 ),
	.shareout(\resq[27]~87 ));
defparam \resq[27]~85 .extended_lut = "off";
defparam \resq[27]~85 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[27]~85 .shared_arith = "on";

arriav_lcell_comb \resq[28]~89 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][28]~q ),
	.datad(!dout_291),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[27]~86 ),
	.sharein(\resq[27]~87 ),
	.combout(),
	.sumout(\resq[28]~89_sumout ),
	.cout(\resq[28]~90 ),
	.shareout(\resq[28]~91 ));
defparam \resq[28]~89 .extended_lut = "off";
defparam \resq[28]~89 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[28]~89 .shared_arith = "on";

arriav_lcell_comb \resq[29]~93 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][29]~q ),
	.datad(!dout_301),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[28]~90 ),
	.sharein(\resq[28]~91 ),
	.combout(),
	.sumout(\resq[29]~93_sumout ),
	.cout(\resq[29]~94 ),
	.shareout(\resq[29]~95 ));
defparam \resq[29]~93 .extended_lut = "off";
defparam \resq[29]~93 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[29]~93 .shared_arith = "on";

arriav_lcell_comb \resq[30]~97 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][30]~q ),
	.datad(!dout_311),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[29]~94 ),
	.sharein(\resq[29]~95 ),
	.combout(),
	.sumout(\resq[30]~97_sumout ),
	.cout(\resq[30]~98 ),
	.shareout(\resq[30]~99 ));
defparam \resq[30]~97 .extended_lut = "off";
defparam \resq[30]~97 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[30]~97 .shared_arith = "on";

arriav_lcell_comb \resq[31]~101 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][31]~q ),
	.datad(!dout_321),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[30]~98 ),
	.sharein(\resq[30]~99 ),
	.combout(),
	.sumout(\resq[31]~101_sumout ),
	.cout(\resq[31]~102 ),
	.shareout(\resq[31]~103 ));
defparam \resq[31]~101 .extended_lut = "off";
defparam \resq[31]~101 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[31]~101 .shared_arith = "on";

arriav_lcell_comb \resq[32]~105 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][32]~q ),
	.datad(!dout_331),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[31]~102 ),
	.sharein(\resq[31]~103 ),
	.combout(),
	.sumout(\resq[32]~105_sumout ),
	.cout(\resq[32]~106 ),
	.shareout(\resq[32]~107 ));
defparam \resq[32]~105 .extended_lut = "off";
defparam \resq[32]~105 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[32]~105 .shared_arith = "on";

arriav_lcell_comb \resq[33]~109 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][33]~q ),
	.datad(!dout_34),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[32]~106 ),
	.sharein(\resq[32]~107 ),
	.combout(),
	.sumout(\resq[33]~109_sumout ),
	.cout(),
	.shareout());
defparam \resq[33]~109 .extended_lut = "off";
defparam \resq[33]~109 .lut_mask = 64'h0000000000000FF0;
defparam \resq[33]~109 .shared_arith = "on";

endmodule

module cic_auk_dspip_delay_3 (
	datain,
	register_fifofifo_data06,
	register_fifofifo_data07,
	register_fifofifo_data08,
	register_fifofifo_data09,
	register_fifofifo_data010,
	register_fifofifo_data011,
	register_fifofifo_data012,
	register_fifofifo_data013,
	register_fifofifo_data014,
	register_fifofifo_data015,
	register_fifofifo_data016,
	register_fifofifo_data017,
	register_fifofifo_data018,
	register_fifofifo_data019,
	register_fifofifo_data020,
	register_fifofifo_data021,
	register_fifofifo_data022,
	register_fifofifo_data023,
	register_fifofifo_data024,
	register_fifofifo_data025,
	register_fifofifo_data026,
	register_fifofifo_data027,
	register_fifofifo_data028,
	register_fifofifo_data029,
	register_fifofifo_data030,
	register_fifofifo_data031,
	register_fifofifo_data032,
	register_fifofifo_data033,
	enable,
	register_fifofifo_data05,
	register_fifofifo_data04,
	register_fifofifo_data03,
	register_fifofifo_data02,
	register_fifofifo_data01,
	register_fifofifo_data00,
	clk,
	reset)/* synthesis synthesis_greybox=1 */;
input 	[46:0] datain;
output 	register_fifofifo_data06;
output 	register_fifofifo_data07;
output 	register_fifofifo_data08;
output 	register_fifofifo_data09;
output 	register_fifofifo_data010;
output 	register_fifofifo_data011;
output 	register_fifofifo_data012;
output 	register_fifofifo_data013;
output 	register_fifofifo_data014;
output 	register_fifofifo_data015;
output 	register_fifofifo_data016;
output 	register_fifofifo_data017;
output 	register_fifofifo_data018;
output 	register_fifofifo_data019;
output 	register_fifofifo_data020;
output 	register_fifofifo_data021;
output 	register_fifofifo_data022;
output 	register_fifofifo_data023;
output 	register_fifofifo_data024;
output 	register_fifofifo_data025;
output 	register_fifofifo_data026;
output 	register_fifofifo_data027;
output 	register_fifofifo_data028;
output 	register_fifofifo_data029;
output 	register_fifofifo_data030;
output 	register_fifofifo_data031;
output 	register_fifofifo_data032;
output 	register_fifofifo_data033;
input 	enable;
output 	register_fifofifo_data05;
output 	register_fifofifo_data04;
output 	register_fifofifo_data03;
output 	register_fifofifo_data02;
output 	register_fifofifo_data01;
output 	register_fifofifo_data00;
input 	clk;
input 	reset;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \register_fifo:fifo_data[0][6] (
	.clk(clk),
	.d(datain[6]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data06),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][6] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][6] .power_up = "low";

dffeas \register_fifo:fifo_data[0][7] (
	.clk(clk),
	.d(datain[7]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data07),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][7] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][7] .power_up = "low";

dffeas \register_fifo:fifo_data[0][8] (
	.clk(clk),
	.d(datain[8]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data08),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][8] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][8] .power_up = "low";

dffeas \register_fifo:fifo_data[0][9] (
	.clk(clk),
	.d(datain[9]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data09),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][9] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][9] .power_up = "low";

dffeas \register_fifo:fifo_data[0][10] (
	.clk(clk),
	.d(datain[10]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data010),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][10] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][10] .power_up = "low";

dffeas \register_fifo:fifo_data[0][11] (
	.clk(clk),
	.d(datain[11]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data011),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][11] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][11] .power_up = "low";

dffeas \register_fifo:fifo_data[0][12] (
	.clk(clk),
	.d(datain[12]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data012),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][12] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][12] .power_up = "low";

dffeas \register_fifo:fifo_data[0][13] (
	.clk(clk),
	.d(datain[13]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data013),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][13] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][13] .power_up = "low";

dffeas \register_fifo:fifo_data[0][14] (
	.clk(clk),
	.d(datain[14]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data014),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][14] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][14] .power_up = "low";

dffeas \register_fifo:fifo_data[0][15] (
	.clk(clk),
	.d(datain[15]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data015),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][15] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][15] .power_up = "low";

dffeas \register_fifo:fifo_data[0][16] (
	.clk(clk),
	.d(datain[16]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data016),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][16] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][16] .power_up = "low";

dffeas \register_fifo:fifo_data[0][17] (
	.clk(clk),
	.d(datain[17]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data017),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][17] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][17] .power_up = "low";

dffeas \register_fifo:fifo_data[0][18] (
	.clk(clk),
	.d(datain[18]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data018),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][18] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][18] .power_up = "low";

dffeas \register_fifo:fifo_data[0][19] (
	.clk(clk),
	.d(datain[19]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data019),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][19] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][19] .power_up = "low";

dffeas \register_fifo:fifo_data[0][20] (
	.clk(clk),
	.d(datain[20]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data020),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][20] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][20] .power_up = "low";

dffeas \register_fifo:fifo_data[0][21] (
	.clk(clk),
	.d(datain[21]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data021),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][21] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][21] .power_up = "low";

dffeas \register_fifo:fifo_data[0][22] (
	.clk(clk),
	.d(datain[22]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data022),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][22] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][22] .power_up = "low";

dffeas \register_fifo:fifo_data[0][23] (
	.clk(clk),
	.d(datain[23]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data023),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][23] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][23] .power_up = "low";

dffeas \register_fifo:fifo_data[0][24] (
	.clk(clk),
	.d(datain[24]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data024),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][24] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][24] .power_up = "low";

dffeas \register_fifo:fifo_data[0][25] (
	.clk(clk),
	.d(datain[25]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data025),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][25] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][25] .power_up = "low";

dffeas \register_fifo:fifo_data[0][26] (
	.clk(clk),
	.d(datain[26]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data026),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][26] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][26] .power_up = "low";

dffeas \register_fifo:fifo_data[0][27] (
	.clk(clk),
	.d(datain[27]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data027),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][27] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][27] .power_up = "low";

dffeas \register_fifo:fifo_data[0][28] (
	.clk(clk),
	.d(datain[28]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data028),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][28] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][28] .power_up = "low";

dffeas \register_fifo:fifo_data[0][29] (
	.clk(clk),
	.d(datain[29]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data029),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][29] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][29] .power_up = "low";

dffeas \register_fifo:fifo_data[0][30] (
	.clk(clk),
	.d(datain[30]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data030),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][30] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][30] .power_up = "low";

dffeas \register_fifo:fifo_data[0][31] (
	.clk(clk),
	.d(datain[31]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data031),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][31] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][31] .power_up = "low";

dffeas \register_fifo:fifo_data[0][32] (
	.clk(clk),
	.d(datain[32]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data032),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][32] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][32] .power_up = "low";

dffeas \register_fifo:fifo_data[0][33] (
	.clk(clk),
	.d(datain[33]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data033),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][33] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][33] .power_up = "low";

dffeas \register_fifo:fifo_data[0][5] (
	.clk(clk),
	.d(datain[5]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data05),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][5] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][5] .power_up = "low";

dffeas \register_fifo:fifo_data[0][4] (
	.clk(clk),
	.d(datain[4]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data04),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][4] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][4] .power_up = "low";

dffeas \register_fifo:fifo_data[0][3] (
	.clk(clk),
	.d(datain[3]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data03),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][3] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][3] .power_up = "low";

dffeas \register_fifo:fifo_data[0][2] (
	.clk(clk),
	.d(datain[2]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data02),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][2] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][2] .power_up = "low";

dffeas \register_fifo:fifo_data[0][1] (
	.clk(clk),
	.d(datain[1]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data01),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][1] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][1] .power_up = "low";

dffeas \register_fifo:fifo_data[0][0] (
	.clk(clk),
	.d(datain[0]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data00),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][0] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][0] .power_up = "low";

endmodule

module cic_auk_dspip_differentiator_4 (
	dout_valid1,
	dout_valid2,
	dout_6,
	dout_7,
	dout_8,
	dout_9,
	dout_10,
	dout_11,
	dout_12,
	dout_13,
	dout_14,
	dout_15,
	dout_16,
	dout_17,
	dout_18,
	dout_19,
	dout_20,
	dout_21,
	dout_22,
	dout_23,
	dout_24,
	dout_25,
	dout_26,
	dout_27,
	dout_28,
	dout_29,
	dout_30,
	dout_31,
	dout_32,
	dout_33,
	dout_5,
	dout_61,
	dout_4,
	dout_71,
	dout_81,
	dout_91,
	dout_101,
	dout_111,
	dout_121,
	dout_131,
	dout_141,
	dout_151,
	dout_161,
	dout_171,
	dout_181,
	dout_191,
	dout_201,
	dout_211,
	dout_221,
	dout_231,
	dout_241,
	dout_251,
	dout_261,
	dout_271,
	dout_281,
	dout_291,
	dout_301,
	dout_311,
	dout_321,
	dout_331,
	dout_51,
	dout_3,
	dout_41,
	dout_2,
	dout_34,
	dout_1,
	dout_210,
	dout_110,
	dout_0,
	stall_reg,
	dout_valid3,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	dout_valid1;
input 	dout_valid2;
output 	dout_6;
output 	dout_7;
output 	dout_8;
output 	dout_9;
output 	dout_10;
output 	dout_11;
output 	dout_12;
output 	dout_13;
output 	dout_14;
output 	dout_15;
output 	dout_16;
output 	dout_17;
output 	dout_18;
output 	dout_19;
output 	dout_20;
output 	dout_21;
output 	dout_22;
output 	dout_23;
output 	dout_24;
output 	dout_25;
output 	dout_26;
output 	dout_27;
output 	dout_28;
output 	dout_29;
output 	dout_30;
output 	dout_31;
output 	dout_32;
output 	dout_33;
output 	dout_5;
input 	dout_61;
output 	dout_4;
input 	dout_71;
input 	dout_81;
input 	dout_91;
input 	dout_101;
input 	dout_111;
input 	dout_121;
input 	dout_131;
input 	dout_141;
input 	dout_151;
input 	dout_161;
input 	dout_171;
input 	dout_181;
input 	dout_191;
input 	dout_201;
input 	dout_211;
input 	dout_221;
input 	dout_231;
input 	dout_241;
input 	dout_251;
input 	dout_261;
input 	dout_271;
input 	dout_281;
input 	dout_291;
input 	dout_301;
input 	dout_311;
input 	dout_321;
input 	dout_331;
input 	dout_51;
output 	dout_3;
input 	dout_41;
output 	dout_2;
input 	dout_34;
output 	dout_1;
input 	dout_210;
input 	dout_110;
input 	dout_0;
input 	stall_reg;
input 	dout_valid3;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \glogic:u0|register_fifo:fifo_data[0][6]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][7]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][8]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][9]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][10]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][11]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][12]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][13]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][14]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][15]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][16]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][17]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][18]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][19]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][20]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][21]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][22]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][23]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][24]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][25]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][26]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][27]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][28]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][29]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][30]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][31]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][32]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][33]~q ;
wire \dout~1_combout ;
wire \glogic:u0|register_fifo:fifo_data[0][5]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][4]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][3]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][2]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][1]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][0]~q ;
wire \resq[0]~134_cout ;
wire \resq[0]~135 ;
wire \resq[1]~130 ;
wire \resq[1]~131 ;
wire \resq[2]~126 ;
wire \resq[2]~127 ;
wire \resq[3]~122 ;
wire \resq[3]~123 ;
wire \resq[4]~118 ;
wire \resq[4]~119 ;
wire \resq[5]~114 ;
wire \resq[5]~115 ;
wire \resq[6]~1_sumout ;
wire \dout[18]~0_combout ;
wire \resq[6]~2 ;
wire \resq[6]~3 ;
wire \resq[7]~5_sumout ;
wire \resq[7]~6 ;
wire \resq[7]~7 ;
wire \resq[8]~9_sumout ;
wire \resq[8]~10 ;
wire \resq[8]~11 ;
wire \resq[9]~13_sumout ;
wire \resq[9]~14 ;
wire \resq[9]~15 ;
wire \resq[10]~17_sumout ;
wire \resq[10]~18 ;
wire \resq[10]~19 ;
wire \resq[11]~21_sumout ;
wire \resq[11]~22 ;
wire \resq[11]~23 ;
wire \resq[12]~25_sumout ;
wire \resq[12]~26 ;
wire \resq[12]~27 ;
wire \resq[13]~29_sumout ;
wire \resq[13]~30 ;
wire \resq[13]~31 ;
wire \resq[14]~33_sumout ;
wire \resq[14]~34 ;
wire \resq[14]~35 ;
wire \resq[15]~37_sumout ;
wire \resq[15]~38 ;
wire \resq[15]~39 ;
wire \resq[16]~41_sumout ;
wire \resq[16]~42 ;
wire \resq[16]~43 ;
wire \resq[17]~45_sumout ;
wire \resq[17]~46 ;
wire \resq[17]~47 ;
wire \resq[18]~49_sumout ;
wire \resq[18]~50 ;
wire \resq[18]~51 ;
wire \resq[19]~53_sumout ;
wire \resq[19]~54 ;
wire \resq[19]~55 ;
wire \resq[20]~57_sumout ;
wire \resq[20]~58 ;
wire \resq[20]~59 ;
wire \resq[21]~61_sumout ;
wire \resq[21]~62 ;
wire \resq[21]~63 ;
wire \resq[22]~65_sumout ;
wire \resq[22]~66 ;
wire \resq[22]~67 ;
wire \resq[23]~69_sumout ;
wire \resq[23]~70 ;
wire \resq[23]~71 ;
wire \resq[24]~73_sumout ;
wire \resq[24]~74 ;
wire \resq[24]~75 ;
wire \resq[25]~77_sumout ;
wire \resq[25]~78 ;
wire \resq[25]~79 ;
wire \resq[26]~81_sumout ;
wire \resq[26]~82 ;
wire \resq[26]~83 ;
wire \resq[27]~85_sumout ;
wire \resq[27]~86 ;
wire \resq[27]~87 ;
wire \resq[28]~89_sumout ;
wire \resq[28]~90 ;
wire \resq[28]~91 ;
wire \resq[29]~93_sumout ;
wire \resq[29]~94 ;
wire \resq[29]~95 ;
wire \resq[30]~97_sumout ;
wire \resq[30]~98 ;
wire \resq[30]~99 ;
wire \resq[31]~101_sumout ;
wire \resq[31]~102 ;
wire \resq[31]~103 ;
wire \resq[32]~105_sumout ;
wire \resq[32]~106 ;
wire \resq[32]~107 ;
wire \resq[33]~109_sumout ;
wire \resq[5]~113_sumout ;
wire \resq[4]~117_sumout ;
wire \resq[3]~121_sumout ;
wire \resq[2]~125_sumout ;
wire \resq[1]~129_sumout ;


cic_auk_dspip_delay_4 \glogic:u0 (
	.datain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,dout_331,dout_321,dout_311,dout_301,dout_291,dout_281,dout_271,dout_261,dout_251,dout_241,dout_231,dout_221,dout_211,dout_201,dout_191,dout_181,dout_171,dout_161,dout_151,dout_141,dout_131,dout_121,dout_111,dout_101,dout_91,dout_81,dout_71,
dout_61,dout_51,dout_41,dout_34,dout_210,dout_110,dout_0}),
	.register_fifofifo_data06(\glogic:u0|register_fifo:fifo_data[0][6]~q ),
	.register_fifofifo_data07(\glogic:u0|register_fifo:fifo_data[0][7]~q ),
	.register_fifofifo_data08(\glogic:u0|register_fifo:fifo_data[0][8]~q ),
	.register_fifofifo_data09(\glogic:u0|register_fifo:fifo_data[0][9]~q ),
	.register_fifofifo_data010(\glogic:u0|register_fifo:fifo_data[0][10]~q ),
	.register_fifofifo_data011(\glogic:u0|register_fifo:fifo_data[0][11]~q ),
	.register_fifofifo_data012(\glogic:u0|register_fifo:fifo_data[0][12]~q ),
	.register_fifofifo_data013(\glogic:u0|register_fifo:fifo_data[0][13]~q ),
	.register_fifofifo_data014(\glogic:u0|register_fifo:fifo_data[0][14]~q ),
	.register_fifofifo_data015(\glogic:u0|register_fifo:fifo_data[0][15]~q ),
	.register_fifofifo_data016(\glogic:u0|register_fifo:fifo_data[0][16]~q ),
	.register_fifofifo_data017(\glogic:u0|register_fifo:fifo_data[0][17]~q ),
	.register_fifofifo_data018(\glogic:u0|register_fifo:fifo_data[0][18]~q ),
	.register_fifofifo_data019(\glogic:u0|register_fifo:fifo_data[0][19]~q ),
	.register_fifofifo_data020(\glogic:u0|register_fifo:fifo_data[0][20]~q ),
	.register_fifofifo_data021(\glogic:u0|register_fifo:fifo_data[0][21]~q ),
	.register_fifofifo_data022(\glogic:u0|register_fifo:fifo_data[0][22]~q ),
	.register_fifofifo_data023(\glogic:u0|register_fifo:fifo_data[0][23]~q ),
	.register_fifofifo_data024(\glogic:u0|register_fifo:fifo_data[0][24]~q ),
	.register_fifofifo_data025(\glogic:u0|register_fifo:fifo_data[0][25]~q ),
	.register_fifofifo_data026(\glogic:u0|register_fifo:fifo_data[0][26]~q ),
	.register_fifofifo_data027(\glogic:u0|register_fifo:fifo_data[0][27]~q ),
	.register_fifofifo_data028(\glogic:u0|register_fifo:fifo_data[0][28]~q ),
	.register_fifofifo_data029(\glogic:u0|register_fifo:fifo_data[0][29]~q ),
	.register_fifofifo_data030(\glogic:u0|register_fifo:fifo_data[0][30]~q ),
	.register_fifofifo_data031(\glogic:u0|register_fifo:fifo_data[0][31]~q ),
	.register_fifofifo_data032(\glogic:u0|register_fifo:fifo_data[0][32]~q ),
	.register_fifofifo_data033(\glogic:u0|register_fifo:fifo_data[0][33]~q ),
	.enable(\dout~1_combout ),
	.register_fifofifo_data05(\glogic:u0|register_fifo:fifo_data[0][5]~q ),
	.register_fifofifo_data04(\glogic:u0|register_fifo:fifo_data[0][4]~q ),
	.register_fifofifo_data03(\glogic:u0|register_fifo:fifo_data[0][3]~q ),
	.register_fifofifo_data02(\glogic:u0|register_fifo:fifo_data[0][2]~q ),
	.register_fifofifo_data01(\glogic:u0|register_fifo:fifo_data[0][1]~q ),
	.register_fifofifo_data00(\glogic:u0|register_fifo:fifo_data[0][0]~q ),
	.clk(clk),
	.reset(reset_n));

arriav_lcell_comb \dout~1 (
	.dataa(!stall_reg),
	.datab(!dout_valid2),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dout~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dout~1 .extended_lut = "off";
defparam \dout~1 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \dout~1 .shared_arith = "off";

dffeas dout_valid(
	.clk(clk),
	.d(dout_valid2),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(dout_valid3),
	.q(dout_valid1),
	.prn(vcc));
defparam dout_valid.is_wysiwyg = "true";
defparam dout_valid.power_up = "low";

dffeas \dout[6] (
	.clk(clk),
	.d(\resq[6]~1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[18]~0_combout ),
	.q(dout_6),
	.prn(vcc));
defparam \dout[6] .is_wysiwyg = "true";
defparam \dout[6] .power_up = "low";

dffeas \dout[7] (
	.clk(clk),
	.d(\resq[7]~5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[18]~0_combout ),
	.q(dout_7),
	.prn(vcc));
defparam \dout[7] .is_wysiwyg = "true";
defparam \dout[7] .power_up = "low";

dffeas \dout[8] (
	.clk(clk),
	.d(\resq[8]~9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[18]~0_combout ),
	.q(dout_8),
	.prn(vcc));
defparam \dout[8] .is_wysiwyg = "true";
defparam \dout[8] .power_up = "low";

dffeas \dout[9] (
	.clk(clk),
	.d(\resq[9]~13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[18]~0_combout ),
	.q(dout_9),
	.prn(vcc));
defparam \dout[9] .is_wysiwyg = "true";
defparam \dout[9] .power_up = "low";

dffeas \dout[10] (
	.clk(clk),
	.d(\resq[10]~17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[18]~0_combout ),
	.q(dout_10),
	.prn(vcc));
defparam \dout[10] .is_wysiwyg = "true";
defparam \dout[10] .power_up = "low";

dffeas \dout[11] (
	.clk(clk),
	.d(\resq[11]~21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[18]~0_combout ),
	.q(dout_11),
	.prn(vcc));
defparam \dout[11] .is_wysiwyg = "true";
defparam \dout[11] .power_up = "low";

dffeas \dout[12] (
	.clk(clk),
	.d(\resq[12]~25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[18]~0_combout ),
	.q(dout_12),
	.prn(vcc));
defparam \dout[12] .is_wysiwyg = "true";
defparam \dout[12] .power_up = "low";

dffeas \dout[13] (
	.clk(clk),
	.d(\resq[13]~29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[18]~0_combout ),
	.q(dout_13),
	.prn(vcc));
defparam \dout[13] .is_wysiwyg = "true";
defparam \dout[13] .power_up = "low";

dffeas \dout[14] (
	.clk(clk),
	.d(\resq[14]~33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[18]~0_combout ),
	.q(dout_14),
	.prn(vcc));
defparam \dout[14] .is_wysiwyg = "true";
defparam \dout[14] .power_up = "low";

dffeas \dout[15] (
	.clk(clk),
	.d(\resq[15]~37_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[18]~0_combout ),
	.q(dout_15),
	.prn(vcc));
defparam \dout[15] .is_wysiwyg = "true";
defparam \dout[15] .power_up = "low";

dffeas \dout[16] (
	.clk(clk),
	.d(\resq[16]~41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[18]~0_combout ),
	.q(dout_16),
	.prn(vcc));
defparam \dout[16] .is_wysiwyg = "true";
defparam \dout[16] .power_up = "low";

dffeas \dout[17] (
	.clk(clk),
	.d(\resq[17]~45_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[18]~0_combout ),
	.q(dout_17),
	.prn(vcc));
defparam \dout[17] .is_wysiwyg = "true";
defparam \dout[17] .power_up = "low";

dffeas \dout[18] (
	.clk(clk),
	.d(\resq[18]~49_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[18]~0_combout ),
	.q(dout_18),
	.prn(vcc));
defparam \dout[18] .is_wysiwyg = "true";
defparam \dout[18] .power_up = "low";

dffeas \dout[19] (
	.clk(clk),
	.d(\resq[19]~53_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[18]~0_combout ),
	.q(dout_19),
	.prn(vcc));
defparam \dout[19] .is_wysiwyg = "true";
defparam \dout[19] .power_up = "low";

dffeas \dout[20] (
	.clk(clk),
	.d(\resq[20]~57_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[18]~0_combout ),
	.q(dout_20),
	.prn(vcc));
defparam \dout[20] .is_wysiwyg = "true";
defparam \dout[20] .power_up = "low";

dffeas \dout[21] (
	.clk(clk),
	.d(\resq[21]~61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[18]~0_combout ),
	.q(dout_21),
	.prn(vcc));
defparam \dout[21] .is_wysiwyg = "true";
defparam \dout[21] .power_up = "low";

dffeas \dout[22] (
	.clk(clk),
	.d(\resq[22]~65_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[18]~0_combout ),
	.q(dout_22),
	.prn(vcc));
defparam \dout[22] .is_wysiwyg = "true";
defparam \dout[22] .power_up = "low";

dffeas \dout[23] (
	.clk(clk),
	.d(\resq[23]~69_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[18]~0_combout ),
	.q(dout_23),
	.prn(vcc));
defparam \dout[23] .is_wysiwyg = "true";
defparam \dout[23] .power_up = "low";

dffeas \dout[24] (
	.clk(clk),
	.d(\resq[24]~73_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[18]~0_combout ),
	.q(dout_24),
	.prn(vcc));
defparam \dout[24] .is_wysiwyg = "true";
defparam \dout[24] .power_up = "low";

dffeas \dout[25] (
	.clk(clk),
	.d(\resq[25]~77_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[18]~0_combout ),
	.q(dout_25),
	.prn(vcc));
defparam \dout[25] .is_wysiwyg = "true";
defparam \dout[25] .power_up = "low";

dffeas \dout[26] (
	.clk(clk),
	.d(\resq[26]~81_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[18]~0_combout ),
	.q(dout_26),
	.prn(vcc));
defparam \dout[26] .is_wysiwyg = "true";
defparam \dout[26] .power_up = "low";

dffeas \dout[27] (
	.clk(clk),
	.d(\resq[27]~85_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[18]~0_combout ),
	.q(dout_27),
	.prn(vcc));
defparam \dout[27] .is_wysiwyg = "true";
defparam \dout[27] .power_up = "low";

dffeas \dout[28] (
	.clk(clk),
	.d(\resq[28]~89_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[18]~0_combout ),
	.q(dout_28),
	.prn(vcc));
defparam \dout[28] .is_wysiwyg = "true";
defparam \dout[28] .power_up = "low";

dffeas \dout[29] (
	.clk(clk),
	.d(\resq[29]~93_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[18]~0_combout ),
	.q(dout_29),
	.prn(vcc));
defparam \dout[29] .is_wysiwyg = "true";
defparam \dout[29] .power_up = "low";

dffeas \dout[30] (
	.clk(clk),
	.d(\resq[30]~97_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[18]~0_combout ),
	.q(dout_30),
	.prn(vcc));
defparam \dout[30] .is_wysiwyg = "true";
defparam \dout[30] .power_up = "low";

dffeas \dout[31] (
	.clk(clk),
	.d(\resq[31]~101_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[18]~0_combout ),
	.q(dout_31),
	.prn(vcc));
defparam \dout[31] .is_wysiwyg = "true";
defparam \dout[31] .power_up = "low";

dffeas \dout[32] (
	.clk(clk),
	.d(\resq[32]~105_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[18]~0_combout ),
	.q(dout_32),
	.prn(vcc));
defparam \dout[32] .is_wysiwyg = "true";
defparam \dout[32] .power_up = "low";

dffeas \dout[33] (
	.clk(clk),
	.d(\resq[33]~109_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[18]~0_combout ),
	.q(dout_33),
	.prn(vcc));
defparam \dout[33] .is_wysiwyg = "true";
defparam \dout[33] .power_up = "low";

dffeas \dout[5] (
	.clk(clk),
	.d(\resq[5]~113_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[18]~0_combout ),
	.q(dout_5),
	.prn(vcc));
defparam \dout[5] .is_wysiwyg = "true";
defparam \dout[5] .power_up = "low";

dffeas \dout[4] (
	.clk(clk),
	.d(\resq[4]~117_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[18]~0_combout ),
	.q(dout_4),
	.prn(vcc));
defparam \dout[4] .is_wysiwyg = "true";
defparam \dout[4] .power_up = "low";

dffeas \dout[3] (
	.clk(clk),
	.d(\resq[3]~121_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[18]~0_combout ),
	.q(dout_3),
	.prn(vcc));
defparam \dout[3] .is_wysiwyg = "true";
defparam \dout[3] .power_up = "low";

dffeas \dout[2] (
	.clk(clk),
	.d(\resq[2]~125_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[18]~0_combout ),
	.q(dout_2),
	.prn(vcc));
defparam \dout[2] .is_wysiwyg = "true";
defparam \dout[2] .power_up = "low";

dffeas \dout[1] (
	.clk(clk),
	.d(\resq[1]~129_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[18]~0_combout ),
	.q(dout_1),
	.prn(vcc));
defparam \dout[1] .is_wysiwyg = "true";
defparam \dout[1] .power_up = "low";

arriav_lcell_comb \resq[0]~134 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][0]~q ),
	.datad(!dout_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\resq[0]~134_cout ),
	.shareout(\resq[0]~135 ));
defparam \resq[0]~134 .extended_lut = "off";
defparam \resq[0]~134 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[0]~134 .shared_arith = "on";

arriav_lcell_comb \resq[1]~129 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][1]~q ),
	.datad(!dout_110),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[0]~134_cout ),
	.sharein(\resq[0]~135 ),
	.combout(),
	.sumout(\resq[1]~129_sumout ),
	.cout(\resq[1]~130 ),
	.shareout(\resq[1]~131 ));
defparam \resq[1]~129 .extended_lut = "off";
defparam \resq[1]~129 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[1]~129 .shared_arith = "on";

arriav_lcell_comb \resq[2]~125 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][2]~q ),
	.datad(!dout_210),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[1]~130 ),
	.sharein(\resq[1]~131 ),
	.combout(),
	.sumout(\resq[2]~125_sumout ),
	.cout(\resq[2]~126 ),
	.shareout(\resq[2]~127 ));
defparam \resq[2]~125 .extended_lut = "off";
defparam \resq[2]~125 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[2]~125 .shared_arith = "on";

arriav_lcell_comb \resq[3]~121 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][3]~q ),
	.datad(!dout_34),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[2]~126 ),
	.sharein(\resq[2]~127 ),
	.combout(),
	.sumout(\resq[3]~121_sumout ),
	.cout(\resq[3]~122 ),
	.shareout(\resq[3]~123 ));
defparam \resq[3]~121 .extended_lut = "off";
defparam \resq[3]~121 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[3]~121 .shared_arith = "on";

arriav_lcell_comb \resq[4]~117 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][4]~q ),
	.datad(!dout_41),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[3]~122 ),
	.sharein(\resq[3]~123 ),
	.combout(),
	.sumout(\resq[4]~117_sumout ),
	.cout(\resq[4]~118 ),
	.shareout(\resq[4]~119 ));
defparam \resq[4]~117 .extended_lut = "off";
defparam \resq[4]~117 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[4]~117 .shared_arith = "on";

arriav_lcell_comb \resq[5]~113 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][5]~q ),
	.datad(!dout_51),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[4]~118 ),
	.sharein(\resq[4]~119 ),
	.combout(),
	.sumout(\resq[5]~113_sumout ),
	.cout(\resq[5]~114 ),
	.shareout(\resq[5]~115 ));
defparam \resq[5]~113 .extended_lut = "off";
defparam \resq[5]~113 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[5]~113 .shared_arith = "on";

arriav_lcell_comb \resq[6]~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][6]~q ),
	.datad(!dout_61),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[5]~114 ),
	.sharein(\resq[5]~115 ),
	.combout(),
	.sumout(\resq[6]~1_sumout ),
	.cout(\resq[6]~2 ),
	.shareout(\resq[6]~3 ));
defparam \resq[6]~1 .extended_lut = "off";
defparam \resq[6]~1 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[6]~1 .shared_arith = "on";

arriav_lcell_comb \dout[18]~0 (
	.dataa(!reset_n),
	.datab(!stall_reg),
	.datac(!dout_valid2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dout[18]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dout[18]~0 .extended_lut = "off";
defparam \dout[18]~0 .lut_mask = 64'hEFEFEFEFEFEFEFEF;
defparam \dout[18]~0 .shared_arith = "off";

arriav_lcell_comb \resq[7]~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][7]~q ),
	.datad(!dout_71),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[6]~2 ),
	.sharein(\resq[6]~3 ),
	.combout(),
	.sumout(\resq[7]~5_sumout ),
	.cout(\resq[7]~6 ),
	.shareout(\resq[7]~7 ));
defparam \resq[7]~5 .extended_lut = "off";
defparam \resq[7]~5 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[7]~5 .shared_arith = "on";

arriav_lcell_comb \resq[8]~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][8]~q ),
	.datad(!dout_81),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[7]~6 ),
	.sharein(\resq[7]~7 ),
	.combout(),
	.sumout(\resq[8]~9_sumout ),
	.cout(\resq[8]~10 ),
	.shareout(\resq[8]~11 ));
defparam \resq[8]~9 .extended_lut = "off";
defparam \resq[8]~9 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[8]~9 .shared_arith = "on";

arriav_lcell_comb \resq[9]~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][9]~q ),
	.datad(!dout_91),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[8]~10 ),
	.sharein(\resq[8]~11 ),
	.combout(),
	.sumout(\resq[9]~13_sumout ),
	.cout(\resq[9]~14 ),
	.shareout(\resq[9]~15 ));
defparam \resq[9]~13 .extended_lut = "off";
defparam \resq[9]~13 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[9]~13 .shared_arith = "on";

arriav_lcell_comb \resq[10]~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][10]~q ),
	.datad(!dout_101),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[9]~14 ),
	.sharein(\resq[9]~15 ),
	.combout(),
	.sumout(\resq[10]~17_sumout ),
	.cout(\resq[10]~18 ),
	.shareout(\resq[10]~19 ));
defparam \resq[10]~17 .extended_lut = "off";
defparam \resq[10]~17 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[10]~17 .shared_arith = "on";

arriav_lcell_comb \resq[11]~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][11]~q ),
	.datad(!dout_111),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[10]~18 ),
	.sharein(\resq[10]~19 ),
	.combout(),
	.sumout(\resq[11]~21_sumout ),
	.cout(\resq[11]~22 ),
	.shareout(\resq[11]~23 ));
defparam \resq[11]~21 .extended_lut = "off";
defparam \resq[11]~21 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[11]~21 .shared_arith = "on";

arriav_lcell_comb \resq[12]~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][12]~q ),
	.datad(!dout_121),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[11]~22 ),
	.sharein(\resq[11]~23 ),
	.combout(),
	.sumout(\resq[12]~25_sumout ),
	.cout(\resq[12]~26 ),
	.shareout(\resq[12]~27 ));
defparam \resq[12]~25 .extended_lut = "off";
defparam \resq[12]~25 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[12]~25 .shared_arith = "on";

arriav_lcell_comb \resq[13]~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][13]~q ),
	.datad(!dout_131),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[12]~26 ),
	.sharein(\resq[12]~27 ),
	.combout(),
	.sumout(\resq[13]~29_sumout ),
	.cout(\resq[13]~30 ),
	.shareout(\resq[13]~31 ));
defparam \resq[13]~29 .extended_lut = "off";
defparam \resq[13]~29 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[13]~29 .shared_arith = "on";

arriav_lcell_comb \resq[14]~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][14]~q ),
	.datad(!dout_141),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[13]~30 ),
	.sharein(\resq[13]~31 ),
	.combout(),
	.sumout(\resq[14]~33_sumout ),
	.cout(\resq[14]~34 ),
	.shareout(\resq[14]~35 ));
defparam \resq[14]~33 .extended_lut = "off";
defparam \resq[14]~33 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[14]~33 .shared_arith = "on";

arriav_lcell_comb \resq[15]~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][15]~q ),
	.datad(!dout_151),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[14]~34 ),
	.sharein(\resq[14]~35 ),
	.combout(),
	.sumout(\resq[15]~37_sumout ),
	.cout(\resq[15]~38 ),
	.shareout(\resq[15]~39 ));
defparam \resq[15]~37 .extended_lut = "off";
defparam \resq[15]~37 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[15]~37 .shared_arith = "on";

arriav_lcell_comb \resq[16]~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][16]~q ),
	.datad(!dout_161),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[15]~38 ),
	.sharein(\resq[15]~39 ),
	.combout(),
	.sumout(\resq[16]~41_sumout ),
	.cout(\resq[16]~42 ),
	.shareout(\resq[16]~43 ));
defparam \resq[16]~41 .extended_lut = "off";
defparam \resq[16]~41 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[16]~41 .shared_arith = "on";

arriav_lcell_comb \resq[17]~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][17]~q ),
	.datad(!dout_171),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[16]~42 ),
	.sharein(\resq[16]~43 ),
	.combout(),
	.sumout(\resq[17]~45_sumout ),
	.cout(\resq[17]~46 ),
	.shareout(\resq[17]~47 ));
defparam \resq[17]~45 .extended_lut = "off";
defparam \resq[17]~45 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[17]~45 .shared_arith = "on";

arriav_lcell_comb \resq[18]~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][18]~q ),
	.datad(!dout_181),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[17]~46 ),
	.sharein(\resq[17]~47 ),
	.combout(),
	.sumout(\resq[18]~49_sumout ),
	.cout(\resq[18]~50 ),
	.shareout(\resq[18]~51 ));
defparam \resq[18]~49 .extended_lut = "off";
defparam \resq[18]~49 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[18]~49 .shared_arith = "on";

arriav_lcell_comb \resq[19]~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][19]~q ),
	.datad(!dout_191),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[18]~50 ),
	.sharein(\resq[18]~51 ),
	.combout(),
	.sumout(\resq[19]~53_sumout ),
	.cout(\resq[19]~54 ),
	.shareout(\resq[19]~55 ));
defparam \resq[19]~53 .extended_lut = "off";
defparam \resq[19]~53 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[19]~53 .shared_arith = "on";

arriav_lcell_comb \resq[20]~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][20]~q ),
	.datad(!dout_201),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[19]~54 ),
	.sharein(\resq[19]~55 ),
	.combout(),
	.sumout(\resq[20]~57_sumout ),
	.cout(\resq[20]~58 ),
	.shareout(\resq[20]~59 ));
defparam \resq[20]~57 .extended_lut = "off";
defparam \resq[20]~57 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[20]~57 .shared_arith = "on";

arriav_lcell_comb \resq[21]~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][21]~q ),
	.datad(!dout_211),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[20]~58 ),
	.sharein(\resq[20]~59 ),
	.combout(),
	.sumout(\resq[21]~61_sumout ),
	.cout(\resq[21]~62 ),
	.shareout(\resq[21]~63 ));
defparam \resq[21]~61 .extended_lut = "off";
defparam \resq[21]~61 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[21]~61 .shared_arith = "on";

arriav_lcell_comb \resq[22]~65 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][22]~q ),
	.datad(!dout_221),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[21]~62 ),
	.sharein(\resq[21]~63 ),
	.combout(),
	.sumout(\resq[22]~65_sumout ),
	.cout(\resq[22]~66 ),
	.shareout(\resq[22]~67 ));
defparam \resq[22]~65 .extended_lut = "off";
defparam \resq[22]~65 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[22]~65 .shared_arith = "on";

arriav_lcell_comb \resq[23]~69 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][23]~q ),
	.datad(!dout_231),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[22]~66 ),
	.sharein(\resq[22]~67 ),
	.combout(),
	.sumout(\resq[23]~69_sumout ),
	.cout(\resq[23]~70 ),
	.shareout(\resq[23]~71 ));
defparam \resq[23]~69 .extended_lut = "off";
defparam \resq[23]~69 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[23]~69 .shared_arith = "on";

arriav_lcell_comb \resq[24]~73 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][24]~q ),
	.datad(!dout_241),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[23]~70 ),
	.sharein(\resq[23]~71 ),
	.combout(),
	.sumout(\resq[24]~73_sumout ),
	.cout(\resq[24]~74 ),
	.shareout(\resq[24]~75 ));
defparam \resq[24]~73 .extended_lut = "off";
defparam \resq[24]~73 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[24]~73 .shared_arith = "on";

arriav_lcell_comb \resq[25]~77 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][25]~q ),
	.datad(!dout_251),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[24]~74 ),
	.sharein(\resq[24]~75 ),
	.combout(),
	.sumout(\resq[25]~77_sumout ),
	.cout(\resq[25]~78 ),
	.shareout(\resq[25]~79 ));
defparam \resq[25]~77 .extended_lut = "off";
defparam \resq[25]~77 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[25]~77 .shared_arith = "on";

arriav_lcell_comb \resq[26]~81 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][26]~q ),
	.datad(!dout_261),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[25]~78 ),
	.sharein(\resq[25]~79 ),
	.combout(),
	.sumout(\resq[26]~81_sumout ),
	.cout(\resq[26]~82 ),
	.shareout(\resq[26]~83 ));
defparam \resq[26]~81 .extended_lut = "off";
defparam \resq[26]~81 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[26]~81 .shared_arith = "on";

arriav_lcell_comb \resq[27]~85 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][27]~q ),
	.datad(!dout_271),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[26]~82 ),
	.sharein(\resq[26]~83 ),
	.combout(),
	.sumout(\resq[27]~85_sumout ),
	.cout(\resq[27]~86 ),
	.shareout(\resq[27]~87 ));
defparam \resq[27]~85 .extended_lut = "off";
defparam \resq[27]~85 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[27]~85 .shared_arith = "on";

arriav_lcell_comb \resq[28]~89 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][28]~q ),
	.datad(!dout_281),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[27]~86 ),
	.sharein(\resq[27]~87 ),
	.combout(),
	.sumout(\resq[28]~89_sumout ),
	.cout(\resq[28]~90 ),
	.shareout(\resq[28]~91 ));
defparam \resq[28]~89 .extended_lut = "off";
defparam \resq[28]~89 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[28]~89 .shared_arith = "on";

arriav_lcell_comb \resq[29]~93 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][29]~q ),
	.datad(!dout_291),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[28]~90 ),
	.sharein(\resq[28]~91 ),
	.combout(),
	.sumout(\resq[29]~93_sumout ),
	.cout(\resq[29]~94 ),
	.shareout(\resq[29]~95 ));
defparam \resq[29]~93 .extended_lut = "off";
defparam \resq[29]~93 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[29]~93 .shared_arith = "on";

arriav_lcell_comb \resq[30]~97 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][30]~q ),
	.datad(!dout_301),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[29]~94 ),
	.sharein(\resq[29]~95 ),
	.combout(),
	.sumout(\resq[30]~97_sumout ),
	.cout(\resq[30]~98 ),
	.shareout(\resq[30]~99 ));
defparam \resq[30]~97 .extended_lut = "off";
defparam \resq[30]~97 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[30]~97 .shared_arith = "on";

arriav_lcell_comb \resq[31]~101 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][31]~q ),
	.datad(!dout_311),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[30]~98 ),
	.sharein(\resq[30]~99 ),
	.combout(),
	.sumout(\resq[31]~101_sumout ),
	.cout(\resq[31]~102 ),
	.shareout(\resq[31]~103 ));
defparam \resq[31]~101 .extended_lut = "off";
defparam \resq[31]~101 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[31]~101 .shared_arith = "on";

arriav_lcell_comb \resq[32]~105 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][32]~q ),
	.datad(!dout_321),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[31]~102 ),
	.sharein(\resq[31]~103 ),
	.combout(),
	.sumout(\resq[32]~105_sumout ),
	.cout(\resq[32]~106 ),
	.shareout(\resq[32]~107 ));
defparam \resq[32]~105 .extended_lut = "off";
defparam \resq[32]~105 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[32]~105 .shared_arith = "on";

arriav_lcell_comb \resq[33]~109 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][33]~q ),
	.datad(!dout_331),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[32]~106 ),
	.sharein(\resq[32]~107 ),
	.combout(),
	.sumout(\resq[33]~109_sumout ),
	.cout(),
	.shareout());
defparam \resq[33]~109 .extended_lut = "off";
defparam \resq[33]~109 .lut_mask = 64'h0000000000000FF0;
defparam \resq[33]~109 .shared_arith = "on";

endmodule

module cic_auk_dspip_delay_4 (
	datain,
	register_fifofifo_data06,
	register_fifofifo_data07,
	register_fifofifo_data08,
	register_fifofifo_data09,
	register_fifofifo_data010,
	register_fifofifo_data011,
	register_fifofifo_data012,
	register_fifofifo_data013,
	register_fifofifo_data014,
	register_fifofifo_data015,
	register_fifofifo_data016,
	register_fifofifo_data017,
	register_fifofifo_data018,
	register_fifofifo_data019,
	register_fifofifo_data020,
	register_fifofifo_data021,
	register_fifofifo_data022,
	register_fifofifo_data023,
	register_fifofifo_data024,
	register_fifofifo_data025,
	register_fifofifo_data026,
	register_fifofifo_data027,
	register_fifofifo_data028,
	register_fifofifo_data029,
	register_fifofifo_data030,
	register_fifofifo_data031,
	register_fifofifo_data032,
	register_fifofifo_data033,
	enable,
	register_fifofifo_data05,
	register_fifofifo_data04,
	register_fifofifo_data03,
	register_fifofifo_data02,
	register_fifofifo_data01,
	register_fifofifo_data00,
	clk,
	reset)/* synthesis synthesis_greybox=1 */;
input 	[46:0] datain;
output 	register_fifofifo_data06;
output 	register_fifofifo_data07;
output 	register_fifofifo_data08;
output 	register_fifofifo_data09;
output 	register_fifofifo_data010;
output 	register_fifofifo_data011;
output 	register_fifofifo_data012;
output 	register_fifofifo_data013;
output 	register_fifofifo_data014;
output 	register_fifofifo_data015;
output 	register_fifofifo_data016;
output 	register_fifofifo_data017;
output 	register_fifofifo_data018;
output 	register_fifofifo_data019;
output 	register_fifofifo_data020;
output 	register_fifofifo_data021;
output 	register_fifofifo_data022;
output 	register_fifofifo_data023;
output 	register_fifofifo_data024;
output 	register_fifofifo_data025;
output 	register_fifofifo_data026;
output 	register_fifofifo_data027;
output 	register_fifofifo_data028;
output 	register_fifofifo_data029;
output 	register_fifofifo_data030;
output 	register_fifofifo_data031;
output 	register_fifofifo_data032;
output 	register_fifofifo_data033;
input 	enable;
output 	register_fifofifo_data05;
output 	register_fifofifo_data04;
output 	register_fifofifo_data03;
output 	register_fifofifo_data02;
output 	register_fifofifo_data01;
output 	register_fifofifo_data00;
input 	clk;
input 	reset;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \register_fifo:fifo_data[0][6] (
	.clk(clk),
	.d(datain[6]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data06),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][6] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][6] .power_up = "low";

dffeas \register_fifo:fifo_data[0][7] (
	.clk(clk),
	.d(datain[7]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data07),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][7] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][7] .power_up = "low";

dffeas \register_fifo:fifo_data[0][8] (
	.clk(clk),
	.d(datain[8]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data08),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][8] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][8] .power_up = "low";

dffeas \register_fifo:fifo_data[0][9] (
	.clk(clk),
	.d(datain[9]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data09),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][9] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][9] .power_up = "low";

dffeas \register_fifo:fifo_data[0][10] (
	.clk(clk),
	.d(datain[10]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data010),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][10] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][10] .power_up = "low";

dffeas \register_fifo:fifo_data[0][11] (
	.clk(clk),
	.d(datain[11]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data011),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][11] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][11] .power_up = "low";

dffeas \register_fifo:fifo_data[0][12] (
	.clk(clk),
	.d(datain[12]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data012),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][12] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][12] .power_up = "low";

dffeas \register_fifo:fifo_data[0][13] (
	.clk(clk),
	.d(datain[13]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data013),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][13] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][13] .power_up = "low";

dffeas \register_fifo:fifo_data[0][14] (
	.clk(clk),
	.d(datain[14]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data014),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][14] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][14] .power_up = "low";

dffeas \register_fifo:fifo_data[0][15] (
	.clk(clk),
	.d(datain[15]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data015),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][15] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][15] .power_up = "low";

dffeas \register_fifo:fifo_data[0][16] (
	.clk(clk),
	.d(datain[16]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data016),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][16] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][16] .power_up = "low";

dffeas \register_fifo:fifo_data[0][17] (
	.clk(clk),
	.d(datain[17]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data017),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][17] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][17] .power_up = "low";

dffeas \register_fifo:fifo_data[0][18] (
	.clk(clk),
	.d(datain[18]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data018),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][18] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][18] .power_up = "low";

dffeas \register_fifo:fifo_data[0][19] (
	.clk(clk),
	.d(datain[19]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data019),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][19] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][19] .power_up = "low";

dffeas \register_fifo:fifo_data[0][20] (
	.clk(clk),
	.d(datain[20]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data020),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][20] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][20] .power_up = "low";

dffeas \register_fifo:fifo_data[0][21] (
	.clk(clk),
	.d(datain[21]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data021),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][21] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][21] .power_up = "low";

dffeas \register_fifo:fifo_data[0][22] (
	.clk(clk),
	.d(datain[22]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data022),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][22] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][22] .power_up = "low";

dffeas \register_fifo:fifo_data[0][23] (
	.clk(clk),
	.d(datain[23]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data023),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][23] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][23] .power_up = "low";

dffeas \register_fifo:fifo_data[0][24] (
	.clk(clk),
	.d(datain[24]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data024),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][24] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][24] .power_up = "low";

dffeas \register_fifo:fifo_data[0][25] (
	.clk(clk),
	.d(datain[25]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data025),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][25] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][25] .power_up = "low";

dffeas \register_fifo:fifo_data[0][26] (
	.clk(clk),
	.d(datain[26]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data026),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][26] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][26] .power_up = "low";

dffeas \register_fifo:fifo_data[0][27] (
	.clk(clk),
	.d(datain[27]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data027),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][27] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][27] .power_up = "low";

dffeas \register_fifo:fifo_data[0][28] (
	.clk(clk),
	.d(datain[28]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data028),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][28] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][28] .power_up = "low";

dffeas \register_fifo:fifo_data[0][29] (
	.clk(clk),
	.d(datain[29]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data029),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][29] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][29] .power_up = "low";

dffeas \register_fifo:fifo_data[0][30] (
	.clk(clk),
	.d(datain[30]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data030),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][30] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][30] .power_up = "low";

dffeas \register_fifo:fifo_data[0][31] (
	.clk(clk),
	.d(datain[31]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data031),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][31] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][31] .power_up = "low";

dffeas \register_fifo:fifo_data[0][32] (
	.clk(clk),
	.d(datain[32]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data032),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][32] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][32] .power_up = "low";

dffeas \register_fifo:fifo_data[0][33] (
	.clk(clk),
	.d(datain[33]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data033),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][33] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][33] .power_up = "low";

dffeas \register_fifo:fifo_data[0][5] (
	.clk(clk),
	.d(datain[5]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data05),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][5] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][5] .power_up = "low";

dffeas \register_fifo:fifo_data[0][4] (
	.clk(clk),
	.d(datain[4]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data04),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][4] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][4] .power_up = "low";

dffeas \register_fifo:fifo_data[0][3] (
	.clk(clk),
	.d(datain[3]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data03),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][3] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][3] .power_up = "low";

dffeas \register_fifo:fifo_data[0][2] (
	.clk(clk),
	.d(datain[2]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data02),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][2] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][2] .power_up = "low";

dffeas \register_fifo:fifo_data[0][1] (
	.clk(clk),
	.d(datain[1]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data01),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][1] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][1] .power_up = "low";

dffeas \register_fifo:fifo_data[0][0] (
	.clk(clk),
	.d(datain[0]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data00),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][0] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][0] .power_up = "low";

endmodule

module cic_auk_dspip_differentiator_5 (
	dout_valid1,
	dout_valid2,
	dout_5,
	dout_6,
	dout_7,
	dout_8,
	dout_9,
	dout_10,
	dout_11,
	dout_12,
	dout_13,
	dout_14,
	dout_15,
	dout_16,
	dout_17,
	dout_18,
	dout_19,
	dout_20,
	dout_21,
	dout_22,
	dout_23,
	dout_24,
	dout_25,
	dout_26,
	dout_27,
	dout_28,
	dout_29,
	dout_30,
	dout_31,
	dout_32,
	dout_4,
	dout_61,
	dout_3,
	dout_71,
	dout_81,
	dout_91,
	dout_101,
	dout_111,
	dout_121,
	dout_131,
	dout_141,
	dout_151,
	dout_161,
	dout_171,
	dout_181,
	dout_191,
	dout_201,
	dout_211,
	dout_221,
	dout_231,
	dout_241,
	dout_251,
	dout_261,
	dout_271,
	dout_281,
	dout_291,
	dout_301,
	dout_311,
	dout_321,
	dout_33,
	dout_51,
	dout_2,
	dout_41,
	dout_1,
	dout_34,
	dout_210,
	dout_110,
	stall_reg,
	dout_valid3,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	dout_valid1;
input 	dout_valid2;
output 	dout_5;
output 	dout_6;
output 	dout_7;
output 	dout_8;
output 	dout_9;
output 	dout_10;
output 	dout_11;
output 	dout_12;
output 	dout_13;
output 	dout_14;
output 	dout_15;
output 	dout_16;
output 	dout_17;
output 	dout_18;
output 	dout_19;
output 	dout_20;
output 	dout_21;
output 	dout_22;
output 	dout_23;
output 	dout_24;
output 	dout_25;
output 	dout_26;
output 	dout_27;
output 	dout_28;
output 	dout_29;
output 	dout_30;
output 	dout_31;
output 	dout_32;
output 	dout_4;
input 	dout_61;
output 	dout_3;
input 	dout_71;
input 	dout_81;
input 	dout_91;
input 	dout_101;
input 	dout_111;
input 	dout_121;
input 	dout_131;
input 	dout_141;
input 	dout_151;
input 	dout_161;
input 	dout_171;
input 	dout_181;
input 	dout_191;
input 	dout_201;
input 	dout_211;
input 	dout_221;
input 	dout_231;
input 	dout_241;
input 	dout_251;
input 	dout_261;
input 	dout_271;
input 	dout_281;
input 	dout_291;
input 	dout_301;
input 	dout_311;
input 	dout_321;
input 	dout_33;
input 	dout_51;
output 	dout_2;
input 	dout_41;
output 	dout_1;
input 	dout_34;
input 	dout_210;
input 	dout_110;
input 	stall_reg;
input 	dout_valid3;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \glogic:u0|register_fifo:fifo_data[0][5]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][6]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][7]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][8]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][9]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][10]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][11]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][12]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][13]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][14]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][15]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][16]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][17]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][18]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][19]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][20]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][21]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][22]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][23]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][24]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][25]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][26]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][27]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][28]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][29]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][30]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][31]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][32]~q ;
wire \dout~1_combout ;
wire \glogic:u0|register_fifo:fifo_data[0][4]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][3]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][2]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][1]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][0]~q ;
wire \resq[0]~130_cout ;
wire \resq[0]~131 ;
wire \resq[1]~126 ;
wire \resq[1]~127 ;
wire \resq[2]~122 ;
wire \resq[2]~123 ;
wire \resq[3]~118 ;
wire \resq[3]~119 ;
wire \resq[4]~114 ;
wire \resq[4]~115 ;
wire \resq[5]~1_sumout ;
wire \dout[29]~0_combout ;
wire \resq[5]~2 ;
wire \resq[5]~3 ;
wire \resq[6]~5_sumout ;
wire \resq[6]~6 ;
wire \resq[6]~7 ;
wire \resq[7]~9_sumout ;
wire \resq[7]~10 ;
wire \resq[7]~11 ;
wire \resq[8]~13_sumout ;
wire \resq[8]~14 ;
wire \resq[8]~15 ;
wire \resq[9]~17_sumout ;
wire \resq[9]~18 ;
wire \resq[9]~19 ;
wire \resq[10]~21_sumout ;
wire \resq[10]~22 ;
wire \resq[10]~23 ;
wire \resq[11]~25_sumout ;
wire \resq[11]~26 ;
wire \resq[11]~27 ;
wire \resq[12]~29_sumout ;
wire \resq[12]~30 ;
wire \resq[12]~31 ;
wire \resq[13]~33_sumout ;
wire \resq[13]~34 ;
wire \resq[13]~35 ;
wire \resq[14]~37_sumout ;
wire \resq[14]~38 ;
wire \resq[14]~39 ;
wire \resq[15]~41_sumout ;
wire \resq[15]~42 ;
wire \resq[15]~43 ;
wire \resq[16]~45_sumout ;
wire \resq[16]~46 ;
wire \resq[16]~47 ;
wire \resq[17]~49_sumout ;
wire \resq[17]~50 ;
wire \resq[17]~51 ;
wire \resq[18]~53_sumout ;
wire \resq[18]~54 ;
wire \resq[18]~55 ;
wire \resq[19]~57_sumout ;
wire \resq[19]~58 ;
wire \resq[19]~59 ;
wire \resq[20]~61_sumout ;
wire \resq[20]~62 ;
wire \resq[20]~63 ;
wire \resq[21]~65_sumout ;
wire \resq[21]~66 ;
wire \resq[21]~67 ;
wire \resq[22]~69_sumout ;
wire \resq[22]~70 ;
wire \resq[22]~71 ;
wire \resq[23]~73_sumout ;
wire \resq[23]~74 ;
wire \resq[23]~75 ;
wire \resq[24]~77_sumout ;
wire \resq[24]~78 ;
wire \resq[24]~79 ;
wire \resq[25]~81_sumout ;
wire \resq[25]~82 ;
wire \resq[25]~83 ;
wire \resq[26]~85_sumout ;
wire \resq[26]~86 ;
wire \resq[26]~87 ;
wire \resq[27]~89_sumout ;
wire \resq[27]~90 ;
wire \resq[27]~91 ;
wire \resq[28]~93_sumout ;
wire \resq[28]~94 ;
wire \resq[28]~95 ;
wire \resq[29]~97_sumout ;
wire \resq[29]~98 ;
wire \resq[29]~99 ;
wire \resq[30]~101_sumout ;
wire \resq[30]~102 ;
wire \resq[30]~103 ;
wire \resq[31]~105_sumout ;
wire \resq[31]~106 ;
wire \resq[31]~107 ;
wire \resq[32]~109_sumout ;
wire \resq[4]~113_sumout ;
wire \resq[3]~117_sumout ;
wire \resq[2]~121_sumout ;
wire \resq[1]~125_sumout ;


cic_auk_dspip_delay_5 \glogic:u0 (
	.datain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,dout_33,dout_321,dout_311,dout_301,dout_291,dout_281,dout_271,dout_261,dout_251,dout_241,dout_231,dout_221,dout_211,dout_201,dout_191,dout_181,dout_171,dout_161,dout_151,dout_141,dout_131,dout_121,dout_111,dout_101,dout_91,dout_81,dout_71,
dout_61,dout_51,dout_41,dout_34,dout_210,dout_110}),
	.register_fifofifo_data05(\glogic:u0|register_fifo:fifo_data[0][5]~q ),
	.register_fifofifo_data06(\glogic:u0|register_fifo:fifo_data[0][6]~q ),
	.register_fifofifo_data07(\glogic:u0|register_fifo:fifo_data[0][7]~q ),
	.register_fifofifo_data08(\glogic:u0|register_fifo:fifo_data[0][8]~q ),
	.register_fifofifo_data09(\glogic:u0|register_fifo:fifo_data[0][9]~q ),
	.register_fifofifo_data010(\glogic:u0|register_fifo:fifo_data[0][10]~q ),
	.register_fifofifo_data011(\glogic:u0|register_fifo:fifo_data[0][11]~q ),
	.register_fifofifo_data012(\glogic:u0|register_fifo:fifo_data[0][12]~q ),
	.register_fifofifo_data013(\glogic:u0|register_fifo:fifo_data[0][13]~q ),
	.register_fifofifo_data014(\glogic:u0|register_fifo:fifo_data[0][14]~q ),
	.register_fifofifo_data015(\glogic:u0|register_fifo:fifo_data[0][15]~q ),
	.register_fifofifo_data016(\glogic:u0|register_fifo:fifo_data[0][16]~q ),
	.register_fifofifo_data017(\glogic:u0|register_fifo:fifo_data[0][17]~q ),
	.register_fifofifo_data018(\glogic:u0|register_fifo:fifo_data[0][18]~q ),
	.register_fifofifo_data019(\glogic:u0|register_fifo:fifo_data[0][19]~q ),
	.register_fifofifo_data020(\glogic:u0|register_fifo:fifo_data[0][20]~q ),
	.register_fifofifo_data021(\glogic:u0|register_fifo:fifo_data[0][21]~q ),
	.register_fifofifo_data022(\glogic:u0|register_fifo:fifo_data[0][22]~q ),
	.register_fifofifo_data023(\glogic:u0|register_fifo:fifo_data[0][23]~q ),
	.register_fifofifo_data024(\glogic:u0|register_fifo:fifo_data[0][24]~q ),
	.register_fifofifo_data025(\glogic:u0|register_fifo:fifo_data[0][25]~q ),
	.register_fifofifo_data026(\glogic:u0|register_fifo:fifo_data[0][26]~q ),
	.register_fifofifo_data027(\glogic:u0|register_fifo:fifo_data[0][27]~q ),
	.register_fifofifo_data028(\glogic:u0|register_fifo:fifo_data[0][28]~q ),
	.register_fifofifo_data029(\glogic:u0|register_fifo:fifo_data[0][29]~q ),
	.register_fifofifo_data030(\glogic:u0|register_fifo:fifo_data[0][30]~q ),
	.register_fifofifo_data031(\glogic:u0|register_fifo:fifo_data[0][31]~q ),
	.register_fifofifo_data032(\glogic:u0|register_fifo:fifo_data[0][32]~q ),
	.enable(\dout~1_combout ),
	.register_fifofifo_data04(\glogic:u0|register_fifo:fifo_data[0][4]~q ),
	.register_fifofifo_data03(\glogic:u0|register_fifo:fifo_data[0][3]~q ),
	.register_fifofifo_data02(\glogic:u0|register_fifo:fifo_data[0][2]~q ),
	.register_fifofifo_data01(\glogic:u0|register_fifo:fifo_data[0][1]~q ),
	.register_fifofifo_data00(\glogic:u0|register_fifo:fifo_data[0][0]~q ),
	.clk(clk),
	.reset(reset_n));

arriav_lcell_comb \dout~1 (
	.dataa(!stall_reg),
	.datab(!dout_valid2),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dout~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dout~1 .extended_lut = "off";
defparam \dout~1 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \dout~1 .shared_arith = "off";

dffeas dout_valid(
	.clk(clk),
	.d(dout_valid2),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(dout_valid3),
	.q(dout_valid1),
	.prn(vcc));
defparam dout_valid.is_wysiwyg = "true";
defparam dout_valid.power_up = "low";

dffeas \dout[5] (
	.clk(clk),
	.d(\resq[5]~1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[29]~0_combout ),
	.q(dout_5),
	.prn(vcc));
defparam \dout[5] .is_wysiwyg = "true";
defparam \dout[5] .power_up = "low";

dffeas \dout[6] (
	.clk(clk),
	.d(\resq[6]~5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[29]~0_combout ),
	.q(dout_6),
	.prn(vcc));
defparam \dout[6] .is_wysiwyg = "true";
defparam \dout[6] .power_up = "low";

dffeas \dout[7] (
	.clk(clk),
	.d(\resq[7]~9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[29]~0_combout ),
	.q(dout_7),
	.prn(vcc));
defparam \dout[7] .is_wysiwyg = "true";
defparam \dout[7] .power_up = "low";

dffeas \dout[8] (
	.clk(clk),
	.d(\resq[8]~13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[29]~0_combout ),
	.q(dout_8),
	.prn(vcc));
defparam \dout[8] .is_wysiwyg = "true";
defparam \dout[8] .power_up = "low";

dffeas \dout[9] (
	.clk(clk),
	.d(\resq[9]~17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[29]~0_combout ),
	.q(dout_9),
	.prn(vcc));
defparam \dout[9] .is_wysiwyg = "true";
defparam \dout[9] .power_up = "low";

dffeas \dout[10] (
	.clk(clk),
	.d(\resq[10]~21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[29]~0_combout ),
	.q(dout_10),
	.prn(vcc));
defparam \dout[10] .is_wysiwyg = "true";
defparam \dout[10] .power_up = "low";

dffeas \dout[11] (
	.clk(clk),
	.d(\resq[11]~25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[29]~0_combout ),
	.q(dout_11),
	.prn(vcc));
defparam \dout[11] .is_wysiwyg = "true";
defparam \dout[11] .power_up = "low";

dffeas \dout[12] (
	.clk(clk),
	.d(\resq[12]~29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[29]~0_combout ),
	.q(dout_12),
	.prn(vcc));
defparam \dout[12] .is_wysiwyg = "true";
defparam \dout[12] .power_up = "low";

dffeas \dout[13] (
	.clk(clk),
	.d(\resq[13]~33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[29]~0_combout ),
	.q(dout_13),
	.prn(vcc));
defparam \dout[13] .is_wysiwyg = "true";
defparam \dout[13] .power_up = "low";

dffeas \dout[14] (
	.clk(clk),
	.d(\resq[14]~37_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[29]~0_combout ),
	.q(dout_14),
	.prn(vcc));
defparam \dout[14] .is_wysiwyg = "true";
defparam \dout[14] .power_up = "low";

dffeas \dout[15] (
	.clk(clk),
	.d(\resq[15]~41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[29]~0_combout ),
	.q(dout_15),
	.prn(vcc));
defparam \dout[15] .is_wysiwyg = "true";
defparam \dout[15] .power_up = "low";

dffeas \dout[16] (
	.clk(clk),
	.d(\resq[16]~45_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[29]~0_combout ),
	.q(dout_16),
	.prn(vcc));
defparam \dout[16] .is_wysiwyg = "true";
defparam \dout[16] .power_up = "low";

dffeas \dout[17] (
	.clk(clk),
	.d(\resq[17]~49_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[29]~0_combout ),
	.q(dout_17),
	.prn(vcc));
defparam \dout[17] .is_wysiwyg = "true";
defparam \dout[17] .power_up = "low";

dffeas \dout[18] (
	.clk(clk),
	.d(\resq[18]~53_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[29]~0_combout ),
	.q(dout_18),
	.prn(vcc));
defparam \dout[18] .is_wysiwyg = "true";
defparam \dout[18] .power_up = "low";

dffeas \dout[19] (
	.clk(clk),
	.d(\resq[19]~57_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[29]~0_combout ),
	.q(dout_19),
	.prn(vcc));
defparam \dout[19] .is_wysiwyg = "true";
defparam \dout[19] .power_up = "low";

dffeas \dout[20] (
	.clk(clk),
	.d(\resq[20]~61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[29]~0_combout ),
	.q(dout_20),
	.prn(vcc));
defparam \dout[20] .is_wysiwyg = "true";
defparam \dout[20] .power_up = "low";

dffeas \dout[21] (
	.clk(clk),
	.d(\resq[21]~65_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[29]~0_combout ),
	.q(dout_21),
	.prn(vcc));
defparam \dout[21] .is_wysiwyg = "true";
defparam \dout[21] .power_up = "low";

dffeas \dout[22] (
	.clk(clk),
	.d(\resq[22]~69_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[29]~0_combout ),
	.q(dout_22),
	.prn(vcc));
defparam \dout[22] .is_wysiwyg = "true";
defparam \dout[22] .power_up = "low";

dffeas \dout[23] (
	.clk(clk),
	.d(\resq[23]~73_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[29]~0_combout ),
	.q(dout_23),
	.prn(vcc));
defparam \dout[23] .is_wysiwyg = "true";
defparam \dout[23] .power_up = "low";

dffeas \dout[24] (
	.clk(clk),
	.d(\resq[24]~77_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[29]~0_combout ),
	.q(dout_24),
	.prn(vcc));
defparam \dout[24] .is_wysiwyg = "true";
defparam \dout[24] .power_up = "low";

dffeas \dout[25] (
	.clk(clk),
	.d(\resq[25]~81_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[29]~0_combout ),
	.q(dout_25),
	.prn(vcc));
defparam \dout[25] .is_wysiwyg = "true";
defparam \dout[25] .power_up = "low";

dffeas \dout[26] (
	.clk(clk),
	.d(\resq[26]~85_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[29]~0_combout ),
	.q(dout_26),
	.prn(vcc));
defparam \dout[26] .is_wysiwyg = "true";
defparam \dout[26] .power_up = "low";

dffeas \dout[27] (
	.clk(clk),
	.d(\resq[27]~89_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[29]~0_combout ),
	.q(dout_27),
	.prn(vcc));
defparam \dout[27] .is_wysiwyg = "true";
defparam \dout[27] .power_up = "low";

dffeas \dout[28] (
	.clk(clk),
	.d(\resq[28]~93_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[29]~0_combout ),
	.q(dout_28),
	.prn(vcc));
defparam \dout[28] .is_wysiwyg = "true";
defparam \dout[28] .power_up = "low";

dffeas \dout[29] (
	.clk(clk),
	.d(\resq[29]~97_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[29]~0_combout ),
	.q(dout_29),
	.prn(vcc));
defparam \dout[29] .is_wysiwyg = "true";
defparam \dout[29] .power_up = "low";

dffeas \dout[30] (
	.clk(clk),
	.d(\resq[30]~101_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[29]~0_combout ),
	.q(dout_30),
	.prn(vcc));
defparam \dout[30] .is_wysiwyg = "true";
defparam \dout[30] .power_up = "low";

dffeas \dout[31] (
	.clk(clk),
	.d(\resq[31]~105_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[29]~0_combout ),
	.q(dout_31),
	.prn(vcc));
defparam \dout[31] .is_wysiwyg = "true";
defparam \dout[31] .power_up = "low";

dffeas \dout[32] (
	.clk(clk),
	.d(\resq[32]~109_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[29]~0_combout ),
	.q(dout_32),
	.prn(vcc));
defparam \dout[32] .is_wysiwyg = "true";
defparam \dout[32] .power_up = "low";

dffeas \dout[4] (
	.clk(clk),
	.d(\resq[4]~113_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[29]~0_combout ),
	.q(dout_4),
	.prn(vcc));
defparam \dout[4] .is_wysiwyg = "true";
defparam \dout[4] .power_up = "low";

dffeas \dout[3] (
	.clk(clk),
	.d(\resq[3]~117_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[29]~0_combout ),
	.q(dout_3),
	.prn(vcc));
defparam \dout[3] .is_wysiwyg = "true";
defparam \dout[3] .power_up = "low";

dffeas \dout[2] (
	.clk(clk),
	.d(\resq[2]~121_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[29]~0_combout ),
	.q(dout_2),
	.prn(vcc));
defparam \dout[2] .is_wysiwyg = "true";
defparam \dout[2] .power_up = "low";

dffeas \dout[1] (
	.clk(clk),
	.d(\resq[1]~125_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[29]~0_combout ),
	.q(dout_1),
	.prn(vcc));
defparam \dout[1] .is_wysiwyg = "true";
defparam \dout[1] .power_up = "low";

arriav_lcell_comb \resq[0]~130 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][0]~q ),
	.datad(!dout_110),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\resq[0]~130_cout ),
	.shareout(\resq[0]~131 ));
defparam \resq[0]~130 .extended_lut = "off";
defparam \resq[0]~130 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[0]~130 .shared_arith = "on";

arriav_lcell_comb \resq[1]~125 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][1]~q ),
	.datad(!dout_210),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[0]~130_cout ),
	.sharein(\resq[0]~131 ),
	.combout(),
	.sumout(\resq[1]~125_sumout ),
	.cout(\resq[1]~126 ),
	.shareout(\resq[1]~127 ));
defparam \resq[1]~125 .extended_lut = "off";
defparam \resq[1]~125 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[1]~125 .shared_arith = "on";

arriav_lcell_comb \resq[2]~121 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][2]~q ),
	.datad(!dout_34),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[1]~126 ),
	.sharein(\resq[1]~127 ),
	.combout(),
	.sumout(\resq[2]~121_sumout ),
	.cout(\resq[2]~122 ),
	.shareout(\resq[2]~123 ));
defparam \resq[2]~121 .extended_lut = "off";
defparam \resq[2]~121 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[2]~121 .shared_arith = "on";

arriav_lcell_comb \resq[3]~117 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][3]~q ),
	.datad(!dout_41),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[2]~122 ),
	.sharein(\resq[2]~123 ),
	.combout(),
	.sumout(\resq[3]~117_sumout ),
	.cout(\resq[3]~118 ),
	.shareout(\resq[3]~119 ));
defparam \resq[3]~117 .extended_lut = "off";
defparam \resq[3]~117 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[3]~117 .shared_arith = "on";

arriav_lcell_comb \resq[4]~113 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][4]~q ),
	.datad(!dout_51),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[3]~118 ),
	.sharein(\resq[3]~119 ),
	.combout(),
	.sumout(\resq[4]~113_sumout ),
	.cout(\resq[4]~114 ),
	.shareout(\resq[4]~115 ));
defparam \resq[4]~113 .extended_lut = "off";
defparam \resq[4]~113 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[4]~113 .shared_arith = "on";

arriav_lcell_comb \resq[5]~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][5]~q ),
	.datad(!dout_61),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[4]~114 ),
	.sharein(\resq[4]~115 ),
	.combout(),
	.sumout(\resq[5]~1_sumout ),
	.cout(\resq[5]~2 ),
	.shareout(\resq[5]~3 ));
defparam \resq[5]~1 .extended_lut = "off";
defparam \resq[5]~1 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[5]~1 .shared_arith = "on";

arriav_lcell_comb \dout[29]~0 (
	.dataa(!reset_n),
	.datab(!stall_reg),
	.datac(!dout_valid2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dout[29]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dout[29]~0 .extended_lut = "off";
defparam \dout[29]~0 .lut_mask = 64'hEFEFEFEFEFEFEFEF;
defparam \dout[29]~0 .shared_arith = "off";

arriav_lcell_comb \resq[6]~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][6]~q ),
	.datad(!dout_71),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[5]~2 ),
	.sharein(\resq[5]~3 ),
	.combout(),
	.sumout(\resq[6]~5_sumout ),
	.cout(\resq[6]~6 ),
	.shareout(\resq[6]~7 ));
defparam \resq[6]~5 .extended_lut = "off";
defparam \resq[6]~5 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[6]~5 .shared_arith = "on";

arriav_lcell_comb \resq[7]~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][7]~q ),
	.datad(!dout_81),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[6]~6 ),
	.sharein(\resq[6]~7 ),
	.combout(),
	.sumout(\resq[7]~9_sumout ),
	.cout(\resq[7]~10 ),
	.shareout(\resq[7]~11 ));
defparam \resq[7]~9 .extended_lut = "off";
defparam \resq[7]~9 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[7]~9 .shared_arith = "on";

arriav_lcell_comb \resq[8]~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][8]~q ),
	.datad(!dout_91),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[7]~10 ),
	.sharein(\resq[7]~11 ),
	.combout(),
	.sumout(\resq[8]~13_sumout ),
	.cout(\resq[8]~14 ),
	.shareout(\resq[8]~15 ));
defparam \resq[8]~13 .extended_lut = "off";
defparam \resq[8]~13 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[8]~13 .shared_arith = "on";

arriav_lcell_comb \resq[9]~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][9]~q ),
	.datad(!dout_101),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[8]~14 ),
	.sharein(\resq[8]~15 ),
	.combout(),
	.sumout(\resq[9]~17_sumout ),
	.cout(\resq[9]~18 ),
	.shareout(\resq[9]~19 ));
defparam \resq[9]~17 .extended_lut = "off";
defparam \resq[9]~17 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[9]~17 .shared_arith = "on";

arriav_lcell_comb \resq[10]~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][10]~q ),
	.datad(!dout_111),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[9]~18 ),
	.sharein(\resq[9]~19 ),
	.combout(),
	.sumout(\resq[10]~21_sumout ),
	.cout(\resq[10]~22 ),
	.shareout(\resq[10]~23 ));
defparam \resq[10]~21 .extended_lut = "off";
defparam \resq[10]~21 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[10]~21 .shared_arith = "on";

arriav_lcell_comb \resq[11]~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][11]~q ),
	.datad(!dout_121),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[10]~22 ),
	.sharein(\resq[10]~23 ),
	.combout(),
	.sumout(\resq[11]~25_sumout ),
	.cout(\resq[11]~26 ),
	.shareout(\resq[11]~27 ));
defparam \resq[11]~25 .extended_lut = "off";
defparam \resq[11]~25 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[11]~25 .shared_arith = "on";

arriav_lcell_comb \resq[12]~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][12]~q ),
	.datad(!dout_131),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[11]~26 ),
	.sharein(\resq[11]~27 ),
	.combout(),
	.sumout(\resq[12]~29_sumout ),
	.cout(\resq[12]~30 ),
	.shareout(\resq[12]~31 ));
defparam \resq[12]~29 .extended_lut = "off";
defparam \resq[12]~29 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[12]~29 .shared_arith = "on";

arriav_lcell_comb \resq[13]~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][13]~q ),
	.datad(!dout_141),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[12]~30 ),
	.sharein(\resq[12]~31 ),
	.combout(),
	.sumout(\resq[13]~33_sumout ),
	.cout(\resq[13]~34 ),
	.shareout(\resq[13]~35 ));
defparam \resq[13]~33 .extended_lut = "off";
defparam \resq[13]~33 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[13]~33 .shared_arith = "on";

arriav_lcell_comb \resq[14]~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][14]~q ),
	.datad(!dout_151),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[13]~34 ),
	.sharein(\resq[13]~35 ),
	.combout(),
	.sumout(\resq[14]~37_sumout ),
	.cout(\resq[14]~38 ),
	.shareout(\resq[14]~39 ));
defparam \resq[14]~37 .extended_lut = "off";
defparam \resq[14]~37 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[14]~37 .shared_arith = "on";

arriav_lcell_comb \resq[15]~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][15]~q ),
	.datad(!dout_161),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[14]~38 ),
	.sharein(\resq[14]~39 ),
	.combout(),
	.sumout(\resq[15]~41_sumout ),
	.cout(\resq[15]~42 ),
	.shareout(\resq[15]~43 ));
defparam \resq[15]~41 .extended_lut = "off";
defparam \resq[15]~41 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[15]~41 .shared_arith = "on";

arriav_lcell_comb \resq[16]~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][16]~q ),
	.datad(!dout_171),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[15]~42 ),
	.sharein(\resq[15]~43 ),
	.combout(),
	.sumout(\resq[16]~45_sumout ),
	.cout(\resq[16]~46 ),
	.shareout(\resq[16]~47 ));
defparam \resq[16]~45 .extended_lut = "off";
defparam \resq[16]~45 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[16]~45 .shared_arith = "on";

arriav_lcell_comb \resq[17]~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][17]~q ),
	.datad(!dout_181),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[16]~46 ),
	.sharein(\resq[16]~47 ),
	.combout(),
	.sumout(\resq[17]~49_sumout ),
	.cout(\resq[17]~50 ),
	.shareout(\resq[17]~51 ));
defparam \resq[17]~49 .extended_lut = "off";
defparam \resq[17]~49 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[17]~49 .shared_arith = "on";

arriav_lcell_comb \resq[18]~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][18]~q ),
	.datad(!dout_191),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[17]~50 ),
	.sharein(\resq[17]~51 ),
	.combout(),
	.sumout(\resq[18]~53_sumout ),
	.cout(\resq[18]~54 ),
	.shareout(\resq[18]~55 ));
defparam \resq[18]~53 .extended_lut = "off";
defparam \resq[18]~53 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[18]~53 .shared_arith = "on";

arriav_lcell_comb \resq[19]~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][19]~q ),
	.datad(!dout_201),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[18]~54 ),
	.sharein(\resq[18]~55 ),
	.combout(),
	.sumout(\resq[19]~57_sumout ),
	.cout(\resq[19]~58 ),
	.shareout(\resq[19]~59 ));
defparam \resq[19]~57 .extended_lut = "off";
defparam \resq[19]~57 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[19]~57 .shared_arith = "on";

arriav_lcell_comb \resq[20]~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][20]~q ),
	.datad(!dout_211),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[19]~58 ),
	.sharein(\resq[19]~59 ),
	.combout(),
	.sumout(\resq[20]~61_sumout ),
	.cout(\resq[20]~62 ),
	.shareout(\resq[20]~63 ));
defparam \resq[20]~61 .extended_lut = "off";
defparam \resq[20]~61 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[20]~61 .shared_arith = "on";

arriav_lcell_comb \resq[21]~65 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][21]~q ),
	.datad(!dout_221),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[20]~62 ),
	.sharein(\resq[20]~63 ),
	.combout(),
	.sumout(\resq[21]~65_sumout ),
	.cout(\resq[21]~66 ),
	.shareout(\resq[21]~67 ));
defparam \resq[21]~65 .extended_lut = "off";
defparam \resq[21]~65 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[21]~65 .shared_arith = "on";

arriav_lcell_comb \resq[22]~69 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][22]~q ),
	.datad(!dout_231),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[21]~66 ),
	.sharein(\resq[21]~67 ),
	.combout(),
	.sumout(\resq[22]~69_sumout ),
	.cout(\resq[22]~70 ),
	.shareout(\resq[22]~71 ));
defparam \resq[22]~69 .extended_lut = "off";
defparam \resq[22]~69 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[22]~69 .shared_arith = "on";

arriav_lcell_comb \resq[23]~73 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][23]~q ),
	.datad(!dout_241),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[22]~70 ),
	.sharein(\resq[22]~71 ),
	.combout(),
	.sumout(\resq[23]~73_sumout ),
	.cout(\resq[23]~74 ),
	.shareout(\resq[23]~75 ));
defparam \resq[23]~73 .extended_lut = "off";
defparam \resq[23]~73 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[23]~73 .shared_arith = "on";

arriav_lcell_comb \resq[24]~77 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][24]~q ),
	.datad(!dout_251),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[23]~74 ),
	.sharein(\resq[23]~75 ),
	.combout(),
	.sumout(\resq[24]~77_sumout ),
	.cout(\resq[24]~78 ),
	.shareout(\resq[24]~79 ));
defparam \resq[24]~77 .extended_lut = "off";
defparam \resq[24]~77 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[24]~77 .shared_arith = "on";

arriav_lcell_comb \resq[25]~81 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][25]~q ),
	.datad(!dout_261),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[24]~78 ),
	.sharein(\resq[24]~79 ),
	.combout(),
	.sumout(\resq[25]~81_sumout ),
	.cout(\resq[25]~82 ),
	.shareout(\resq[25]~83 ));
defparam \resq[25]~81 .extended_lut = "off";
defparam \resq[25]~81 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[25]~81 .shared_arith = "on";

arriav_lcell_comb \resq[26]~85 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][26]~q ),
	.datad(!dout_271),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[25]~82 ),
	.sharein(\resq[25]~83 ),
	.combout(),
	.sumout(\resq[26]~85_sumout ),
	.cout(\resq[26]~86 ),
	.shareout(\resq[26]~87 ));
defparam \resq[26]~85 .extended_lut = "off";
defparam \resq[26]~85 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[26]~85 .shared_arith = "on";

arriav_lcell_comb \resq[27]~89 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][27]~q ),
	.datad(!dout_281),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[26]~86 ),
	.sharein(\resq[26]~87 ),
	.combout(),
	.sumout(\resq[27]~89_sumout ),
	.cout(\resq[27]~90 ),
	.shareout(\resq[27]~91 ));
defparam \resq[27]~89 .extended_lut = "off";
defparam \resq[27]~89 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[27]~89 .shared_arith = "on";

arriav_lcell_comb \resq[28]~93 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][28]~q ),
	.datad(!dout_291),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[27]~90 ),
	.sharein(\resq[27]~91 ),
	.combout(),
	.sumout(\resq[28]~93_sumout ),
	.cout(\resq[28]~94 ),
	.shareout(\resq[28]~95 ));
defparam \resq[28]~93 .extended_lut = "off";
defparam \resq[28]~93 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[28]~93 .shared_arith = "on";

arriav_lcell_comb \resq[29]~97 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][29]~q ),
	.datad(!dout_301),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[28]~94 ),
	.sharein(\resq[28]~95 ),
	.combout(),
	.sumout(\resq[29]~97_sumout ),
	.cout(\resq[29]~98 ),
	.shareout(\resq[29]~99 ));
defparam \resq[29]~97 .extended_lut = "off";
defparam \resq[29]~97 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[29]~97 .shared_arith = "on";

arriav_lcell_comb \resq[30]~101 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][30]~q ),
	.datad(!dout_311),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[29]~98 ),
	.sharein(\resq[29]~99 ),
	.combout(),
	.sumout(\resq[30]~101_sumout ),
	.cout(\resq[30]~102 ),
	.shareout(\resq[30]~103 ));
defparam \resq[30]~101 .extended_lut = "off";
defparam \resq[30]~101 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[30]~101 .shared_arith = "on";

arriav_lcell_comb \resq[31]~105 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][31]~q ),
	.datad(!dout_321),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[30]~102 ),
	.sharein(\resq[30]~103 ),
	.combout(),
	.sumout(\resq[31]~105_sumout ),
	.cout(\resq[31]~106 ),
	.shareout(\resq[31]~107 ));
defparam \resq[31]~105 .extended_lut = "off";
defparam \resq[31]~105 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[31]~105 .shared_arith = "on";

arriav_lcell_comb \resq[32]~109 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][32]~q ),
	.datad(!dout_33),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[31]~106 ),
	.sharein(\resq[31]~107 ),
	.combout(),
	.sumout(\resq[32]~109_sumout ),
	.cout(),
	.shareout());
defparam \resq[32]~109 .extended_lut = "off";
defparam \resq[32]~109 .lut_mask = 64'h0000000000000FF0;
defparam \resq[32]~109 .shared_arith = "on";

endmodule

module cic_auk_dspip_delay_5 (
	datain,
	register_fifofifo_data05,
	register_fifofifo_data06,
	register_fifofifo_data07,
	register_fifofifo_data08,
	register_fifofifo_data09,
	register_fifofifo_data010,
	register_fifofifo_data011,
	register_fifofifo_data012,
	register_fifofifo_data013,
	register_fifofifo_data014,
	register_fifofifo_data015,
	register_fifofifo_data016,
	register_fifofifo_data017,
	register_fifofifo_data018,
	register_fifofifo_data019,
	register_fifofifo_data020,
	register_fifofifo_data021,
	register_fifofifo_data022,
	register_fifofifo_data023,
	register_fifofifo_data024,
	register_fifofifo_data025,
	register_fifofifo_data026,
	register_fifofifo_data027,
	register_fifofifo_data028,
	register_fifofifo_data029,
	register_fifofifo_data030,
	register_fifofifo_data031,
	register_fifofifo_data032,
	enable,
	register_fifofifo_data04,
	register_fifofifo_data03,
	register_fifofifo_data02,
	register_fifofifo_data01,
	register_fifofifo_data00,
	clk,
	reset)/* synthesis synthesis_greybox=1 */;
input 	[46:0] datain;
output 	register_fifofifo_data05;
output 	register_fifofifo_data06;
output 	register_fifofifo_data07;
output 	register_fifofifo_data08;
output 	register_fifofifo_data09;
output 	register_fifofifo_data010;
output 	register_fifofifo_data011;
output 	register_fifofifo_data012;
output 	register_fifofifo_data013;
output 	register_fifofifo_data014;
output 	register_fifofifo_data015;
output 	register_fifofifo_data016;
output 	register_fifofifo_data017;
output 	register_fifofifo_data018;
output 	register_fifofifo_data019;
output 	register_fifofifo_data020;
output 	register_fifofifo_data021;
output 	register_fifofifo_data022;
output 	register_fifofifo_data023;
output 	register_fifofifo_data024;
output 	register_fifofifo_data025;
output 	register_fifofifo_data026;
output 	register_fifofifo_data027;
output 	register_fifofifo_data028;
output 	register_fifofifo_data029;
output 	register_fifofifo_data030;
output 	register_fifofifo_data031;
output 	register_fifofifo_data032;
input 	enable;
output 	register_fifofifo_data04;
output 	register_fifofifo_data03;
output 	register_fifofifo_data02;
output 	register_fifofifo_data01;
output 	register_fifofifo_data00;
input 	clk;
input 	reset;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \register_fifo:fifo_data[0][5] (
	.clk(clk),
	.d(datain[5]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data05),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][5] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][5] .power_up = "low";

dffeas \register_fifo:fifo_data[0][6] (
	.clk(clk),
	.d(datain[6]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data06),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][6] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][6] .power_up = "low";

dffeas \register_fifo:fifo_data[0][7] (
	.clk(clk),
	.d(datain[7]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data07),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][7] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][7] .power_up = "low";

dffeas \register_fifo:fifo_data[0][8] (
	.clk(clk),
	.d(datain[8]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data08),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][8] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][8] .power_up = "low";

dffeas \register_fifo:fifo_data[0][9] (
	.clk(clk),
	.d(datain[9]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data09),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][9] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][9] .power_up = "low";

dffeas \register_fifo:fifo_data[0][10] (
	.clk(clk),
	.d(datain[10]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data010),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][10] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][10] .power_up = "low";

dffeas \register_fifo:fifo_data[0][11] (
	.clk(clk),
	.d(datain[11]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data011),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][11] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][11] .power_up = "low";

dffeas \register_fifo:fifo_data[0][12] (
	.clk(clk),
	.d(datain[12]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data012),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][12] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][12] .power_up = "low";

dffeas \register_fifo:fifo_data[0][13] (
	.clk(clk),
	.d(datain[13]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data013),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][13] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][13] .power_up = "low";

dffeas \register_fifo:fifo_data[0][14] (
	.clk(clk),
	.d(datain[14]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data014),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][14] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][14] .power_up = "low";

dffeas \register_fifo:fifo_data[0][15] (
	.clk(clk),
	.d(datain[15]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data015),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][15] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][15] .power_up = "low";

dffeas \register_fifo:fifo_data[0][16] (
	.clk(clk),
	.d(datain[16]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data016),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][16] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][16] .power_up = "low";

dffeas \register_fifo:fifo_data[0][17] (
	.clk(clk),
	.d(datain[17]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data017),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][17] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][17] .power_up = "low";

dffeas \register_fifo:fifo_data[0][18] (
	.clk(clk),
	.d(datain[18]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data018),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][18] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][18] .power_up = "low";

dffeas \register_fifo:fifo_data[0][19] (
	.clk(clk),
	.d(datain[19]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data019),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][19] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][19] .power_up = "low";

dffeas \register_fifo:fifo_data[0][20] (
	.clk(clk),
	.d(datain[20]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data020),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][20] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][20] .power_up = "low";

dffeas \register_fifo:fifo_data[0][21] (
	.clk(clk),
	.d(datain[21]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data021),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][21] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][21] .power_up = "low";

dffeas \register_fifo:fifo_data[0][22] (
	.clk(clk),
	.d(datain[22]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data022),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][22] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][22] .power_up = "low";

dffeas \register_fifo:fifo_data[0][23] (
	.clk(clk),
	.d(datain[23]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data023),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][23] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][23] .power_up = "low";

dffeas \register_fifo:fifo_data[0][24] (
	.clk(clk),
	.d(datain[24]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data024),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][24] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][24] .power_up = "low";

dffeas \register_fifo:fifo_data[0][25] (
	.clk(clk),
	.d(datain[25]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data025),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][25] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][25] .power_up = "low";

dffeas \register_fifo:fifo_data[0][26] (
	.clk(clk),
	.d(datain[26]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data026),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][26] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][26] .power_up = "low";

dffeas \register_fifo:fifo_data[0][27] (
	.clk(clk),
	.d(datain[27]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data027),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][27] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][27] .power_up = "low";

dffeas \register_fifo:fifo_data[0][28] (
	.clk(clk),
	.d(datain[28]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data028),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][28] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][28] .power_up = "low";

dffeas \register_fifo:fifo_data[0][29] (
	.clk(clk),
	.d(datain[29]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data029),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][29] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][29] .power_up = "low";

dffeas \register_fifo:fifo_data[0][30] (
	.clk(clk),
	.d(datain[30]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data030),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][30] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][30] .power_up = "low";

dffeas \register_fifo:fifo_data[0][31] (
	.clk(clk),
	.d(datain[31]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data031),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][31] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][31] .power_up = "low";

dffeas \register_fifo:fifo_data[0][32] (
	.clk(clk),
	.d(datain[32]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data032),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][32] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][32] .power_up = "low";

dffeas \register_fifo:fifo_data[0][4] (
	.clk(clk),
	.d(datain[4]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data04),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][4] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][4] .power_up = "low";

dffeas \register_fifo:fifo_data[0][3] (
	.clk(clk),
	.d(datain[3]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data03),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][3] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][3] .power_up = "low";

dffeas \register_fifo:fifo_data[0][2] (
	.clk(clk),
	.d(datain[2]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data02),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][2] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][2] .power_up = "low";

dffeas \register_fifo:fifo_data[0][1] (
	.clk(clk),
	.d(datain[1]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data01),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][1] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][1] .power_up = "low";

dffeas \register_fifo:fifo_data[0][0] (
	.clk(clk),
	.d(datain[0]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data00),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][0] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][0] .power_up = "low";

endmodule

module cic_auk_dspip_differentiator_6 (
	dout_valid1,
	dout_valid2,
	dout_4,
	dout_5,
	dout_6,
	dout_7,
	dout_8,
	dout_9,
	dout_10,
	dout_11,
	dout_12,
	dout_13,
	dout_14,
	dout_15,
	dout_16,
	dout_17,
	dout_18,
	dout_19,
	dout_20,
	dout_21,
	dout_22,
	dout_23,
	dout_24,
	dout_25,
	dout_26,
	dout_27,
	dout_28,
	dout_29,
	dout_30,
	dout_31,
	dout_3,
	dout_51,
	dout_2,
	dout_61,
	dout_71,
	dout_81,
	dout_91,
	dout_101,
	dout_111,
	dout_121,
	dout_131,
	dout_141,
	dout_151,
	dout_161,
	dout_171,
	dout_181,
	dout_191,
	dout_201,
	dout_211,
	dout_221,
	dout_231,
	dout_241,
	dout_251,
	dout_261,
	dout_271,
	dout_281,
	dout_291,
	dout_301,
	dout_311,
	dout_32,
	dout_41,
	dout_1,
	dout_33,
	dout_210,
	dout_110,
	stall_reg,
	dout_valid3,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	dout_valid1;
input 	dout_valid2;
output 	dout_4;
output 	dout_5;
output 	dout_6;
output 	dout_7;
output 	dout_8;
output 	dout_9;
output 	dout_10;
output 	dout_11;
output 	dout_12;
output 	dout_13;
output 	dout_14;
output 	dout_15;
output 	dout_16;
output 	dout_17;
output 	dout_18;
output 	dout_19;
output 	dout_20;
output 	dout_21;
output 	dout_22;
output 	dout_23;
output 	dout_24;
output 	dout_25;
output 	dout_26;
output 	dout_27;
output 	dout_28;
output 	dout_29;
output 	dout_30;
output 	dout_31;
output 	dout_3;
input 	dout_51;
output 	dout_2;
input 	dout_61;
input 	dout_71;
input 	dout_81;
input 	dout_91;
input 	dout_101;
input 	dout_111;
input 	dout_121;
input 	dout_131;
input 	dout_141;
input 	dout_151;
input 	dout_161;
input 	dout_171;
input 	dout_181;
input 	dout_191;
input 	dout_201;
input 	dout_211;
input 	dout_221;
input 	dout_231;
input 	dout_241;
input 	dout_251;
input 	dout_261;
input 	dout_271;
input 	dout_281;
input 	dout_291;
input 	dout_301;
input 	dout_311;
input 	dout_32;
input 	dout_41;
output 	dout_1;
input 	dout_33;
input 	dout_210;
input 	dout_110;
input 	stall_reg;
input 	dout_valid3;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \glogic:u0|register_fifo:fifo_data[0][4]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][5]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][6]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][7]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][8]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][9]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][10]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][11]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][12]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][13]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][14]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][15]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][16]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][17]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][18]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][19]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][20]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][21]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][22]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][23]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][24]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][25]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][26]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][27]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][28]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][29]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][30]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][31]~q ;
wire \dout~1_combout ;
wire \glogic:u0|register_fifo:fifo_data[0][3]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][2]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][1]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][0]~q ;
wire \resq[0]~126_cout ;
wire \resq[0]~127 ;
wire \resq[1]~122 ;
wire \resq[1]~123 ;
wire \resq[2]~118 ;
wire \resq[2]~119 ;
wire \resq[3]~114 ;
wire \resq[3]~115 ;
wire \resq[4]~1_sumout ;
wire \dout[20]~0_combout ;
wire \resq[4]~2 ;
wire \resq[4]~3 ;
wire \resq[5]~5_sumout ;
wire \resq[5]~6 ;
wire \resq[5]~7 ;
wire \resq[6]~9_sumout ;
wire \resq[6]~10 ;
wire \resq[6]~11 ;
wire \resq[7]~13_sumout ;
wire \resq[7]~14 ;
wire \resq[7]~15 ;
wire \resq[8]~17_sumout ;
wire \resq[8]~18 ;
wire \resq[8]~19 ;
wire \resq[9]~21_sumout ;
wire \resq[9]~22 ;
wire \resq[9]~23 ;
wire \resq[10]~25_sumout ;
wire \resq[10]~26 ;
wire \resq[10]~27 ;
wire \resq[11]~29_sumout ;
wire \resq[11]~30 ;
wire \resq[11]~31 ;
wire \resq[12]~33_sumout ;
wire \resq[12]~34 ;
wire \resq[12]~35 ;
wire \resq[13]~37_sumout ;
wire \resq[13]~38 ;
wire \resq[13]~39 ;
wire \resq[14]~41_sumout ;
wire \resq[14]~42 ;
wire \resq[14]~43 ;
wire \resq[15]~45_sumout ;
wire \resq[15]~46 ;
wire \resq[15]~47 ;
wire \resq[16]~49_sumout ;
wire \resq[16]~50 ;
wire \resq[16]~51 ;
wire \resq[17]~53_sumout ;
wire \resq[17]~54 ;
wire \resq[17]~55 ;
wire \resq[18]~57_sumout ;
wire \resq[18]~58 ;
wire \resq[18]~59 ;
wire \resq[19]~61_sumout ;
wire \resq[19]~62 ;
wire \resq[19]~63 ;
wire \resq[20]~65_sumout ;
wire \resq[20]~66 ;
wire \resq[20]~67 ;
wire \resq[21]~69_sumout ;
wire \resq[21]~70 ;
wire \resq[21]~71 ;
wire \resq[22]~73_sumout ;
wire \resq[22]~74 ;
wire \resq[22]~75 ;
wire \resq[23]~77_sumout ;
wire \resq[23]~78 ;
wire \resq[23]~79 ;
wire \resq[24]~81_sumout ;
wire \resq[24]~82 ;
wire \resq[24]~83 ;
wire \resq[25]~85_sumout ;
wire \resq[25]~86 ;
wire \resq[25]~87 ;
wire \resq[26]~89_sumout ;
wire \resq[26]~90 ;
wire \resq[26]~91 ;
wire \resq[27]~93_sumout ;
wire \resq[27]~94 ;
wire \resq[27]~95 ;
wire \resq[28]~97_sumout ;
wire \resq[28]~98 ;
wire \resq[28]~99 ;
wire \resq[29]~101_sumout ;
wire \resq[29]~102 ;
wire \resq[29]~103 ;
wire \resq[30]~105_sumout ;
wire \resq[30]~106 ;
wire \resq[30]~107 ;
wire \resq[31]~109_sumout ;
wire \resq[3]~113_sumout ;
wire \resq[2]~117_sumout ;
wire \resq[1]~121_sumout ;


cic_auk_dspip_delay_6 \glogic:u0 (
	.datain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,dout_32,dout_311,dout_301,dout_291,dout_281,dout_271,dout_261,dout_251,dout_241,dout_231,dout_221,dout_211,dout_201,dout_191,dout_181,dout_171,dout_161,dout_151,dout_141,dout_131,dout_121,dout_111,dout_101,dout_91,dout_81,dout_71,dout_61,
dout_51,dout_41,dout_33,dout_210,dout_110}),
	.register_fifofifo_data04(\glogic:u0|register_fifo:fifo_data[0][4]~q ),
	.register_fifofifo_data05(\glogic:u0|register_fifo:fifo_data[0][5]~q ),
	.register_fifofifo_data06(\glogic:u0|register_fifo:fifo_data[0][6]~q ),
	.register_fifofifo_data07(\glogic:u0|register_fifo:fifo_data[0][7]~q ),
	.register_fifofifo_data08(\glogic:u0|register_fifo:fifo_data[0][8]~q ),
	.register_fifofifo_data09(\glogic:u0|register_fifo:fifo_data[0][9]~q ),
	.register_fifofifo_data010(\glogic:u0|register_fifo:fifo_data[0][10]~q ),
	.register_fifofifo_data011(\glogic:u0|register_fifo:fifo_data[0][11]~q ),
	.register_fifofifo_data012(\glogic:u0|register_fifo:fifo_data[0][12]~q ),
	.register_fifofifo_data013(\glogic:u0|register_fifo:fifo_data[0][13]~q ),
	.register_fifofifo_data014(\glogic:u0|register_fifo:fifo_data[0][14]~q ),
	.register_fifofifo_data015(\glogic:u0|register_fifo:fifo_data[0][15]~q ),
	.register_fifofifo_data016(\glogic:u0|register_fifo:fifo_data[0][16]~q ),
	.register_fifofifo_data017(\glogic:u0|register_fifo:fifo_data[0][17]~q ),
	.register_fifofifo_data018(\glogic:u0|register_fifo:fifo_data[0][18]~q ),
	.register_fifofifo_data019(\glogic:u0|register_fifo:fifo_data[0][19]~q ),
	.register_fifofifo_data020(\glogic:u0|register_fifo:fifo_data[0][20]~q ),
	.register_fifofifo_data021(\glogic:u0|register_fifo:fifo_data[0][21]~q ),
	.register_fifofifo_data022(\glogic:u0|register_fifo:fifo_data[0][22]~q ),
	.register_fifofifo_data023(\glogic:u0|register_fifo:fifo_data[0][23]~q ),
	.register_fifofifo_data024(\glogic:u0|register_fifo:fifo_data[0][24]~q ),
	.register_fifofifo_data025(\glogic:u0|register_fifo:fifo_data[0][25]~q ),
	.register_fifofifo_data026(\glogic:u0|register_fifo:fifo_data[0][26]~q ),
	.register_fifofifo_data027(\glogic:u0|register_fifo:fifo_data[0][27]~q ),
	.register_fifofifo_data028(\glogic:u0|register_fifo:fifo_data[0][28]~q ),
	.register_fifofifo_data029(\glogic:u0|register_fifo:fifo_data[0][29]~q ),
	.register_fifofifo_data030(\glogic:u0|register_fifo:fifo_data[0][30]~q ),
	.register_fifofifo_data031(\glogic:u0|register_fifo:fifo_data[0][31]~q ),
	.enable(\dout~1_combout ),
	.register_fifofifo_data03(\glogic:u0|register_fifo:fifo_data[0][3]~q ),
	.register_fifofifo_data02(\glogic:u0|register_fifo:fifo_data[0][2]~q ),
	.register_fifofifo_data01(\glogic:u0|register_fifo:fifo_data[0][1]~q ),
	.register_fifofifo_data00(\glogic:u0|register_fifo:fifo_data[0][0]~q ),
	.clk(clk),
	.reset(reset_n));

arriav_lcell_comb \dout~1 (
	.dataa(!stall_reg),
	.datab(!dout_valid2),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dout~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dout~1 .extended_lut = "off";
defparam \dout~1 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \dout~1 .shared_arith = "off";

dffeas dout_valid(
	.clk(clk),
	.d(dout_valid2),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(dout_valid3),
	.q(dout_valid1),
	.prn(vcc));
defparam dout_valid.is_wysiwyg = "true";
defparam dout_valid.power_up = "low";

dffeas \dout[4] (
	.clk(clk),
	.d(\resq[4]~1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[20]~0_combout ),
	.q(dout_4),
	.prn(vcc));
defparam \dout[4] .is_wysiwyg = "true";
defparam \dout[4] .power_up = "low";

dffeas \dout[5] (
	.clk(clk),
	.d(\resq[5]~5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[20]~0_combout ),
	.q(dout_5),
	.prn(vcc));
defparam \dout[5] .is_wysiwyg = "true";
defparam \dout[5] .power_up = "low";

dffeas \dout[6] (
	.clk(clk),
	.d(\resq[6]~9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[20]~0_combout ),
	.q(dout_6),
	.prn(vcc));
defparam \dout[6] .is_wysiwyg = "true";
defparam \dout[6] .power_up = "low";

dffeas \dout[7] (
	.clk(clk),
	.d(\resq[7]~13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[20]~0_combout ),
	.q(dout_7),
	.prn(vcc));
defparam \dout[7] .is_wysiwyg = "true";
defparam \dout[7] .power_up = "low";

dffeas \dout[8] (
	.clk(clk),
	.d(\resq[8]~17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[20]~0_combout ),
	.q(dout_8),
	.prn(vcc));
defparam \dout[8] .is_wysiwyg = "true";
defparam \dout[8] .power_up = "low";

dffeas \dout[9] (
	.clk(clk),
	.d(\resq[9]~21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[20]~0_combout ),
	.q(dout_9),
	.prn(vcc));
defparam \dout[9] .is_wysiwyg = "true";
defparam \dout[9] .power_up = "low";

dffeas \dout[10] (
	.clk(clk),
	.d(\resq[10]~25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[20]~0_combout ),
	.q(dout_10),
	.prn(vcc));
defparam \dout[10] .is_wysiwyg = "true";
defparam \dout[10] .power_up = "low";

dffeas \dout[11] (
	.clk(clk),
	.d(\resq[11]~29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[20]~0_combout ),
	.q(dout_11),
	.prn(vcc));
defparam \dout[11] .is_wysiwyg = "true";
defparam \dout[11] .power_up = "low";

dffeas \dout[12] (
	.clk(clk),
	.d(\resq[12]~33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[20]~0_combout ),
	.q(dout_12),
	.prn(vcc));
defparam \dout[12] .is_wysiwyg = "true";
defparam \dout[12] .power_up = "low";

dffeas \dout[13] (
	.clk(clk),
	.d(\resq[13]~37_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[20]~0_combout ),
	.q(dout_13),
	.prn(vcc));
defparam \dout[13] .is_wysiwyg = "true";
defparam \dout[13] .power_up = "low";

dffeas \dout[14] (
	.clk(clk),
	.d(\resq[14]~41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[20]~0_combout ),
	.q(dout_14),
	.prn(vcc));
defparam \dout[14] .is_wysiwyg = "true";
defparam \dout[14] .power_up = "low";

dffeas \dout[15] (
	.clk(clk),
	.d(\resq[15]~45_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[20]~0_combout ),
	.q(dout_15),
	.prn(vcc));
defparam \dout[15] .is_wysiwyg = "true";
defparam \dout[15] .power_up = "low";

dffeas \dout[16] (
	.clk(clk),
	.d(\resq[16]~49_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[20]~0_combout ),
	.q(dout_16),
	.prn(vcc));
defparam \dout[16] .is_wysiwyg = "true";
defparam \dout[16] .power_up = "low";

dffeas \dout[17] (
	.clk(clk),
	.d(\resq[17]~53_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[20]~0_combout ),
	.q(dout_17),
	.prn(vcc));
defparam \dout[17] .is_wysiwyg = "true";
defparam \dout[17] .power_up = "low";

dffeas \dout[18] (
	.clk(clk),
	.d(\resq[18]~57_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[20]~0_combout ),
	.q(dout_18),
	.prn(vcc));
defparam \dout[18] .is_wysiwyg = "true";
defparam \dout[18] .power_up = "low";

dffeas \dout[19] (
	.clk(clk),
	.d(\resq[19]~61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[20]~0_combout ),
	.q(dout_19),
	.prn(vcc));
defparam \dout[19] .is_wysiwyg = "true";
defparam \dout[19] .power_up = "low";

dffeas \dout[20] (
	.clk(clk),
	.d(\resq[20]~65_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[20]~0_combout ),
	.q(dout_20),
	.prn(vcc));
defparam \dout[20] .is_wysiwyg = "true";
defparam \dout[20] .power_up = "low";

dffeas \dout[21] (
	.clk(clk),
	.d(\resq[21]~69_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[20]~0_combout ),
	.q(dout_21),
	.prn(vcc));
defparam \dout[21] .is_wysiwyg = "true";
defparam \dout[21] .power_up = "low";

dffeas \dout[22] (
	.clk(clk),
	.d(\resq[22]~73_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[20]~0_combout ),
	.q(dout_22),
	.prn(vcc));
defparam \dout[22] .is_wysiwyg = "true";
defparam \dout[22] .power_up = "low";

dffeas \dout[23] (
	.clk(clk),
	.d(\resq[23]~77_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[20]~0_combout ),
	.q(dout_23),
	.prn(vcc));
defparam \dout[23] .is_wysiwyg = "true";
defparam \dout[23] .power_up = "low";

dffeas \dout[24] (
	.clk(clk),
	.d(\resq[24]~81_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[20]~0_combout ),
	.q(dout_24),
	.prn(vcc));
defparam \dout[24] .is_wysiwyg = "true";
defparam \dout[24] .power_up = "low";

dffeas \dout[25] (
	.clk(clk),
	.d(\resq[25]~85_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[20]~0_combout ),
	.q(dout_25),
	.prn(vcc));
defparam \dout[25] .is_wysiwyg = "true";
defparam \dout[25] .power_up = "low";

dffeas \dout[26] (
	.clk(clk),
	.d(\resq[26]~89_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[20]~0_combout ),
	.q(dout_26),
	.prn(vcc));
defparam \dout[26] .is_wysiwyg = "true";
defparam \dout[26] .power_up = "low";

dffeas \dout[27] (
	.clk(clk),
	.d(\resq[27]~93_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[20]~0_combout ),
	.q(dout_27),
	.prn(vcc));
defparam \dout[27] .is_wysiwyg = "true";
defparam \dout[27] .power_up = "low";

dffeas \dout[28] (
	.clk(clk),
	.d(\resq[28]~97_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[20]~0_combout ),
	.q(dout_28),
	.prn(vcc));
defparam \dout[28] .is_wysiwyg = "true";
defparam \dout[28] .power_up = "low";

dffeas \dout[29] (
	.clk(clk),
	.d(\resq[29]~101_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[20]~0_combout ),
	.q(dout_29),
	.prn(vcc));
defparam \dout[29] .is_wysiwyg = "true";
defparam \dout[29] .power_up = "low";

dffeas \dout[30] (
	.clk(clk),
	.d(\resq[30]~105_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[20]~0_combout ),
	.q(dout_30),
	.prn(vcc));
defparam \dout[30] .is_wysiwyg = "true";
defparam \dout[30] .power_up = "low";

dffeas \dout[31] (
	.clk(clk),
	.d(\resq[31]~109_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[20]~0_combout ),
	.q(dout_31),
	.prn(vcc));
defparam \dout[31] .is_wysiwyg = "true";
defparam \dout[31] .power_up = "low";

dffeas \dout[3] (
	.clk(clk),
	.d(\resq[3]~113_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[20]~0_combout ),
	.q(dout_3),
	.prn(vcc));
defparam \dout[3] .is_wysiwyg = "true";
defparam \dout[3] .power_up = "low";

dffeas \dout[2] (
	.clk(clk),
	.d(\resq[2]~117_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[20]~0_combout ),
	.q(dout_2),
	.prn(vcc));
defparam \dout[2] .is_wysiwyg = "true";
defparam \dout[2] .power_up = "low";

dffeas \dout[1] (
	.clk(clk),
	.d(\resq[1]~121_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[20]~0_combout ),
	.q(dout_1),
	.prn(vcc));
defparam \dout[1] .is_wysiwyg = "true";
defparam \dout[1] .power_up = "low";

arriav_lcell_comb \resq[0]~126 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][0]~q ),
	.datad(!dout_110),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\resq[0]~126_cout ),
	.shareout(\resq[0]~127 ));
defparam \resq[0]~126 .extended_lut = "off";
defparam \resq[0]~126 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[0]~126 .shared_arith = "on";

arriav_lcell_comb \resq[1]~121 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][1]~q ),
	.datad(!dout_210),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[0]~126_cout ),
	.sharein(\resq[0]~127 ),
	.combout(),
	.sumout(\resq[1]~121_sumout ),
	.cout(\resq[1]~122 ),
	.shareout(\resq[1]~123 ));
defparam \resq[1]~121 .extended_lut = "off";
defparam \resq[1]~121 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[1]~121 .shared_arith = "on";

arriav_lcell_comb \resq[2]~117 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][2]~q ),
	.datad(!dout_33),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[1]~122 ),
	.sharein(\resq[1]~123 ),
	.combout(),
	.sumout(\resq[2]~117_sumout ),
	.cout(\resq[2]~118 ),
	.shareout(\resq[2]~119 ));
defparam \resq[2]~117 .extended_lut = "off";
defparam \resq[2]~117 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[2]~117 .shared_arith = "on";

arriav_lcell_comb \resq[3]~113 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][3]~q ),
	.datad(!dout_41),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[2]~118 ),
	.sharein(\resq[2]~119 ),
	.combout(),
	.sumout(\resq[3]~113_sumout ),
	.cout(\resq[3]~114 ),
	.shareout(\resq[3]~115 ));
defparam \resq[3]~113 .extended_lut = "off";
defparam \resq[3]~113 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[3]~113 .shared_arith = "on";

arriav_lcell_comb \resq[4]~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][4]~q ),
	.datad(!dout_51),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[3]~114 ),
	.sharein(\resq[3]~115 ),
	.combout(),
	.sumout(\resq[4]~1_sumout ),
	.cout(\resq[4]~2 ),
	.shareout(\resq[4]~3 ));
defparam \resq[4]~1 .extended_lut = "off";
defparam \resq[4]~1 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[4]~1 .shared_arith = "on";

arriav_lcell_comb \dout[20]~0 (
	.dataa(!reset_n),
	.datab(!stall_reg),
	.datac(!dout_valid2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dout[20]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dout[20]~0 .extended_lut = "off";
defparam \dout[20]~0 .lut_mask = 64'hEFEFEFEFEFEFEFEF;
defparam \dout[20]~0 .shared_arith = "off";

arriav_lcell_comb \resq[5]~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][5]~q ),
	.datad(!dout_61),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[4]~2 ),
	.sharein(\resq[4]~3 ),
	.combout(),
	.sumout(\resq[5]~5_sumout ),
	.cout(\resq[5]~6 ),
	.shareout(\resq[5]~7 ));
defparam \resq[5]~5 .extended_lut = "off";
defparam \resq[5]~5 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[5]~5 .shared_arith = "on";

arriav_lcell_comb \resq[6]~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][6]~q ),
	.datad(!dout_71),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[5]~6 ),
	.sharein(\resq[5]~7 ),
	.combout(),
	.sumout(\resq[6]~9_sumout ),
	.cout(\resq[6]~10 ),
	.shareout(\resq[6]~11 ));
defparam \resq[6]~9 .extended_lut = "off";
defparam \resq[6]~9 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[6]~9 .shared_arith = "on";

arriav_lcell_comb \resq[7]~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][7]~q ),
	.datad(!dout_81),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[6]~10 ),
	.sharein(\resq[6]~11 ),
	.combout(),
	.sumout(\resq[7]~13_sumout ),
	.cout(\resq[7]~14 ),
	.shareout(\resq[7]~15 ));
defparam \resq[7]~13 .extended_lut = "off";
defparam \resq[7]~13 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[7]~13 .shared_arith = "on";

arriav_lcell_comb \resq[8]~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][8]~q ),
	.datad(!dout_91),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[7]~14 ),
	.sharein(\resq[7]~15 ),
	.combout(),
	.sumout(\resq[8]~17_sumout ),
	.cout(\resq[8]~18 ),
	.shareout(\resq[8]~19 ));
defparam \resq[8]~17 .extended_lut = "off";
defparam \resq[8]~17 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[8]~17 .shared_arith = "on";

arriav_lcell_comb \resq[9]~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][9]~q ),
	.datad(!dout_101),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[8]~18 ),
	.sharein(\resq[8]~19 ),
	.combout(),
	.sumout(\resq[9]~21_sumout ),
	.cout(\resq[9]~22 ),
	.shareout(\resq[9]~23 ));
defparam \resq[9]~21 .extended_lut = "off";
defparam \resq[9]~21 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[9]~21 .shared_arith = "on";

arriav_lcell_comb \resq[10]~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][10]~q ),
	.datad(!dout_111),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[9]~22 ),
	.sharein(\resq[9]~23 ),
	.combout(),
	.sumout(\resq[10]~25_sumout ),
	.cout(\resq[10]~26 ),
	.shareout(\resq[10]~27 ));
defparam \resq[10]~25 .extended_lut = "off";
defparam \resq[10]~25 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[10]~25 .shared_arith = "on";

arriav_lcell_comb \resq[11]~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][11]~q ),
	.datad(!dout_121),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[10]~26 ),
	.sharein(\resq[10]~27 ),
	.combout(),
	.sumout(\resq[11]~29_sumout ),
	.cout(\resq[11]~30 ),
	.shareout(\resq[11]~31 ));
defparam \resq[11]~29 .extended_lut = "off";
defparam \resq[11]~29 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[11]~29 .shared_arith = "on";

arriav_lcell_comb \resq[12]~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][12]~q ),
	.datad(!dout_131),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[11]~30 ),
	.sharein(\resq[11]~31 ),
	.combout(),
	.sumout(\resq[12]~33_sumout ),
	.cout(\resq[12]~34 ),
	.shareout(\resq[12]~35 ));
defparam \resq[12]~33 .extended_lut = "off";
defparam \resq[12]~33 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[12]~33 .shared_arith = "on";

arriav_lcell_comb \resq[13]~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][13]~q ),
	.datad(!dout_141),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[12]~34 ),
	.sharein(\resq[12]~35 ),
	.combout(),
	.sumout(\resq[13]~37_sumout ),
	.cout(\resq[13]~38 ),
	.shareout(\resq[13]~39 ));
defparam \resq[13]~37 .extended_lut = "off";
defparam \resq[13]~37 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[13]~37 .shared_arith = "on";

arriav_lcell_comb \resq[14]~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][14]~q ),
	.datad(!dout_151),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[13]~38 ),
	.sharein(\resq[13]~39 ),
	.combout(),
	.sumout(\resq[14]~41_sumout ),
	.cout(\resq[14]~42 ),
	.shareout(\resq[14]~43 ));
defparam \resq[14]~41 .extended_lut = "off";
defparam \resq[14]~41 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[14]~41 .shared_arith = "on";

arriav_lcell_comb \resq[15]~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][15]~q ),
	.datad(!dout_161),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[14]~42 ),
	.sharein(\resq[14]~43 ),
	.combout(),
	.sumout(\resq[15]~45_sumout ),
	.cout(\resq[15]~46 ),
	.shareout(\resq[15]~47 ));
defparam \resq[15]~45 .extended_lut = "off";
defparam \resq[15]~45 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[15]~45 .shared_arith = "on";

arriav_lcell_comb \resq[16]~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][16]~q ),
	.datad(!dout_171),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[15]~46 ),
	.sharein(\resq[15]~47 ),
	.combout(),
	.sumout(\resq[16]~49_sumout ),
	.cout(\resq[16]~50 ),
	.shareout(\resq[16]~51 ));
defparam \resq[16]~49 .extended_lut = "off";
defparam \resq[16]~49 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[16]~49 .shared_arith = "on";

arriav_lcell_comb \resq[17]~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][17]~q ),
	.datad(!dout_181),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[16]~50 ),
	.sharein(\resq[16]~51 ),
	.combout(),
	.sumout(\resq[17]~53_sumout ),
	.cout(\resq[17]~54 ),
	.shareout(\resq[17]~55 ));
defparam \resq[17]~53 .extended_lut = "off";
defparam \resq[17]~53 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[17]~53 .shared_arith = "on";

arriav_lcell_comb \resq[18]~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][18]~q ),
	.datad(!dout_191),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[17]~54 ),
	.sharein(\resq[17]~55 ),
	.combout(),
	.sumout(\resq[18]~57_sumout ),
	.cout(\resq[18]~58 ),
	.shareout(\resq[18]~59 ));
defparam \resq[18]~57 .extended_lut = "off";
defparam \resq[18]~57 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[18]~57 .shared_arith = "on";

arriav_lcell_comb \resq[19]~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][19]~q ),
	.datad(!dout_201),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[18]~58 ),
	.sharein(\resq[18]~59 ),
	.combout(),
	.sumout(\resq[19]~61_sumout ),
	.cout(\resq[19]~62 ),
	.shareout(\resq[19]~63 ));
defparam \resq[19]~61 .extended_lut = "off";
defparam \resq[19]~61 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[19]~61 .shared_arith = "on";

arriav_lcell_comb \resq[20]~65 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][20]~q ),
	.datad(!dout_211),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[19]~62 ),
	.sharein(\resq[19]~63 ),
	.combout(),
	.sumout(\resq[20]~65_sumout ),
	.cout(\resq[20]~66 ),
	.shareout(\resq[20]~67 ));
defparam \resq[20]~65 .extended_lut = "off";
defparam \resq[20]~65 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[20]~65 .shared_arith = "on";

arriav_lcell_comb \resq[21]~69 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][21]~q ),
	.datad(!dout_221),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[20]~66 ),
	.sharein(\resq[20]~67 ),
	.combout(),
	.sumout(\resq[21]~69_sumout ),
	.cout(\resq[21]~70 ),
	.shareout(\resq[21]~71 ));
defparam \resq[21]~69 .extended_lut = "off";
defparam \resq[21]~69 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[21]~69 .shared_arith = "on";

arriav_lcell_comb \resq[22]~73 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][22]~q ),
	.datad(!dout_231),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[21]~70 ),
	.sharein(\resq[21]~71 ),
	.combout(),
	.sumout(\resq[22]~73_sumout ),
	.cout(\resq[22]~74 ),
	.shareout(\resq[22]~75 ));
defparam \resq[22]~73 .extended_lut = "off";
defparam \resq[22]~73 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[22]~73 .shared_arith = "on";

arriav_lcell_comb \resq[23]~77 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][23]~q ),
	.datad(!dout_241),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[22]~74 ),
	.sharein(\resq[22]~75 ),
	.combout(),
	.sumout(\resq[23]~77_sumout ),
	.cout(\resq[23]~78 ),
	.shareout(\resq[23]~79 ));
defparam \resq[23]~77 .extended_lut = "off";
defparam \resq[23]~77 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[23]~77 .shared_arith = "on";

arriav_lcell_comb \resq[24]~81 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][24]~q ),
	.datad(!dout_251),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[23]~78 ),
	.sharein(\resq[23]~79 ),
	.combout(),
	.sumout(\resq[24]~81_sumout ),
	.cout(\resq[24]~82 ),
	.shareout(\resq[24]~83 ));
defparam \resq[24]~81 .extended_lut = "off";
defparam \resq[24]~81 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[24]~81 .shared_arith = "on";

arriav_lcell_comb \resq[25]~85 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][25]~q ),
	.datad(!dout_261),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[24]~82 ),
	.sharein(\resq[24]~83 ),
	.combout(),
	.sumout(\resq[25]~85_sumout ),
	.cout(\resq[25]~86 ),
	.shareout(\resq[25]~87 ));
defparam \resq[25]~85 .extended_lut = "off";
defparam \resq[25]~85 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[25]~85 .shared_arith = "on";

arriav_lcell_comb \resq[26]~89 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][26]~q ),
	.datad(!dout_271),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[25]~86 ),
	.sharein(\resq[25]~87 ),
	.combout(),
	.sumout(\resq[26]~89_sumout ),
	.cout(\resq[26]~90 ),
	.shareout(\resq[26]~91 ));
defparam \resq[26]~89 .extended_lut = "off";
defparam \resq[26]~89 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[26]~89 .shared_arith = "on";

arriav_lcell_comb \resq[27]~93 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][27]~q ),
	.datad(!dout_281),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[26]~90 ),
	.sharein(\resq[26]~91 ),
	.combout(),
	.sumout(\resq[27]~93_sumout ),
	.cout(\resq[27]~94 ),
	.shareout(\resq[27]~95 ));
defparam \resq[27]~93 .extended_lut = "off";
defparam \resq[27]~93 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[27]~93 .shared_arith = "on";

arriav_lcell_comb \resq[28]~97 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][28]~q ),
	.datad(!dout_291),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[27]~94 ),
	.sharein(\resq[27]~95 ),
	.combout(),
	.sumout(\resq[28]~97_sumout ),
	.cout(\resq[28]~98 ),
	.shareout(\resq[28]~99 ));
defparam \resq[28]~97 .extended_lut = "off";
defparam \resq[28]~97 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[28]~97 .shared_arith = "on";

arriav_lcell_comb \resq[29]~101 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][29]~q ),
	.datad(!dout_301),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[28]~98 ),
	.sharein(\resq[28]~99 ),
	.combout(),
	.sumout(\resq[29]~101_sumout ),
	.cout(\resq[29]~102 ),
	.shareout(\resq[29]~103 ));
defparam \resq[29]~101 .extended_lut = "off";
defparam \resq[29]~101 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[29]~101 .shared_arith = "on";

arriav_lcell_comb \resq[30]~105 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][30]~q ),
	.datad(!dout_311),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[29]~102 ),
	.sharein(\resq[29]~103 ),
	.combout(),
	.sumout(\resq[30]~105_sumout ),
	.cout(\resq[30]~106 ),
	.shareout(\resq[30]~107 ));
defparam \resq[30]~105 .extended_lut = "off";
defparam \resq[30]~105 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[30]~105 .shared_arith = "on";

arriav_lcell_comb \resq[31]~109 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][31]~q ),
	.datad(!dout_32),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[30]~106 ),
	.sharein(\resq[30]~107 ),
	.combout(),
	.sumout(\resq[31]~109_sumout ),
	.cout(),
	.shareout());
defparam \resq[31]~109 .extended_lut = "off";
defparam \resq[31]~109 .lut_mask = 64'h0000000000000FF0;
defparam \resq[31]~109 .shared_arith = "on";

endmodule

module cic_auk_dspip_delay_6 (
	datain,
	register_fifofifo_data04,
	register_fifofifo_data05,
	register_fifofifo_data06,
	register_fifofifo_data07,
	register_fifofifo_data08,
	register_fifofifo_data09,
	register_fifofifo_data010,
	register_fifofifo_data011,
	register_fifofifo_data012,
	register_fifofifo_data013,
	register_fifofifo_data014,
	register_fifofifo_data015,
	register_fifofifo_data016,
	register_fifofifo_data017,
	register_fifofifo_data018,
	register_fifofifo_data019,
	register_fifofifo_data020,
	register_fifofifo_data021,
	register_fifofifo_data022,
	register_fifofifo_data023,
	register_fifofifo_data024,
	register_fifofifo_data025,
	register_fifofifo_data026,
	register_fifofifo_data027,
	register_fifofifo_data028,
	register_fifofifo_data029,
	register_fifofifo_data030,
	register_fifofifo_data031,
	enable,
	register_fifofifo_data03,
	register_fifofifo_data02,
	register_fifofifo_data01,
	register_fifofifo_data00,
	clk,
	reset)/* synthesis synthesis_greybox=1 */;
input 	[46:0] datain;
output 	register_fifofifo_data04;
output 	register_fifofifo_data05;
output 	register_fifofifo_data06;
output 	register_fifofifo_data07;
output 	register_fifofifo_data08;
output 	register_fifofifo_data09;
output 	register_fifofifo_data010;
output 	register_fifofifo_data011;
output 	register_fifofifo_data012;
output 	register_fifofifo_data013;
output 	register_fifofifo_data014;
output 	register_fifofifo_data015;
output 	register_fifofifo_data016;
output 	register_fifofifo_data017;
output 	register_fifofifo_data018;
output 	register_fifofifo_data019;
output 	register_fifofifo_data020;
output 	register_fifofifo_data021;
output 	register_fifofifo_data022;
output 	register_fifofifo_data023;
output 	register_fifofifo_data024;
output 	register_fifofifo_data025;
output 	register_fifofifo_data026;
output 	register_fifofifo_data027;
output 	register_fifofifo_data028;
output 	register_fifofifo_data029;
output 	register_fifofifo_data030;
output 	register_fifofifo_data031;
input 	enable;
output 	register_fifofifo_data03;
output 	register_fifofifo_data02;
output 	register_fifofifo_data01;
output 	register_fifofifo_data00;
input 	clk;
input 	reset;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \register_fifo:fifo_data[0][4] (
	.clk(clk),
	.d(datain[4]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data04),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][4] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][4] .power_up = "low";

dffeas \register_fifo:fifo_data[0][5] (
	.clk(clk),
	.d(datain[5]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data05),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][5] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][5] .power_up = "low";

dffeas \register_fifo:fifo_data[0][6] (
	.clk(clk),
	.d(datain[6]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data06),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][6] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][6] .power_up = "low";

dffeas \register_fifo:fifo_data[0][7] (
	.clk(clk),
	.d(datain[7]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data07),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][7] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][7] .power_up = "low";

dffeas \register_fifo:fifo_data[0][8] (
	.clk(clk),
	.d(datain[8]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data08),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][8] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][8] .power_up = "low";

dffeas \register_fifo:fifo_data[0][9] (
	.clk(clk),
	.d(datain[9]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data09),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][9] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][9] .power_up = "low";

dffeas \register_fifo:fifo_data[0][10] (
	.clk(clk),
	.d(datain[10]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data010),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][10] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][10] .power_up = "low";

dffeas \register_fifo:fifo_data[0][11] (
	.clk(clk),
	.d(datain[11]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data011),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][11] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][11] .power_up = "low";

dffeas \register_fifo:fifo_data[0][12] (
	.clk(clk),
	.d(datain[12]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data012),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][12] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][12] .power_up = "low";

dffeas \register_fifo:fifo_data[0][13] (
	.clk(clk),
	.d(datain[13]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data013),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][13] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][13] .power_up = "low";

dffeas \register_fifo:fifo_data[0][14] (
	.clk(clk),
	.d(datain[14]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data014),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][14] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][14] .power_up = "low";

dffeas \register_fifo:fifo_data[0][15] (
	.clk(clk),
	.d(datain[15]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data015),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][15] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][15] .power_up = "low";

dffeas \register_fifo:fifo_data[0][16] (
	.clk(clk),
	.d(datain[16]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data016),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][16] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][16] .power_up = "low";

dffeas \register_fifo:fifo_data[0][17] (
	.clk(clk),
	.d(datain[17]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data017),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][17] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][17] .power_up = "low";

dffeas \register_fifo:fifo_data[0][18] (
	.clk(clk),
	.d(datain[18]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data018),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][18] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][18] .power_up = "low";

dffeas \register_fifo:fifo_data[0][19] (
	.clk(clk),
	.d(datain[19]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data019),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][19] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][19] .power_up = "low";

dffeas \register_fifo:fifo_data[0][20] (
	.clk(clk),
	.d(datain[20]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data020),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][20] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][20] .power_up = "low";

dffeas \register_fifo:fifo_data[0][21] (
	.clk(clk),
	.d(datain[21]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data021),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][21] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][21] .power_up = "low";

dffeas \register_fifo:fifo_data[0][22] (
	.clk(clk),
	.d(datain[22]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data022),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][22] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][22] .power_up = "low";

dffeas \register_fifo:fifo_data[0][23] (
	.clk(clk),
	.d(datain[23]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data023),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][23] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][23] .power_up = "low";

dffeas \register_fifo:fifo_data[0][24] (
	.clk(clk),
	.d(datain[24]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data024),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][24] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][24] .power_up = "low";

dffeas \register_fifo:fifo_data[0][25] (
	.clk(clk),
	.d(datain[25]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data025),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][25] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][25] .power_up = "low";

dffeas \register_fifo:fifo_data[0][26] (
	.clk(clk),
	.d(datain[26]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data026),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][26] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][26] .power_up = "low";

dffeas \register_fifo:fifo_data[0][27] (
	.clk(clk),
	.d(datain[27]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data027),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][27] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][27] .power_up = "low";

dffeas \register_fifo:fifo_data[0][28] (
	.clk(clk),
	.d(datain[28]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data028),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][28] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][28] .power_up = "low";

dffeas \register_fifo:fifo_data[0][29] (
	.clk(clk),
	.d(datain[29]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data029),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][29] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][29] .power_up = "low";

dffeas \register_fifo:fifo_data[0][30] (
	.clk(clk),
	.d(datain[30]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data030),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][30] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][30] .power_up = "low";

dffeas \register_fifo:fifo_data[0][31] (
	.clk(clk),
	.d(datain[31]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data031),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][31] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][31] .power_up = "low";

dffeas \register_fifo:fifo_data[0][3] (
	.clk(clk),
	.d(datain[3]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data03),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][3] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][3] .power_up = "low";

dffeas \register_fifo:fifo_data[0][2] (
	.clk(clk),
	.d(datain[2]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data02),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][2] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][2] .power_up = "low";

dffeas \register_fifo:fifo_data[0][1] (
	.clk(clk),
	.d(datain[1]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data01),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][1] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][1] .power_up = "low";

dffeas \register_fifo:fifo_data[0][0] (
	.clk(clk),
	.d(datain[0]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data00),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][0] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][0] .power_up = "low";

endmodule

module cic_auk_dspip_differentiator_7 (
	dout_valid1,
	dout_3,
	dout_4,
	dout_5,
	dout_6,
	dout_7,
	dout_8,
	dout_9,
	dout_10,
	dout_11,
	dout_12,
	dout_13,
	dout_14,
	dout_15,
	dout_16,
	dout_17,
	dout_18,
	dout_19,
	dout_20,
	dout_21,
	dout_22,
	dout_23,
	dout_24,
	dout_25,
	dout_26,
	dout_27,
	dout_28,
	dout_29,
	dout_30,
	dout_valid2,
	dout_41,
	dout_51,
	dout_61,
	dout_71,
	dout_81,
	dout_91,
	dout_101,
	dout_111,
	dout_121,
	dout_131,
	dout_141,
	dout_151,
	dout_161,
	dout_171,
	dout_181,
	dout_191,
	dout_201,
	dout_211,
	dout_221,
	dout_231,
	dout_241,
	dout_251,
	dout_261,
	dout_271,
	dout_281,
	dout_291,
	dout_301,
	dout_31,
	dout_32,
	dout_2,
	dout_1,
	stall_reg,
	dout_valid3,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	dout_valid1;
output 	dout_3;
output 	dout_4;
output 	dout_5;
output 	dout_6;
output 	dout_7;
output 	dout_8;
output 	dout_9;
output 	dout_10;
output 	dout_11;
output 	dout_12;
output 	dout_13;
output 	dout_14;
output 	dout_15;
output 	dout_16;
output 	dout_17;
output 	dout_18;
output 	dout_19;
output 	dout_20;
output 	dout_21;
output 	dout_22;
output 	dout_23;
output 	dout_24;
output 	dout_25;
output 	dout_26;
output 	dout_27;
output 	dout_28;
output 	dout_29;
output 	dout_30;
input 	dout_valid2;
input 	dout_41;
input 	dout_51;
input 	dout_61;
input 	dout_71;
input 	dout_81;
input 	dout_91;
input 	dout_101;
input 	dout_111;
input 	dout_121;
input 	dout_131;
input 	dout_141;
input 	dout_151;
input 	dout_161;
input 	dout_171;
input 	dout_181;
input 	dout_191;
input 	dout_201;
input 	dout_211;
input 	dout_221;
input 	dout_231;
input 	dout_241;
input 	dout_251;
input 	dout_261;
input 	dout_271;
input 	dout_281;
input 	dout_291;
input 	dout_301;
input 	dout_31;
input 	dout_32;
input 	dout_2;
input 	dout_1;
input 	stall_reg;
output 	dout_valid3;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \glogic:u0|register_fifo:fifo_data[0][3]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][4]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][5]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][6]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][7]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][8]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][9]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][10]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][11]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][12]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][13]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][14]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][15]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][16]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][17]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][18]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][19]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][20]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][21]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][22]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][23]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][24]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][25]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][26]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][27]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][28]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][29]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][30]~q ;
wire \dout~1_combout ;
wire \glogic:u0|register_fifo:fifo_data[0][2]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][1]~q ;
wire \glogic:u0|register_fifo:fifo_data[0][0]~q ;
wire \resq[0]~122_cout ;
wire \resq[0]~123 ;
wire \resq[1]~118_cout ;
wire \resq[1]~119 ;
wire \resq[2]~114_cout ;
wire \resq[2]~115 ;
wire \resq[3]~1_sumout ;
wire \dout[20]~0_combout ;
wire \resq[3]~2 ;
wire \resq[3]~3 ;
wire \resq[4]~5_sumout ;
wire \resq[4]~6 ;
wire \resq[4]~7 ;
wire \resq[5]~9_sumout ;
wire \resq[5]~10 ;
wire \resq[5]~11 ;
wire \resq[6]~13_sumout ;
wire \resq[6]~14 ;
wire \resq[6]~15 ;
wire \resq[7]~17_sumout ;
wire \resq[7]~18 ;
wire \resq[7]~19 ;
wire \resq[8]~21_sumout ;
wire \resq[8]~22 ;
wire \resq[8]~23 ;
wire \resq[9]~25_sumout ;
wire \resq[9]~26 ;
wire \resq[9]~27 ;
wire \resq[10]~29_sumout ;
wire \resq[10]~30 ;
wire \resq[10]~31 ;
wire \resq[11]~33_sumout ;
wire \resq[11]~34 ;
wire \resq[11]~35 ;
wire \resq[12]~37_sumout ;
wire \resq[12]~38 ;
wire \resq[12]~39 ;
wire \resq[13]~41_sumout ;
wire \resq[13]~42 ;
wire \resq[13]~43 ;
wire \resq[14]~45_sumout ;
wire \resq[14]~46 ;
wire \resq[14]~47 ;
wire \resq[15]~49_sumout ;
wire \resq[15]~50 ;
wire \resq[15]~51 ;
wire \resq[16]~53_sumout ;
wire \resq[16]~54 ;
wire \resq[16]~55 ;
wire \resq[17]~57_sumout ;
wire \resq[17]~58 ;
wire \resq[17]~59 ;
wire \resq[18]~61_sumout ;
wire \resq[18]~62 ;
wire \resq[18]~63 ;
wire \resq[19]~65_sumout ;
wire \resq[19]~66 ;
wire \resq[19]~67 ;
wire \resq[20]~69_sumout ;
wire \resq[20]~70 ;
wire \resq[20]~71 ;
wire \resq[21]~73_sumout ;
wire \resq[21]~74 ;
wire \resq[21]~75 ;
wire \resq[22]~77_sumout ;
wire \resq[22]~78 ;
wire \resq[22]~79 ;
wire \resq[23]~81_sumout ;
wire \resq[23]~82 ;
wire \resq[23]~83 ;
wire \resq[24]~85_sumout ;
wire \resq[24]~86 ;
wire \resq[24]~87 ;
wire \resq[25]~89_sumout ;
wire \resq[25]~90 ;
wire \resq[25]~91 ;
wire \resq[26]~93_sumout ;
wire \resq[26]~94 ;
wire \resq[26]~95 ;
wire \resq[27]~97_sumout ;
wire \resq[27]~98 ;
wire \resq[27]~99 ;
wire \resq[28]~101_sumout ;
wire \resq[28]~102 ;
wire \resq[28]~103 ;
wire \resq[29]~105_sumout ;
wire \resq[29]~106 ;
wire \resq[29]~107 ;
wire \resq[30]~109_sumout ;


cic_auk_dspip_delay_7 \glogic:u0 (
	.datain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,dout_31,dout_301,dout_291,dout_281,dout_271,dout_261,dout_251,dout_241,dout_231,dout_221,dout_211,dout_201,dout_191,dout_181,dout_171,dout_161,dout_151,dout_141,dout_131,dout_121,dout_111,dout_101,dout_91,dout_81,dout_71,dout_61,
dout_51,dout_41,dout_32,dout_2,dout_1}),
	.register_fifofifo_data03(\glogic:u0|register_fifo:fifo_data[0][3]~q ),
	.register_fifofifo_data04(\glogic:u0|register_fifo:fifo_data[0][4]~q ),
	.register_fifofifo_data05(\glogic:u0|register_fifo:fifo_data[0][5]~q ),
	.register_fifofifo_data06(\glogic:u0|register_fifo:fifo_data[0][6]~q ),
	.register_fifofifo_data07(\glogic:u0|register_fifo:fifo_data[0][7]~q ),
	.register_fifofifo_data08(\glogic:u0|register_fifo:fifo_data[0][8]~q ),
	.register_fifofifo_data09(\glogic:u0|register_fifo:fifo_data[0][9]~q ),
	.register_fifofifo_data010(\glogic:u0|register_fifo:fifo_data[0][10]~q ),
	.register_fifofifo_data011(\glogic:u0|register_fifo:fifo_data[0][11]~q ),
	.register_fifofifo_data012(\glogic:u0|register_fifo:fifo_data[0][12]~q ),
	.register_fifofifo_data013(\glogic:u0|register_fifo:fifo_data[0][13]~q ),
	.register_fifofifo_data014(\glogic:u0|register_fifo:fifo_data[0][14]~q ),
	.register_fifofifo_data015(\glogic:u0|register_fifo:fifo_data[0][15]~q ),
	.register_fifofifo_data016(\glogic:u0|register_fifo:fifo_data[0][16]~q ),
	.register_fifofifo_data017(\glogic:u0|register_fifo:fifo_data[0][17]~q ),
	.register_fifofifo_data018(\glogic:u0|register_fifo:fifo_data[0][18]~q ),
	.register_fifofifo_data019(\glogic:u0|register_fifo:fifo_data[0][19]~q ),
	.register_fifofifo_data020(\glogic:u0|register_fifo:fifo_data[0][20]~q ),
	.register_fifofifo_data021(\glogic:u0|register_fifo:fifo_data[0][21]~q ),
	.register_fifofifo_data022(\glogic:u0|register_fifo:fifo_data[0][22]~q ),
	.register_fifofifo_data023(\glogic:u0|register_fifo:fifo_data[0][23]~q ),
	.register_fifofifo_data024(\glogic:u0|register_fifo:fifo_data[0][24]~q ),
	.register_fifofifo_data025(\glogic:u0|register_fifo:fifo_data[0][25]~q ),
	.register_fifofifo_data026(\glogic:u0|register_fifo:fifo_data[0][26]~q ),
	.register_fifofifo_data027(\glogic:u0|register_fifo:fifo_data[0][27]~q ),
	.register_fifofifo_data028(\glogic:u0|register_fifo:fifo_data[0][28]~q ),
	.register_fifofifo_data029(\glogic:u0|register_fifo:fifo_data[0][29]~q ),
	.register_fifofifo_data030(\glogic:u0|register_fifo:fifo_data[0][30]~q ),
	.enable(\dout~1_combout ),
	.register_fifofifo_data02(\glogic:u0|register_fifo:fifo_data[0][2]~q ),
	.register_fifofifo_data01(\glogic:u0|register_fifo:fifo_data[0][1]~q ),
	.register_fifofifo_data00(\glogic:u0|register_fifo:fifo_data[0][0]~q ),
	.clk(clk),
	.reset(reset_n));

arriav_lcell_comb \dout~1 (
	.dataa(!stall_reg),
	.datab(!dout_valid2),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dout~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dout~1 .extended_lut = "off";
defparam \dout~1 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \dout~1 .shared_arith = "off";

dffeas dout_valid(
	.clk(clk),
	.d(dout_valid2),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(dout_valid3),
	.q(dout_valid1),
	.prn(vcc));
defparam dout_valid.is_wysiwyg = "true";
defparam dout_valid.power_up = "low";

dffeas \dout[3] (
	.clk(clk),
	.d(\resq[3]~1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[20]~0_combout ),
	.q(dout_3),
	.prn(vcc));
defparam \dout[3] .is_wysiwyg = "true";
defparam \dout[3] .power_up = "low";

dffeas \dout[4] (
	.clk(clk),
	.d(\resq[4]~5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[20]~0_combout ),
	.q(dout_4),
	.prn(vcc));
defparam \dout[4] .is_wysiwyg = "true";
defparam \dout[4] .power_up = "low";

dffeas \dout[5] (
	.clk(clk),
	.d(\resq[5]~9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[20]~0_combout ),
	.q(dout_5),
	.prn(vcc));
defparam \dout[5] .is_wysiwyg = "true";
defparam \dout[5] .power_up = "low";

dffeas \dout[6] (
	.clk(clk),
	.d(\resq[6]~13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[20]~0_combout ),
	.q(dout_6),
	.prn(vcc));
defparam \dout[6] .is_wysiwyg = "true";
defparam \dout[6] .power_up = "low";

dffeas \dout[7] (
	.clk(clk),
	.d(\resq[7]~17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[20]~0_combout ),
	.q(dout_7),
	.prn(vcc));
defparam \dout[7] .is_wysiwyg = "true";
defparam \dout[7] .power_up = "low";

dffeas \dout[8] (
	.clk(clk),
	.d(\resq[8]~21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[20]~0_combout ),
	.q(dout_8),
	.prn(vcc));
defparam \dout[8] .is_wysiwyg = "true";
defparam \dout[8] .power_up = "low";

dffeas \dout[9] (
	.clk(clk),
	.d(\resq[9]~25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[20]~0_combout ),
	.q(dout_9),
	.prn(vcc));
defparam \dout[9] .is_wysiwyg = "true";
defparam \dout[9] .power_up = "low";

dffeas \dout[10] (
	.clk(clk),
	.d(\resq[10]~29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[20]~0_combout ),
	.q(dout_10),
	.prn(vcc));
defparam \dout[10] .is_wysiwyg = "true";
defparam \dout[10] .power_up = "low";

dffeas \dout[11] (
	.clk(clk),
	.d(\resq[11]~33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[20]~0_combout ),
	.q(dout_11),
	.prn(vcc));
defparam \dout[11] .is_wysiwyg = "true";
defparam \dout[11] .power_up = "low";

dffeas \dout[12] (
	.clk(clk),
	.d(\resq[12]~37_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[20]~0_combout ),
	.q(dout_12),
	.prn(vcc));
defparam \dout[12] .is_wysiwyg = "true";
defparam \dout[12] .power_up = "low";

dffeas \dout[13] (
	.clk(clk),
	.d(\resq[13]~41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[20]~0_combout ),
	.q(dout_13),
	.prn(vcc));
defparam \dout[13] .is_wysiwyg = "true";
defparam \dout[13] .power_up = "low";

dffeas \dout[14] (
	.clk(clk),
	.d(\resq[14]~45_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[20]~0_combout ),
	.q(dout_14),
	.prn(vcc));
defparam \dout[14] .is_wysiwyg = "true";
defparam \dout[14] .power_up = "low";

dffeas \dout[15] (
	.clk(clk),
	.d(\resq[15]~49_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[20]~0_combout ),
	.q(dout_15),
	.prn(vcc));
defparam \dout[15] .is_wysiwyg = "true";
defparam \dout[15] .power_up = "low";

dffeas \dout[16] (
	.clk(clk),
	.d(\resq[16]~53_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[20]~0_combout ),
	.q(dout_16),
	.prn(vcc));
defparam \dout[16] .is_wysiwyg = "true";
defparam \dout[16] .power_up = "low";

dffeas \dout[17] (
	.clk(clk),
	.d(\resq[17]~57_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[20]~0_combout ),
	.q(dout_17),
	.prn(vcc));
defparam \dout[17] .is_wysiwyg = "true";
defparam \dout[17] .power_up = "low";

dffeas \dout[18] (
	.clk(clk),
	.d(\resq[18]~61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[20]~0_combout ),
	.q(dout_18),
	.prn(vcc));
defparam \dout[18] .is_wysiwyg = "true";
defparam \dout[18] .power_up = "low";

dffeas \dout[19] (
	.clk(clk),
	.d(\resq[19]~65_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[20]~0_combout ),
	.q(dout_19),
	.prn(vcc));
defparam \dout[19] .is_wysiwyg = "true";
defparam \dout[19] .power_up = "low";

dffeas \dout[20] (
	.clk(clk),
	.d(\resq[20]~69_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[20]~0_combout ),
	.q(dout_20),
	.prn(vcc));
defparam \dout[20] .is_wysiwyg = "true";
defparam \dout[20] .power_up = "low";

dffeas \dout[21] (
	.clk(clk),
	.d(\resq[21]~73_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[20]~0_combout ),
	.q(dout_21),
	.prn(vcc));
defparam \dout[21] .is_wysiwyg = "true";
defparam \dout[21] .power_up = "low";

dffeas \dout[22] (
	.clk(clk),
	.d(\resq[22]~77_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[20]~0_combout ),
	.q(dout_22),
	.prn(vcc));
defparam \dout[22] .is_wysiwyg = "true";
defparam \dout[22] .power_up = "low";

dffeas \dout[23] (
	.clk(clk),
	.d(\resq[23]~81_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[20]~0_combout ),
	.q(dout_23),
	.prn(vcc));
defparam \dout[23] .is_wysiwyg = "true";
defparam \dout[23] .power_up = "low";

dffeas \dout[24] (
	.clk(clk),
	.d(\resq[24]~85_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[20]~0_combout ),
	.q(dout_24),
	.prn(vcc));
defparam \dout[24] .is_wysiwyg = "true";
defparam \dout[24] .power_up = "low";

dffeas \dout[25] (
	.clk(clk),
	.d(\resq[25]~89_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[20]~0_combout ),
	.q(dout_25),
	.prn(vcc));
defparam \dout[25] .is_wysiwyg = "true";
defparam \dout[25] .power_up = "low";

dffeas \dout[26] (
	.clk(clk),
	.d(\resq[26]~93_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[20]~0_combout ),
	.q(dout_26),
	.prn(vcc));
defparam \dout[26] .is_wysiwyg = "true";
defparam \dout[26] .power_up = "low";

dffeas \dout[27] (
	.clk(clk),
	.d(\resq[27]~97_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[20]~0_combout ),
	.q(dout_27),
	.prn(vcc));
defparam \dout[27] .is_wysiwyg = "true";
defparam \dout[27] .power_up = "low";

dffeas \dout[28] (
	.clk(clk),
	.d(\resq[28]~101_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[20]~0_combout ),
	.q(dout_28),
	.prn(vcc));
defparam \dout[28] .is_wysiwyg = "true";
defparam \dout[28] .power_up = "low";

dffeas \dout[29] (
	.clk(clk),
	.d(\resq[29]~105_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[20]~0_combout ),
	.q(dout_29),
	.prn(vcc));
defparam \dout[29] .is_wysiwyg = "true";
defparam \dout[29] .power_up = "low";

dffeas \dout[30] (
	.clk(clk),
	.d(\resq[30]~109_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[20]~0_combout ),
	.q(dout_30),
	.prn(vcc));
defparam \dout[30] .is_wysiwyg = "true";
defparam \dout[30] .power_up = "low";

arriav_lcell_comb \dout_valid~0 (
	.dataa(!reset_n),
	.datab(!stall_reg),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(dout_valid3),
	.sumout(),
	.cout(),
	.shareout());
defparam \dout_valid~0 .extended_lut = "off";
defparam \dout_valid~0 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \dout_valid~0 .shared_arith = "off";

arriav_lcell_comb \resq[0]~122 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][0]~q ),
	.datad(!dout_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\resq[0]~122_cout ),
	.shareout(\resq[0]~123 ));
defparam \resq[0]~122 .extended_lut = "off";
defparam \resq[0]~122 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[0]~122 .shared_arith = "on";

arriav_lcell_comb \resq[1]~118 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][1]~q ),
	.datad(!dout_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[0]~122_cout ),
	.sharein(\resq[0]~123 ),
	.combout(),
	.sumout(),
	.cout(\resq[1]~118_cout ),
	.shareout(\resq[1]~119 ));
defparam \resq[1]~118 .extended_lut = "off";
defparam \resq[1]~118 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[1]~118 .shared_arith = "on";

arriav_lcell_comb \resq[2]~114 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][2]~q ),
	.datad(!dout_32),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[1]~118_cout ),
	.sharein(\resq[1]~119 ),
	.combout(),
	.sumout(),
	.cout(\resq[2]~114_cout ),
	.shareout(\resq[2]~115 ));
defparam \resq[2]~114 .extended_lut = "off";
defparam \resq[2]~114 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[2]~114 .shared_arith = "on";

arriav_lcell_comb \resq[3]~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][3]~q ),
	.datad(!dout_41),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[2]~114_cout ),
	.sharein(\resq[2]~115 ),
	.combout(),
	.sumout(\resq[3]~1_sumout ),
	.cout(\resq[3]~2 ),
	.shareout(\resq[3]~3 ));
defparam \resq[3]~1 .extended_lut = "off";
defparam \resq[3]~1 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[3]~1 .shared_arith = "on";

arriav_lcell_comb \dout[20]~0 (
	.dataa(!reset_n),
	.datab(!stall_reg),
	.datac(!dout_valid2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dout[20]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dout[20]~0 .extended_lut = "off";
defparam \dout[20]~0 .lut_mask = 64'hEFEFEFEFEFEFEFEF;
defparam \dout[20]~0 .shared_arith = "off";

arriav_lcell_comb \resq[4]~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][4]~q ),
	.datad(!dout_51),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[3]~2 ),
	.sharein(\resq[3]~3 ),
	.combout(),
	.sumout(\resq[4]~5_sumout ),
	.cout(\resq[4]~6 ),
	.shareout(\resq[4]~7 ));
defparam \resq[4]~5 .extended_lut = "off";
defparam \resq[4]~5 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[4]~5 .shared_arith = "on";

arriav_lcell_comb \resq[5]~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][5]~q ),
	.datad(!dout_61),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[4]~6 ),
	.sharein(\resq[4]~7 ),
	.combout(),
	.sumout(\resq[5]~9_sumout ),
	.cout(\resq[5]~10 ),
	.shareout(\resq[5]~11 ));
defparam \resq[5]~9 .extended_lut = "off";
defparam \resq[5]~9 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[5]~9 .shared_arith = "on";

arriav_lcell_comb \resq[6]~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][6]~q ),
	.datad(!dout_71),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[5]~10 ),
	.sharein(\resq[5]~11 ),
	.combout(),
	.sumout(\resq[6]~13_sumout ),
	.cout(\resq[6]~14 ),
	.shareout(\resq[6]~15 ));
defparam \resq[6]~13 .extended_lut = "off";
defparam \resq[6]~13 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[6]~13 .shared_arith = "on";

arriav_lcell_comb \resq[7]~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][7]~q ),
	.datad(!dout_81),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[6]~14 ),
	.sharein(\resq[6]~15 ),
	.combout(),
	.sumout(\resq[7]~17_sumout ),
	.cout(\resq[7]~18 ),
	.shareout(\resq[7]~19 ));
defparam \resq[7]~17 .extended_lut = "off";
defparam \resq[7]~17 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[7]~17 .shared_arith = "on";

arriav_lcell_comb \resq[8]~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][8]~q ),
	.datad(!dout_91),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[7]~18 ),
	.sharein(\resq[7]~19 ),
	.combout(),
	.sumout(\resq[8]~21_sumout ),
	.cout(\resq[8]~22 ),
	.shareout(\resq[8]~23 ));
defparam \resq[8]~21 .extended_lut = "off";
defparam \resq[8]~21 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[8]~21 .shared_arith = "on";

arriav_lcell_comb \resq[9]~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][9]~q ),
	.datad(!dout_101),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[8]~22 ),
	.sharein(\resq[8]~23 ),
	.combout(),
	.sumout(\resq[9]~25_sumout ),
	.cout(\resq[9]~26 ),
	.shareout(\resq[9]~27 ));
defparam \resq[9]~25 .extended_lut = "off";
defparam \resq[9]~25 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[9]~25 .shared_arith = "on";

arriav_lcell_comb \resq[10]~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][10]~q ),
	.datad(!dout_111),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[9]~26 ),
	.sharein(\resq[9]~27 ),
	.combout(),
	.sumout(\resq[10]~29_sumout ),
	.cout(\resq[10]~30 ),
	.shareout(\resq[10]~31 ));
defparam \resq[10]~29 .extended_lut = "off";
defparam \resq[10]~29 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[10]~29 .shared_arith = "on";

arriav_lcell_comb \resq[11]~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][11]~q ),
	.datad(!dout_121),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[10]~30 ),
	.sharein(\resq[10]~31 ),
	.combout(),
	.sumout(\resq[11]~33_sumout ),
	.cout(\resq[11]~34 ),
	.shareout(\resq[11]~35 ));
defparam \resq[11]~33 .extended_lut = "off";
defparam \resq[11]~33 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[11]~33 .shared_arith = "on";

arriav_lcell_comb \resq[12]~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][12]~q ),
	.datad(!dout_131),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[11]~34 ),
	.sharein(\resq[11]~35 ),
	.combout(),
	.sumout(\resq[12]~37_sumout ),
	.cout(\resq[12]~38 ),
	.shareout(\resq[12]~39 ));
defparam \resq[12]~37 .extended_lut = "off";
defparam \resq[12]~37 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[12]~37 .shared_arith = "on";

arriav_lcell_comb \resq[13]~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][13]~q ),
	.datad(!dout_141),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[12]~38 ),
	.sharein(\resq[12]~39 ),
	.combout(),
	.sumout(\resq[13]~41_sumout ),
	.cout(\resq[13]~42 ),
	.shareout(\resq[13]~43 ));
defparam \resq[13]~41 .extended_lut = "off";
defparam \resq[13]~41 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[13]~41 .shared_arith = "on";

arriav_lcell_comb \resq[14]~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][14]~q ),
	.datad(!dout_151),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[13]~42 ),
	.sharein(\resq[13]~43 ),
	.combout(),
	.sumout(\resq[14]~45_sumout ),
	.cout(\resq[14]~46 ),
	.shareout(\resq[14]~47 ));
defparam \resq[14]~45 .extended_lut = "off";
defparam \resq[14]~45 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[14]~45 .shared_arith = "on";

arriav_lcell_comb \resq[15]~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][15]~q ),
	.datad(!dout_161),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[14]~46 ),
	.sharein(\resq[14]~47 ),
	.combout(),
	.sumout(\resq[15]~49_sumout ),
	.cout(\resq[15]~50 ),
	.shareout(\resq[15]~51 ));
defparam \resq[15]~49 .extended_lut = "off";
defparam \resq[15]~49 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[15]~49 .shared_arith = "on";

arriav_lcell_comb \resq[16]~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][16]~q ),
	.datad(!dout_171),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[15]~50 ),
	.sharein(\resq[15]~51 ),
	.combout(),
	.sumout(\resq[16]~53_sumout ),
	.cout(\resq[16]~54 ),
	.shareout(\resq[16]~55 ));
defparam \resq[16]~53 .extended_lut = "off";
defparam \resq[16]~53 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[16]~53 .shared_arith = "on";

arriav_lcell_comb \resq[17]~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][17]~q ),
	.datad(!dout_181),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[16]~54 ),
	.sharein(\resq[16]~55 ),
	.combout(),
	.sumout(\resq[17]~57_sumout ),
	.cout(\resq[17]~58 ),
	.shareout(\resq[17]~59 ));
defparam \resq[17]~57 .extended_lut = "off";
defparam \resq[17]~57 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[17]~57 .shared_arith = "on";

arriav_lcell_comb \resq[18]~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][18]~q ),
	.datad(!dout_191),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[17]~58 ),
	.sharein(\resq[17]~59 ),
	.combout(),
	.sumout(\resq[18]~61_sumout ),
	.cout(\resq[18]~62 ),
	.shareout(\resq[18]~63 ));
defparam \resq[18]~61 .extended_lut = "off";
defparam \resq[18]~61 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[18]~61 .shared_arith = "on";

arriav_lcell_comb \resq[19]~65 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][19]~q ),
	.datad(!dout_201),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[18]~62 ),
	.sharein(\resq[18]~63 ),
	.combout(),
	.sumout(\resq[19]~65_sumout ),
	.cout(\resq[19]~66 ),
	.shareout(\resq[19]~67 ));
defparam \resq[19]~65 .extended_lut = "off";
defparam \resq[19]~65 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[19]~65 .shared_arith = "on";

arriav_lcell_comb \resq[20]~69 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][20]~q ),
	.datad(!dout_211),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[19]~66 ),
	.sharein(\resq[19]~67 ),
	.combout(),
	.sumout(\resq[20]~69_sumout ),
	.cout(\resq[20]~70 ),
	.shareout(\resq[20]~71 ));
defparam \resq[20]~69 .extended_lut = "off";
defparam \resq[20]~69 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[20]~69 .shared_arith = "on";

arriav_lcell_comb \resq[21]~73 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][21]~q ),
	.datad(!dout_221),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[20]~70 ),
	.sharein(\resq[20]~71 ),
	.combout(),
	.sumout(\resq[21]~73_sumout ),
	.cout(\resq[21]~74 ),
	.shareout(\resq[21]~75 ));
defparam \resq[21]~73 .extended_lut = "off";
defparam \resq[21]~73 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[21]~73 .shared_arith = "on";

arriav_lcell_comb \resq[22]~77 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][22]~q ),
	.datad(!dout_231),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[21]~74 ),
	.sharein(\resq[21]~75 ),
	.combout(),
	.sumout(\resq[22]~77_sumout ),
	.cout(\resq[22]~78 ),
	.shareout(\resq[22]~79 ));
defparam \resq[22]~77 .extended_lut = "off";
defparam \resq[22]~77 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[22]~77 .shared_arith = "on";

arriav_lcell_comb \resq[23]~81 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][23]~q ),
	.datad(!dout_241),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[22]~78 ),
	.sharein(\resq[22]~79 ),
	.combout(),
	.sumout(\resq[23]~81_sumout ),
	.cout(\resq[23]~82 ),
	.shareout(\resq[23]~83 ));
defparam \resq[23]~81 .extended_lut = "off";
defparam \resq[23]~81 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[23]~81 .shared_arith = "on";

arriav_lcell_comb \resq[24]~85 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][24]~q ),
	.datad(!dout_251),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[23]~82 ),
	.sharein(\resq[23]~83 ),
	.combout(),
	.sumout(\resq[24]~85_sumout ),
	.cout(\resq[24]~86 ),
	.shareout(\resq[24]~87 ));
defparam \resq[24]~85 .extended_lut = "off";
defparam \resq[24]~85 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[24]~85 .shared_arith = "on";

arriav_lcell_comb \resq[25]~89 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][25]~q ),
	.datad(!dout_261),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[24]~86 ),
	.sharein(\resq[24]~87 ),
	.combout(),
	.sumout(\resq[25]~89_sumout ),
	.cout(\resq[25]~90 ),
	.shareout(\resq[25]~91 ));
defparam \resq[25]~89 .extended_lut = "off";
defparam \resq[25]~89 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[25]~89 .shared_arith = "on";

arriav_lcell_comb \resq[26]~93 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][26]~q ),
	.datad(!dout_271),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[25]~90 ),
	.sharein(\resq[25]~91 ),
	.combout(),
	.sumout(\resq[26]~93_sumout ),
	.cout(\resq[26]~94 ),
	.shareout(\resq[26]~95 ));
defparam \resq[26]~93 .extended_lut = "off";
defparam \resq[26]~93 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[26]~93 .shared_arith = "on";

arriav_lcell_comb \resq[27]~97 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][27]~q ),
	.datad(!dout_281),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[26]~94 ),
	.sharein(\resq[26]~95 ),
	.combout(),
	.sumout(\resq[27]~97_sumout ),
	.cout(\resq[27]~98 ),
	.shareout(\resq[27]~99 ));
defparam \resq[27]~97 .extended_lut = "off";
defparam \resq[27]~97 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[27]~97 .shared_arith = "on";

arriav_lcell_comb \resq[28]~101 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][28]~q ),
	.datad(!dout_291),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[27]~98 ),
	.sharein(\resq[27]~99 ),
	.combout(),
	.sumout(\resq[28]~101_sumout ),
	.cout(\resq[28]~102 ),
	.shareout(\resq[28]~103 ));
defparam \resq[28]~101 .extended_lut = "off";
defparam \resq[28]~101 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[28]~101 .shared_arith = "on";

arriav_lcell_comb \resq[29]~105 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][29]~q ),
	.datad(!dout_301),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[28]~102 ),
	.sharein(\resq[28]~103 ),
	.combout(),
	.sumout(\resq[29]~105_sumout ),
	.cout(\resq[29]~106 ),
	.shareout(\resq[29]~107 ));
defparam \resq[29]~105 .extended_lut = "off";
defparam \resq[29]~105 .lut_mask = 64'h0000F0FF00000FF0;
defparam \resq[29]~105 .shared_arith = "on";

arriav_lcell_comb \resq[30]~109 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\glogic:u0|register_fifo:fifo_data[0][30]~q ),
	.datad(!dout_31),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\resq[29]~106 ),
	.sharein(\resq[29]~107 ),
	.combout(),
	.sumout(\resq[30]~109_sumout ),
	.cout(),
	.shareout());
defparam \resq[30]~109 .extended_lut = "off";
defparam \resq[30]~109 .lut_mask = 64'h0000000000000FF0;
defparam \resq[30]~109 .shared_arith = "on";

endmodule

module cic_auk_dspip_delay_7 (
	datain,
	register_fifofifo_data03,
	register_fifofifo_data04,
	register_fifofifo_data05,
	register_fifofifo_data06,
	register_fifofifo_data07,
	register_fifofifo_data08,
	register_fifofifo_data09,
	register_fifofifo_data010,
	register_fifofifo_data011,
	register_fifofifo_data012,
	register_fifofifo_data013,
	register_fifofifo_data014,
	register_fifofifo_data015,
	register_fifofifo_data016,
	register_fifofifo_data017,
	register_fifofifo_data018,
	register_fifofifo_data019,
	register_fifofifo_data020,
	register_fifofifo_data021,
	register_fifofifo_data022,
	register_fifofifo_data023,
	register_fifofifo_data024,
	register_fifofifo_data025,
	register_fifofifo_data026,
	register_fifofifo_data027,
	register_fifofifo_data028,
	register_fifofifo_data029,
	register_fifofifo_data030,
	enable,
	register_fifofifo_data02,
	register_fifofifo_data01,
	register_fifofifo_data00,
	clk,
	reset)/* synthesis synthesis_greybox=1 */;
input 	[46:0] datain;
output 	register_fifofifo_data03;
output 	register_fifofifo_data04;
output 	register_fifofifo_data05;
output 	register_fifofifo_data06;
output 	register_fifofifo_data07;
output 	register_fifofifo_data08;
output 	register_fifofifo_data09;
output 	register_fifofifo_data010;
output 	register_fifofifo_data011;
output 	register_fifofifo_data012;
output 	register_fifofifo_data013;
output 	register_fifofifo_data014;
output 	register_fifofifo_data015;
output 	register_fifofifo_data016;
output 	register_fifofifo_data017;
output 	register_fifofifo_data018;
output 	register_fifofifo_data019;
output 	register_fifofifo_data020;
output 	register_fifofifo_data021;
output 	register_fifofifo_data022;
output 	register_fifofifo_data023;
output 	register_fifofifo_data024;
output 	register_fifofifo_data025;
output 	register_fifofifo_data026;
output 	register_fifofifo_data027;
output 	register_fifofifo_data028;
output 	register_fifofifo_data029;
output 	register_fifofifo_data030;
input 	enable;
output 	register_fifofifo_data02;
output 	register_fifofifo_data01;
output 	register_fifofifo_data00;
input 	clk;
input 	reset;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \register_fifo:fifo_data[0][3] (
	.clk(clk),
	.d(datain[3]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data03),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][3] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][3] .power_up = "low";

dffeas \register_fifo:fifo_data[0][4] (
	.clk(clk),
	.d(datain[4]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data04),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][4] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][4] .power_up = "low";

dffeas \register_fifo:fifo_data[0][5] (
	.clk(clk),
	.d(datain[5]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data05),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][5] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][5] .power_up = "low";

dffeas \register_fifo:fifo_data[0][6] (
	.clk(clk),
	.d(datain[6]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data06),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][6] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][6] .power_up = "low";

dffeas \register_fifo:fifo_data[0][7] (
	.clk(clk),
	.d(datain[7]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data07),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][7] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][7] .power_up = "low";

dffeas \register_fifo:fifo_data[0][8] (
	.clk(clk),
	.d(datain[8]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data08),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][8] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][8] .power_up = "low";

dffeas \register_fifo:fifo_data[0][9] (
	.clk(clk),
	.d(datain[9]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data09),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][9] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][9] .power_up = "low";

dffeas \register_fifo:fifo_data[0][10] (
	.clk(clk),
	.d(datain[10]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data010),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][10] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][10] .power_up = "low";

dffeas \register_fifo:fifo_data[0][11] (
	.clk(clk),
	.d(datain[11]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data011),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][11] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][11] .power_up = "low";

dffeas \register_fifo:fifo_data[0][12] (
	.clk(clk),
	.d(datain[12]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data012),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][12] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][12] .power_up = "low";

dffeas \register_fifo:fifo_data[0][13] (
	.clk(clk),
	.d(datain[13]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data013),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][13] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][13] .power_up = "low";

dffeas \register_fifo:fifo_data[0][14] (
	.clk(clk),
	.d(datain[14]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data014),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][14] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][14] .power_up = "low";

dffeas \register_fifo:fifo_data[0][15] (
	.clk(clk),
	.d(datain[15]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data015),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][15] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][15] .power_up = "low";

dffeas \register_fifo:fifo_data[0][16] (
	.clk(clk),
	.d(datain[16]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data016),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][16] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][16] .power_up = "low";

dffeas \register_fifo:fifo_data[0][17] (
	.clk(clk),
	.d(datain[17]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data017),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][17] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][17] .power_up = "low";

dffeas \register_fifo:fifo_data[0][18] (
	.clk(clk),
	.d(datain[18]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data018),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][18] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][18] .power_up = "low";

dffeas \register_fifo:fifo_data[0][19] (
	.clk(clk),
	.d(datain[19]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data019),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][19] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][19] .power_up = "low";

dffeas \register_fifo:fifo_data[0][20] (
	.clk(clk),
	.d(datain[20]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data020),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][20] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][20] .power_up = "low";

dffeas \register_fifo:fifo_data[0][21] (
	.clk(clk),
	.d(datain[21]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data021),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][21] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][21] .power_up = "low";

dffeas \register_fifo:fifo_data[0][22] (
	.clk(clk),
	.d(datain[22]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data022),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][22] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][22] .power_up = "low";

dffeas \register_fifo:fifo_data[0][23] (
	.clk(clk),
	.d(datain[23]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data023),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][23] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][23] .power_up = "low";

dffeas \register_fifo:fifo_data[0][24] (
	.clk(clk),
	.d(datain[24]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data024),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][24] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][24] .power_up = "low";

dffeas \register_fifo:fifo_data[0][25] (
	.clk(clk),
	.d(datain[25]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data025),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][25] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][25] .power_up = "low";

dffeas \register_fifo:fifo_data[0][26] (
	.clk(clk),
	.d(datain[26]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data026),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][26] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][26] .power_up = "low";

dffeas \register_fifo:fifo_data[0][27] (
	.clk(clk),
	.d(datain[27]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data027),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][27] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][27] .power_up = "low";

dffeas \register_fifo:fifo_data[0][28] (
	.clk(clk),
	.d(datain[28]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data028),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][28] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][28] .power_up = "low";

dffeas \register_fifo:fifo_data[0][29] (
	.clk(clk),
	.d(datain[29]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data029),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][29] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][29] .power_up = "low";

dffeas \register_fifo:fifo_data[0][30] (
	.clk(clk),
	.d(datain[30]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data030),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][30] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][30] .power_up = "low";

dffeas \register_fifo:fifo_data[0][2] (
	.clk(clk),
	.d(datain[2]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data02),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][2] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][2] .power_up = "low";

dffeas \register_fifo:fifo_data[0][1] (
	.clk(clk),
	.d(datain[1]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data01),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][1] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][1] .power_up = "low";

dffeas \register_fifo:fifo_data[0][0] (
	.clk(clk),
	.d(datain[0]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(register_fifofifo_data00),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][0] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][0] .power_up = "low";

endmodule

module cic_auk_dspip_downsample (
	sample_state_0,
	stall_reg,
	count_0,
	count_3,
	count_1,
	count_2,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	sample_state_0;
input 	stall_reg;
output 	count_0;
output 	count_3;
output 	count_1;
output 	count_2;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cic_counter_module_1 counter_fs_inst(
	.sample_state_0(sample_state_0),
	.stall_reg(stall_reg),
	.count_0(count_0),
	.count_3(count_3),
	.count_1(count_1),
	.count_2(count_2),
	.clk(clk),
	.reset_n(reset_n));

endmodule

module cic_counter_module_1 (
	sample_state_0,
	stall_reg,
	count_0,
	count_3,
	count_1,
	count_2,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	sample_state_0;
input 	stall_reg;
output 	count_0;
output 	count_3;
output 	count_1;
output 	count_2;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \count~0_combout ;
wire \count[1]~1_combout ;
wire \count~2_combout ;
wire \count~3_combout ;
wire \count~4_combout ;


dffeas \count[0] (
	.clk(clk),
	.d(\count~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\count[1]~1_combout ),
	.q(count_0),
	.prn(vcc));
defparam \count[0] .is_wysiwyg = "true";
defparam \count[0] .power_up = "low";

dffeas \count[3] (
	.clk(clk),
	.d(\count~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\count[1]~1_combout ),
	.q(count_3),
	.prn(vcc));
defparam \count[3] .is_wysiwyg = "true";
defparam \count[3] .power_up = "low";

dffeas \count[1] (
	.clk(clk),
	.d(\count~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\count[1]~1_combout ),
	.q(count_1),
	.prn(vcc));
defparam \count[1] .is_wysiwyg = "true";
defparam \count[1] .power_up = "low";

dffeas \count[2] (
	.clk(clk),
	.d(\count~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\count[1]~1_combout ),
	.q(count_2),
	.prn(vcc));
defparam \count[2] .is_wysiwyg = "true";
defparam \count[2] .power_up = "low";

arriav_lcell_comb \count~0 (
	.dataa(!reset_n),
	.datab(!count_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\count~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \count~0 .extended_lut = "off";
defparam \count~0 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \count~0 .shared_arith = "off";

arriav_lcell_comb \count[1]~1 (
	.dataa(!reset_n),
	.datab(!stall_reg),
	.datac(!sample_state_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\count[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \count[1]~1 .extended_lut = "off";
defparam \count[1]~1 .lut_mask = 64'hEFEFEFEFEFEFEFEF;
defparam \count[1]~1 .shared_arith = "off";

arriav_lcell_comb \count~2 (
	.dataa(!reset_n),
	.datab(!count_0),
	.datac(!count_3),
	.datad(!count_1),
	.datae(!count_2),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\count~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \count~2 .extended_lut = "off";
defparam \count~2 .lut_mask = 64'h7DD7D77D7DD7D77D;
defparam \count~2 .shared_arith = "off";

arriav_lcell_comb \count~3 (
	.dataa(!reset_n),
	.datab(!count_0),
	.datac(!count_3),
	.datad(!count_1),
	.datae(!count_2),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\count~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \count~3 .extended_lut = "off";
defparam \count~3 .lut_mask = 64'hF7FDFFFFF7FDFFFF;
defparam \count~3 .shared_arith = "off";

arriav_lcell_comb \count~4 (
	.dataa(!reset_n),
	.datab(!count_0),
	.datac(gnd),
	.datad(!count_1),
	.datae(!count_2),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\count~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \count~4 .extended_lut = "off";
defparam \count~4 .lut_mask = 64'hDD7777DDDD7777DD;
defparam \count~4 .shared_arith = "off";

endmodule

module cic_auk_dspip_integrator (
	q_b_19,
	q_b_18,
	q_b_17,
	q_b_16,
	q_b_15,
	q_b_14,
	q_b_13,
	q_b_12,
	q_b_11,
	q_b_10,
	q_b_9,
	q_b_8,
	q_b_7,
	q_b_6,
	q_b_5,
	q_b_4,
	q_b_3,
	q_b_2,
	q_b_1,
	q_b_0,
	stall_reg,
	register_fifofifo_data019,
	register_fifofifo_data020,
	register_fifofifo_data021,
	register_fifofifo_data022,
	register_fifofifo_data023,
	register_fifofifo_data024,
	register_fifofifo_data025,
	register_fifofifo_data026,
	register_fifofifo_data027,
	register_fifofifo_data028,
	register_fifofifo_data029,
	register_fifofifo_data030,
	register_fifofifo_data031,
	register_fifofifo_data032,
	register_fifofifo_data033,
	register_fifofifo_data034,
	register_fifofifo_data035,
	register_fifofifo_data036,
	register_fifofifo_data037,
	register_fifofifo_data038,
	register_fifofifo_data039,
	register_fifofifo_data040,
	register_fifofifo_data041,
	register_fifofifo_data042,
	register_fifofifo_data043,
	register_fifofifo_data044,
	register_fifofifo_data045,
	register_fifofifo_data046,
	register_fifofifo_data018,
	register_fifofifo_data017,
	register_fifofifo_data016,
	register_fifofifo_data015,
	register_fifofifo_data014,
	register_fifofifo_data013,
	register_fifofifo_data012,
	register_fifofifo_data011,
	register_fifofifo_data010,
	register_fifofifo_data09,
	register_fifofifo_data08,
	register_fifofifo_data07,
	register_fifofifo_data06,
	register_fifofifo_data05,
	register_fifofifo_data04,
	register_fifofifo_data03,
	register_fifofifo_data02,
	register_fifofifo_data01,
	register_fifofifo_data00,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	q_b_19;
input 	q_b_18;
input 	q_b_17;
input 	q_b_16;
input 	q_b_15;
input 	q_b_14;
input 	q_b_13;
input 	q_b_12;
input 	q_b_11;
input 	q_b_10;
input 	q_b_9;
input 	q_b_8;
input 	q_b_7;
input 	q_b_6;
input 	q_b_5;
input 	q_b_4;
input 	q_b_3;
input 	q_b_2;
input 	q_b_1;
input 	q_b_0;
input 	stall_reg;
output 	register_fifofifo_data019;
output 	register_fifofifo_data020;
output 	register_fifofifo_data021;
output 	register_fifofifo_data022;
output 	register_fifofifo_data023;
output 	register_fifofifo_data024;
output 	register_fifofifo_data025;
output 	register_fifofifo_data026;
output 	register_fifofifo_data027;
output 	register_fifofifo_data028;
output 	register_fifofifo_data029;
output 	register_fifofifo_data030;
output 	register_fifofifo_data031;
output 	register_fifofifo_data032;
output 	register_fifofifo_data033;
output 	register_fifofifo_data034;
output 	register_fifofifo_data035;
output 	register_fifofifo_data036;
output 	register_fifofifo_data037;
output 	register_fifofifo_data038;
output 	register_fifofifo_data039;
output 	register_fifofifo_data040;
output 	register_fifofifo_data041;
output 	register_fifofifo_data042;
output 	register_fifofifo_data043;
output 	register_fifofifo_data044;
output 	register_fifofifo_data045;
output 	register_fifofifo_data046;
output 	register_fifofifo_data018;
output 	register_fifofifo_data017;
output 	register_fifofifo_data016;
output 	register_fifofifo_data015;
output 	register_fifofifo_data014;
output 	register_fifofifo_data013;
output 	register_fifofifo_data012;
output 	register_fifofifo_data011;
output 	register_fifofifo_data010;
output 	register_fifofifo_data09;
output 	register_fifofifo_data08;
output 	register_fifofifo_data07;
output 	register_fifofifo_data06;
output 	register_fifofifo_data05;
output 	register_fifofifo_data04;
output 	register_fifofifo_data03;
output 	register_fifofifo_data02;
output 	register_fifofifo_data01;
output 	register_fifofifo_data00;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Add0~1_sumout ;
wire \Add0~2 ;
wire \Add0~5_sumout ;
wire \Add0~6 ;
wire \Add0~9_sumout ;
wire \Add0~10 ;
wire \Add0~13_sumout ;
wire \Add0~14 ;
wire \Add0~17_sumout ;
wire \Add0~18 ;
wire \Add0~21_sumout ;
wire \Add0~22 ;
wire \Add0~25_sumout ;
wire \Add0~26 ;
wire \Add0~29_sumout ;
wire \Add0~30 ;
wire \Add0~33_sumout ;
wire \Add0~34 ;
wire \Add0~37_sumout ;
wire \Add0~38 ;
wire \Add0~41_sumout ;
wire \Add0~42 ;
wire \Add0~45_sumout ;
wire \Add0~46 ;
wire \Add0~49_sumout ;
wire \Add0~50 ;
wire \Add0~53_sumout ;
wire \Add0~54 ;
wire \Add0~57_sumout ;
wire \Add0~58 ;
wire \Add0~61_sumout ;
wire \Add0~62 ;
wire \Add0~65_sumout ;
wire \Add0~66 ;
wire \Add0~69_sumout ;
wire \Add0~70 ;
wire \Add0~73_sumout ;
wire \Add0~74 ;
wire \Add0~77_sumout ;
wire \Add0~78 ;
wire \Add0~81_sumout ;
wire \Add0~82 ;
wire \Add0~85_sumout ;
wire \Add0~86 ;
wire \Add0~89_sumout ;
wire \Add0~90 ;
wire \Add0~93_sumout ;
wire \Add0~94 ;
wire \Add0~97_sumout ;
wire \Add0~98 ;
wire \Add0~101_sumout ;
wire \Add0~102 ;
wire \Add0~105_sumout ;
wire \Add0~106 ;
wire \Add0~109_sumout ;
wire \Add0~113_sumout ;
wire \Add0~114 ;
wire \Add0~117_sumout ;
wire \Add0~118 ;
wire \Add0~121_sumout ;
wire \Add0~122 ;
wire \Add0~125_sumout ;
wire \Add0~126 ;
wire \Add0~129_sumout ;
wire \Add0~130 ;
wire \Add0~133_sumout ;
wire \Add0~134 ;
wire \Add0~137_sumout ;
wire \Add0~138 ;
wire \Add0~141_sumout ;
wire \Add0~142 ;
wire \Add0~145_sumout ;
wire \Add0~146 ;
wire \Add0~149_sumout ;
wire \Add0~150 ;
wire \Add0~153_sumout ;
wire \Add0~154 ;
wire \Add0~157_sumout ;
wire \Add0~158 ;
wire \Add0~161_sumout ;
wire \Add0~162 ;
wire \Add0~165_sumout ;
wire \Add0~166 ;
wire \Add0~169_sumout ;
wire \Add0~170 ;
wire \Add0~173_sumout ;
wire \Add0~174 ;
wire \Add0~177_sumout ;
wire \Add0~178 ;
wire \Add0~181_sumout ;
wire \Add0~182 ;
wire \Add0~185_sumout ;
wire \Add0~186 ;


cic_auk_dspip_delay_8 \glogic:integrator_pipeline_0_generate:u1 (
	.datain({\Add0~109_sumout ,\Add0~105_sumout ,\Add0~101_sumout ,\Add0~97_sumout ,\Add0~93_sumout ,\Add0~89_sumout ,\Add0~85_sumout ,\Add0~81_sumout ,\Add0~77_sumout ,\Add0~73_sumout ,\Add0~69_sumout ,\Add0~65_sumout ,\Add0~61_sumout ,\Add0~57_sumout ,\Add0~53_sumout ,
\Add0~49_sumout ,\Add0~45_sumout ,\Add0~41_sumout ,\Add0~37_sumout ,\Add0~33_sumout ,\Add0~29_sumout ,\Add0~25_sumout ,\Add0~21_sumout ,\Add0~17_sumout ,\Add0~13_sumout ,\Add0~9_sumout ,\Add0~5_sumout ,\Add0~1_sumout ,\Add0~113_sumout ,\Add0~117_sumout ,\Add0~121_sumout ,
\Add0~125_sumout ,\Add0~129_sumout ,\Add0~133_sumout ,\Add0~137_sumout ,\Add0~141_sumout ,\Add0~145_sumout ,\Add0~149_sumout ,\Add0~153_sumout ,\Add0~157_sumout ,\Add0~161_sumout ,\Add0~165_sumout ,\Add0~169_sumout ,\Add0~173_sumout ,\Add0~177_sumout ,\Add0~181_sumout ,
\Add0~185_sumout }),
	.enable(stall_reg),
	.register_fifofifo_data019(register_fifofifo_data019),
	.register_fifofifo_data020(register_fifofifo_data020),
	.register_fifofifo_data021(register_fifofifo_data021),
	.register_fifofifo_data022(register_fifofifo_data022),
	.register_fifofifo_data023(register_fifofifo_data023),
	.register_fifofifo_data024(register_fifofifo_data024),
	.register_fifofifo_data025(register_fifofifo_data025),
	.register_fifofifo_data026(register_fifofifo_data026),
	.register_fifofifo_data027(register_fifofifo_data027),
	.register_fifofifo_data028(register_fifofifo_data028),
	.register_fifofifo_data029(register_fifofifo_data029),
	.register_fifofifo_data030(register_fifofifo_data030),
	.register_fifofifo_data031(register_fifofifo_data031),
	.register_fifofifo_data032(register_fifofifo_data032),
	.register_fifofifo_data033(register_fifofifo_data033),
	.register_fifofifo_data034(register_fifofifo_data034),
	.register_fifofifo_data035(register_fifofifo_data035),
	.register_fifofifo_data036(register_fifofifo_data036),
	.register_fifofifo_data037(register_fifofifo_data037),
	.register_fifofifo_data038(register_fifofifo_data038),
	.register_fifofifo_data039(register_fifofifo_data039),
	.register_fifofifo_data040(register_fifofifo_data040),
	.register_fifofifo_data041(register_fifofifo_data041),
	.register_fifofifo_data042(register_fifofifo_data042),
	.register_fifofifo_data043(register_fifofifo_data043),
	.register_fifofifo_data044(register_fifofifo_data044),
	.register_fifofifo_data045(register_fifofifo_data045),
	.register_fifofifo_data046(register_fifofifo_data046),
	.register_fifofifo_data018(register_fifofifo_data018),
	.register_fifofifo_data017(register_fifofifo_data017),
	.register_fifofifo_data016(register_fifofifo_data016),
	.register_fifofifo_data015(register_fifofifo_data015),
	.register_fifofifo_data014(register_fifofifo_data014),
	.register_fifofifo_data013(register_fifofifo_data013),
	.register_fifofifo_data012(register_fifofifo_data012),
	.register_fifofifo_data011(register_fifofifo_data011),
	.register_fifofifo_data010(register_fifofifo_data010),
	.register_fifofifo_data09(register_fifofifo_data09),
	.register_fifofifo_data08(register_fifofifo_data08),
	.register_fifofifo_data07(register_fifofifo_data07),
	.register_fifofifo_data06(register_fifofifo_data06),
	.register_fifofifo_data05(register_fifofifo_data05),
	.register_fifofifo_data04(register_fifofifo_data04),
	.register_fifofifo_data03(register_fifofifo_data03),
	.register_fifofifo_data02(register_fifofifo_data02),
	.register_fifofifo_data01(register_fifofifo_data01),
	.register_fifofifo_data00(register_fifofifo_data00),
	.clk(clk),
	.reset(reset_n));

arriav_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data019),
	.datae(gnd),
	.dataf(!q_b_19),
	.datag(gnd),
	.cin(\Add0~114 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(\Add0~2 ),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~1 .shared_arith = "off";

arriav_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data020),
	.datae(gnd),
	.dataf(!q_b_19),
	.datag(gnd),
	.cin(\Add0~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~5 .shared_arith = "off";

arriav_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data021),
	.datae(gnd),
	.dataf(!q_b_19),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~9 .shared_arith = "off";

arriav_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data022),
	.datae(gnd),
	.dataf(!q_b_19),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~13 .shared_arith = "off";

arriav_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data023),
	.datae(gnd),
	.dataf(!q_b_19),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout());
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~17 .shared_arith = "off";

arriav_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data024),
	.datae(gnd),
	.dataf(!q_b_19),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout());
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~21 .shared_arith = "off";

arriav_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data025),
	.datae(gnd),
	.dataf(!q_b_19),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout());
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~25 .shared_arith = "off";

arriav_lcell_comb \Add0~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data026),
	.datae(gnd),
	.dataf(!q_b_19),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout());
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~29 .shared_arith = "off";

arriav_lcell_comb \Add0~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data027),
	.datae(gnd),
	.dataf(!q_b_19),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~33_sumout ),
	.cout(\Add0~34 ),
	.shareout());
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~33 .shared_arith = "off";

arriav_lcell_comb \Add0~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data028),
	.datae(gnd),
	.dataf(!q_b_19),
	.datag(gnd),
	.cin(\Add0~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~37_sumout ),
	.cout(\Add0~38 ),
	.shareout());
defparam \Add0~37 .extended_lut = "off";
defparam \Add0~37 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~37 .shared_arith = "off";

arriav_lcell_comb \Add0~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data029),
	.datae(gnd),
	.dataf(!q_b_19),
	.datag(gnd),
	.cin(\Add0~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~41_sumout ),
	.cout(\Add0~42 ),
	.shareout());
defparam \Add0~41 .extended_lut = "off";
defparam \Add0~41 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~41 .shared_arith = "off";

arriav_lcell_comb \Add0~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data030),
	.datae(gnd),
	.dataf(!q_b_19),
	.datag(gnd),
	.cin(\Add0~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~45_sumout ),
	.cout(\Add0~46 ),
	.shareout());
defparam \Add0~45 .extended_lut = "off";
defparam \Add0~45 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~45 .shared_arith = "off";

arriav_lcell_comb \Add0~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data031),
	.datae(gnd),
	.dataf(!q_b_19),
	.datag(gnd),
	.cin(\Add0~46 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~49_sumout ),
	.cout(\Add0~50 ),
	.shareout());
defparam \Add0~49 .extended_lut = "off";
defparam \Add0~49 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~49 .shared_arith = "off";

arriav_lcell_comb \Add0~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data032),
	.datae(gnd),
	.dataf(!q_b_19),
	.datag(gnd),
	.cin(\Add0~50 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~53_sumout ),
	.cout(\Add0~54 ),
	.shareout());
defparam \Add0~53 .extended_lut = "off";
defparam \Add0~53 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~53 .shared_arith = "off";

arriav_lcell_comb \Add0~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data033),
	.datae(gnd),
	.dataf(!q_b_19),
	.datag(gnd),
	.cin(\Add0~54 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~57_sumout ),
	.cout(\Add0~58 ),
	.shareout());
defparam \Add0~57 .extended_lut = "off";
defparam \Add0~57 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~57 .shared_arith = "off";

arriav_lcell_comb \Add0~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data034),
	.datae(gnd),
	.dataf(!q_b_19),
	.datag(gnd),
	.cin(\Add0~58 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~61_sumout ),
	.cout(\Add0~62 ),
	.shareout());
defparam \Add0~61 .extended_lut = "off";
defparam \Add0~61 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~61 .shared_arith = "off";

arriav_lcell_comb \Add0~65 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data035),
	.datae(gnd),
	.dataf(!q_b_19),
	.datag(gnd),
	.cin(\Add0~62 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~65_sumout ),
	.cout(\Add0~66 ),
	.shareout());
defparam \Add0~65 .extended_lut = "off";
defparam \Add0~65 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~65 .shared_arith = "off";

arriav_lcell_comb \Add0~69 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data036),
	.datae(gnd),
	.dataf(!q_b_19),
	.datag(gnd),
	.cin(\Add0~66 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~69_sumout ),
	.cout(\Add0~70 ),
	.shareout());
defparam \Add0~69 .extended_lut = "off";
defparam \Add0~69 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~69 .shared_arith = "off";

arriav_lcell_comb \Add0~73 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data037),
	.datae(gnd),
	.dataf(!q_b_19),
	.datag(gnd),
	.cin(\Add0~70 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~73_sumout ),
	.cout(\Add0~74 ),
	.shareout());
defparam \Add0~73 .extended_lut = "off";
defparam \Add0~73 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~73 .shared_arith = "off";

arriav_lcell_comb \Add0~77 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data038),
	.datae(gnd),
	.dataf(!q_b_19),
	.datag(gnd),
	.cin(\Add0~74 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~77_sumout ),
	.cout(\Add0~78 ),
	.shareout());
defparam \Add0~77 .extended_lut = "off";
defparam \Add0~77 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~77 .shared_arith = "off";

arriav_lcell_comb \Add0~81 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data039),
	.datae(gnd),
	.dataf(!q_b_19),
	.datag(gnd),
	.cin(\Add0~78 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~81_sumout ),
	.cout(\Add0~82 ),
	.shareout());
defparam \Add0~81 .extended_lut = "off";
defparam \Add0~81 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~81 .shared_arith = "off";

arriav_lcell_comb \Add0~85 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data040),
	.datae(gnd),
	.dataf(!q_b_19),
	.datag(gnd),
	.cin(\Add0~82 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~85_sumout ),
	.cout(\Add0~86 ),
	.shareout());
defparam \Add0~85 .extended_lut = "off";
defparam \Add0~85 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~85 .shared_arith = "off";

arriav_lcell_comb \Add0~89 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data041),
	.datae(gnd),
	.dataf(!q_b_19),
	.datag(gnd),
	.cin(\Add0~86 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~89_sumout ),
	.cout(\Add0~90 ),
	.shareout());
defparam \Add0~89 .extended_lut = "off";
defparam \Add0~89 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~89 .shared_arith = "off";

arriav_lcell_comb \Add0~93 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data042),
	.datae(gnd),
	.dataf(!q_b_19),
	.datag(gnd),
	.cin(\Add0~90 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~93_sumout ),
	.cout(\Add0~94 ),
	.shareout());
defparam \Add0~93 .extended_lut = "off";
defparam \Add0~93 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~93 .shared_arith = "off";

arriav_lcell_comb \Add0~97 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data043),
	.datae(gnd),
	.dataf(!q_b_19),
	.datag(gnd),
	.cin(\Add0~94 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~97_sumout ),
	.cout(\Add0~98 ),
	.shareout());
defparam \Add0~97 .extended_lut = "off";
defparam \Add0~97 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~97 .shared_arith = "off";

arriav_lcell_comb \Add0~101 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data044),
	.datae(gnd),
	.dataf(!q_b_19),
	.datag(gnd),
	.cin(\Add0~98 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~101_sumout ),
	.cout(\Add0~102 ),
	.shareout());
defparam \Add0~101 .extended_lut = "off";
defparam \Add0~101 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~101 .shared_arith = "off";

arriav_lcell_comb \Add0~105 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data045),
	.datae(gnd),
	.dataf(!q_b_19),
	.datag(gnd),
	.cin(\Add0~102 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~105_sumout ),
	.cout(\Add0~106 ),
	.shareout());
defparam \Add0~105 .extended_lut = "off";
defparam \Add0~105 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~105 .shared_arith = "off";

arriav_lcell_comb \Add0~109 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data046),
	.datae(gnd),
	.dataf(!q_b_19),
	.datag(gnd),
	.cin(\Add0~106 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~109_sumout ),
	.cout(),
	.shareout());
defparam \Add0~109 .extended_lut = "off";
defparam \Add0~109 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~109 .shared_arith = "off";

arriav_lcell_comb \Add0~113 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data018),
	.datae(gnd),
	.dataf(!q_b_18),
	.datag(gnd),
	.cin(\Add0~118 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~113_sumout ),
	.cout(\Add0~114 ),
	.shareout());
defparam \Add0~113 .extended_lut = "off";
defparam \Add0~113 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~113 .shared_arith = "off";

arriav_lcell_comb \Add0~117 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data017),
	.datae(gnd),
	.dataf(!q_b_17),
	.datag(gnd),
	.cin(\Add0~122 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~117_sumout ),
	.cout(\Add0~118 ),
	.shareout());
defparam \Add0~117 .extended_lut = "off";
defparam \Add0~117 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~117 .shared_arith = "off";

arriav_lcell_comb \Add0~121 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data016),
	.datae(gnd),
	.dataf(!q_b_16),
	.datag(gnd),
	.cin(\Add0~126 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~121_sumout ),
	.cout(\Add0~122 ),
	.shareout());
defparam \Add0~121 .extended_lut = "off";
defparam \Add0~121 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~121 .shared_arith = "off";

arriav_lcell_comb \Add0~125 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data015),
	.datae(gnd),
	.dataf(!q_b_15),
	.datag(gnd),
	.cin(\Add0~130 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~125_sumout ),
	.cout(\Add0~126 ),
	.shareout());
defparam \Add0~125 .extended_lut = "off";
defparam \Add0~125 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~125 .shared_arith = "off";

arriav_lcell_comb \Add0~129 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data014),
	.datae(gnd),
	.dataf(!q_b_14),
	.datag(gnd),
	.cin(\Add0~134 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~129_sumout ),
	.cout(\Add0~130 ),
	.shareout());
defparam \Add0~129 .extended_lut = "off";
defparam \Add0~129 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~129 .shared_arith = "off";

arriav_lcell_comb \Add0~133 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data013),
	.datae(gnd),
	.dataf(!q_b_13),
	.datag(gnd),
	.cin(\Add0~138 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~133_sumout ),
	.cout(\Add0~134 ),
	.shareout());
defparam \Add0~133 .extended_lut = "off";
defparam \Add0~133 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~133 .shared_arith = "off";

arriav_lcell_comb \Add0~137 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data012),
	.datae(gnd),
	.dataf(!q_b_12),
	.datag(gnd),
	.cin(\Add0~142 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~137_sumout ),
	.cout(\Add0~138 ),
	.shareout());
defparam \Add0~137 .extended_lut = "off";
defparam \Add0~137 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~137 .shared_arith = "off";

arriav_lcell_comb \Add0~141 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data011),
	.datae(gnd),
	.dataf(!q_b_11),
	.datag(gnd),
	.cin(\Add0~146 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~141_sumout ),
	.cout(\Add0~142 ),
	.shareout());
defparam \Add0~141 .extended_lut = "off";
defparam \Add0~141 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~141 .shared_arith = "off";

arriav_lcell_comb \Add0~145 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data010),
	.datae(gnd),
	.dataf(!q_b_10),
	.datag(gnd),
	.cin(\Add0~150 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~145_sumout ),
	.cout(\Add0~146 ),
	.shareout());
defparam \Add0~145 .extended_lut = "off";
defparam \Add0~145 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~145 .shared_arith = "off";

arriav_lcell_comb \Add0~149 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data09),
	.datae(gnd),
	.dataf(!q_b_9),
	.datag(gnd),
	.cin(\Add0~154 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~149_sumout ),
	.cout(\Add0~150 ),
	.shareout());
defparam \Add0~149 .extended_lut = "off";
defparam \Add0~149 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~149 .shared_arith = "off";

arriav_lcell_comb \Add0~153 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data08),
	.datae(gnd),
	.dataf(!q_b_8),
	.datag(gnd),
	.cin(\Add0~158 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~153_sumout ),
	.cout(\Add0~154 ),
	.shareout());
defparam \Add0~153 .extended_lut = "off";
defparam \Add0~153 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~153 .shared_arith = "off";

arriav_lcell_comb \Add0~157 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data07),
	.datae(gnd),
	.dataf(!q_b_7),
	.datag(gnd),
	.cin(\Add0~162 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~157_sumout ),
	.cout(\Add0~158 ),
	.shareout());
defparam \Add0~157 .extended_lut = "off";
defparam \Add0~157 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~157 .shared_arith = "off";

arriav_lcell_comb \Add0~161 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data06),
	.datae(gnd),
	.dataf(!q_b_6),
	.datag(gnd),
	.cin(\Add0~166 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~161_sumout ),
	.cout(\Add0~162 ),
	.shareout());
defparam \Add0~161 .extended_lut = "off";
defparam \Add0~161 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~161 .shared_arith = "off";

arriav_lcell_comb \Add0~165 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data05),
	.datae(gnd),
	.dataf(!q_b_5),
	.datag(gnd),
	.cin(\Add0~170 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~165_sumout ),
	.cout(\Add0~166 ),
	.shareout());
defparam \Add0~165 .extended_lut = "off";
defparam \Add0~165 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~165 .shared_arith = "off";

arriav_lcell_comb \Add0~169 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data04),
	.datae(gnd),
	.dataf(!q_b_4),
	.datag(gnd),
	.cin(\Add0~174 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~169_sumout ),
	.cout(\Add0~170 ),
	.shareout());
defparam \Add0~169 .extended_lut = "off";
defparam \Add0~169 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~169 .shared_arith = "off";

arriav_lcell_comb \Add0~173 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data03),
	.datae(gnd),
	.dataf(!q_b_3),
	.datag(gnd),
	.cin(\Add0~178 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~173_sumout ),
	.cout(\Add0~174 ),
	.shareout());
defparam \Add0~173 .extended_lut = "off";
defparam \Add0~173 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~173 .shared_arith = "off";

arriav_lcell_comb \Add0~177 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data02),
	.datae(gnd),
	.dataf(!q_b_2),
	.datag(gnd),
	.cin(\Add0~182 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~177_sumout ),
	.cout(\Add0~178 ),
	.shareout());
defparam \Add0~177 .extended_lut = "off";
defparam \Add0~177 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~177 .shared_arith = "off";

arriav_lcell_comb \Add0~181 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data01),
	.datae(gnd),
	.dataf(!q_b_1),
	.datag(gnd),
	.cin(\Add0~186 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~181_sumout ),
	.cout(\Add0~182 ),
	.shareout());
defparam \Add0~181 .extended_lut = "off";
defparam \Add0~181 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~181 .shared_arith = "off";

arriav_lcell_comb \Add0~185 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data00),
	.datae(gnd),
	.dataf(!q_b_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~185_sumout ),
	.cout(\Add0~186 ),
	.shareout());
defparam \Add0~185 .extended_lut = "off";
defparam \Add0~185 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~185 .shared_arith = "off";

endmodule

module cic_auk_dspip_delay_8 (
	datain,
	enable,
	register_fifofifo_data019,
	register_fifofifo_data020,
	register_fifofifo_data021,
	register_fifofifo_data022,
	register_fifofifo_data023,
	register_fifofifo_data024,
	register_fifofifo_data025,
	register_fifofifo_data026,
	register_fifofifo_data027,
	register_fifofifo_data028,
	register_fifofifo_data029,
	register_fifofifo_data030,
	register_fifofifo_data031,
	register_fifofifo_data032,
	register_fifofifo_data033,
	register_fifofifo_data034,
	register_fifofifo_data035,
	register_fifofifo_data036,
	register_fifofifo_data037,
	register_fifofifo_data038,
	register_fifofifo_data039,
	register_fifofifo_data040,
	register_fifofifo_data041,
	register_fifofifo_data042,
	register_fifofifo_data043,
	register_fifofifo_data044,
	register_fifofifo_data045,
	register_fifofifo_data046,
	register_fifofifo_data018,
	register_fifofifo_data017,
	register_fifofifo_data016,
	register_fifofifo_data015,
	register_fifofifo_data014,
	register_fifofifo_data013,
	register_fifofifo_data012,
	register_fifofifo_data011,
	register_fifofifo_data010,
	register_fifofifo_data09,
	register_fifofifo_data08,
	register_fifofifo_data07,
	register_fifofifo_data06,
	register_fifofifo_data05,
	register_fifofifo_data04,
	register_fifofifo_data03,
	register_fifofifo_data02,
	register_fifofifo_data01,
	register_fifofifo_data00,
	clk,
	reset)/* synthesis synthesis_greybox=1 */;
input 	[46:0] datain;
input 	enable;
output 	register_fifofifo_data019;
output 	register_fifofifo_data020;
output 	register_fifofifo_data021;
output 	register_fifofifo_data022;
output 	register_fifofifo_data023;
output 	register_fifofifo_data024;
output 	register_fifofifo_data025;
output 	register_fifofifo_data026;
output 	register_fifofifo_data027;
output 	register_fifofifo_data028;
output 	register_fifofifo_data029;
output 	register_fifofifo_data030;
output 	register_fifofifo_data031;
output 	register_fifofifo_data032;
output 	register_fifofifo_data033;
output 	register_fifofifo_data034;
output 	register_fifofifo_data035;
output 	register_fifofifo_data036;
output 	register_fifofifo_data037;
output 	register_fifofifo_data038;
output 	register_fifofifo_data039;
output 	register_fifofifo_data040;
output 	register_fifofifo_data041;
output 	register_fifofifo_data042;
output 	register_fifofifo_data043;
output 	register_fifofifo_data044;
output 	register_fifofifo_data045;
output 	register_fifofifo_data046;
output 	register_fifofifo_data018;
output 	register_fifofifo_data017;
output 	register_fifofifo_data016;
output 	register_fifofifo_data015;
output 	register_fifofifo_data014;
output 	register_fifofifo_data013;
output 	register_fifofifo_data012;
output 	register_fifofifo_data011;
output 	register_fifofifo_data010;
output 	register_fifofifo_data09;
output 	register_fifofifo_data08;
output 	register_fifofifo_data07;
output 	register_fifofifo_data06;
output 	register_fifofifo_data05;
output 	register_fifofifo_data04;
output 	register_fifofifo_data03;
output 	register_fifofifo_data02;
output 	register_fifofifo_data01;
output 	register_fifofifo_data00;
input 	clk;
input 	reset;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \register_fifo:fifo_data[0][19] (
	.clk(clk),
	.d(datain[19]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data019),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][19] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][19] .power_up = "low";

dffeas \register_fifo:fifo_data[0][20] (
	.clk(clk),
	.d(datain[20]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data020),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][20] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][20] .power_up = "low";

dffeas \register_fifo:fifo_data[0][21] (
	.clk(clk),
	.d(datain[21]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data021),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][21] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][21] .power_up = "low";

dffeas \register_fifo:fifo_data[0][22] (
	.clk(clk),
	.d(datain[22]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data022),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][22] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][22] .power_up = "low";

dffeas \register_fifo:fifo_data[0][23] (
	.clk(clk),
	.d(datain[23]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data023),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][23] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][23] .power_up = "low";

dffeas \register_fifo:fifo_data[0][24] (
	.clk(clk),
	.d(datain[24]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data024),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][24] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][24] .power_up = "low";

dffeas \register_fifo:fifo_data[0][25] (
	.clk(clk),
	.d(datain[25]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data025),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][25] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][25] .power_up = "low";

dffeas \register_fifo:fifo_data[0][26] (
	.clk(clk),
	.d(datain[26]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data026),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][26] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][26] .power_up = "low";

dffeas \register_fifo:fifo_data[0][27] (
	.clk(clk),
	.d(datain[27]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data027),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][27] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][27] .power_up = "low";

dffeas \register_fifo:fifo_data[0][28] (
	.clk(clk),
	.d(datain[28]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data028),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][28] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][28] .power_up = "low";

dffeas \register_fifo:fifo_data[0][29] (
	.clk(clk),
	.d(datain[29]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data029),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][29] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][29] .power_up = "low";

dffeas \register_fifo:fifo_data[0][30] (
	.clk(clk),
	.d(datain[30]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data030),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][30] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][30] .power_up = "low";

dffeas \register_fifo:fifo_data[0][31] (
	.clk(clk),
	.d(datain[31]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data031),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][31] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][31] .power_up = "low";

dffeas \register_fifo:fifo_data[0][32] (
	.clk(clk),
	.d(datain[32]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data032),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][32] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][32] .power_up = "low";

dffeas \register_fifo:fifo_data[0][33] (
	.clk(clk),
	.d(datain[33]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data033),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][33] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][33] .power_up = "low";

dffeas \register_fifo:fifo_data[0][34] (
	.clk(clk),
	.d(datain[34]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data034),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][34] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][34] .power_up = "low";

dffeas \register_fifo:fifo_data[0][35] (
	.clk(clk),
	.d(datain[35]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data035),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][35] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][35] .power_up = "low";

dffeas \register_fifo:fifo_data[0][36] (
	.clk(clk),
	.d(datain[36]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data036),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][36] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][36] .power_up = "low";

dffeas \register_fifo:fifo_data[0][37] (
	.clk(clk),
	.d(datain[37]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data037),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][37] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][37] .power_up = "low";

dffeas \register_fifo:fifo_data[0][38] (
	.clk(clk),
	.d(datain[38]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data038),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][38] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][38] .power_up = "low";

dffeas \register_fifo:fifo_data[0][39] (
	.clk(clk),
	.d(datain[39]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data039),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][39] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][39] .power_up = "low";

dffeas \register_fifo:fifo_data[0][40] (
	.clk(clk),
	.d(datain[40]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data040),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][40] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][40] .power_up = "low";

dffeas \register_fifo:fifo_data[0][41] (
	.clk(clk),
	.d(datain[41]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data041),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][41] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][41] .power_up = "low";

dffeas \register_fifo:fifo_data[0][42] (
	.clk(clk),
	.d(datain[42]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data042),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][42] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][42] .power_up = "low";

dffeas \register_fifo:fifo_data[0][43] (
	.clk(clk),
	.d(datain[43]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data043),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][43] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][43] .power_up = "low";

dffeas \register_fifo:fifo_data[0][44] (
	.clk(clk),
	.d(datain[44]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data044),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][44] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][44] .power_up = "low";

dffeas \register_fifo:fifo_data[0][45] (
	.clk(clk),
	.d(datain[45]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data045),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][45] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][45] .power_up = "low";

dffeas \register_fifo:fifo_data[0][46] (
	.clk(clk),
	.d(datain[46]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data046),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][46] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][46] .power_up = "low";

dffeas \register_fifo:fifo_data[0][18] (
	.clk(clk),
	.d(datain[18]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data018),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][18] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][18] .power_up = "low";

dffeas \register_fifo:fifo_data[0][17] (
	.clk(clk),
	.d(datain[17]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data017),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][17] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][17] .power_up = "low";

dffeas \register_fifo:fifo_data[0][16] (
	.clk(clk),
	.d(datain[16]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data016),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][16] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][16] .power_up = "low";

dffeas \register_fifo:fifo_data[0][15] (
	.clk(clk),
	.d(datain[15]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data015),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][15] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][15] .power_up = "low";

dffeas \register_fifo:fifo_data[0][14] (
	.clk(clk),
	.d(datain[14]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data014),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][14] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][14] .power_up = "low";

dffeas \register_fifo:fifo_data[0][13] (
	.clk(clk),
	.d(datain[13]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data013),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][13] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][13] .power_up = "low";

dffeas \register_fifo:fifo_data[0][12] (
	.clk(clk),
	.d(datain[12]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data012),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][12] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][12] .power_up = "low";

dffeas \register_fifo:fifo_data[0][11] (
	.clk(clk),
	.d(datain[11]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data011),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][11] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][11] .power_up = "low";

dffeas \register_fifo:fifo_data[0][10] (
	.clk(clk),
	.d(datain[10]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data010),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][10] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][10] .power_up = "low";

dffeas \register_fifo:fifo_data[0][9] (
	.clk(clk),
	.d(datain[9]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data09),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][9] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][9] .power_up = "low";

dffeas \register_fifo:fifo_data[0][8] (
	.clk(clk),
	.d(datain[8]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data08),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][8] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][8] .power_up = "low";

dffeas \register_fifo:fifo_data[0][7] (
	.clk(clk),
	.d(datain[7]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data07),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][7] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][7] .power_up = "low";

dffeas \register_fifo:fifo_data[0][6] (
	.clk(clk),
	.d(datain[6]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data06),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][6] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][6] .power_up = "low";

dffeas \register_fifo:fifo_data[0][5] (
	.clk(clk),
	.d(datain[5]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data05),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][5] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][5] .power_up = "low";

dffeas \register_fifo:fifo_data[0][4] (
	.clk(clk),
	.d(datain[4]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data04),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][4] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][4] .power_up = "low";

dffeas \register_fifo:fifo_data[0][3] (
	.clk(clk),
	.d(datain[3]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data03),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][3] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][3] .power_up = "low";

dffeas \register_fifo:fifo_data[0][2] (
	.clk(clk),
	.d(datain[2]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data02),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][2] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][2] .power_up = "low";

dffeas \register_fifo:fifo_data[0][1] (
	.clk(clk),
	.d(datain[1]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data01),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][1] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][1] .power_up = "low";

dffeas \register_fifo:fifo_data[0][0] (
	.clk(clk),
	.d(datain[0]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data00),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][0] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][0] .power_up = "low";

endmodule

module cic_auk_dspip_integrator_1 (
	stall_reg,
	register_fifofifo_data019,
	register_fifofifo_data020,
	register_fifofifo_data021,
	register_fifofifo_data022,
	register_fifofifo_data023,
	register_fifofifo_data024,
	register_fifofifo_data025,
	register_fifofifo_data026,
	register_fifofifo_data027,
	register_fifofifo_data028,
	register_fifofifo_data029,
	register_fifofifo_data030,
	register_fifofifo_data031,
	register_fifofifo_data032,
	register_fifofifo_data033,
	register_fifofifo_data034,
	register_fifofifo_data035,
	register_fifofifo_data036,
	register_fifofifo_data037,
	register_fifofifo_data038,
	register_fifofifo_data039,
	register_fifofifo_data040,
	register_fifofifo_data041,
	register_fifofifo_data042,
	register_fifofifo_data043,
	register_fifofifo_data044,
	register_fifofifo_data045,
	register_fifofifo_data046,
	register_fifofifo_data018,
	register_fifofifo_data0191,
	register_fifofifo_data017,
	register_fifofifo_data0201,
	register_fifofifo_data0211,
	register_fifofifo_data0221,
	register_fifofifo_data0231,
	register_fifofifo_data0241,
	register_fifofifo_data0251,
	register_fifofifo_data0261,
	register_fifofifo_data0271,
	register_fifofifo_data0281,
	register_fifofifo_data0291,
	register_fifofifo_data0301,
	register_fifofifo_data0311,
	register_fifofifo_data0321,
	register_fifofifo_data0331,
	register_fifofifo_data0341,
	register_fifofifo_data0351,
	register_fifofifo_data0361,
	register_fifofifo_data0371,
	register_fifofifo_data0381,
	register_fifofifo_data0391,
	register_fifofifo_data0401,
	register_fifofifo_data0411,
	register_fifofifo_data0421,
	register_fifofifo_data0431,
	register_fifofifo_data0441,
	register_fifofifo_data0451,
	register_fifofifo_data0461,
	register_fifofifo_data0181,
	register_fifofifo_data016,
	register_fifofifo_data0171,
	register_fifofifo_data015,
	register_fifofifo_data0161,
	register_fifofifo_data014,
	register_fifofifo_data0151,
	register_fifofifo_data013,
	register_fifofifo_data0141,
	register_fifofifo_data012,
	register_fifofifo_data0131,
	register_fifofifo_data011,
	register_fifofifo_data0121,
	register_fifofifo_data010,
	register_fifofifo_data0111,
	register_fifofifo_data09,
	register_fifofifo_data0101,
	register_fifofifo_data08,
	register_fifofifo_data091,
	register_fifofifo_data07,
	register_fifofifo_data081,
	register_fifofifo_data06,
	register_fifofifo_data071,
	register_fifofifo_data05,
	register_fifofifo_data061,
	register_fifofifo_data04,
	register_fifofifo_data051,
	register_fifofifo_data03,
	register_fifofifo_data047,
	register_fifofifo_data02,
	register_fifofifo_data0310,
	register_fifofifo_data01,
	register_fifofifo_data0210,
	register_fifofifo_data00,
	register_fifofifo_data0110,
	register_fifofifo_data001,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	stall_reg;
output 	register_fifofifo_data019;
output 	register_fifofifo_data020;
output 	register_fifofifo_data021;
output 	register_fifofifo_data022;
output 	register_fifofifo_data023;
output 	register_fifofifo_data024;
output 	register_fifofifo_data025;
output 	register_fifofifo_data026;
output 	register_fifofifo_data027;
output 	register_fifofifo_data028;
output 	register_fifofifo_data029;
output 	register_fifofifo_data030;
output 	register_fifofifo_data031;
output 	register_fifofifo_data032;
output 	register_fifofifo_data033;
output 	register_fifofifo_data034;
output 	register_fifofifo_data035;
output 	register_fifofifo_data036;
output 	register_fifofifo_data037;
output 	register_fifofifo_data038;
output 	register_fifofifo_data039;
output 	register_fifofifo_data040;
output 	register_fifofifo_data041;
output 	register_fifofifo_data042;
output 	register_fifofifo_data043;
output 	register_fifofifo_data044;
output 	register_fifofifo_data045;
output 	register_fifofifo_data046;
output 	register_fifofifo_data018;
input 	register_fifofifo_data0191;
output 	register_fifofifo_data017;
input 	register_fifofifo_data0201;
input 	register_fifofifo_data0211;
input 	register_fifofifo_data0221;
input 	register_fifofifo_data0231;
input 	register_fifofifo_data0241;
input 	register_fifofifo_data0251;
input 	register_fifofifo_data0261;
input 	register_fifofifo_data0271;
input 	register_fifofifo_data0281;
input 	register_fifofifo_data0291;
input 	register_fifofifo_data0301;
input 	register_fifofifo_data0311;
input 	register_fifofifo_data0321;
input 	register_fifofifo_data0331;
input 	register_fifofifo_data0341;
input 	register_fifofifo_data0351;
input 	register_fifofifo_data0361;
input 	register_fifofifo_data0371;
input 	register_fifofifo_data0381;
input 	register_fifofifo_data0391;
input 	register_fifofifo_data0401;
input 	register_fifofifo_data0411;
input 	register_fifofifo_data0421;
input 	register_fifofifo_data0431;
input 	register_fifofifo_data0441;
input 	register_fifofifo_data0451;
input 	register_fifofifo_data0461;
input 	register_fifofifo_data0181;
output 	register_fifofifo_data016;
input 	register_fifofifo_data0171;
output 	register_fifofifo_data015;
input 	register_fifofifo_data0161;
output 	register_fifofifo_data014;
input 	register_fifofifo_data0151;
output 	register_fifofifo_data013;
input 	register_fifofifo_data0141;
output 	register_fifofifo_data012;
input 	register_fifofifo_data0131;
output 	register_fifofifo_data011;
input 	register_fifofifo_data0121;
output 	register_fifofifo_data010;
input 	register_fifofifo_data0111;
output 	register_fifofifo_data09;
input 	register_fifofifo_data0101;
output 	register_fifofifo_data08;
input 	register_fifofifo_data091;
output 	register_fifofifo_data07;
input 	register_fifofifo_data081;
output 	register_fifofifo_data06;
input 	register_fifofifo_data071;
output 	register_fifofifo_data05;
input 	register_fifofifo_data061;
output 	register_fifofifo_data04;
input 	register_fifofifo_data051;
output 	register_fifofifo_data03;
input 	register_fifofifo_data047;
output 	register_fifofifo_data02;
input 	register_fifofifo_data0310;
output 	register_fifofifo_data01;
input 	register_fifofifo_data0210;
output 	register_fifofifo_data00;
input 	register_fifofifo_data0110;
input 	register_fifofifo_data001;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Add0~1_sumout ;
wire \Add0~2 ;
wire \Add0~5_sumout ;
wire \Add0~6 ;
wire \Add0~9_sumout ;
wire \Add0~10 ;
wire \Add0~13_sumout ;
wire \Add0~14 ;
wire \Add0~17_sumout ;
wire \Add0~18 ;
wire \Add0~21_sumout ;
wire \Add0~22 ;
wire \Add0~25_sumout ;
wire \Add0~26 ;
wire \Add0~29_sumout ;
wire \Add0~30 ;
wire \Add0~33_sumout ;
wire \Add0~34 ;
wire \Add0~37_sumout ;
wire \Add0~38 ;
wire \Add0~41_sumout ;
wire \Add0~42 ;
wire \Add0~45_sumout ;
wire \Add0~46 ;
wire \Add0~49_sumout ;
wire \Add0~50 ;
wire \Add0~53_sumout ;
wire \Add0~54 ;
wire \Add0~57_sumout ;
wire \Add0~58 ;
wire \Add0~61_sumout ;
wire \Add0~62 ;
wire \Add0~65_sumout ;
wire \Add0~66 ;
wire \Add0~69_sumout ;
wire \Add0~70 ;
wire \Add0~73_sumout ;
wire \Add0~74 ;
wire \Add0~77_sumout ;
wire \Add0~78 ;
wire \Add0~81_sumout ;
wire \Add0~82 ;
wire \Add0~85_sumout ;
wire \Add0~86 ;
wire \Add0~89_sumout ;
wire \Add0~90 ;
wire \Add0~93_sumout ;
wire \Add0~94 ;
wire \Add0~97_sumout ;
wire \Add0~98 ;
wire \Add0~101_sumout ;
wire \Add0~102 ;
wire \Add0~105_sumout ;
wire \Add0~106 ;
wire \Add0~109_sumout ;
wire \Add0~113_sumout ;
wire \Add0~114 ;
wire \Add0~117_sumout ;
wire \Add0~118 ;
wire \Add0~121_sumout ;
wire \Add0~122 ;
wire \Add0~125_sumout ;
wire \Add0~126 ;
wire \Add0~129_sumout ;
wire \Add0~130 ;
wire \Add0~133_sumout ;
wire \Add0~134 ;
wire \Add0~137_sumout ;
wire \Add0~138 ;
wire \Add0~141_sumout ;
wire \Add0~142 ;
wire \Add0~145_sumout ;
wire \Add0~146 ;
wire \Add0~149_sumout ;
wire \Add0~150 ;
wire \Add0~153_sumout ;
wire \Add0~154 ;
wire \Add0~157_sumout ;
wire \Add0~158 ;
wire \Add0~161_sumout ;
wire \Add0~162 ;
wire \Add0~165_sumout ;
wire \Add0~166 ;
wire \Add0~169_sumout ;
wire \Add0~170 ;
wire \Add0~173_sumout ;
wire \Add0~174 ;
wire \Add0~177_sumout ;
wire \Add0~178 ;
wire \Add0~181_sumout ;
wire \Add0~182 ;
wire \Add0~185_sumout ;
wire \Add0~186 ;


cic_auk_dspip_delay_9 \glogic:integrator_pipeline_0_generate:u1 (
	.datain({\Add0~109_sumout ,\Add0~105_sumout ,\Add0~101_sumout ,\Add0~97_sumout ,\Add0~93_sumout ,\Add0~89_sumout ,\Add0~85_sumout ,\Add0~81_sumout ,\Add0~77_sumout ,\Add0~73_sumout ,\Add0~69_sumout ,\Add0~65_sumout ,\Add0~61_sumout ,\Add0~57_sumout ,\Add0~53_sumout ,
\Add0~49_sumout ,\Add0~45_sumout ,\Add0~41_sumout ,\Add0~37_sumout ,\Add0~33_sumout ,\Add0~29_sumout ,\Add0~25_sumout ,\Add0~21_sumout ,\Add0~17_sumout ,\Add0~13_sumout ,\Add0~9_sumout ,\Add0~5_sumout ,\Add0~1_sumout ,\Add0~113_sumout ,\Add0~117_sumout ,\Add0~121_sumout ,
\Add0~125_sumout ,\Add0~129_sumout ,\Add0~133_sumout ,\Add0~137_sumout ,\Add0~141_sumout ,\Add0~145_sumout ,\Add0~149_sumout ,\Add0~153_sumout ,\Add0~157_sumout ,\Add0~161_sumout ,\Add0~165_sumout ,\Add0~169_sumout ,\Add0~173_sumout ,\Add0~177_sumout ,\Add0~181_sumout ,
\Add0~185_sumout }),
	.enable(stall_reg),
	.register_fifofifo_data019(register_fifofifo_data019),
	.register_fifofifo_data020(register_fifofifo_data020),
	.register_fifofifo_data021(register_fifofifo_data021),
	.register_fifofifo_data022(register_fifofifo_data022),
	.register_fifofifo_data023(register_fifofifo_data023),
	.register_fifofifo_data024(register_fifofifo_data024),
	.register_fifofifo_data025(register_fifofifo_data025),
	.register_fifofifo_data026(register_fifofifo_data026),
	.register_fifofifo_data027(register_fifofifo_data027),
	.register_fifofifo_data028(register_fifofifo_data028),
	.register_fifofifo_data029(register_fifofifo_data029),
	.register_fifofifo_data030(register_fifofifo_data030),
	.register_fifofifo_data031(register_fifofifo_data031),
	.register_fifofifo_data032(register_fifofifo_data032),
	.register_fifofifo_data033(register_fifofifo_data033),
	.register_fifofifo_data034(register_fifofifo_data034),
	.register_fifofifo_data035(register_fifofifo_data035),
	.register_fifofifo_data036(register_fifofifo_data036),
	.register_fifofifo_data037(register_fifofifo_data037),
	.register_fifofifo_data038(register_fifofifo_data038),
	.register_fifofifo_data039(register_fifofifo_data039),
	.register_fifofifo_data040(register_fifofifo_data040),
	.register_fifofifo_data041(register_fifofifo_data041),
	.register_fifofifo_data042(register_fifofifo_data042),
	.register_fifofifo_data043(register_fifofifo_data043),
	.register_fifofifo_data044(register_fifofifo_data044),
	.register_fifofifo_data045(register_fifofifo_data045),
	.register_fifofifo_data046(register_fifofifo_data046),
	.register_fifofifo_data018(register_fifofifo_data018),
	.register_fifofifo_data017(register_fifofifo_data017),
	.register_fifofifo_data016(register_fifofifo_data016),
	.register_fifofifo_data015(register_fifofifo_data015),
	.register_fifofifo_data014(register_fifofifo_data014),
	.register_fifofifo_data013(register_fifofifo_data013),
	.register_fifofifo_data012(register_fifofifo_data012),
	.register_fifofifo_data011(register_fifofifo_data011),
	.register_fifofifo_data010(register_fifofifo_data010),
	.register_fifofifo_data09(register_fifofifo_data09),
	.register_fifofifo_data08(register_fifofifo_data08),
	.register_fifofifo_data07(register_fifofifo_data07),
	.register_fifofifo_data06(register_fifofifo_data06),
	.register_fifofifo_data05(register_fifofifo_data05),
	.register_fifofifo_data04(register_fifofifo_data04),
	.register_fifofifo_data03(register_fifofifo_data03),
	.register_fifofifo_data02(register_fifofifo_data02),
	.register_fifofifo_data01(register_fifofifo_data01),
	.register_fifofifo_data00(register_fifofifo_data00),
	.clk(clk),
	.reset(reset_n));

arriav_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data019),
	.datae(gnd),
	.dataf(!register_fifofifo_data0191),
	.datag(gnd),
	.cin(\Add0~114 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(\Add0~2 ),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~1 .shared_arith = "off";

arriav_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data020),
	.datae(gnd),
	.dataf(!register_fifofifo_data0201),
	.datag(gnd),
	.cin(\Add0~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~5 .shared_arith = "off";

arriav_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data021),
	.datae(gnd),
	.dataf(!register_fifofifo_data0211),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~9 .shared_arith = "off";

arriav_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data022),
	.datae(gnd),
	.dataf(!register_fifofifo_data0221),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~13 .shared_arith = "off";

arriav_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data023),
	.datae(gnd),
	.dataf(!register_fifofifo_data0231),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout());
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~17 .shared_arith = "off";

arriav_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data024),
	.datae(gnd),
	.dataf(!register_fifofifo_data0241),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout());
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~21 .shared_arith = "off";

arriav_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data025),
	.datae(gnd),
	.dataf(!register_fifofifo_data0251),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout());
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~25 .shared_arith = "off";

arriav_lcell_comb \Add0~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data026),
	.datae(gnd),
	.dataf(!register_fifofifo_data0261),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout());
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~29 .shared_arith = "off";

arriav_lcell_comb \Add0~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data027),
	.datae(gnd),
	.dataf(!register_fifofifo_data0271),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~33_sumout ),
	.cout(\Add0~34 ),
	.shareout());
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~33 .shared_arith = "off";

arriav_lcell_comb \Add0~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data028),
	.datae(gnd),
	.dataf(!register_fifofifo_data0281),
	.datag(gnd),
	.cin(\Add0~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~37_sumout ),
	.cout(\Add0~38 ),
	.shareout());
defparam \Add0~37 .extended_lut = "off";
defparam \Add0~37 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~37 .shared_arith = "off";

arriav_lcell_comb \Add0~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data029),
	.datae(gnd),
	.dataf(!register_fifofifo_data0291),
	.datag(gnd),
	.cin(\Add0~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~41_sumout ),
	.cout(\Add0~42 ),
	.shareout());
defparam \Add0~41 .extended_lut = "off";
defparam \Add0~41 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~41 .shared_arith = "off";

arriav_lcell_comb \Add0~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data030),
	.datae(gnd),
	.dataf(!register_fifofifo_data0301),
	.datag(gnd),
	.cin(\Add0~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~45_sumout ),
	.cout(\Add0~46 ),
	.shareout());
defparam \Add0~45 .extended_lut = "off";
defparam \Add0~45 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~45 .shared_arith = "off";

arriav_lcell_comb \Add0~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data031),
	.datae(gnd),
	.dataf(!register_fifofifo_data0311),
	.datag(gnd),
	.cin(\Add0~46 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~49_sumout ),
	.cout(\Add0~50 ),
	.shareout());
defparam \Add0~49 .extended_lut = "off";
defparam \Add0~49 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~49 .shared_arith = "off";

arriav_lcell_comb \Add0~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data032),
	.datae(gnd),
	.dataf(!register_fifofifo_data0321),
	.datag(gnd),
	.cin(\Add0~50 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~53_sumout ),
	.cout(\Add0~54 ),
	.shareout());
defparam \Add0~53 .extended_lut = "off";
defparam \Add0~53 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~53 .shared_arith = "off";

arriav_lcell_comb \Add0~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data033),
	.datae(gnd),
	.dataf(!register_fifofifo_data0331),
	.datag(gnd),
	.cin(\Add0~54 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~57_sumout ),
	.cout(\Add0~58 ),
	.shareout());
defparam \Add0~57 .extended_lut = "off";
defparam \Add0~57 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~57 .shared_arith = "off";

arriav_lcell_comb \Add0~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data034),
	.datae(gnd),
	.dataf(!register_fifofifo_data0341),
	.datag(gnd),
	.cin(\Add0~58 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~61_sumout ),
	.cout(\Add0~62 ),
	.shareout());
defparam \Add0~61 .extended_lut = "off";
defparam \Add0~61 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~61 .shared_arith = "off";

arriav_lcell_comb \Add0~65 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data035),
	.datae(gnd),
	.dataf(!register_fifofifo_data0351),
	.datag(gnd),
	.cin(\Add0~62 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~65_sumout ),
	.cout(\Add0~66 ),
	.shareout());
defparam \Add0~65 .extended_lut = "off";
defparam \Add0~65 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~65 .shared_arith = "off";

arriav_lcell_comb \Add0~69 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data036),
	.datae(gnd),
	.dataf(!register_fifofifo_data0361),
	.datag(gnd),
	.cin(\Add0~66 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~69_sumout ),
	.cout(\Add0~70 ),
	.shareout());
defparam \Add0~69 .extended_lut = "off";
defparam \Add0~69 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~69 .shared_arith = "off";

arriav_lcell_comb \Add0~73 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data037),
	.datae(gnd),
	.dataf(!register_fifofifo_data0371),
	.datag(gnd),
	.cin(\Add0~70 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~73_sumout ),
	.cout(\Add0~74 ),
	.shareout());
defparam \Add0~73 .extended_lut = "off";
defparam \Add0~73 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~73 .shared_arith = "off";

arriav_lcell_comb \Add0~77 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data038),
	.datae(gnd),
	.dataf(!register_fifofifo_data0381),
	.datag(gnd),
	.cin(\Add0~74 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~77_sumout ),
	.cout(\Add0~78 ),
	.shareout());
defparam \Add0~77 .extended_lut = "off";
defparam \Add0~77 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~77 .shared_arith = "off";

arriav_lcell_comb \Add0~81 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data039),
	.datae(gnd),
	.dataf(!register_fifofifo_data0391),
	.datag(gnd),
	.cin(\Add0~78 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~81_sumout ),
	.cout(\Add0~82 ),
	.shareout());
defparam \Add0~81 .extended_lut = "off";
defparam \Add0~81 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~81 .shared_arith = "off";

arriav_lcell_comb \Add0~85 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data040),
	.datae(gnd),
	.dataf(!register_fifofifo_data0401),
	.datag(gnd),
	.cin(\Add0~82 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~85_sumout ),
	.cout(\Add0~86 ),
	.shareout());
defparam \Add0~85 .extended_lut = "off";
defparam \Add0~85 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~85 .shared_arith = "off";

arriav_lcell_comb \Add0~89 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data041),
	.datae(gnd),
	.dataf(!register_fifofifo_data0411),
	.datag(gnd),
	.cin(\Add0~86 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~89_sumout ),
	.cout(\Add0~90 ),
	.shareout());
defparam \Add0~89 .extended_lut = "off";
defparam \Add0~89 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~89 .shared_arith = "off";

arriav_lcell_comb \Add0~93 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data042),
	.datae(gnd),
	.dataf(!register_fifofifo_data0421),
	.datag(gnd),
	.cin(\Add0~90 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~93_sumout ),
	.cout(\Add0~94 ),
	.shareout());
defparam \Add0~93 .extended_lut = "off";
defparam \Add0~93 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~93 .shared_arith = "off";

arriav_lcell_comb \Add0~97 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data043),
	.datae(gnd),
	.dataf(!register_fifofifo_data0431),
	.datag(gnd),
	.cin(\Add0~94 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~97_sumout ),
	.cout(\Add0~98 ),
	.shareout());
defparam \Add0~97 .extended_lut = "off";
defparam \Add0~97 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~97 .shared_arith = "off";

arriav_lcell_comb \Add0~101 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data044),
	.datae(gnd),
	.dataf(!register_fifofifo_data0441),
	.datag(gnd),
	.cin(\Add0~98 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~101_sumout ),
	.cout(\Add0~102 ),
	.shareout());
defparam \Add0~101 .extended_lut = "off";
defparam \Add0~101 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~101 .shared_arith = "off";

arriav_lcell_comb \Add0~105 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data045),
	.datae(gnd),
	.dataf(!register_fifofifo_data0451),
	.datag(gnd),
	.cin(\Add0~102 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~105_sumout ),
	.cout(\Add0~106 ),
	.shareout());
defparam \Add0~105 .extended_lut = "off";
defparam \Add0~105 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~105 .shared_arith = "off";

arriav_lcell_comb \Add0~109 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data046),
	.datae(gnd),
	.dataf(!register_fifofifo_data0461),
	.datag(gnd),
	.cin(\Add0~106 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~109_sumout ),
	.cout(),
	.shareout());
defparam \Add0~109 .extended_lut = "off";
defparam \Add0~109 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~109 .shared_arith = "off";

arriav_lcell_comb \Add0~113 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data018),
	.datae(gnd),
	.dataf(!register_fifofifo_data0181),
	.datag(gnd),
	.cin(\Add0~118 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~113_sumout ),
	.cout(\Add0~114 ),
	.shareout());
defparam \Add0~113 .extended_lut = "off";
defparam \Add0~113 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~113 .shared_arith = "off";

arriav_lcell_comb \Add0~117 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data017),
	.datae(gnd),
	.dataf(!register_fifofifo_data0171),
	.datag(gnd),
	.cin(\Add0~122 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~117_sumout ),
	.cout(\Add0~118 ),
	.shareout());
defparam \Add0~117 .extended_lut = "off";
defparam \Add0~117 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~117 .shared_arith = "off";

arriav_lcell_comb \Add0~121 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data016),
	.datae(gnd),
	.dataf(!register_fifofifo_data0161),
	.datag(gnd),
	.cin(\Add0~126 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~121_sumout ),
	.cout(\Add0~122 ),
	.shareout());
defparam \Add0~121 .extended_lut = "off";
defparam \Add0~121 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~121 .shared_arith = "off";

arriav_lcell_comb \Add0~125 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data015),
	.datae(gnd),
	.dataf(!register_fifofifo_data0151),
	.datag(gnd),
	.cin(\Add0~130 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~125_sumout ),
	.cout(\Add0~126 ),
	.shareout());
defparam \Add0~125 .extended_lut = "off";
defparam \Add0~125 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~125 .shared_arith = "off";

arriav_lcell_comb \Add0~129 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data014),
	.datae(gnd),
	.dataf(!register_fifofifo_data0141),
	.datag(gnd),
	.cin(\Add0~134 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~129_sumout ),
	.cout(\Add0~130 ),
	.shareout());
defparam \Add0~129 .extended_lut = "off";
defparam \Add0~129 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~129 .shared_arith = "off";

arriav_lcell_comb \Add0~133 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data013),
	.datae(gnd),
	.dataf(!register_fifofifo_data0131),
	.datag(gnd),
	.cin(\Add0~138 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~133_sumout ),
	.cout(\Add0~134 ),
	.shareout());
defparam \Add0~133 .extended_lut = "off";
defparam \Add0~133 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~133 .shared_arith = "off";

arriav_lcell_comb \Add0~137 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data012),
	.datae(gnd),
	.dataf(!register_fifofifo_data0121),
	.datag(gnd),
	.cin(\Add0~142 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~137_sumout ),
	.cout(\Add0~138 ),
	.shareout());
defparam \Add0~137 .extended_lut = "off";
defparam \Add0~137 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~137 .shared_arith = "off";

arriav_lcell_comb \Add0~141 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data011),
	.datae(gnd),
	.dataf(!register_fifofifo_data0111),
	.datag(gnd),
	.cin(\Add0~146 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~141_sumout ),
	.cout(\Add0~142 ),
	.shareout());
defparam \Add0~141 .extended_lut = "off";
defparam \Add0~141 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~141 .shared_arith = "off";

arriav_lcell_comb \Add0~145 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data010),
	.datae(gnd),
	.dataf(!register_fifofifo_data0101),
	.datag(gnd),
	.cin(\Add0~150 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~145_sumout ),
	.cout(\Add0~146 ),
	.shareout());
defparam \Add0~145 .extended_lut = "off";
defparam \Add0~145 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~145 .shared_arith = "off";

arriav_lcell_comb \Add0~149 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data09),
	.datae(gnd),
	.dataf(!register_fifofifo_data091),
	.datag(gnd),
	.cin(\Add0~154 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~149_sumout ),
	.cout(\Add0~150 ),
	.shareout());
defparam \Add0~149 .extended_lut = "off";
defparam \Add0~149 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~149 .shared_arith = "off";

arriav_lcell_comb \Add0~153 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data08),
	.datae(gnd),
	.dataf(!register_fifofifo_data081),
	.datag(gnd),
	.cin(\Add0~158 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~153_sumout ),
	.cout(\Add0~154 ),
	.shareout());
defparam \Add0~153 .extended_lut = "off";
defparam \Add0~153 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~153 .shared_arith = "off";

arriav_lcell_comb \Add0~157 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data07),
	.datae(gnd),
	.dataf(!register_fifofifo_data071),
	.datag(gnd),
	.cin(\Add0~162 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~157_sumout ),
	.cout(\Add0~158 ),
	.shareout());
defparam \Add0~157 .extended_lut = "off";
defparam \Add0~157 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~157 .shared_arith = "off";

arriav_lcell_comb \Add0~161 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data06),
	.datae(gnd),
	.dataf(!register_fifofifo_data061),
	.datag(gnd),
	.cin(\Add0~166 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~161_sumout ),
	.cout(\Add0~162 ),
	.shareout());
defparam \Add0~161 .extended_lut = "off";
defparam \Add0~161 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~161 .shared_arith = "off";

arriav_lcell_comb \Add0~165 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data05),
	.datae(gnd),
	.dataf(!register_fifofifo_data051),
	.datag(gnd),
	.cin(\Add0~170 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~165_sumout ),
	.cout(\Add0~166 ),
	.shareout());
defparam \Add0~165 .extended_lut = "off";
defparam \Add0~165 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~165 .shared_arith = "off";

arriav_lcell_comb \Add0~169 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data04),
	.datae(gnd),
	.dataf(!register_fifofifo_data047),
	.datag(gnd),
	.cin(\Add0~174 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~169_sumout ),
	.cout(\Add0~170 ),
	.shareout());
defparam \Add0~169 .extended_lut = "off";
defparam \Add0~169 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~169 .shared_arith = "off";

arriav_lcell_comb \Add0~173 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data03),
	.datae(gnd),
	.dataf(!register_fifofifo_data0310),
	.datag(gnd),
	.cin(\Add0~178 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~173_sumout ),
	.cout(\Add0~174 ),
	.shareout());
defparam \Add0~173 .extended_lut = "off";
defparam \Add0~173 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~173 .shared_arith = "off";

arriav_lcell_comb \Add0~177 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data02),
	.datae(gnd),
	.dataf(!register_fifofifo_data0210),
	.datag(gnd),
	.cin(\Add0~182 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~177_sumout ),
	.cout(\Add0~178 ),
	.shareout());
defparam \Add0~177 .extended_lut = "off";
defparam \Add0~177 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~177 .shared_arith = "off";

arriav_lcell_comb \Add0~181 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data01),
	.datae(gnd),
	.dataf(!register_fifofifo_data0110),
	.datag(gnd),
	.cin(\Add0~186 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~181_sumout ),
	.cout(\Add0~182 ),
	.shareout());
defparam \Add0~181 .extended_lut = "off";
defparam \Add0~181 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~181 .shared_arith = "off";

arriav_lcell_comb \Add0~185 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data00),
	.datae(gnd),
	.dataf(!register_fifofifo_data001),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~185_sumout ),
	.cout(\Add0~186 ),
	.shareout());
defparam \Add0~185 .extended_lut = "off";
defparam \Add0~185 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~185 .shared_arith = "off";

endmodule

module cic_auk_dspip_delay_9 (
	datain,
	enable,
	register_fifofifo_data019,
	register_fifofifo_data020,
	register_fifofifo_data021,
	register_fifofifo_data022,
	register_fifofifo_data023,
	register_fifofifo_data024,
	register_fifofifo_data025,
	register_fifofifo_data026,
	register_fifofifo_data027,
	register_fifofifo_data028,
	register_fifofifo_data029,
	register_fifofifo_data030,
	register_fifofifo_data031,
	register_fifofifo_data032,
	register_fifofifo_data033,
	register_fifofifo_data034,
	register_fifofifo_data035,
	register_fifofifo_data036,
	register_fifofifo_data037,
	register_fifofifo_data038,
	register_fifofifo_data039,
	register_fifofifo_data040,
	register_fifofifo_data041,
	register_fifofifo_data042,
	register_fifofifo_data043,
	register_fifofifo_data044,
	register_fifofifo_data045,
	register_fifofifo_data046,
	register_fifofifo_data018,
	register_fifofifo_data017,
	register_fifofifo_data016,
	register_fifofifo_data015,
	register_fifofifo_data014,
	register_fifofifo_data013,
	register_fifofifo_data012,
	register_fifofifo_data011,
	register_fifofifo_data010,
	register_fifofifo_data09,
	register_fifofifo_data08,
	register_fifofifo_data07,
	register_fifofifo_data06,
	register_fifofifo_data05,
	register_fifofifo_data04,
	register_fifofifo_data03,
	register_fifofifo_data02,
	register_fifofifo_data01,
	register_fifofifo_data00,
	clk,
	reset)/* synthesis synthesis_greybox=1 */;
input 	[46:0] datain;
input 	enable;
output 	register_fifofifo_data019;
output 	register_fifofifo_data020;
output 	register_fifofifo_data021;
output 	register_fifofifo_data022;
output 	register_fifofifo_data023;
output 	register_fifofifo_data024;
output 	register_fifofifo_data025;
output 	register_fifofifo_data026;
output 	register_fifofifo_data027;
output 	register_fifofifo_data028;
output 	register_fifofifo_data029;
output 	register_fifofifo_data030;
output 	register_fifofifo_data031;
output 	register_fifofifo_data032;
output 	register_fifofifo_data033;
output 	register_fifofifo_data034;
output 	register_fifofifo_data035;
output 	register_fifofifo_data036;
output 	register_fifofifo_data037;
output 	register_fifofifo_data038;
output 	register_fifofifo_data039;
output 	register_fifofifo_data040;
output 	register_fifofifo_data041;
output 	register_fifofifo_data042;
output 	register_fifofifo_data043;
output 	register_fifofifo_data044;
output 	register_fifofifo_data045;
output 	register_fifofifo_data046;
output 	register_fifofifo_data018;
output 	register_fifofifo_data017;
output 	register_fifofifo_data016;
output 	register_fifofifo_data015;
output 	register_fifofifo_data014;
output 	register_fifofifo_data013;
output 	register_fifofifo_data012;
output 	register_fifofifo_data011;
output 	register_fifofifo_data010;
output 	register_fifofifo_data09;
output 	register_fifofifo_data08;
output 	register_fifofifo_data07;
output 	register_fifofifo_data06;
output 	register_fifofifo_data05;
output 	register_fifofifo_data04;
output 	register_fifofifo_data03;
output 	register_fifofifo_data02;
output 	register_fifofifo_data01;
output 	register_fifofifo_data00;
input 	clk;
input 	reset;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \register_fifo:fifo_data[0][19] (
	.clk(clk),
	.d(datain[19]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data019),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][19] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][19] .power_up = "low";

dffeas \register_fifo:fifo_data[0][20] (
	.clk(clk),
	.d(datain[20]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data020),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][20] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][20] .power_up = "low";

dffeas \register_fifo:fifo_data[0][21] (
	.clk(clk),
	.d(datain[21]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data021),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][21] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][21] .power_up = "low";

dffeas \register_fifo:fifo_data[0][22] (
	.clk(clk),
	.d(datain[22]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data022),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][22] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][22] .power_up = "low";

dffeas \register_fifo:fifo_data[0][23] (
	.clk(clk),
	.d(datain[23]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data023),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][23] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][23] .power_up = "low";

dffeas \register_fifo:fifo_data[0][24] (
	.clk(clk),
	.d(datain[24]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data024),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][24] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][24] .power_up = "low";

dffeas \register_fifo:fifo_data[0][25] (
	.clk(clk),
	.d(datain[25]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data025),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][25] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][25] .power_up = "low";

dffeas \register_fifo:fifo_data[0][26] (
	.clk(clk),
	.d(datain[26]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data026),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][26] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][26] .power_up = "low";

dffeas \register_fifo:fifo_data[0][27] (
	.clk(clk),
	.d(datain[27]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data027),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][27] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][27] .power_up = "low";

dffeas \register_fifo:fifo_data[0][28] (
	.clk(clk),
	.d(datain[28]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data028),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][28] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][28] .power_up = "low";

dffeas \register_fifo:fifo_data[0][29] (
	.clk(clk),
	.d(datain[29]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data029),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][29] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][29] .power_up = "low";

dffeas \register_fifo:fifo_data[0][30] (
	.clk(clk),
	.d(datain[30]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data030),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][30] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][30] .power_up = "low";

dffeas \register_fifo:fifo_data[0][31] (
	.clk(clk),
	.d(datain[31]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data031),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][31] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][31] .power_up = "low";

dffeas \register_fifo:fifo_data[0][32] (
	.clk(clk),
	.d(datain[32]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data032),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][32] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][32] .power_up = "low";

dffeas \register_fifo:fifo_data[0][33] (
	.clk(clk),
	.d(datain[33]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data033),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][33] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][33] .power_up = "low";

dffeas \register_fifo:fifo_data[0][34] (
	.clk(clk),
	.d(datain[34]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data034),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][34] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][34] .power_up = "low";

dffeas \register_fifo:fifo_data[0][35] (
	.clk(clk),
	.d(datain[35]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data035),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][35] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][35] .power_up = "low";

dffeas \register_fifo:fifo_data[0][36] (
	.clk(clk),
	.d(datain[36]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data036),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][36] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][36] .power_up = "low";

dffeas \register_fifo:fifo_data[0][37] (
	.clk(clk),
	.d(datain[37]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data037),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][37] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][37] .power_up = "low";

dffeas \register_fifo:fifo_data[0][38] (
	.clk(clk),
	.d(datain[38]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data038),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][38] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][38] .power_up = "low";

dffeas \register_fifo:fifo_data[0][39] (
	.clk(clk),
	.d(datain[39]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data039),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][39] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][39] .power_up = "low";

dffeas \register_fifo:fifo_data[0][40] (
	.clk(clk),
	.d(datain[40]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data040),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][40] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][40] .power_up = "low";

dffeas \register_fifo:fifo_data[0][41] (
	.clk(clk),
	.d(datain[41]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data041),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][41] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][41] .power_up = "low";

dffeas \register_fifo:fifo_data[0][42] (
	.clk(clk),
	.d(datain[42]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data042),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][42] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][42] .power_up = "low";

dffeas \register_fifo:fifo_data[0][43] (
	.clk(clk),
	.d(datain[43]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data043),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][43] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][43] .power_up = "low";

dffeas \register_fifo:fifo_data[0][44] (
	.clk(clk),
	.d(datain[44]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data044),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][44] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][44] .power_up = "low";

dffeas \register_fifo:fifo_data[0][45] (
	.clk(clk),
	.d(datain[45]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data045),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][45] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][45] .power_up = "low";

dffeas \register_fifo:fifo_data[0][46] (
	.clk(clk),
	.d(datain[46]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data046),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][46] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][46] .power_up = "low";

dffeas \register_fifo:fifo_data[0][18] (
	.clk(clk),
	.d(datain[18]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data018),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][18] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][18] .power_up = "low";

dffeas \register_fifo:fifo_data[0][17] (
	.clk(clk),
	.d(datain[17]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data017),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][17] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][17] .power_up = "low";

dffeas \register_fifo:fifo_data[0][16] (
	.clk(clk),
	.d(datain[16]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data016),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][16] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][16] .power_up = "low";

dffeas \register_fifo:fifo_data[0][15] (
	.clk(clk),
	.d(datain[15]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data015),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][15] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][15] .power_up = "low";

dffeas \register_fifo:fifo_data[0][14] (
	.clk(clk),
	.d(datain[14]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data014),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][14] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][14] .power_up = "low";

dffeas \register_fifo:fifo_data[0][13] (
	.clk(clk),
	.d(datain[13]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data013),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][13] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][13] .power_up = "low";

dffeas \register_fifo:fifo_data[0][12] (
	.clk(clk),
	.d(datain[12]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data012),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][12] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][12] .power_up = "low";

dffeas \register_fifo:fifo_data[0][11] (
	.clk(clk),
	.d(datain[11]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data011),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][11] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][11] .power_up = "low";

dffeas \register_fifo:fifo_data[0][10] (
	.clk(clk),
	.d(datain[10]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data010),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][10] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][10] .power_up = "low";

dffeas \register_fifo:fifo_data[0][9] (
	.clk(clk),
	.d(datain[9]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data09),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][9] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][9] .power_up = "low";

dffeas \register_fifo:fifo_data[0][8] (
	.clk(clk),
	.d(datain[8]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data08),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][8] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][8] .power_up = "low";

dffeas \register_fifo:fifo_data[0][7] (
	.clk(clk),
	.d(datain[7]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data07),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][7] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][7] .power_up = "low";

dffeas \register_fifo:fifo_data[0][6] (
	.clk(clk),
	.d(datain[6]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data06),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][6] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][6] .power_up = "low";

dffeas \register_fifo:fifo_data[0][5] (
	.clk(clk),
	.d(datain[5]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data05),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][5] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][5] .power_up = "low";

dffeas \register_fifo:fifo_data[0][4] (
	.clk(clk),
	.d(datain[4]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data04),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][4] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][4] .power_up = "low";

dffeas \register_fifo:fifo_data[0][3] (
	.clk(clk),
	.d(datain[3]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data03),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][3] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][3] .power_up = "low";

dffeas \register_fifo:fifo_data[0][2] (
	.clk(clk),
	.d(datain[2]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data02),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][2] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][2] .power_up = "low";

dffeas \register_fifo:fifo_data[0][1] (
	.clk(clk),
	.d(datain[1]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data01),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][1] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][1] .power_up = "low";

dffeas \register_fifo:fifo_data[0][0] (
	.clk(clk),
	.d(datain[0]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data00),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][0] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][0] .power_up = "low";

endmodule

module cic_auk_dspip_integrator_2 (
	stall_reg,
	register_fifofifo_data019,
	register_fifofifo_data020,
	register_fifofifo_data021,
	register_fifofifo_data022,
	register_fifofifo_data023,
	register_fifofifo_data024,
	register_fifofifo_data025,
	register_fifofifo_data026,
	register_fifofifo_data027,
	register_fifofifo_data028,
	register_fifofifo_data029,
	register_fifofifo_data030,
	register_fifofifo_data031,
	register_fifofifo_data032,
	register_fifofifo_data033,
	register_fifofifo_data034,
	register_fifofifo_data035,
	register_fifofifo_data036,
	register_fifofifo_data037,
	register_fifofifo_data038,
	register_fifofifo_data039,
	register_fifofifo_data040,
	register_fifofifo_data041,
	register_fifofifo_data042,
	register_fifofifo_data043,
	register_fifofifo_data044,
	register_fifofifo_data045,
	register_fifofifo_data046,
	register_fifofifo_data018,
	register_fifofifo_data0191,
	register_fifofifo_data017,
	register_fifofifo_data0201,
	register_fifofifo_data0211,
	register_fifofifo_data0221,
	register_fifofifo_data0231,
	register_fifofifo_data0241,
	register_fifofifo_data0251,
	register_fifofifo_data0261,
	register_fifofifo_data0271,
	register_fifofifo_data0281,
	register_fifofifo_data0291,
	register_fifofifo_data0301,
	register_fifofifo_data0311,
	register_fifofifo_data0321,
	register_fifofifo_data0331,
	register_fifofifo_data0341,
	register_fifofifo_data0351,
	register_fifofifo_data0361,
	register_fifofifo_data0371,
	register_fifofifo_data0381,
	register_fifofifo_data0391,
	register_fifofifo_data0401,
	register_fifofifo_data0411,
	register_fifofifo_data0421,
	register_fifofifo_data0431,
	register_fifofifo_data0441,
	register_fifofifo_data0451,
	register_fifofifo_data0461,
	register_fifofifo_data0181,
	register_fifofifo_data016,
	register_fifofifo_data0171,
	register_fifofifo_data015,
	register_fifofifo_data0161,
	register_fifofifo_data014,
	register_fifofifo_data0151,
	register_fifofifo_data013,
	register_fifofifo_data0141,
	register_fifofifo_data012,
	register_fifofifo_data0131,
	register_fifofifo_data011,
	register_fifofifo_data0121,
	register_fifofifo_data010,
	register_fifofifo_data0111,
	register_fifofifo_data09,
	register_fifofifo_data0101,
	register_fifofifo_data08,
	register_fifofifo_data091,
	register_fifofifo_data07,
	register_fifofifo_data081,
	register_fifofifo_data06,
	register_fifofifo_data071,
	register_fifofifo_data05,
	register_fifofifo_data061,
	register_fifofifo_data04,
	register_fifofifo_data051,
	register_fifofifo_data03,
	register_fifofifo_data047,
	register_fifofifo_data02,
	register_fifofifo_data0310,
	register_fifofifo_data01,
	register_fifofifo_data0210,
	register_fifofifo_data0110,
	register_fifofifo_data00,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	stall_reg;
output 	register_fifofifo_data019;
output 	register_fifofifo_data020;
output 	register_fifofifo_data021;
output 	register_fifofifo_data022;
output 	register_fifofifo_data023;
output 	register_fifofifo_data024;
output 	register_fifofifo_data025;
output 	register_fifofifo_data026;
output 	register_fifofifo_data027;
output 	register_fifofifo_data028;
output 	register_fifofifo_data029;
output 	register_fifofifo_data030;
output 	register_fifofifo_data031;
output 	register_fifofifo_data032;
output 	register_fifofifo_data033;
output 	register_fifofifo_data034;
output 	register_fifofifo_data035;
output 	register_fifofifo_data036;
output 	register_fifofifo_data037;
output 	register_fifofifo_data038;
output 	register_fifofifo_data039;
output 	register_fifofifo_data040;
output 	register_fifofifo_data041;
output 	register_fifofifo_data042;
output 	register_fifofifo_data043;
output 	register_fifofifo_data044;
output 	register_fifofifo_data045;
output 	register_fifofifo_data046;
output 	register_fifofifo_data018;
input 	register_fifofifo_data0191;
output 	register_fifofifo_data017;
input 	register_fifofifo_data0201;
input 	register_fifofifo_data0211;
input 	register_fifofifo_data0221;
input 	register_fifofifo_data0231;
input 	register_fifofifo_data0241;
input 	register_fifofifo_data0251;
input 	register_fifofifo_data0261;
input 	register_fifofifo_data0271;
input 	register_fifofifo_data0281;
input 	register_fifofifo_data0291;
input 	register_fifofifo_data0301;
input 	register_fifofifo_data0311;
input 	register_fifofifo_data0321;
input 	register_fifofifo_data0331;
input 	register_fifofifo_data0341;
input 	register_fifofifo_data0351;
input 	register_fifofifo_data0361;
input 	register_fifofifo_data0371;
input 	register_fifofifo_data0381;
input 	register_fifofifo_data0391;
input 	register_fifofifo_data0401;
input 	register_fifofifo_data0411;
input 	register_fifofifo_data0421;
input 	register_fifofifo_data0431;
input 	register_fifofifo_data0441;
input 	register_fifofifo_data0451;
input 	register_fifofifo_data0461;
input 	register_fifofifo_data0181;
output 	register_fifofifo_data016;
input 	register_fifofifo_data0171;
output 	register_fifofifo_data015;
input 	register_fifofifo_data0161;
output 	register_fifofifo_data014;
input 	register_fifofifo_data0151;
output 	register_fifofifo_data013;
input 	register_fifofifo_data0141;
output 	register_fifofifo_data012;
input 	register_fifofifo_data0131;
output 	register_fifofifo_data011;
input 	register_fifofifo_data0121;
output 	register_fifofifo_data010;
input 	register_fifofifo_data0111;
output 	register_fifofifo_data09;
input 	register_fifofifo_data0101;
output 	register_fifofifo_data08;
input 	register_fifofifo_data091;
output 	register_fifofifo_data07;
input 	register_fifofifo_data081;
output 	register_fifofifo_data06;
input 	register_fifofifo_data071;
output 	register_fifofifo_data05;
input 	register_fifofifo_data061;
output 	register_fifofifo_data04;
input 	register_fifofifo_data051;
output 	register_fifofifo_data03;
input 	register_fifofifo_data047;
output 	register_fifofifo_data02;
input 	register_fifofifo_data0310;
output 	register_fifofifo_data01;
input 	register_fifofifo_data0210;
input 	register_fifofifo_data0110;
input 	register_fifofifo_data00;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Add0~1_sumout ;
wire \Add0~2 ;
wire \Add0~5_sumout ;
wire \Add0~6 ;
wire \Add0~9_sumout ;
wire \Add0~10 ;
wire \Add0~13_sumout ;
wire \Add0~14 ;
wire \Add0~17_sumout ;
wire \Add0~18 ;
wire \Add0~21_sumout ;
wire \Add0~22 ;
wire \Add0~25_sumout ;
wire \Add0~26 ;
wire \Add0~29_sumout ;
wire \Add0~30 ;
wire \Add0~33_sumout ;
wire \Add0~34 ;
wire \Add0~37_sumout ;
wire \Add0~38 ;
wire \Add0~41_sumout ;
wire \Add0~42 ;
wire \Add0~45_sumout ;
wire \Add0~46 ;
wire \Add0~49_sumout ;
wire \Add0~50 ;
wire \Add0~53_sumout ;
wire \Add0~54 ;
wire \Add0~57_sumout ;
wire \Add0~58 ;
wire \Add0~61_sumout ;
wire \Add0~62 ;
wire \Add0~65_sumout ;
wire \Add0~66 ;
wire \Add0~69_sumout ;
wire \Add0~70 ;
wire \Add0~73_sumout ;
wire \Add0~74 ;
wire \Add0~77_sumout ;
wire \Add0~78 ;
wire \Add0~81_sumout ;
wire \Add0~82 ;
wire \Add0~85_sumout ;
wire \Add0~86 ;
wire \Add0~89_sumout ;
wire \Add0~90 ;
wire \Add0~93_sumout ;
wire \Add0~94 ;
wire \Add0~97_sumout ;
wire \Add0~98 ;
wire \Add0~101_sumout ;
wire \Add0~102 ;
wire \Add0~105_sumout ;
wire \Add0~106 ;
wire \Add0~109_sumout ;
wire \Add0~113_sumout ;
wire \Add0~114 ;
wire \Add0~117_sumout ;
wire \Add0~118 ;
wire \Add0~121_sumout ;
wire \Add0~122 ;
wire \Add0~125_sumout ;
wire \Add0~126 ;
wire \Add0~129_sumout ;
wire \Add0~130 ;
wire \Add0~133_sumout ;
wire \Add0~134 ;
wire \Add0~137_sumout ;
wire \Add0~138 ;
wire \Add0~141_sumout ;
wire \Add0~142 ;
wire \Add0~145_sumout ;
wire \Add0~146 ;
wire \Add0~149_sumout ;
wire \Add0~150 ;
wire \Add0~153_sumout ;
wire \Add0~154 ;
wire \Add0~157_sumout ;
wire \Add0~158 ;
wire \Add0~161_sumout ;
wire \Add0~162 ;
wire \Add0~165_sumout ;
wire \Add0~166 ;
wire \Add0~169_sumout ;
wire \Add0~170 ;
wire \Add0~173_sumout ;
wire \Add0~174 ;
wire \Add0~177_sumout ;
wire \Add0~178 ;
wire \Add0~181_sumout ;
wire \Add0~182 ;
wire \Add0~185_sumout ;
wire \Add0~186 ;
wire \glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][0]~q ;


cic_auk_dspip_delay_10 \glogic:integrator_pipeline_0_generate:u1 (
	.datain({\Add0~109_sumout ,\Add0~105_sumout ,\Add0~101_sumout ,\Add0~97_sumout ,\Add0~93_sumout ,\Add0~89_sumout ,\Add0~85_sumout ,\Add0~81_sumout ,\Add0~77_sumout ,\Add0~73_sumout ,\Add0~69_sumout ,\Add0~65_sumout ,\Add0~61_sumout ,\Add0~57_sumout ,\Add0~53_sumout ,
\Add0~49_sumout ,\Add0~45_sumout ,\Add0~41_sumout ,\Add0~37_sumout ,\Add0~33_sumout ,\Add0~29_sumout ,\Add0~25_sumout ,\Add0~21_sumout ,\Add0~17_sumout ,\Add0~13_sumout ,\Add0~9_sumout ,\Add0~5_sumout ,\Add0~1_sumout ,\Add0~113_sumout ,\Add0~117_sumout ,\Add0~121_sumout ,
\Add0~125_sumout ,\Add0~129_sumout ,\Add0~133_sumout ,\Add0~137_sumout ,\Add0~141_sumout ,\Add0~145_sumout ,\Add0~149_sumout ,\Add0~153_sumout ,\Add0~157_sumout ,\Add0~161_sumout ,\Add0~165_sumout ,\Add0~169_sumout ,\Add0~173_sumout ,\Add0~177_sumout ,\Add0~181_sumout ,
\Add0~185_sumout }),
	.enable(stall_reg),
	.register_fifofifo_data019(register_fifofifo_data019),
	.register_fifofifo_data020(register_fifofifo_data020),
	.register_fifofifo_data021(register_fifofifo_data021),
	.register_fifofifo_data022(register_fifofifo_data022),
	.register_fifofifo_data023(register_fifofifo_data023),
	.register_fifofifo_data024(register_fifofifo_data024),
	.register_fifofifo_data025(register_fifofifo_data025),
	.register_fifofifo_data026(register_fifofifo_data026),
	.register_fifofifo_data027(register_fifofifo_data027),
	.register_fifofifo_data028(register_fifofifo_data028),
	.register_fifofifo_data029(register_fifofifo_data029),
	.register_fifofifo_data030(register_fifofifo_data030),
	.register_fifofifo_data031(register_fifofifo_data031),
	.register_fifofifo_data032(register_fifofifo_data032),
	.register_fifofifo_data033(register_fifofifo_data033),
	.register_fifofifo_data034(register_fifofifo_data034),
	.register_fifofifo_data035(register_fifofifo_data035),
	.register_fifofifo_data036(register_fifofifo_data036),
	.register_fifofifo_data037(register_fifofifo_data037),
	.register_fifofifo_data038(register_fifofifo_data038),
	.register_fifofifo_data039(register_fifofifo_data039),
	.register_fifofifo_data040(register_fifofifo_data040),
	.register_fifofifo_data041(register_fifofifo_data041),
	.register_fifofifo_data042(register_fifofifo_data042),
	.register_fifofifo_data043(register_fifofifo_data043),
	.register_fifofifo_data044(register_fifofifo_data044),
	.register_fifofifo_data045(register_fifofifo_data045),
	.register_fifofifo_data046(register_fifofifo_data046),
	.register_fifofifo_data018(register_fifofifo_data018),
	.register_fifofifo_data017(register_fifofifo_data017),
	.register_fifofifo_data016(register_fifofifo_data016),
	.register_fifofifo_data015(register_fifofifo_data015),
	.register_fifofifo_data014(register_fifofifo_data014),
	.register_fifofifo_data013(register_fifofifo_data013),
	.register_fifofifo_data012(register_fifofifo_data012),
	.register_fifofifo_data011(register_fifofifo_data011),
	.register_fifofifo_data010(register_fifofifo_data010),
	.register_fifofifo_data09(register_fifofifo_data09),
	.register_fifofifo_data08(register_fifofifo_data08),
	.register_fifofifo_data07(register_fifofifo_data07),
	.register_fifofifo_data06(register_fifofifo_data06),
	.register_fifofifo_data05(register_fifofifo_data05),
	.register_fifofifo_data04(register_fifofifo_data04),
	.register_fifofifo_data03(register_fifofifo_data03),
	.register_fifofifo_data02(register_fifofifo_data02),
	.register_fifofifo_data01(register_fifofifo_data01),
	.register_fifofifo_data00(\glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][0]~q ),
	.clk(clk),
	.reset(reset_n));

arriav_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data019),
	.datae(gnd),
	.dataf(!register_fifofifo_data0191),
	.datag(gnd),
	.cin(\Add0~114 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(\Add0~2 ),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~1 .shared_arith = "off";

arriav_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data020),
	.datae(gnd),
	.dataf(!register_fifofifo_data0201),
	.datag(gnd),
	.cin(\Add0~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~5 .shared_arith = "off";

arriav_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data021),
	.datae(gnd),
	.dataf(!register_fifofifo_data0211),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~9 .shared_arith = "off";

arriav_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data022),
	.datae(gnd),
	.dataf(!register_fifofifo_data0221),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~13 .shared_arith = "off";

arriav_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data023),
	.datae(gnd),
	.dataf(!register_fifofifo_data0231),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout());
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~17 .shared_arith = "off";

arriav_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data024),
	.datae(gnd),
	.dataf(!register_fifofifo_data0241),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout());
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~21 .shared_arith = "off";

arriav_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data025),
	.datae(gnd),
	.dataf(!register_fifofifo_data0251),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout());
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~25 .shared_arith = "off";

arriav_lcell_comb \Add0~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data026),
	.datae(gnd),
	.dataf(!register_fifofifo_data0261),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout());
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~29 .shared_arith = "off";

arriav_lcell_comb \Add0~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data027),
	.datae(gnd),
	.dataf(!register_fifofifo_data0271),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~33_sumout ),
	.cout(\Add0~34 ),
	.shareout());
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~33 .shared_arith = "off";

arriav_lcell_comb \Add0~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data028),
	.datae(gnd),
	.dataf(!register_fifofifo_data0281),
	.datag(gnd),
	.cin(\Add0~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~37_sumout ),
	.cout(\Add0~38 ),
	.shareout());
defparam \Add0~37 .extended_lut = "off";
defparam \Add0~37 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~37 .shared_arith = "off";

arriav_lcell_comb \Add0~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data029),
	.datae(gnd),
	.dataf(!register_fifofifo_data0291),
	.datag(gnd),
	.cin(\Add0~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~41_sumout ),
	.cout(\Add0~42 ),
	.shareout());
defparam \Add0~41 .extended_lut = "off";
defparam \Add0~41 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~41 .shared_arith = "off";

arriav_lcell_comb \Add0~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data030),
	.datae(gnd),
	.dataf(!register_fifofifo_data0301),
	.datag(gnd),
	.cin(\Add0~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~45_sumout ),
	.cout(\Add0~46 ),
	.shareout());
defparam \Add0~45 .extended_lut = "off";
defparam \Add0~45 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~45 .shared_arith = "off";

arriav_lcell_comb \Add0~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data031),
	.datae(gnd),
	.dataf(!register_fifofifo_data0311),
	.datag(gnd),
	.cin(\Add0~46 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~49_sumout ),
	.cout(\Add0~50 ),
	.shareout());
defparam \Add0~49 .extended_lut = "off";
defparam \Add0~49 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~49 .shared_arith = "off";

arriav_lcell_comb \Add0~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data032),
	.datae(gnd),
	.dataf(!register_fifofifo_data0321),
	.datag(gnd),
	.cin(\Add0~50 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~53_sumout ),
	.cout(\Add0~54 ),
	.shareout());
defparam \Add0~53 .extended_lut = "off";
defparam \Add0~53 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~53 .shared_arith = "off";

arriav_lcell_comb \Add0~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data033),
	.datae(gnd),
	.dataf(!register_fifofifo_data0331),
	.datag(gnd),
	.cin(\Add0~54 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~57_sumout ),
	.cout(\Add0~58 ),
	.shareout());
defparam \Add0~57 .extended_lut = "off";
defparam \Add0~57 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~57 .shared_arith = "off";

arriav_lcell_comb \Add0~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data034),
	.datae(gnd),
	.dataf(!register_fifofifo_data0341),
	.datag(gnd),
	.cin(\Add0~58 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~61_sumout ),
	.cout(\Add0~62 ),
	.shareout());
defparam \Add0~61 .extended_lut = "off";
defparam \Add0~61 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~61 .shared_arith = "off";

arriav_lcell_comb \Add0~65 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data035),
	.datae(gnd),
	.dataf(!register_fifofifo_data0351),
	.datag(gnd),
	.cin(\Add0~62 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~65_sumout ),
	.cout(\Add0~66 ),
	.shareout());
defparam \Add0~65 .extended_lut = "off";
defparam \Add0~65 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~65 .shared_arith = "off";

arriav_lcell_comb \Add0~69 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data036),
	.datae(gnd),
	.dataf(!register_fifofifo_data0361),
	.datag(gnd),
	.cin(\Add0~66 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~69_sumout ),
	.cout(\Add0~70 ),
	.shareout());
defparam \Add0~69 .extended_lut = "off";
defparam \Add0~69 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~69 .shared_arith = "off";

arriav_lcell_comb \Add0~73 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data037),
	.datae(gnd),
	.dataf(!register_fifofifo_data0371),
	.datag(gnd),
	.cin(\Add0~70 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~73_sumout ),
	.cout(\Add0~74 ),
	.shareout());
defparam \Add0~73 .extended_lut = "off";
defparam \Add0~73 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~73 .shared_arith = "off";

arriav_lcell_comb \Add0~77 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data038),
	.datae(gnd),
	.dataf(!register_fifofifo_data0381),
	.datag(gnd),
	.cin(\Add0~74 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~77_sumout ),
	.cout(\Add0~78 ),
	.shareout());
defparam \Add0~77 .extended_lut = "off";
defparam \Add0~77 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~77 .shared_arith = "off";

arriav_lcell_comb \Add0~81 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data039),
	.datae(gnd),
	.dataf(!register_fifofifo_data0391),
	.datag(gnd),
	.cin(\Add0~78 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~81_sumout ),
	.cout(\Add0~82 ),
	.shareout());
defparam \Add0~81 .extended_lut = "off";
defparam \Add0~81 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~81 .shared_arith = "off";

arriav_lcell_comb \Add0~85 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data040),
	.datae(gnd),
	.dataf(!register_fifofifo_data0401),
	.datag(gnd),
	.cin(\Add0~82 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~85_sumout ),
	.cout(\Add0~86 ),
	.shareout());
defparam \Add0~85 .extended_lut = "off";
defparam \Add0~85 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~85 .shared_arith = "off";

arriav_lcell_comb \Add0~89 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data041),
	.datae(gnd),
	.dataf(!register_fifofifo_data0411),
	.datag(gnd),
	.cin(\Add0~86 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~89_sumout ),
	.cout(\Add0~90 ),
	.shareout());
defparam \Add0~89 .extended_lut = "off";
defparam \Add0~89 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~89 .shared_arith = "off";

arriav_lcell_comb \Add0~93 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data042),
	.datae(gnd),
	.dataf(!register_fifofifo_data0421),
	.datag(gnd),
	.cin(\Add0~90 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~93_sumout ),
	.cout(\Add0~94 ),
	.shareout());
defparam \Add0~93 .extended_lut = "off";
defparam \Add0~93 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~93 .shared_arith = "off";

arriav_lcell_comb \Add0~97 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data043),
	.datae(gnd),
	.dataf(!register_fifofifo_data0431),
	.datag(gnd),
	.cin(\Add0~94 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~97_sumout ),
	.cout(\Add0~98 ),
	.shareout());
defparam \Add0~97 .extended_lut = "off";
defparam \Add0~97 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~97 .shared_arith = "off";

arriav_lcell_comb \Add0~101 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data044),
	.datae(gnd),
	.dataf(!register_fifofifo_data0441),
	.datag(gnd),
	.cin(\Add0~98 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~101_sumout ),
	.cout(\Add0~102 ),
	.shareout());
defparam \Add0~101 .extended_lut = "off";
defparam \Add0~101 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~101 .shared_arith = "off";

arriav_lcell_comb \Add0~105 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data045),
	.datae(gnd),
	.dataf(!register_fifofifo_data0451),
	.datag(gnd),
	.cin(\Add0~102 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~105_sumout ),
	.cout(\Add0~106 ),
	.shareout());
defparam \Add0~105 .extended_lut = "off";
defparam \Add0~105 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~105 .shared_arith = "off";

arriav_lcell_comb \Add0~109 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data046),
	.datae(gnd),
	.dataf(!register_fifofifo_data0461),
	.datag(gnd),
	.cin(\Add0~106 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~109_sumout ),
	.cout(),
	.shareout());
defparam \Add0~109 .extended_lut = "off";
defparam \Add0~109 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~109 .shared_arith = "off";

arriav_lcell_comb \Add0~113 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data018),
	.datae(gnd),
	.dataf(!register_fifofifo_data0181),
	.datag(gnd),
	.cin(\Add0~118 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~113_sumout ),
	.cout(\Add0~114 ),
	.shareout());
defparam \Add0~113 .extended_lut = "off";
defparam \Add0~113 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~113 .shared_arith = "off";

arriav_lcell_comb \Add0~117 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data017),
	.datae(gnd),
	.dataf(!register_fifofifo_data0171),
	.datag(gnd),
	.cin(\Add0~122 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~117_sumout ),
	.cout(\Add0~118 ),
	.shareout());
defparam \Add0~117 .extended_lut = "off";
defparam \Add0~117 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~117 .shared_arith = "off";

arriav_lcell_comb \Add0~121 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data016),
	.datae(gnd),
	.dataf(!register_fifofifo_data0161),
	.datag(gnd),
	.cin(\Add0~126 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~121_sumout ),
	.cout(\Add0~122 ),
	.shareout());
defparam \Add0~121 .extended_lut = "off";
defparam \Add0~121 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~121 .shared_arith = "off";

arriav_lcell_comb \Add0~125 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data015),
	.datae(gnd),
	.dataf(!register_fifofifo_data0151),
	.datag(gnd),
	.cin(\Add0~130 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~125_sumout ),
	.cout(\Add0~126 ),
	.shareout());
defparam \Add0~125 .extended_lut = "off";
defparam \Add0~125 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~125 .shared_arith = "off";

arriav_lcell_comb \Add0~129 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data014),
	.datae(gnd),
	.dataf(!register_fifofifo_data0141),
	.datag(gnd),
	.cin(\Add0~134 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~129_sumout ),
	.cout(\Add0~130 ),
	.shareout());
defparam \Add0~129 .extended_lut = "off";
defparam \Add0~129 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~129 .shared_arith = "off";

arriav_lcell_comb \Add0~133 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data013),
	.datae(gnd),
	.dataf(!register_fifofifo_data0131),
	.datag(gnd),
	.cin(\Add0~138 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~133_sumout ),
	.cout(\Add0~134 ),
	.shareout());
defparam \Add0~133 .extended_lut = "off";
defparam \Add0~133 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~133 .shared_arith = "off";

arriav_lcell_comb \Add0~137 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data012),
	.datae(gnd),
	.dataf(!register_fifofifo_data0121),
	.datag(gnd),
	.cin(\Add0~142 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~137_sumout ),
	.cout(\Add0~138 ),
	.shareout());
defparam \Add0~137 .extended_lut = "off";
defparam \Add0~137 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~137 .shared_arith = "off";

arriav_lcell_comb \Add0~141 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data011),
	.datae(gnd),
	.dataf(!register_fifofifo_data0111),
	.datag(gnd),
	.cin(\Add0~146 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~141_sumout ),
	.cout(\Add0~142 ),
	.shareout());
defparam \Add0~141 .extended_lut = "off";
defparam \Add0~141 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~141 .shared_arith = "off";

arriav_lcell_comb \Add0~145 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data010),
	.datae(gnd),
	.dataf(!register_fifofifo_data0101),
	.datag(gnd),
	.cin(\Add0~150 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~145_sumout ),
	.cout(\Add0~146 ),
	.shareout());
defparam \Add0~145 .extended_lut = "off";
defparam \Add0~145 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~145 .shared_arith = "off";

arriav_lcell_comb \Add0~149 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data09),
	.datae(gnd),
	.dataf(!register_fifofifo_data091),
	.datag(gnd),
	.cin(\Add0~154 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~149_sumout ),
	.cout(\Add0~150 ),
	.shareout());
defparam \Add0~149 .extended_lut = "off";
defparam \Add0~149 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~149 .shared_arith = "off";

arriav_lcell_comb \Add0~153 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data08),
	.datae(gnd),
	.dataf(!register_fifofifo_data081),
	.datag(gnd),
	.cin(\Add0~158 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~153_sumout ),
	.cout(\Add0~154 ),
	.shareout());
defparam \Add0~153 .extended_lut = "off";
defparam \Add0~153 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~153 .shared_arith = "off";

arriav_lcell_comb \Add0~157 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data07),
	.datae(gnd),
	.dataf(!register_fifofifo_data071),
	.datag(gnd),
	.cin(\Add0~162 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~157_sumout ),
	.cout(\Add0~158 ),
	.shareout());
defparam \Add0~157 .extended_lut = "off";
defparam \Add0~157 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~157 .shared_arith = "off";

arriav_lcell_comb \Add0~161 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data06),
	.datae(gnd),
	.dataf(!register_fifofifo_data061),
	.datag(gnd),
	.cin(\Add0~166 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~161_sumout ),
	.cout(\Add0~162 ),
	.shareout());
defparam \Add0~161 .extended_lut = "off";
defparam \Add0~161 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~161 .shared_arith = "off";

arriav_lcell_comb \Add0~165 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data05),
	.datae(gnd),
	.dataf(!register_fifofifo_data051),
	.datag(gnd),
	.cin(\Add0~170 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~165_sumout ),
	.cout(\Add0~166 ),
	.shareout());
defparam \Add0~165 .extended_lut = "off";
defparam \Add0~165 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~165 .shared_arith = "off";

arriav_lcell_comb \Add0~169 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data04),
	.datae(gnd),
	.dataf(!register_fifofifo_data047),
	.datag(gnd),
	.cin(\Add0~174 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~169_sumout ),
	.cout(\Add0~170 ),
	.shareout());
defparam \Add0~169 .extended_lut = "off";
defparam \Add0~169 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~169 .shared_arith = "off";

arriav_lcell_comb \Add0~173 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data03),
	.datae(gnd),
	.dataf(!register_fifofifo_data0310),
	.datag(gnd),
	.cin(\Add0~178 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~173_sumout ),
	.cout(\Add0~174 ),
	.shareout());
defparam \Add0~173 .extended_lut = "off";
defparam \Add0~173 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~173 .shared_arith = "off";

arriav_lcell_comb \Add0~177 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data02),
	.datae(gnd),
	.dataf(!register_fifofifo_data0210),
	.datag(gnd),
	.cin(\Add0~182 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~177_sumout ),
	.cout(\Add0~178 ),
	.shareout());
defparam \Add0~177 .extended_lut = "off";
defparam \Add0~177 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~177 .shared_arith = "off";

arriav_lcell_comb \Add0~181 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data01),
	.datae(gnd),
	.dataf(!register_fifofifo_data0110),
	.datag(gnd),
	.cin(\Add0~186 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~181_sumout ),
	.cout(\Add0~182 ),
	.shareout());
defparam \Add0~181 .extended_lut = "off";
defparam \Add0~181 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~181 .shared_arith = "off";

arriav_lcell_comb \Add0~185 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][0]~q ),
	.datae(gnd),
	.dataf(!register_fifofifo_data00),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~185_sumout ),
	.cout(\Add0~186 ),
	.shareout());
defparam \Add0~185 .extended_lut = "off";
defparam \Add0~185 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~185 .shared_arith = "off";

endmodule

module cic_auk_dspip_delay_10 (
	datain,
	enable,
	register_fifofifo_data019,
	register_fifofifo_data020,
	register_fifofifo_data021,
	register_fifofifo_data022,
	register_fifofifo_data023,
	register_fifofifo_data024,
	register_fifofifo_data025,
	register_fifofifo_data026,
	register_fifofifo_data027,
	register_fifofifo_data028,
	register_fifofifo_data029,
	register_fifofifo_data030,
	register_fifofifo_data031,
	register_fifofifo_data032,
	register_fifofifo_data033,
	register_fifofifo_data034,
	register_fifofifo_data035,
	register_fifofifo_data036,
	register_fifofifo_data037,
	register_fifofifo_data038,
	register_fifofifo_data039,
	register_fifofifo_data040,
	register_fifofifo_data041,
	register_fifofifo_data042,
	register_fifofifo_data043,
	register_fifofifo_data044,
	register_fifofifo_data045,
	register_fifofifo_data046,
	register_fifofifo_data018,
	register_fifofifo_data017,
	register_fifofifo_data016,
	register_fifofifo_data015,
	register_fifofifo_data014,
	register_fifofifo_data013,
	register_fifofifo_data012,
	register_fifofifo_data011,
	register_fifofifo_data010,
	register_fifofifo_data09,
	register_fifofifo_data08,
	register_fifofifo_data07,
	register_fifofifo_data06,
	register_fifofifo_data05,
	register_fifofifo_data04,
	register_fifofifo_data03,
	register_fifofifo_data02,
	register_fifofifo_data01,
	register_fifofifo_data00,
	clk,
	reset)/* synthesis synthesis_greybox=1 */;
input 	[46:0] datain;
input 	enable;
output 	register_fifofifo_data019;
output 	register_fifofifo_data020;
output 	register_fifofifo_data021;
output 	register_fifofifo_data022;
output 	register_fifofifo_data023;
output 	register_fifofifo_data024;
output 	register_fifofifo_data025;
output 	register_fifofifo_data026;
output 	register_fifofifo_data027;
output 	register_fifofifo_data028;
output 	register_fifofifo_data029;
output 	register_fifofifo_data030;
output 	register_fifofifo_data031;
output 	register_fifofifo_data032;
output 	register_fifofifo_data033;
output 	register_fifofifo_data034;
output 	register_fifofifo_data035;
output 	register_fifofifo_data036;
output 	register_fifofifo_data037;
output 	register_fifofifo_data038;
output 	register_fifofifo_data039;
output 	register_fifofifo_data040;
output 	register_fifofifo_data041;
output 	register_fifofifo_data042;
output 	register_fifofifo_data043;
output 	register_fifofifo_data044;
output 	register_fifofifo_data045;
output 	register_fifofifo_data046;
output 	register_fifofifo_data018;
output 	register_fifofifo_data017;
output 	register_fifofifo_data016;
output 	register_fifofifo_data015;
output 	register_fifofifo_data014;
output 	register_fifofifo_data013;
output 	register_fifofifo_data012;
output 	register_fifofifo_data011;
output 	register_fifofifo_data010;
output 	register_fifofifo_data09;
output 	register_fifofifo_data08;
output 	register_fifofifo_data07;
output 	register_fifofifo_data06;
output 	register_fifofifo_data05;
output 	register_fifofifo_data04;
output 	register_fifofifo_data03;
output 	register_fifofifo_data02;
output 	register_fifofifo_data01;
output 	register_fifofifo_data00;
input 	clk;
input 	reset;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \register_fifo:fifo_data[0][19] (
	.clk(clk),
	.d(datain[19]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data019),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][19] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][19] .power_up = "low";

dffeas \register_fifo:fifo_data[0][20] (
	.clk(clk),
	.d(datain[20]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data020),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][20] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][20] .power_up = "low";

dffeas \register_fifo:fifo_data[0][21] (
	.clk(clk),
	.d(datain[21]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data021),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][21] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][21] .power_up = "low";

dffeas \register_fifo:fifo_data[0][22] (
	.clk(clk),
	.d(datain[22]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data022),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][22] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][22] .power_up = "low";

dffeas \register_fifo:fifo_data[0][23] (
	.clk(clk),
	.d(datain[23]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data023),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][23] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][23] .power_up = "low";

dffeas \register_fifo:fifo_data[0][24] (
	.clk(clk),
	.d(datain[24]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data024),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][24] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][24] .power_up = "low";

dffeas \register_fifo:fifo_data[0][25] (
	.clk(clk),
	.d(datain[25]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data025),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][25] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][25] .power_up = "low";

dffeas \register_fifo:fifo_data[0][26] (
	.clk(clk),
	.d(datain[26]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data026),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][26] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][26] .power_up = "low";

dffeas \register_fifo:fifo_data[0][27] (
	.clk(clk),
	.d(datain[27]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data027),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][27] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][27] .power_up = "low";

dffeas \register_fifo:fifo_data[0][28] (
	.clk(clk),
	.d(datain[28]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data028),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][28] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][28] .power_up = "low";

dffeas \register_fifo:fifo_data[0][29] (
	.clk(clk),
	.d(datain[29]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data029),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][29] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][29] .power_up = "low";

dffeas \register_fifo:fifo_data[0][30] (
	.clk(clk),
	.d(datain[30]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data030),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][30] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][30] .power_up = "low";

dffeas \register_fifo:fifo_data[0][31] (
	.clk(clk),
	.d(datain[31]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data031),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][31] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][31] .power_up = "low";

dffeas \register_fifo:fifo_data[0][32] (
	.clk(clk),
	.d(datain[32]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data032),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][32] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][32] .power_up = "low";

dffeas \register_fifo:fifo_data[0][33] (
	.clk(clk),
	.d(datain[33]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data033),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][33] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][33] .power_up = "low";

dffeas \register_fifo:fifo_data[0][34] (
	.clk(clk),
	.d(datain[34]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data034),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][34] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][34] .power_up = "low";

dffeas \register_fifo:fifo_data[0][35] (
	.clk(clk),
	.d(datain[35]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data035),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][35] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][35] .power_up = "low";

dffeas \register_fifo:fifo_data[0][36] (
	.clk(clk),
	.d(datain[36]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data036),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][36] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][36] .power_up = "low";

dffeas \register_fifo:fifo_data[0][37] (
	.clk(clk),
	.d(datain[37]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data037),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][37] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][37] .power_up = "low";

dffeas \register_fifo:fifo_data[0][38] (
	.clk(clk),
	.d(datain[38]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data038),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][38] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][38] .power_up = "low";

dffeas \register_fifo:fifo_data[0][39] (
	.clk(clk),
	.d(datain[39]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data039),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][39] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][39] .power_up = "low";

dffeas \register_fifo:fifo_data[0][40] (
	.clk(clk),
	.d(datain[40]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data040),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][40] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][40] .power_up = "low";

dffeas \register_fifo:fifo_data[0][41] (
	.clk(clk),
	.d(datain[41]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data041),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][41] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][41] .power_up = "low";

dffeas \register_fifo:fifo_data[0][42] (
	.clk(clk),
	.d(datain[42]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data042),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][42] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][42] .power_up = "low";

dffeas \register_fifo:fifo_data[0][43] (
	.clk(clk),
	.d(datain[43]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data043),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][43] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][43] .power_up = "low";

dffeas \register_fifo:fifo_data[0][44] (
	.clk(clk),
	.d(datain[44]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data044),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][44] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][44] .power_up = "low";

dffeas \register_fifo:fifo_data[0][45] (
	.clk(clk),
	.d(datain[45]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data045),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][45] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][45] .power_up = "low";

dffeas \register_fifo:fifo_data[0][46] (
	.clk(clk),
	.d(datain[46]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data046),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][46] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][46] .power_up = "low";

dffeas \register_fifo:fifo_data[0][18] (
	.clk(clk),
	.d(datain[18]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data018),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][18] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][18] .power_up = "low";

dffeas \register_fifo:fifo_data[0][17] (
	.clk(clk),
	.d(datain[17]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data017),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][17] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][17] .power_up = "low";

dffeas \register_fifo:fifo_data[0][16] (
	.clk(clk),
	.d(datain[16]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data016),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][16] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][16] .power_up = "low";

dffeas \register_fifo:fifo_data[0][15] (
	.clk(clk),
	.d(datain[15]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data015),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][15] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][15] .power_up = "low";

dffeas \register_fifo:fifo_data[0][14] (
	.clk(clk),
	.d(datain[14]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data014),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][14] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][14] .power_up = "low";

dffeas \register_fifo:fifo_data[0][13] (
	.clk(clk),
	.d(datain[13]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data013),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][13] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][13] .power_up = "low";

dffeas \register_fifo:fifo_data[0][12] (
	.clk(clk),
	.d(datain[12]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data012),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][12] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][12] .power_up = "low";

dffeas \register_fifo:fifo_data[0][11] (
	.clk(clk),
	.d(datain[11]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data011),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][11] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][11] .power_up = "low";

dffeas \register_fifo:fifo_data[0][10] (
	.clk(clk),
	.d(datain[10]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data010),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][10] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][10] .power_up = "low";

dffeas \register_fifo:fifo_data[0][9] (
	.clk(clk),
	.d(datain[9]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data09),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][9] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][9] .power_up = "low";

dffeas \register_fifo:fifo_data[0][8] (
	.clk(clk),
	.d(datain[8]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data08),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][8] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][8] .power_up = "low";

dffeas \register_fifo:fifo_data[0][7] (
	.clk(clk),
	.d(datain[7]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data07),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][7] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][7] .power_up = "low";

dffeas \register_fifo:fifo_data[0][6] (
	.clk(clk),
	.d(datain[6]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data06),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][6] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][6] .power_up = "low";

dffeas \register_fifo:fifo_data[0][5] (
	.clk(clk),
	.d(datain[5]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data05),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][5] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][5] .power_up = "low";

dffeas \register_fifo:fifo_data[0][4] (
	.clk(clk),
	.d(datain[4]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data04),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][4] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][4] .power_up = "low";

dffeas \register_fifo:fifo_data[0][3] (
	.clk(clk),
	.d(datain[3]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data03),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][3] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][3] .power_up = "low";

dffeas \register_fifo:fifo_data[0][2] (
	.clk(clk),
	.d(datain[2]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data02),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][2] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][2] .power_up = "low";

dffeas \register_fifo:fifo_data[0][1] (
	.clk(clk),
	.d(datain[1]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data01),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][1] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][1] .power_up = "low";

dffeas \register_fifo:fifo_data[0][0] (
	.clk(clk),
	.d(datain[0]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data00),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][0] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][0] .power_up = "low";

endmodule

module cic_auk_dspip_integrator_3 (
	stall_reg,
	register_fifofifo_data018,
	register_fifofifo_data019,
	register_fifofifo_data020,
	register_fifofifo_data021,
	register_fifofifo_data022,
	register_fifofifo_data023,
	register_fifofifo_data024,
	register_fifofifo_data025,
	register_fifofifo_data026,
	register_fifofifo_data027,
	register_fifofifo_data028,
	register_fifofifo_data029,
	register_fifofifo_data030,
	register_fifofifo_data031,
	register_fifofifo_data032,
	register_fifofifo_data033,
	register_fifofifo_data034,
	register_fifofifo_data035,
	register_fifofifo_data036,
	register_fifofifo_data037,
	register_fifofifo_data038,
	register_fifofifo_data039,
	register_fifofifo_data040,
	register_fifofifo_data041,
	register_fifofifo_data042,
	register_fifofifo_data043,
	register_fifofifo_data044,
	register_fifofifo_data045,
	register_fifofifo_data017,
	register_fifofifo_data0191,
	register_fifofifo_data016,
	register_fifofifo_data0201,
	register_fifofifo_data0211,
	register_fifofifo_data0221,
	register_fifofifo_data0231,
	register_fifofifo_data0241,
	register_fifofifo_data0251,
	register_fifofifo_data0261,
	register_fifofifo_data0271,
	register_fifofifo_data0281,
	register_fifofifo_data0291,
	register_fifofifo_data0301,
	register_fifofifo_data0311,
	register_fifofifo_data0321,
	register_fifofifo_data0331,
	register_fifofifo_data0341,
	register_fifofifo_data0351,
	register_fifofifo_data0361,
	register_fifofifo_data0371,
	register_fifofifo_data0381,
	register_fifofifo_data0391,
	register_fifofifo_data0401,
	register_fifofifo_data0411,
	register_fifofifo_data0421,
	register_fifofifo_data0431,
	register_fifofifo_data0441,
	register_fifofifo_data0451,
	register_fifofifo_data046,
	register_fifofifo_data0181,
	register_fifofifo_data015,
	register_fifofifo_data0171,
	register_fifofifo_data014,
	register_fifofifo_data0161,
	register_fifofifo_data013,
	register_fifofifo_data0151,
	register_fifofifo_data012,
	register_fifofifo_data0141,
	register_fifofifo_data011,
	register_fifofifo_data0131,
	register_fifofifo_data010,
	register_fifofifo_data0121,
	register_fifofifo_data09,
	register_fifofifo_data0111,
	register_fifofifo_data08,
	register_fifofifo_data0101,
	register_fifofifo_data07,
	register_fifofifo_data091,
	register_fifofifo_data06,
	register_fifofifo_data081,
	register_fifofifo_data05,
	register_fifofifo_data071,
	register_fifofifo_data04,
	register_fifofifo_data061,
	register_fifofifo_data03,
	register_fifofifo_data051,
	register_fifofifo_data02,
	register_fifofifo_data047,
	register_fifofifo_data0310,
	register_fifofifo_data0210,
	register_fifofifo_data01,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	stall_reg;
output 	register_fifofifo_data018;
output 	register_fifofifo_data019;
output 	register_fifofifo_data020;
output 	register_fifofifo_data021;
output 	register_fifofifo_data022;
output 	register_fifofifo_data023;
output 	register_fifofifo_data024;
output 	register_fifofifo_data025;
output 	register_fifofifo_data026;
output 	register_fifofifo_data027;
output 	register_fifofifo_data028;
output 	register_fifofifo_data029;
output 	register_fifofifo_data030;
output 	register_fifofifo_data031;
output 	register_fifofifo_data032;
output 	register_fifofifo_data033;
output 	register_fifofifo_data034;
output 	register_fifofifo_data035;
output 	register_fifofifo_data036;
output 	register_fifofifo_data037;
output 	register_fifofifo_data038;
output 	register_fifofifo_data039;
output 	register_fifofifo_data040;
output 	register_fifofifo_data041;
output 	register_fifofifo_data042;
output 	register_fifofifo_data043;
output 	register_fifofifo_data044;
output 	register_fifofifo_data045;
output 	register_fifofifo_data017;
input 	register_fifofifo_data0191;
output 	register_fifofifo_data016;
input 	register_fifofifo_data0201;
input 	register_fifofifo_data0211;
input 	register_fifofifo_data0221;
input 	register_fifofifo_data0231;
input 	register_fifofifo_data0241;
input 	register_fifofifo_data0251;
input 	register_fifofifo_data0261;
input 	register_fifofifo_data0271;
input 	register_fifofifo_data0281;
input 	register_fifofifo_data0291;
input 	register_fifofifo_data0301;
input 	register_fifofifo_data0311;
input 	register_fifofifo_data0321;
input 	register_fifofifo_data0331;
input 	register_fifofifo_data0341;
input 	register_fifofifo_data0351;
input 	register_fifofifo_data0361;
input 	register_fifofifo_data0371;
input 	register_fifofifo_data0381;
input 	register_fifofifo_data0391;
input 	register_fifofifo_data0401;
input 	register_fifofifo_data0411;
input 	register_fifofifo_data0421;
input 	register_fifofifo_data0431;
input 	register_fifofifo_data0441;
input 	register_fifofifo_data0451;
input 	register_fifofifo_data046;
input 	register_fifofifo_data0181;
output 	register_fifofifo_data015;
input 	register_fifofifo_data0171;
output 	register_fifofifo_data014;
input 	register_fifofifo_data0161;
output 	register_fifofifo_data013;
input 	register_fifofifo_data0151;
output 	register_fifofifo_data012;
input 	register_fifofifo_data0141;
output 	register_fifofifo_data011;
input 	register_fifofifo_data0131;
output 	register_fifofifo_data010;
input 	register_fifofifo_data0121;
output 	register_fifofifo_data09;
input 	register_fifofifo_data0111;
output 	register_fifofifo_data08;
input 	register_fifofifo_data0101;
output 	register_fifofifo_data07;
input 	register_fifofifo_data091;
output 	register_fifofifo_data06;
input 	register_fifofifo_data081;
output 	register_fifofifo_data05;
input 	register_fifofifo_data071;
output 	register_fifofifo_data04;
input 	register_fifofifo_data061;
output 	register_fifofifo_data03;
input 	register_fifofifo_data051;
output 	register_fifofifo_data02;
input 	register_fifofifo_data047;
input 	register_fifofifo_data0310;
input 	register_fifofifo_data0210;
input 	register_fifofifo_data01;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Add0~1_sumout ;
wire \Add0~2 ;
wire \Add0~5_sumout ;
wire \Add0~6 ;
wire \Add0~9_sumout ;
wire \Add0~10 ;
wire \Add0~13_sumout ;
wire \Add0~14 ;
wire \Add0~17_sumout ;
wire \Add0~18 ;
wire \Add0~21_sumout ;
wire \Add0~22 ;
wire \Add0~25_sumout ;
wire \Add0~26 ;
wire \Add0~29_sumout ;
wire \Add0~30 ;
wire \Add0~33_sumout ;
wire \Add0~34 ;
wire \Add0~37_sumout ;
wire \Add0~38 ;
wire \Add0~41_sumout ;
wire \Add0~42 ;
wire \Add0~45_sumout ;
wire \Add0~46 ;
wire \Add0~49_sumout ;
wire \Add0~50 ;
wire \Add0~53_sumout ;
wire \Add0~54 ;
wire \Add0~57_sumout ;
wire \Add0~58 ;
wire \Add0~61_sumout ;
wire \Add0~62 ;
wire \Add0~65_sumout ;
wire \Add0~66 ;
wire \Add0~69_sumout ;
wire \Add0~70 ;
wire \Add0~73_sumout ;
wire \Add0~74 ;
wire \Add0~77_sumout ;
wire \Add0~78 ;
wire \Add0~81_sumout ;
wire \Add0~82 ;
wire \Add0~85_sumout ;
wire \Add0~86 ;
wire \Add0~89_sumout ;
wire \Add0~90 ;
wire \Add0~93_sumout ;
wire \Add0~94 ;
wire \Add0~97_sumout ;
wire \Add0~98 ;
wire \Add0~101_sumout ;
wire \Add0~102 ;
wire \Add0~105_sumout ;
wire \Add0~106 ;
wire \Add0~109_sumout ;
wire \Add0~113_sumout ;
wire \Add0~114 ;
wire \Add0~117_sumout ;
wire \Add0~118 ;
wire \Add0~121_sumout ;
wire \Add0~122 ;
wire \Add0~125_sumout ;
wire \Add0~126 ;
wire \Add0~129_sumout ;
wire \Add0~130 ;
wire \Add0~133_sumout ;
wire \Add0~134 ;
wire \Add0~137_sumout ;
wire \Add0~138 ;
wire \Add0~141_sumout ;
wire \Add0~142 ;
wire \Add0~145_sumout ;
wire \Add0~146 ;
wire \Add0~149_sumout ;
wire \Add0~150 ;
wire \Add0~153_sumout ;
wire \Add0~154 ;
wire \Add0~157_sumout ;
wire \Add0~158 ;
wire \Add0~161_sumout ;
wire \Add0~162 ;
wire \Add0~165_sumout ;
wire \Add0~166 ;
wire \Add0~169_sumout ;
wire \Add0~170 ;
wire \Add0~173_sumout ;
wire \Add0~174 ;
wire \Add0~177_sumout ;
wire \Add0~178 ;
wire \Add0~181_sumout ;
wire \Add0~182 ;
wire \glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][1]~q ;
wire \glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][0]~q ;


cic_auk_dspip_delay_11 \glogic:integrator_pipeline_0_generate:u1 (
	.datain({gnd,\Add0~109_sumout ,\Add0~105_sumout ,\Add0~101_sumout ,\Add0~97_sumout ,\Add0~93_sumout ,\Add0~89_sumout ,\Add0~85_sumout ,\Add0~81_sumout ,\Add0~77_sumout ,\Add0~73_sumout ,\Add0~69_sumout ,\Add0~65_sumout ,\Add0~61_sumout ,\Add0~57_sumout ,\Add0~53_sumout ,
\Add0~49_sumout ,\Add0~45_sumout ,\Add0~41_sumout ,\Add0~37_sumout ,\Add0~33_sumout ,\Add0~29_sumout ,\Add0~25_sumout ,\Add0~21_sumout ,\Add0~17_sumout ,\Add0~13_sumout ,\Add0~9_sumout ,\Add0~5_sumout ,\Add0~1_sumout ,\Add0~113_sumout ,\Add0~117_sumout ,\Add0~121_sumout ,
\Add0~125_sumout ,\Add0~129_sumout ,\Add0~133_sumout ,\Add0~137_sumout ,\Add0~141_sumout ,\Add0~145_sumout ,\Add0~149_sumout ,\Add0~153_sumout ,\Add0~157_sumout ,\Add0~161_sumout ,\Add0~165_sumout ,\Add0~169_sumout ,\Add0~173_sumout ,\Add0~177_sumout ,\Add0~181_sumout }),
	.enable(stall_reg),
	.register_fifofifo_data018(register_fifofifo_data018),
	.register_fifofifo_data019(register_fifofifo_data019),
	.register_fifofifo_data020(register_fifofifo_data020),
	.register_fifofifo_data021(register_fifofifo_data021),
	.register_fifofifo_data022(register_fifofifo_data022),
	.register_fifofifo_data023(register_fifofifo_data023),
	.register_fifofifo_data024(register_fifofifo_data024),
	.register_fifofifo_data025(register_fifofifo_data025),
	.register_fifofifo_data026(register_fifofifo_data026),
	.register_fifofifo_data027(register_fifofifo_data027),
	.register_fifofifo_data028(register_fifofifo_data028),
	.register_fifofifo_data029(register_fifofifo_data029),
	.register_fifofifo_data030(register_fifofifo_data030),
	.register_fifofifo_data031(register_fifofifo_data031),
	.register_fifofifo_data032(register_fifofifo_data032),
	.register_fifofifo_data033(register_fifofifo_data033),
	.register_fifofifo_data034(register_fifofifo_data034),
	.register_fifofifo_data035(register_fifofifo_data035),
	.register_fifofifo_data036(register_fifofifo_data036),
	.register_fifofifo_data037(register_fifofifo_data037),
	.register_fifofifo_data038(register_fifofifo_data038),
	.register_fifofifo_data039(register_fifofifo_data039),
	.register_fifofifo_data040(register_fifofifo_data040),
	.register_fifofifo_data041(register_fifofifo_data041),
	.register_fifofifo_data042(register_fifofifo_data042),
	.register_fifofifo_data043(register_fifofifo_data043),
	.register_fifofifo_data044(register_fifofifo_data044),
	.register_fifofifo_data045(register_fifofifo_data045),
	.register_fifofifo_data017(register_fifofifo_data017),
	.register_fifofifo_data016(register_fifofifo_data016),
	.register_fifofifo_data015(register_fifofifo_data015),
	.register_fifofifo_data014(register_fifofifo_data014),
	.register_fifofifo_data013(register_fifofifo_data013),
	.register_fifofifo_data012(register_fifofifo_data012),
	.register_fifofifo_data011(register_fifofifo_data011),
	.register_fifofifo_data010(register_fifofifo_data010),
	.register_fifofifo_data09(register_fifofifo_data09),
	.register_fifofifo_data08(register_fifofifo_data08),
	.register_fifofifo_data07(register_fifofifo_data07),
	.register_fifofifo_data06(register_fifofifo_data06),
	.register_fifofifo_data05(register_fifofifo_data05),
	.register_fifofifo_data04(register_fifofifo_data04),
	.register_fifofifo_data03(register_fifofifo_data03),
	.register_fifofifo_data02(register_fifofifo_data02),
	.register_fifofifo_data01(\glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][1]~q ),
	.register_fifofifo_data00(\glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][0]~q ),
	.clk(clk),
	.reset(reset_n));

arriav_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data018),
	.datae(gnd),
	.dataf(!register_fifofifo_data0191),
	.datag(gnd),
	.cin(\Add0~114 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(\Add0~2 ),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~1 .shared_arith = "off";

arriav_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data019),
	.datae(gnd),
	.dataf(!register_fifofifo_data0201),
	.datag(gnd),
	.cin(\Add0~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~5 .shared_arith = "off";

arriav_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data020),
	.datae(gnd),
	.dataf(!register_fifofifo_data0211),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~9 .shared_arith = "off";

arriav_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data021),
	.datae(gnd),
	.dataf(!register_fifofifo_data0221),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~13 .shared_arith = "off";

arriav_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data022),
	.datae(gnd),
	.dataf(!register_fifofifo_data0231),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout());
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~17 .shared_arith = "off";

arriav_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data023),
	.datae(gnd),
	.dataf(!register_fifofifo_data0241),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout());
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~21 .shared_arith = "off";

arriav_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data024),
	.datae(gnd),
	.dataf(!register_fifofifo_data0251),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout());
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~25 .shared_arith = "off";

arriav_lcell_comb \Add0~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data025),
	.datae(gnd),
	.dataf(!register_fifofifo_data0261),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout());
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~29 .shared_arith = "off";

arriav_lcell_comb \Add0~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data026),
	.datae(gnd),
	.dataf(!register_fifofifo_data0271),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~33_sumout ),
	.cout(\Add0~34 ),
	.shareout());
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~33 .shared_arith = "off";

arriav_lcell_comb \Add0~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data027),
	.datae(gnd),
	.dataf(!register_fifofifo_data0281),
	.datag(gnd),
	.cin(\Add0~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~37_sumout ),
	.cout(\Add0~38 ),
	.shareout());
defparam \Add0~37 .extended_lut = "off";
defparam \Add0~37 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~37 .shared_arith = "off";

arriav_lcell_comb \Add0~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data028),
	.datae(gnd),
	.dataf(!register_fifofifo_data0291),
	.datag(gnd),
	.cin(\Add0~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~41_sumout ),
	.cout(\Add0~42 ),
	.shareout());
defparam \Add0~41 .extended_lut = "off";
defparam \Add0~41 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~41 .shared_arith = "off";

arriav_lcell_comb \Add0~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data029),
	.datae(gnd),
	.dataf(!register_fifofifo_data0301),
	.datag(gnd),
	.cin(\Add0~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~45_sumout ),
	.cout(\Add0~46 ),
	.shareout());
defparam \Add0~45 .extended_lut = "off";
defparam \Add0~45 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~45 .shared_arith = "off";

arriav_lcell_comb \Add0~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data030),
	.datae(gnd),
	.dataf(!register_fifofifo_data0311),
	.datag(gnd),
	.cin(\Add0~46 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~49_sumout ),
	.cout(\Add0~50 ),
	.shareout());
defparam \Add0~49 .extended_lut = "off";
defparam \Add0~49 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~49 .shared_arith = "off";

arriav_lcell_comb \Add0~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data031),
	.datae(gnd),
	.dataf(!register_fifofifo_data0321),
	.datag(gnd),
	.cin(\Add0~50 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~53_sumout ),
	.cout(\Add0~54 ),
	.shareout());
defparam \Add0~53 .extended_lut = "off";
defparam \Add0~53 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~53 .shared_arith = "off";

arriav_lcell_comb \Add0~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data032),
	.datae(gnd),
	.dataf(!register_fifofifo_data0331),
	.datag(gnd),
	.cin(\Add0~54 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~57_sumout ),
	.cout(\Add0~58 ),
	.shareout());
defparam \Add0~57 .extended_lut = "off";
defparam \Add0~57 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~57 .shared_arith = "off";

arriav_lcell_comb \Add0~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data033),
	.datae(gnd),
	.dataf(!register_fifofifo_data0341),
	.datag(gnd),
	.cin(\Add0~58 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~61_sumout ),
	.cout(\Add0~62 ),
	.shareout());
defparam \Add0~61 .extended_lut = "off";
defparam \Add0~61 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~61 .shared_arith = "off";

arriav_lcell_comb \Add0~65 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data034),
	.datae(gnd),
	.dataf(!register_fifofifo_data0351),
	.datag(gnd),
	.cin(\Add0~62 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~65_sumout ),
	.cout(\Add0~66 ),
	.shareout());
defparam \Add0~65 .extended_lut = "off";
defparam \Add0~65 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~65 .shared_arith = "off";

arriav_lcell_comb \Add0~69 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data035),
	.datae(gnd),
	.dataf(!register_fifofifo_data0361),
	.datag(gnd),
	.cin(\Add0~66 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~69_sumout ),
	.cout(\Add0~70 ),
	.shareout());
defparam \Add0~69 .extended_lut = "off";
defparam \Add0~69 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~69 .shared_arith = "off";

arriav_lcell_comb \Add0~73 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data036),
	.datae(gnd),
	.dataf(!register_fifofifo_data0371),
	.datag(gnd),
	.cin(\Add0~70 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~73_sumout ),
	.cout(\Add0~74 ),
	.shareout());
defparam \Add0~73 .extended_lut = "off";
defparam \Add0~73 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~73 .shared_arith = "off";

arriav_lcell_comb \Add0~77 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data037),
	.datae(gnd),
	.dataf(!register_fifofifo_data0381),
	.datag(gnd),
	.cin(\Add0~74 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~77_sumout ),
	.cout(\Add0~78 ),
	.shareout());
defparam \Add0~77 .extended_lut = "off";
defparam \Add0~77 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~77 .shared_arith = "off";

arriav_lcell_comb \Add0~81 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data038),
	.datae(gnd),
	.dataf(!register_fifofifo_data0391),
	.datag(gnd),
	.cin(\Add0~78 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~81_sumout ),
	.cout(\Add0~82 ),
	.shareout());
defparam \Add0~81 .extended_lut = "off";
defparam \Add0~81 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~81 .shared_arith = "off";

arriav_lcell_comb \Add0~85 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data039),
	.datae(gnd),
	.dataf(!register_fifofifo_data0401),
	.datag(gnd),
	.cin(\Add0~82 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~85_sumout ),
	.cout(\Add0~86 ),
	.shareout());
defparam \Add0~85 .extended_lut = "off";
defparam \Add0~85 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~85 .shared_arith = "off";

arriav_lcell_comb \Add0~89 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data040),
	.datae(gnd),
	.dataf(!register_fifofifo_data0411),
	.datag(gnd),
	.cin(\Add0~86 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~89_sumout ),
	.cout(\Add0~90 ),
	.shareout());
defparam \Add0~89 .extended_lut = "off";
defparam \Add0~89 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~89 .shared_arith = "off";

arriav_lcell_comb \Add0~93 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data041),
	.datae(gnd),
	.dataf(!register_fifofifo_data0421),
	.datag(gnd),
	.cin(\Add0~90 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~93_sumout ),
	.cout(\Add0~94 ),
	.shareout());
defparam \Add0~93 .extended_lut = "off";
defparam \Add0~93 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~93 .shared_arith = "off";

arriav_lcell_comb \Add0~97 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data042),
	.datae(gnd),
	.dataf(!register_fifofifo_data0431),
	.datag(gnd),
	.cin(\Add0~94 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~97_sumout ),
	.cout(\Add0~98 ),
	.shareout());
defparam \Add0~97 .extended_lut = "off";
defparam \Add0~97 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~97 .shared_arith = "off";

arriav_lcell_comb \Add0~101 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data043),
	.datae(gnd),
	.dataf(!register_fifofifo_data0441),
	.datag(gnd),
	.cin(\Add0~98 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~101_sumout ),
	.cout(\Add0~102 ),
	.shareout());
defparam \Add0~101 .extended_lut = "off";
defparam \Add0~101 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~101 .shared_arith = "off";

arriav_lcell_comb \Add0~105 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data044),
	.datae(gnd),
	.dataf(!register_fifofifo_data0451),
	.datag(gnd),
	.cin(\Add0~102 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~105_sumout ),
	.cout(\Add0~106 ),
	.shareout());
defparam \Add0~105 .extended_lut = "off";
defparam \Add0~105 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~105 .shared_arith = "off";

arriav_lcell_comb \Add0~109 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data045),
	.datae(gnd),
	.dataf(!register_fifofifo_data046),
	.datag(gnd),
	.cin(\Add0~106 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~109_sumout ),
	.cout(),
	.shareout());
defparam \Add0~109 .extended_lut = "off";
defparam \Add0~109 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~109 .shared_arith = "off";

arriav_lcell_comb \Add0~113 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data017),
	.datae(gnd),
	.dataf(!register_fifofifo_data0181),
	.datag(gnd),
	.cin(\Add0~118 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~113_sumout ),
	.cout(\Add0~114 ),
	.shareout());
defparam \Add0~113 .extended_lut = "off";
defparam \Add0~113 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~113 .shared_arith = "off";

arriav_lcell_comb \Add0~117 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data016),
	.datae(gnd),
	.dataf(!register_fifofifo_data0171),
	.datag(gnd),
	.cin(\Add0~122 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~117_sumout ),
	.cout(\Add0~118 ),
	.shareout());
defparam \Add0~117 .extended_lut = "off";
defparam \Add0~117 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~117 .shared_arith = "off";

arriav_lcell_comb \Add0~121 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data015),
	.datae(gnd),
	.dataf(!register_fifofifo_data0161),
	.datag(gnd),
	.cin(\Add0~126 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~121_sumout ),
	.cout(\Add0~122 ),
	.shareout());
defparam \Add0~121 .extended_lut = "off";
defparam \Add0~121 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~121 .shared_arith = "off";

arriav_lcell_comb \Add0~125 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data014),
	.datae(gnd),
	.dataf(!register_fifofifo_data0151),
	.datag(gnd),
	.cin(\Add0~130 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~125_sumout ),
	.cout(\Add0~126 ),
	.shareout());
defparam \Add0~125 .extended_lut = "off";
defparam \Add0~125 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~125 .shared_arith = "off";

arriav_lcell_comb \Add0~129 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data013),
	.datae(gnd),
	.dataf(!register_fifofifo_data0141),
	.datag(gnd),
	.cin(\Add0~134 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~129_sumout ),
	.cout(\Add0~130 ),
	.shareout());
defparam \Add0~129 .extended_lut = "off";
defparam \Add0~129 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~129 .shared_arith = "off";

arriav_lcell_comb \Add0~133 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data012),
	.datae(gnd),
	.dataf(!register_fifofifo_data0131),
	.datag(gnd),
	.cin(\Add0~138 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~133_sumout ),
	.cout(\Add0~134 ),
	.shareout());
defparam \Add0~133 .extended_lut = "off";
defparam \Add0~133 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~133 .shared_arith = "off";

arriav_lcell_comb \Add0~137 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data011),
	.datae(gnd),
	.dataf(!register_fifofifo_data0121),
	.datag(gnd),
	.cin(\Add0~142 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~137_sumout ),
	.cout(\Add0~138 ),
	.shareout());
defparam \Add0~137 .extended_lut = "off";
defparam \Add0~137 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~137 .shared_arith = "off";

arriav_lcell_comb \Add0~141 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data010),
	.datae(gnd),
	.dataf(!register_fifofifo_data0111),
	.datag(gnd),
	.cin(\Add0~146 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~141_sumout ),
	.cout(\Add0~142 ),
	.shareout());
defparam \Add0~141 .extended_lut = "off";
defparam \Add0~141 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~141 .shared_arith = "off";

arriav_lcell_comb \Add0~145 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data09),
	.datae(gnd),
	.dataf(!register_fifofifo_data0101),
	.datag(gnd),
	.cin(\Add0~150 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~145_sumout ),
	.cout(\Add0~146 ),
	.shareout());
defparam \Add0~145 .extended_lut = "off";
defparam \Add0~145 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~145 .shared_arith = "off";

arriav_lcell_comb \Add0~149 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data08),
	.datae(gnd),
	.dataf(!register_fifofifo_data091),
	.datag(gnd),
	.cin(\Add0~154 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~149_sumout ),
	.cout(\Add0~150 ),
	.shareout());
defparam \Add0~149 .extended_lut = "off";
defparam \Add0~149 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~149 .shared_arith = "off";

arriav_lcell_comb \Add0~153 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data07),
	.datae(gnd),
	.dataf(!register_fifofifo_data081),
	.datag(gnd),
	.cin(\Add0~158 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~153_sumout ),
	.cout(\Add0~154 ),
	.shareout());
defparam \Add0~153 .extended_lut = "off";
defparam \Add0~153 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~153 .shared_arith = "off";

arriav_lcell_comb \Add0~157 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data06),
	.datae(gnd),
	.dataf(!register_fifofifo_data071),
	.datag(gnd),
	.cin(\Add0~162 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~157_sumout ),
	.cout(\Add0~158 ),
	.shareout());
defparam \Add0~157 .extended_lut = "off";
defparam \Add0~157 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~157 .shared_arith = "off";

arriav_lcell_comb \Add0~161 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data05),
	.datae(gnd),
	.dataf(!register_fifofifo_data061),
	.datag(gnd),
	.cin(\Add0~166 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~161_sumout ),
	.cout(\Add0~162 ),
	.shareout());
defparam \Add0~161 .extended_lut = "off";
defparam \Add0~161 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~161 .shared_arith = "off";

arriav_lcell_comb \Add0~165 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data04),
	.datae(gnd),
	.dataf(!register_fifofifo_data051),
	.datag(gnd),
	.cin(\Add0~170 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~165_sumout ),
	.cout(\Add0~166 ),
	.shareout());
defparam \Add0~165 .extended_lut = "off";
defparam \Add0~165 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~165 .shared_arith = "off";

arriav_lcell_comb \Add0~169 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data03),
	.datae(gnd),
	.dataf(!register_fifofifo_data047),
	.datag(gnd),
	.cin(\Add0~174 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~169_sumout ),
	.cout(\Add0~170 ),
	.shareout());
defparam \Add0~169 .extended_lut = "off";
defparam \Add0~169 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~169 .shared_arith = "off";

arriav_lcell_comb \Add0~173 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data02),
	.datae(gnd),
	.dataf(!register_fifofifo_data0310),
	.datag(gnd),
	.cin(\Add0~178 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~173_sumout ),
	.cout(\Add0~174 ),
	.shareout());
defparam \Add0~173 .extended_lut = "off";
defparam \Add0~173 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~173 .shared_arith = "off";

arriav_lcell_comb \Add0~177 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][1]~q ),
	.datae(gnd),
	.dataf(!register_fifofifo_data0210),
	.datag(gnd),
	.cin(\Add0~182 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~177_sumout ),
	.cout(\Add0~178 ),
	.shareout());
defparam \Add0~177 .extended_lut = "off";
defparam \Add0~177 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~177 .shared_arith = "off";

arriav_lcell_comb \Add0~181 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][0]~q ),
	.datae(gnd),
	.dataf(!register_fifofifo_data01),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~181_sumout ),
	.cout(\Add0~182 ),
	.shareout());
defparam \Add0~181 .extended_lut = "off";
defparam \Add0~181 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~181 .shared_arith = "off";

endmodule

module cic_auk_dspip_delay_11 (
	datain,
	enable,
	register_fifofifo_data018,
	register_fifofifo_data019,
	register_fifofifo_data020,
	register_fifofifo_data021,
	register_fifofifo_data022,
	register_fifofifo_data023,
	register_fifofifo_data024,
	register_fifofifo_data025,
	register_fifofifo_data026,
	register_fifofifo_data027,
	register_fifofifo_data028,
	register_fifofifo_data029,
	register_fifofifo_data030,
	register_fifofifo_data031,
	register_fifofifo_data032,
	register_fifofifo_data033,
	register_fifofifo_data034,
	register_fifofifo_data035,
	register_fifofifo_data036,
	register_fifofifo_data037,
	register_fifofifo_data038,
	register_fifofifo_data039,
	register_fifofifo_data040,
	register_fifofifo_data041,
	register_fifofifo_data042,
	register_fifofifo_data043,
	register_fifofifo_data044,
	register_fifofifo_data045,
	register_fifofifo_data017,
	register_fifofifo_data016,
	register_fifofifo_data015,
	register_fifofifo_data014,
	register_fifofifo_data013,
	register_fifofifo_data012,
	register_fifofifo_data011,
	register_fifofifo_data010,
	register_fifofifo_data09,
	register_fifofifo_data08,
	register_fifofifo_data07,
	register_fifofifo_data06,
	register_fifofifo_data05,
	register_fifofifo_data04,
	register_fifofifo_data03,
	register_fifofifo_data02,
	register_fifofifo_data01,
	register_fifofifo_data00,
	clk,
	reset)/* synthesis synthesis_greybox=1 */;
input 	[46:0] datain;
input 	enable;
output 	register_fifofifo_data018;
output 	register_fifofifo_data019;
output 	register_fifofifo_data020;
output 	register_fifofifo_data021;
output 	register_fifofifo_data022;
output 	register_fifofifo_data023;
output 	register_fifofifo_data024;
output 	register_fifofifo_data025;
output 	register_fifofifo_data026;
output 	register_fifofifo_data027;
output 	register_fifofifo_data028;
output 	register_fifofifo_data029;
output 	register_fifofifo_data030;
output 	register_fifofifo_data031;
output 	register_fifofifo_data032;
output 	register_fifofifo_data033;
output 	register_fifofifo_data034;
output 	register_fifofifo_data035;
output 	register_fifofifo_data036;
output 	register_fifofifo_data037;
output 	register_fifofifo_data038;
output 	register_fifofifo_data039;
output 	register_fifofifo_data040;
output 	register_fifofifo_data041;
output 	register_fifofifo_data042;
output 	register_fifofifo_data043;
output 	register_fifofifo_data044;
output 	register_fifofifo_data045;
output 	register_fifofifo_data017;
output 	register_fifofifo_data016;
output 	register_fifofifo_data015;
output 	register_fifofifo_data014;
output 	register_fifofifo_data013;
output 	register_fifofifo_data012;
output 	register_fifofifo_data011;
output 	register_fifofifo_data010;
output 	register_fifofifo_data09;
output 	register_fifofifo_data08;
output 	register_fifofifo_data07;
output 	register_fifofifo_data06;
output 	register_fifofifo_data05;
output 	register_fifofifo_data04;
output 	register_fifofifo_data03;
output 	register_fifofifo_data02;
output 	register_fifofifo_data01;
output 	register_fifofifo_data00;
input 	clk;
input 	reset;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \register_fifo:fifo_data[0][18] (
	.clk(clk),
	.d(datain[18]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data018),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][18] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][18] .power_up = "low";

dffeas \register_fifo:fifo_data[0][19] (
	.clk(clk),
	.d(datain[19]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data019),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][19] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][19] .power_up = "low";

dffeas \register_fifo:fifo_data[0][20] (
	.clk(clk),
	.d(datain[20]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data020),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][20] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][20] .power_up = "low";

dffeas \register_fifo:fifo_data[0][21] (
	.clk(clk),
	.d(datain[21]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data021),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][21] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][21] .power_up = "low";

dffeas \register_fifo:fifo_data[0][22] (
	.clk(clk),
	.d(datain[22]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data022),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][22] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][22] .power_up = "low";

dffeas \register_fifo:fifo_data[0][23] (
	.clk(clk),
	.d(datain[23]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data023),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][23] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][23] .power_up = "low";

dffeas \register_fifo:fifo_data[0][24] (
	.clk(clk),
	.d(datain[24]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data024),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][24] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][24] .power_up = "low";

dffeas \register_fifo:fifo_data[0][25] (
	.clk(clk),
	.d(datain[25]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data025),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][25] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][25] .power_up = "low";

dffeas \register_fifo:fifo_data[0][26] (
	.clk(clk),
	.d(datain[26]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data026),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][26] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][26] .power_up = "low";

dffeas \register_fifo:fifo_data[0][27] (
	.clk(clk),
	.d(datain[27]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data027),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][27] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][27] .power_up = "low";

dffeas \register_fifo:fifo_data[0][28] (
	.clk(clk),
	.d(datain[28]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data028),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][28] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][28] .power_up = "low";

dffeas \register_fifo:fifo_data[0][29] (
	.clk(clk),
	.d(datain[29]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data029),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][29] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][29] .power_up = "low";

dffeas \register_fifo:fifo_data[0][30] (
	.clk(clk),
	.d(datain[30]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data030),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][30] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][30] .power_up = "low";

dffeas \register_fifo:fifo_data[0][31] (
	.clk(clk),
	.d(datain[31]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data031),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][31] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][31] .power_up = "low";

dffeas \register_fifo:fifo_data[0][32] (
	.clk(clk),
	.d(datain[32]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data032),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][32] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][32] .power_up = "low";

dffeas \register_fifo:fifo_data[0][33] (
	.clk(clk),
	.d(datain[33]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data033),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][33] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][33] .power_up = "low";

dffeas \register_fifo:fifo_data[0][34] (
	.clk(clk),
	.d(datain[34]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data034),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][34] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][34] .power_up = "low";

dffeas \register_fifo:fifo_data[0][35] (
	.clk(clk),
	.d(datain[35]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data035),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][35] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][35] .power_up = "low";

dffeas \register_fifo:fifo_data[0][36] (
	.clk(clk),
	.d(datain[36]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data036),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][36] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][36] .power_up = "low";

dffeas \register_fifo:fifo_data[0][37] (
	.clk(clk),
	.d(datain[37]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data037),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][37] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][37] .power_up = "low";

dffeas \register_fifo:fifo_data[0][38] (
	.clk(clk),
	.d(datain[38]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data038),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][38] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][38] .power_up = "low";

dffeas \register_fifo:fifo_data[0][39] (
	.clk(clk),
	.d(datain[39]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data039),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][39] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][39] .power_up = "low";

dffeas \register_fifo:fifo_data[0][40] (
	.clk(clk),
	.d(datain[40]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data040),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][40] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][40] .power_up = "low";

dffeas \register_fifo:fifo_data[0][41] (
	.clk(clk),
	.d(datain[41]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data041),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][41] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][41] .power_up = "low";

dffeas \register_fifo:fifo_data[0][42] (
	.clk(clk),
	.d(datain[42]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data042),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][42] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][42] .power_up = "low";

dffeas \register_fifo:fifo_data[0][43] (
	.clk(clk),
	.d(datain[43]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data043),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][43] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][43] .power_up = "low";

dffeas \register_fifo:fifo_data[0][44] (
	.clk(clk),
	.d(datain[44]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data044),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][44] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][44] .power_up = "low";

dffeas \register_fifo:fifo_data[0][45] (
	.clk(clk),
	.d(datain[45]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data045),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][45] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][45] .power_up = "low";

dffeas \register_fifo:fifo_data[0][17] (
	.clk(clk),
	.d(datain[17]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data017),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][17] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][17] .power_up = "low";

dffeas \register_fifo:fifo_data[0][16] (
	.clk(clk),
	.d(datain[16]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data016),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][16] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][16] .power_up = "low";

dffeas \register_fifo:fifo_data[0][15] (
	.clk(clk),
	.d(datain[15]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data015),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][15] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][15] .power_up = "low";

dffeas \register_fifo:fifo_data[0][14] (
	.clk(clk),
	.d(datain[14]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data014),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][14] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][14] .power_up = "low";

dffeas \register_fifo:fifo_data[0][13] (
	.clk(clk),
	.d(datain[13]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data013),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][13] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][13] .power_up = "low";

dffeas \register_fifo:fifo_data[0][12] (
	.clk(clk),
	.d(datain[12]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data012),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][12] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][12] .power_up = "low";

dffeas \register_fifo:fifo_data[0][11] (
	.clk(clk),
	.d(datain[11]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data011),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][11] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][11] .power_up = "low";

dffeas \register_fifo:fifo_data[0][10] (
	.clk(clk),
	.d(datain[10]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data010),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][10] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][10] .power_up = "low";

dffeas \register_fifo:fifo_data[0][9] (
	.clk(clk),
	.d(datain[9]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data09),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][9] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][9] .power_up = "low";

dffeas \register_fifo:fifo_data[0][8] (
	.clk(clk),
	.d(datain[8]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data08),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][8] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][8] .power_up = "low";

dffeas \register_fifo:fifo_data[0][7] (
	.clk(clk),
	.d(datain[7]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data07),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][7] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][7] .power_up = "low";

dffeas \register_fifo:fifo_data[0][6] (
	.clk(clk),
	.d(datain[6]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data06),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][6] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][6] .power_up = "low";

dffeas \register_fifo:fifo_data[0][5] (
	.clk(clk),
	.d(datain[5]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data05),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][5] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][5] .power_up = "low";

dffeas \register_fifo:fifo_data[0][4] (
	.clk(clk),
	.d(datain[4]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data04),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][4] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][4] .power_up = "low";

dffeas \register_fifo:fifo_data[0][3] (
	.clk(clk),
	.d(datain[3]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data03),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][3] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][3] .power_up = "low";

dffeas \register_fifo:fifo_data[0][2] (
	.clk(clk),
	.d(datain[2]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data02),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][2] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][2] .power_up = "low";

dffeas \register_fifo:fifo_data[0][1] (
	.clk(clk),
	.d(datain[1]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data01),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][1] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][1] .power_up = "low";

dffeas \register_fifo:fifo_data[0][0] (
	.clk(clk),
	.d(datain[0]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data00),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][0] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][0] .power_up = "low";

endmodule

module cic_auk_dspip_integrator_4 (
	stall_reg,
	register_fifofifo_data016,
	register_fifofifo_data017,
	register_fifofifo_data018,
	register_fifofifo_data019,
	register_fifofifo_data020,
	register_fifofifo_data021,
	register_fifofifo_data022,
	register_fifofifo_data023,
	register_fifofifo_data024,
	register_fifofifo_data025,
	register_fifofifo_data026,
	register_fifofifo_data027,
	register_fifofifo_data028,
	register_fifofifo_data029,
	register_fifofifo_data030,
	register_fifofifo_data031,
	register_fifofifo_data032,
	register_fifofifo_data033,
	register_fifofifo_data034,
	register_fifofifo_data035,
	register_fifofifo_data036,
	register_fifofifo_data037,
	register_fifofifo_data038,
	register_fifofifo_data039,
	register_fifofifo_data040,
	register_fifofifo_data041,
	register_fifofifo_data042,
	register_fifofifo_data043,
	register_fifofifo_data015,
	register_fifofifo_data0181,
	register_fifofifo_data014,
	register_fifofifo_data0191,
	register_fifofifo_data0201,
	register_fifofifo_data0211,
	register_fifofifo_data0221,
	register_fifofifo_data0231,
	register_fifofifo_data0241,
	register_fifofifo_data0251,
	register_fifofifo_data0261,
	register_fifofifo_data0271,
	register_fifofifo_data0281,
	register_fifofifo_data0291,
	register_fifofifo_data0301,
	register_fifofifo_data0311,
	register_fifofifo_data0321,
	register_fifofifo_data0331,
	register_fifofifo_data0341,
	register_fifofifo_data0351,
	register_fifofifo_data0361,
	register_fifofifo_data0371,
	register_fifofifo_data0381,
	register_fifofifo_data0391,
	register_fifofifo_data0401,
	register_fifofifo_data0411,
	register_fifofifo_data0421,
	register_fifofifo_data0431,
	register_fifofifo_data044,
	register_fifofifo_data045,
	register_fifofifo_data0171,
	register_fifofifo_data013,
	register_fifofifo_data0161,
	register_fifofifo_data012,
	register_fifofifo_data0151,
	register_fifofifo_data011,
	register_fifofifo_data0141,
	register_fifofifo_data010,
	register_fifofifo_data0131,
	register_fifofifo_data09,
	register_fifofifo_data0121,
	register_fifofifo_data08,
	register_fifofifo_data0111,
	register_fifofifo_data07,
	register_fifofifo_data0101,
	register_fifofifo_data06,
	register_fifofifo_data091,
	register_fifofifo_data05,
	register_fifofifo_data081,
	register_fifofifo_data04,
	register_fifofifo_data071,
	register_fifofifo_data03,
	register_fifofifo_data061,
	register_fifofifo_data02,
	register_fifofifo_data051,
	register_fifofifo_data046,
	register_fifofifo_data0310,
	register_fifofifo_data0210,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	stall_reg;
output 	register_fifofifo_data016;
output 	register_fifofifo_data017;
output 	register_fifofifo_data018;
output 	register_fifofifo_data019;
output 	register_fifofifo_data020;
output 	register_fifofifo_data021;
output 	register_fifofifo_data022;
output 	register_fifofifo_data023;
output 	register_fifofifo_data024;
output 	register_fifofifo_data025;
output 	register_fifofifo_data026;
output 	register_fifofifo_data027;
output 	register_fifofifo_data028;
output 	register_fifofifo_data029;
output 	register_fifofifo_data030;
output 	register_fifofifo_data031;
output 	register_fifofifo_data032;
output 	register_fifofifo_data033;
output 	register_fifofifo_data034;
output 	register_fifofifo_data035;
output 	register_fifofifo_data036;
output 	register_fifofifo_data037;
output 	register_fifofifo_data038;
output 	register_fifofifo_data039;
output 	register_fifofifo_data040;
output 	register_fifofifo_data041;
output 	register_fifofifo_data042;
output 	register_fifofifo_data043;
output 	register_fifofifo_data015;
input 	register_fifofifo_data0181;
output 	register_fifofifo_data014;
input 	register_fifofifo_data0191;
input 	register_fifofifo_data0201;
input 	register_fifofifo_data0211;
input 	register_fifofifo_data0221;
input 	register_fifofifo_data0231;
input 	register_fifofifo_data0241;
input 	register_fifofifo_data0251;
input 	register_fifofifo_data0261;
input 	register_fifofifo_data0271;
input 	register_fifofifo_data0281;
input 	register_fifofifo_data0291;
input 	register_fifofifo_data0301;
input 	register_fifofifo_data0311;
input 	register_fifofifo_data0321;
input 	register_fifofifo_data0331;
input 	register_fifofifo_data0341;
input 	register_fifofifo_data0351;
input 	register_fifofifo_data0361;
input 	register_fifofifo_data0371;
input 	register_fifofifo_data0381;
input 	register_fifofifo_data0391;
input 	register_fifofifo_data0401;
input 	register_fifofifo_data0411;
input 	register_fifofifo_data0421;
input 	register_fifofifo_data0431;
input 	register_fifofifo_data044;
input 	register_fifofifo_data045;
input 	register_fifofifo_data0171;
output 	register_fifofifo_data013;
input 	register_fifofifo_data0161;
output 	register_fifofifo_data012;
input 	register_fifofifo_data0151;
output 	register_fifofifo_data011;
input 	register_fifofifo_data0141;
output 	register_fifofifo_data010;
input 	register_fifofifo_data0131;
output 	register_fifofifo_data09;
input 	register_fifofifo_data0121;
output 	register_fifofifo_data08;
input 	register_fifofifo_data0111;
output 	register_fifofifo_data07;
input 	register_fifofifo_data0101;
output 	register_fifofifo_data06;
input 	register_fifofifo_data091;
output 	register_fifofifo_data05;
input 	register_fifofifo_data081;
output 	register_fifofifo_data04;
input 	register_fifofifo_data071;
output 	register_fifofifo_data03;
input 	register_fifofifo_data061;
output 	register_fifofifo_data02;
input 	register_fifofifo_data051;
input 	register_fifofifo_data046;
input 	register_fifofifo_data0310;
input 	register_fifofifo_data0210;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Add0~1_sumout ;
wire \Add0~2 ;
wire \Add0~5_sumout ;
wire \Add0~6 ;
wire \Add0~9_sumout ;
wire \Add0~10 ;
wire \Add0~13_sumout ;
wire \Add0~14 ;
wire \Add0~17_sumout ;
wire \Add0~18 ;
wire \Add0~21_sumout ;
wire \Add0~22 ;
wire \Add0~25_sumout ;
wire \Add0~26 ;
wire \Add0~29_sumout ;
wire \Add0~30 ;
wire \Add0~33_sumout ;
wire \Add0~34 ;
wire \Add0~37_sumout ;
wire \Add0~38 ;
wire \Add0~41_sumout ;
wire \Add0~42 ;
wire \Add0~45_sumout ;
wire \Add0~46 ;
wire \Add0~49_sumout ;
wire \Add0~50 ;
wire \Add0~53_sumout ;
wire \Add0~54 ;
wire \Add0~57_sumout ;
wire \Add0~58 ;
wire \Add0~61_sumout ;
wire \Add0~62 ;
wire \Add0~65_sumout ;
wire \Add0~66 ;
wire \Add0~69_sumout ;
wire \Add0~70 ;
wire \Add0~73_sumout ;
wire \Add0~74 ;
wire \Add0~77_sumout ;
wire \Add0~78 ;
wire \Add0~81_sumout ;
wire \Add0~82 ;
wire \Add0~85_sumout ;
wire \Add0~86 ;
wire \Add0~89_sumout ;
wire \Add0~90 ;
wire \Add0~93_sumout ;
wire \Add0~94 ;
wire \Add0~97_sumout ;
wire \Add0~98 ;
wire \Add0~101_sumout ;
wire \Add0~102 ;
wire \Add0~105_sumout ;
wire \Add0~106 ;
wire \Add0~109_sumout ;
wire \Add0~113_sumout ;
wire \Add0~114 ;
wire \Add0~117_sumout ;
wire \Add0~118 ;
wire \Add0~121_sumout ;
wire \Add0~122 ;
wire \Add0~125_sumout ;
wire \Add0~126 ;
wire \Add0~129_sumout ;
wire \Add0~130 ;
wire \Add0~133_sumout ;
wire \Add0~134 ;
wire \Add0~137_sumout ;
wire \Add0~138 ;
wire \Add0~141_sumout ;
wire \Add0~142 ;
wire \Add0~145_sumout ;
wire \Add0~146 ;
wire \Add0~149_sumout ;
wire \Add0~150 ;
wire \Add0~153_sumout ;
wire \Add0~154 ;
wire \Add0~157_sumout ;
wire \Add0~158 ;
wire \Add0~161_sumout ;
wire \Add0~162 ;
wire \Add0~165_sumout ;
wire \Add0~166 ;
wire \Add0~169_sumout ;
wire \Add0~170 ;
wire \Add0~173_sumout ;
wire \Add0~174 ;
wire \glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][1]~q ;
wire \glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][0]~q ;


cic_auk_dspip_delay_12 \glogic:integrator_pipeline_0_generate:u1 (
	.datain({gnd,gnd,gnd,\Add0~109_sumout ,\Add0~105_sumout ,\Add0~101_sumout ,\Add0~97_sumout ,\Add0~93_sumout ,\Add0~89_sumout ,\Add0~85_sumout ,\Add0~81_sumout ,\Add0~77_sumout ,\Add0~73_sumout ,\Add0~69_sumout ,\Add0~65_sumout ,\Add0~61_sumout ,\Add0~57_sumout ,\Add0~53_sumout ,
\Add0~49_sumout ,\Add0~45_sumout ,\Add0~41_sumout ,\Add0~37_sumout ,\Add0~33_sumout ,\Add0~29_sumout ,\Add0~25_sumout ,\Add0~21_sumout ,\Add0~17_sumout ,\Add0~13_sumout ,\Add0~9_sumout ,\Add0~5_sumout ,\Add0~1_sumout ,\Add0~113_sumout ,\Add0~117_sumout ,\Add0~121_sumout ,
\Add0~125_sumout ,\Add0~129_sumout ,\Add0~133_sumout ,\Add0~137_sumout ,\Add0~141_sumout ,\Add0~145_sumout ,\Add0~149_sumout ,\Add0~153_sumout ,\Add0~157_sumout ,\Add0~161_sumout ,\Add0~165_sumout ,\Add0~169_sumout ,\Add0~173_sumout }),
	.enable(stall_reg),
	.register_fifofifo_data016(register_fifofifo_data016),
	.register_fifofifo_data017(register_fifofifo_data017),
	.register_fifofifo_data018(register_fifofifo_data018),
	.register_fifofifo_data019(register_fifofifo_data019),
	.register_fifofifo_data020(register_fifofifo_data020),
	.register_fifofifo_data021(register_fifofifo_data021),
	.register_fifofifo_data022(register_fifofifo_data022),
	.register_fifofifo_data023(register_fifofifo_data023),
	.register_fifofifo_data024(register_fifofifo_data024),
	.register_fifofifo_data025(register_fifofifo_data025),
	.register_fifofifo_data026(register_fifofifo_data026),
	.register_fifofifo_data027(register_fifofifo_data027),
	.register_fifofifo_data028(register_fifofifo_data028),
	.register_fifofifo_data029(register_fifofifo_data029),
	.register_fifofifo_data030(register_fifofifo_data030),
	.register_fifofifo_data031(register_fifofifo_data031),
	.register_fifofifo_data032(register_fifofifo_data032),
	.register_fifofifo_data033(register_fifofifo_data033),
	.register_fifofifo_data034(register_fifofifo_data034),
	.register_fifofifo_data035(register_fifofifo_data035),
	.register_fifofifo_data036(register_fifofifo_data036),
	.register_fifofifo_data037(register_fifofifo_data037),
	.register_fifofifo_data038(register_fifofifo_data038),
	.register_fifofifo_data039(register_fifofifo_data039),
	.register_fifofifo_data040(register_fifofifo_data040),
	.register_fifofifo_data041(register_fifofifo_data041),
	.register_fifofifo_data042(register_fifofifo_data042),
	.register_fifofifo_data043(register_fifofifo_data043),
	.register_fifofifo_data015(register_fifofifo_data015),
	.register_fifofifo_data014(register_fifofifo_data014),
	.register_fifofifo_data013(register_fifofifo_data013),
	.register_fifofifo_data012(register_fifofifo_data012),
	.register_fifofifo_data011(register_fifofifo_data011),
	.register_fifofifo_data010(register_fifofifo_data010),
	.register_fifofifo_data09(register_fifofifo_data09),
	.register_fifofifo_data08(register_fifofifo_data08),
	.register_fifofifo_data07(register_fifofifo_data07),
	.register_fifofifo_data06(register_fifofifo_data06),
	.register_fifofifo_data05(register_fifofifo_data05),
	.register_fifofifo_data04(register_fifofifo_data04),
	.register_fifofifo_data03(register_fifofifo_data03),
	.register_fifofifo_data02(register_fifofifo_data02),
	.register_fifofifo_data01(\glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][1]~q ),
	.register_fifofifo_data00(\glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][0]~q ),
	.clk(clk),
	.reset(reset_n));

arriav_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data016),
	.datae(gnd),
	.dataf(!register_fifofifo_data0181),
	.datag(gnd),
	.cin(\Add0~114 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(\Add0~2 ),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~1 .shared_arith = "off";

arriav_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data017),
	.datae(gnd),
	.dataf(!register_fifofifo_data0191),
	.datag(gnd),
	.cin(\Add0~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~5 .shared_arith = "off";

arriav_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data018),
	.datae(gnd),
	.dataf(!register_fifofifo_data0201),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~9 .shared_arith = "off";

arriav_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data019),
	.datae(gnd),
	.dataf(!register_fifofifo_data0211),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~13 .shared_arith = "off";

arriav_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data020),
	.datae(gnd),
	.dataf(!register_fifofifo_data0221),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout());
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~17 .shared_arith = "off";

arriav_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data021),
	.datae(gnd),
	.dataf(!register_fifofifo_data0231),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout());
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~21 .shared_arith = "off";

arriav_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data022),
	.datae(gnd),
	.dataf(!register_fifofifo_data0241),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout());
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~25 .shared_arith = "off";

arriav_lcell_comb \Add0~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data023),
	.datae(gnd),
	.dataf(!register_fifofifo_data0251),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout());
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~29 .shared_arith = "off";

arriav_lcell_comb \Add0~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data024),
	.datae(gnd),
	.dataf(!register_fifofifo_data0261),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~33_sumout ),
	.cout(\Add0~34 ),
	.shareout());
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~33 .shared_arith = "off";

arriav_lcell_comb \Add0~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data025),
	.datae(gnd),
	.dataf(!register_fifofifo_data0271),
	.datag(gnd),
	.cin(\Add0~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~37_sumout ),
	.cout(\Add0~38 ),
	.shareout());
defparam \Add0~37 .extended_lut = "off";
defparam \Add0~37 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~37 .shared_arith = "off";

arriav_lcell_comb \Add0~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data026),
	.datae(gnd),
	.dataf(!register_fifofifo_data0281),
	.datag(gnd),
	.cin(\Add0~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~41_sumout ),
	.cout(\Add0~42 ),
	.shareout());
defparam \Add0~41 .extended_lut = "off";
defparam \Add0~41 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~41 .shared_arith = "off";

arriav_lcell_comb \Add0~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data027),
	.datae(gnd),
	.dataf(!register_fifofifo_data0291),
	.datag(gnd),
	.cin(\Add0~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~45_sumout ),
	.cout(\Add0~46 ),
	.shareout());
defparam \Add0~45 .extended_lut = "off";
defparam \Add0~45 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~45 .shared_arith = "off";

arriav_lcell_comb \Add0~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data028),
	.datae(gnd),
	.dataf(!register_fifofifo_data0301),
	.datag(gnd),
	.cin(\Add0~46 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~49_sumout ),
	.cout(\Add0~50 ),
	.shareout());
defparam \Add0~49 .extended_lut = "off";
defparam \Add0~49 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~49 .shared_arith = "off";

arriav_lcell_comb \Add0~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data029),
	.datae(gnd),
	.dataf(!register_fifofifo_data0311),
	.datag(gnd),
	.cin(\Add0~50 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~53_sumout ),
	.cout(\Add0~54 ),
	.shareout());
defparam \Add0~53 .extended_lut = "off";
defparam \Add0~53 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~53 .shared_arith = "off";

arriav_lcell_comb \Add0~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data030),
	.datae(gnd),
	.dataf(!register_fifofifo_data0321),
	.datag(gnd),
	.cin(\Add0~54 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~57_sumout ),
	.cout(\Add0~58 ),
	.shareout());
defparam \Add0~57 .extended_lut = "off";
defparam \Add0~57 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~57 .shared_arith = "off";

arriav_lcell_comb \Add0~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data031),
	.datae(gnd),
	.dataf(!register_fifofifo_data0331),
	.datag(gnd),
	.cin(\Add0~58 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~61_sumout ),
	.cout(\Add0~62 ),
	.shareout());
defparam \Add0~61 .extended_lut = "off";
defparam \Add0~61 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~61 .shared_arith = "off";

arriav_lcell_comb \Add0~65 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data032),
	.datae(gnd),
	.dataf(!register_fifofifo_data0341),
	.datag(gnd),
	.cin(\Add0~62 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~65_sumout ),
	.cout(\Add0~66 ),
	.shareout());
defparam \Add0~65 .extended_lut = "off";
defparam \Add0~65 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~65 .shared_arith = "off";

arriav_lcell_comb \Add0~69 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data033),
	.datae(gnd),
	.dataf(!register_fifofifo_data0351),
	.datag(gnd),
	.cin(\Add0~66 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~69_sumout ),
	.cout(\Add0~70 ),
	.shareout());
defparam \Add0~69 .extended_lut = "off";
defparam \Add0~69 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~69 .shared_arith = "off";

arriav_lcell_comb \Add0~73 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data034),
	.datae(gnd),
	.dataf(!register_fifofifo_data0361),
	.datag(gnd),
	.cin(\Add0~70 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~73_sumout ),
	.cout(\Add0~74 ),
	.shareout());
defparam \Add0~73 .extended_lut = "off";
defparam \Add0~73 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~73 .shared_arith = "off";

arriav_lcell_comb \Add0~77 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data035),
	.datae(gnd),
	.dataf(!register_fifofifo_data0371),
	.datag(gnd),
	.cin(\Add0~74 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~77_sumout ),
	.cout(\Add0~78 ),
	.shareout());
defparam \Add0~77 .extended_lut = "off";
defparam \Add0~77 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~77 .shared_arith = "off";

arriav_lcell_comb \Add0~81 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data036),
	.datae(gnd),
	.dataf(!register_fifofifo_data0381),
	.datag(gnd),
	.cin(\Add0~78 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~81_sumout ),
	.cout(\Add0~82 ),
	.shareout());
defparam \Add0~81 .extended_lut = "off";
defparam \Add0~81 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~81 .shared_arith = "off";

arriav_lcell_comb \Add0~85 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data037),
	.datae(gnd),
	.dataf(!register_fifofifo_data0391),
	.datag(gnd),
	.cin(\Add0~82 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~85_sumout ),
	.cout(\Add0~86 ),
	.shareout());
defparam \Add0~85 .extended_lut = "off";
defparam \Add0~85 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~85 .shared_arith = "off";

arriav_lcell_comb \Add0~89 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data038),
	.datae(gnd),
	.dataf(!register_fifofifo_data0401),
	.datag(gnd),
	.cin(\Add0~86 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~89_sumout ),
	.cout(\Add0~90 ),
	.shareout());
defparam \Add0~89 .extended_lut = "off";
defparam \Add0~89 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~89 .shared_arith = "off";

arriav_lcell_comb \Add0~93 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data039),
	.datae(gnd),
	.dataf(!register_fifofifo_data0411),
	.datag(gnd),
	.cin(\Add0~90 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~93_sumout ),
	.cout(\Add0~94 ),
	.shareout());
defparam \Add0~93 .extended_lut = "off";
defparam \Add0~93 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~93 .shared_arith = "off";

arriav_lcell_comb \Add0~97 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data040),
	.datae(gnd),
	.dataf(!register_fifofifo_data0421),
	.datag(gnd),
	.cin(\Add0~94 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~97_sumout ),
	.cout(\Add0~98 ),
	.shareout());
defparam \Add0~97 .extended_lut = "off";
defparam \Add0~97 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~97 .shared_arith = "off";

arriav_lcell_comb \Add0~101 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data041),
	.datae(gnd),
	.dataf(!register_fifofifo_data0431),
	.datag(gnd),
	.cin(\Add0~98 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~101_sumout ),
	.cout(\Add0~102 ),
	.shareout());
defparam \Add0~101 .extended_lut = "off";
defparam \Add0~101 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~101 .shared_arith = "off";

arriav_lcell_comb \Add0~105 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data042),
	.datae(gnd),
	.dataf(!register_fifofifo_data044),
	.datag(gnd),
	.cin(\Add0~102 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~105_sumout ),
	.cout(\Add0~106 ),
	.shareout());
defparam \Add0~105 .extended_lut = "off";
defparam \Add0~105 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~105 .shared_arith = "off";

arriav_lcell_comb \Add0~109 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data043),
	.datae(gnd),
	.dataf(!register_fifofifo_data045),
	.datag(gnd),
	.cin(\Add0~106 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~109_sumout ),
	.cout(),
	.shareout());
defparam \Add0~109 .extended_lut = "off";
defparam \Add0~109 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~109 .shared_arith = "off";

arriav_lcell_comb \Add0~113 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data015),
	.datae(gnd),
	.dataf(!register_fifofifo_data0171),
	.datag(gnd),
	.cin(\Add0~118 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~113_sumout ),
	.cout(\Add0~114 ),
	.shareout());
defparam \Add0~113 .extended_lut = "off";
defparam \Add0~113 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~113 .shared_arith = "off";

arriav_lcell_comb \Add0~117 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data014),
	.datae(gnd),
	.dataf(!register_fifofifo_data0161),
	.datag(gnd),
	.cin(\Add0~122 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~117_sumout ),
	.cout(\Add0~118 ),
	.shareout());
defparam \Add0~117 .extended_lut = "off";
defparam \Add0~117 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~117 .shared_arith = "off";

arriav_lcell_comb \Add0~121 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data013),
	.datae(gnd),
	.dataf(!register_fifofifo_data0151),
	.datag(gnd),
	.cin(\Add0~126 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~121_sumout ),
	.cout(\Add0~122 ),
	.shareout());
defparam \Add0~121 .extended_lut = "off";
defparam \Add0~121 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~121 .shared_arith = "off";

arriav_lcell_comb \Add0~125 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data012),
	.datae(gnd),
	.dataf(!register_fifofifo_data0141),
	.datag(gnd),
	.cin(\Add0~130 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~125_sumout ),
	.cout(\Add0~126 ),
	.shareout());
defparam \Add0~125 .extended_lut = "off";
defparam \Add0~125 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~125 .shared_arith = "off";

arriav_lcell_comb \Add0~129 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data011),
	.datae(gnd),
	.dataf(!register_fifofifo_data0131),
	.datag(gnd),
	.cin(\Add0~134 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~129_sumout ),
	.cout(\Add0~130 ),
	.shareout());
defparam \Add0~129 .extended_lut = "off";
defparam \Add0~129 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~129 .shared_arith = "off";

arriav_lcell_comb \Add0~133 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data010),
	.datae(gnd),
	.dataf(!register_fifofifo_data0121),
	.datag(gnd),
	.cin(\Add0~138 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~133_sumout ),
	.cout(\Add0~134 ),
	.shareout());
defparam \Add0~133 .extended_lut = "off";
defparam \Add0~133 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~133 .shared_arith = "off";

arriav_lcell_comb \Add0~137 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data09),
	.datae(gnd),
	.dataf(!register_fifofifo_data0111),
	.datag(gnd),
	.cin(\Add0~142 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~137_sumout ),
	.cout(\Add0~138 ),
	.shareout());
defparam \Add0~137 .extended_lut = "off";
defparam \Add0~137 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~137 .shared_arith = "off";

arriav_lcell_comb \Add0~141 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data08),
	.datae(gnd),
	.dataf(!register_fifofifo_data0101),
	.datag(gnd),
	.cin(\Add0~146 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~141_sumout ),
	.cout(\Add0~142 ),
	.shareout());
defparam \Add0~141 .extended_lut = "off";
defparam \Add0~141 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~141 .shared_arith = "off";

arriav_lcell_comb \Add0~145 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data07),
	.datae(gnd),
	.dataf(!register_fifofifo_data091),
	.datag(gnd),
	.cin(\Add0~150 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~145_sumout ),
	.cout(\Add0~146 ),
	.shareout());
defparam \Add0~145 .extended_lut = "off";
defparam \Add0~145 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~145 .shared_arith = "off";

arriav_lcell_comb \Add0~149 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data06),
	.datae(gnd),
	.dataf(!register_fifofifo_data081),
	.datag(gnd),
	.cin(\Add0~154 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~149_sumout ),
	.cout(\Add0~150 ),
	.shareout());
defparam \Add0~149 .extended_lut = "off";
defparam \Add0~149 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~149 .shared_arith = "off";

arriav_lcell_comb \Add0~153 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data05),
	.datae(gnd),
	.dataf(!register_fifofifo_data071),
	.datag(gnd),
	.cin(\Add0~158 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~153_sumout ),
	.cout(\Add0~154 ),
	.shareout());
defparam \Add0~153 .extended_lut = "off";
defparam \Add0~153 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~153 .shared_arith = "off";

arriav_lcell_comb \Add0~157 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data04),
	.datae(gnd),
	.dataf(!register_fifofifo_data061),
	.datag(gnd),
	.cin(\Add0~162 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~157_sumout ),
	.cout(\Add0~158 ),
	.shareout());
defparam \Add0~157 .extended_lut = "off";
defparam \Add0~157 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~157 .shared_arith = "off";

arriav_lcell_comb \Add0~161 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data03),
	.datae(gnd),
	.dataf(!register_fifofifo_data051),
	.datag(gnd),
	.cin(\Add0~166 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~161_sumout ),
	.cout(\Add0~162 ),
	.shareout());
defparam \Add0~161 .extended_lut = "off";
defparam \Add0~161 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~161 .shared_arith = "off";

arriav_lcell_comb \Add0~165 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data02),
	.datae(gnd),
	.dataf(!register_fifofifo_data046),
	.datag(gnd),
	.cin(\Add0~170 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~165_sumout ),
	.cout(\Add0~166 ),
	.shareout());
defparam \Add0~165 .extended_lut = "off";
defparam \Add0~165 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~165 .shared_arith = "off";

arriav_lcell_comb \Add0~169 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][1]~q ),
	.datae(gnd),
	.dataf(!register_fifofifo_data0310),
	.datag(gnd),
	.cin(\Add0~174 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~169_sumout ),
	.cout(\Add0~170 ),
	.shareout());
defparam \Add0~169 .extended_lut = "off";
defparam \Add0~169 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~169 .shared_arith = "off";

arriav_lcell_comb \Add0~173 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][0]~q ),
	.datae(gnd),
	.dataf(!register_fifofifo_data0210),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~173_sumout ),
	.cout(\Add0~174 ),
	.shareout());
defparam \Add0~173 .extended_lut = "off";
defparam \Add0~173 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~173 .shared_arith = "off";

endmodule

module cic_auk_dspip_delay_12 (
	datain,
	enable,
	register_fifofifo_data016,
	register_fifofifo_data017,
	register_fifofifo_data018,
	register_fifofifo_data019,
	register_fifofifo_data020,
	register_fifofifo_data021,
	register_fifofifo_data022,
	register_fifofifo_data023,
	register_fifofifo_data024,
	register_fifofifo_data025,
	register_fifofifo_data026,
	register_fifofifo_data027,
	register_fifofifo_data028,
	register_fifofifo_data029,
	register_fifofifo_data030,
	register_fifofifo_data031,
	register_fifofifo_data032,
	register_fifofifo_data033,
	register_fifofifo_data034,
	register_fifofifo_data035,
	register_fifofifo_data036,
	register_fifofifo_data037,
	register_fifofifo_data038,
	register_fifofifo_data039,
	register_fifofifo_data040,
	register_fifofifo_data041,
	register_fifofifo_data042,
	register_fifofifo_data043,
	register_fifofifo_data015,
	register_fifofifo_data014,
	register_fifofifo_data013,
	register_fifofifo_data012,
	register_fifofifo_data011,
	register_fifofifo_data010,
	register_fifofifo_data09,
	register_fifofifo_data08,
	register_fifofifo_data07,
	register_fifofifo_data06,
	register_fifofifo_data05,
	register_fifofifo_data04,
	register_fifofifo_data03,
	register_fifofifo_data02,
	register_fifofifo_data01,
	register_fifofifo_data00,
	clk,
	reset)/* synthesis synthesis_greybox=1 */;
input 	[46:0] datain;
input 	enable;
output 	register_fifofifo_data016;
output 	register_fifofifo_data017;
output 	register_fifofifo_data018;
output 	register_fifofifo_data019;
output 	register_fifofifo_data020;
output 	register_fifofifo_data021;
output 	register_fifofifo_data022;
output 	register_fifofifo_data023;
output 	register_fifofifo_data024;
output 	register_fifofifo_data025;
output 	register_fifofifo_data026;
output 	register_fifofifo_data027;
output 	register_fifofifo_data028;
output 	register_fifofifo_data029;
output 	register_fifofifo_data030;
output 	register_fifofifo_data031;
output 	register_fifofifo_data032;
output 	register_fifofifo_data033;
output 	register_fifofifo_data034;
output 	register_fifofifo_data035;
output 	register_fifofifo_data036;
output 	register_fifofifo_data037;
output 	register_fifofifo_data038;
output 	register_fifofifo_data039;
output 	register_fifofifo_data040;
output 	register_fifofifo_data041;
output 	register_fifofifo_data042;
output 	register_fifofifo_data043;
output 	register_fifofifo_data015;
output 	register_fifofifo_data014;
output 	register_fifofifo_data013;
output 	register_fifofifo_data012;
output 	register_fifofifo_data011;
output 	register_fifofifo_data010;
output 	register_fifofifo_data09;
output 	register_fifofifo_data08;
output 	register_fifofifo_data07;
output 	register_fifofifo_data06;
output 	register_fifofifo_data05;
output 	register_fifofifo_data04;
output 	register_fifofifo_data03;
output 	register_fifofifo_data02;
output 	register_fifofifo_data01;
output 	register_fifofifo_data00;
input 	clk;
input 	reset;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \register_fifo:fifo_data[0][16] (
	.clk(clk),
	.d(datain[16]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data016),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][16] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][16] .power_up = "low";

dffeas \register_fifo:fifo_data[0][17] (
	.clk(clk),
	.d(datain[17]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data017),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][17] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][17] .power_up = "low";

dffeas \register_fifo:fifo_data[0][18] (
	.clk(clk),
	.d(datain[18]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data018),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][18] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][18] .power_up = "low";

dffeas \register_fifo:fifo_data[0][19] (
	.clk(clk),
	.d(datain[19]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data019),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][19] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][19] .power_up = "low";

dffeas \register_fifo:fifo_data[0][20] (
	.clk(clk),
	.d(datain[20]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data020),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][20] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][20] .power_up = "low";

dffeas \register_fifo:fifo_data[0][21] (
	.clk(clk),
	.d(datain[21]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data021),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][21] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][21] .power_up = "low";

dffeas \register_fifo:fifo_data[0][22] (
	.clk(clk),
	.d(datain[22]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data022),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][22] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][22] .power_up = "low";

dffeas \register_fifo:fifo_data[0][23] (
	.clk(clk),
	.d(datain[23]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data023),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][23] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][23] .power_up = "low";

dffeas \register_fifo:fifo_data[0][24] (
	.clk(clk),
	.d(datain[24]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data024),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][24] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][24] .power_up = "low";

dffeas \register_fifo:fifo_data[0][25] (
	.clk(clk),
	.d(datain[25]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data025),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][25] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][25] .power_up = "low";

dffeas \register_fifo:fifo_data[0][26] (
	.clk(clk),
	.d(datain[26]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data026),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][26] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][26] .power_up = "low";

dffeas \register_fifo:fifo_data[0][27] (
	.clk(clk),
	.d(datain[27]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data027),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][27] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][27] .power_up = "low";

dffeas \register_fifo:fifo_data[0][28] (
	.clk(clk),
	.d(datain[28]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data028),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][28] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][28] .power_up = "low";

dffeas \register_fifo:fifo_data[0][29] (
	.clk(clk),
	.d(datain[29]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data029),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][29] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][29] .power_up = "low";

dffeas \register_fifo:fifo_data[0][30] (
	.clk(clk),
	.d(datain[30]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data030),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][30] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][30] .power_up = "low";

dffeas \register_fifo:fifo_data[0][31] (
	.clk(clk),
	.d(datain[31]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data031),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][31] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][31] .power_up = "low";

dffeas \register_fifo:fifo_data[0][32] (
	.clk(clk),
	.d(datain[32]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data032),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][32] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][32] .power_up = "low";

dffeas \register_fifo:fifo_data[0][33] (
	.clk(clk),
	.d(datain[33]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data033),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][33] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][33] .power_up = "low";

dffeas \register_fifo:fifo_data[0][34] (
	.clk(clk),
	.d(datain[34]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data034),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][34] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][34] .power_up = "low";

dffeas \register_fifo:fifo_data[0][35] (
	.clk(clk),
	.d(datain[35]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data035),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][35] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][35] .power_up = "low";

dffeas \register_fifo:fifo_data[0][36] (
	.clk(clk),
	.d(datain[36]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data036),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][36] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][36] .power_up = "low";

dffeas \register_fifo:fifo_data[0][37] (
	.clk(clk),
	.d(datain[37]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data037),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][37] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][37] .power_up = "low";

dffeas \register_fifo:fifo_data[0][38] (
	.clk(clk),
	.d(datain[38]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data038),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][38] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][38] .power_up = "low";

dffeas \register_fifo:fifo_data[0][39] (
	.clk(clk),
	.d(datain[39]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data039),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][39] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][39] .power_up = "low";

dffeas \register_fifo:fifo_data[0][40] (
	.clk(clk),
	.d(datain[40]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data040),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][40] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][40] .power_up = "low";

dffeas \register_fifo:fifo_data[0][41] (
	.clk(clk),
	.d(datain[41]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data041),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][41] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][41] .power_up = "low";

dffeas \register_fifo:fifo_data[0][42] (
	.clk(clk),
	.d(datain[42]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data042),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][42] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][42] .power_up = "low";

dffeas \register_fifo:fifo_data[0][43] (
	.clk(clk),
	.d(datain[43]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data043),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][43] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][43] .power_up = "low";

dffeas \register_fifo:fifo_data[0][15] (
	.clk(clk),
	.d(datain[15]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data015),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][15] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][15] .power_up = "low";

dffeas \register_fifo:fifo_data[0][14] (
	.clk(clk),
	.d(datain[14]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data014),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][14] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][14] .power_up = "low";

dffeas \register_fifo:fifo_data[0][13] (
	.clk(clk),
	.d(datain[13]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data013),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][13] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][13] .power_up = "low";

dffeas \register_fifo:fifo_data[0][12] (
	.clk(clk),
	.d(datain[12]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data012),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][12] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][12] .power_up = "low";

dffeas \register_fifo:fifo_data[0][11] (
	.clk(clk),
	.d(datain[11]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data011),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][11] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][11] .power_up = "low";

dffeas \register_fifo:fifo_data[0][10] (
	.clk(clk),
	.d(datain[10]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data010),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][10] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][10] .power_up = "low";

dffeas \register_fifo:fifo_data[0][9] (
	.clk(clk),
	.d(datain[9]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data09),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][9] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][9] .power_up = "low";

dffeas \register_fifo:fifo_data[0][8] (
	.clk(clk),
	.d(datain[8]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data08),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][8] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][8] .power_up = "low";

dffeas \register_fifo:fifo_data[0][7] (
	.clk(clk),
	.d(datain[7]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data07),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][7] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][7] .power_up = "low";

dffeas \register_fifo:fifo_data[0][6] (
	.clk(clk),
	.d(datain[6]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data06),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][6] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][6] .power_up = "low";

dffeas \register_fifo:fifo_data[0][5] (
	.clk(clk),
	.d(datain[5]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data05),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][5] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][5] .power_up = "low";

dffeas \register_fifo:fifo_data[0][4] (
	.clk(clk),
	.d(datain[4]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data04),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][4] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][4] .power_up = "low";

dffeas \register_fifo:fifo_data[0][3] (
	.clk(clk),
	.d(datain[3]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data03),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][3] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][3] .power_up = "low";

dffeas \register_fifo:fifo_data[0][2] (
	.clk(clk),
	.d(datain[2]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data02),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][2] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][2] .power_up = "low";

dffeas \register_fifo:fifo_data[0][1] (
	.clk(clk),
	.d(datain[1]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data01),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][1] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][1] .power_up = "low";

dffeas \register_fifo:fifo_data[0][0] (
	.clk(clk),
	.d(datain[0]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data00),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][0] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][0] .power_up = "low";

endmodule

module cic_auk_dspip_integrator_5 (
	stall_reg,
	register_fifofifo_data014,
	register_fifofifo_data015,
	register_fifofifo_data016,
	register_fifofifo_data017,
	register_fifofifo_data018,
	register_fifofifo_data019,
	register_fifofifo_data020,
	register_fifofifo_data021,
	register_fifofifo_data022,
	register_fifofifo_data023,
	register_fifofifo_data024,
	register_fifofifo_data025,
	register_fifofifo_data026,
	register_fifofifo_data027,
	register_fifofifo_data028,
	register_fifofifo_data029,
	register_fifofifo_data030,
	register_fifofifo_data031,
	register_fifofifo_data032,
	register_fifofifo_data033,
	register_fifofifo_data034,
	register_fifofifo_data035,
	register_fifofifo_data036,
	register_fifofifo_data037,
	register_fifofifo_data038,
	register_fifofifo_data039,
	register_fifofifo_data040,
	register_fifofifo_data041,
	register_fifofifo_data013,
	register_fifofifo_data0161,
	register_fifofifo_data012,
	register_fifofifo_data0171,
	register_fifofifo_data0181,
	register_fifofifo_data0191,
	register_fifofifo_data0201,
	register_fifofifo_data0211,
	register_fifofifo_data0221,
	register_fifofifo_data0231,
	register_fifofifo_data0241,
	register_fifofifo_data0251,
	register_fifofifo_data0261,
	register_fifofifo_data0271,
	register_fifofifo_data0281,
	register_fifofifo_data0291,
	register_fifofifo_data0301,
	register_fifofifo_data0311,
	register_fifofifo_data0321,
	register_fifofifo_data0331,
	register_fifofifo_data0341,
	register_fifofifo_data0351,
	register_fifofifo_data0361,
	register_fifofifo_data0371,
	register_fifofifo_data0381,
	register_fifofifo_data0391,
	register_fifofifo_data0401,
	register_fifofifo_data0411,
	register_fifofifo_data042,
	register_fifofifo_data043,
	register_fifofifo_data0151,
	register_fifofifo_data011,
	register_fifofifo_data0141,
	register_fifofifo_data010,
	register_fifofifo_data0131,
	register_fifofifo_data09,
	register_fifofifo_data0121,
	register_fifofifo_data08,
	register_fifofifo_data0111,
	register_fifofifo_data07,
	register_fifofifo_data0101,
	register_fifofifo_data06,
	register_fifofifo_data091,
	register_fifofifo_data05,
	register_fifofifo_data081,
	register_fifofifo_data04,
	register_fifofifo_data071,
	register_fifofifo_data03,
	register_fifofifo_data061,
	register_fifofifo_data02,
	register_fifofifo_data051,
	register_fifofifo_data044,
	register_fifofifo_data0310,
	register_fifofifo_data0210,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	stall_reg;
output 	register_fifofifo_data014;
output 	register_fifofifo_data015;
output 	register_fifofifo_data016;
output 	register_fifofifo_data017;
output 	register_fifofifo_data018;
output 	register_fifofifo_data019;
output 	register_fifofifo_data020;
output 	register_fifofifo_data021;
output 	register_fifofifo_data022;
output 	register_fifofifo_data023;
output 	register_fifofifo_data024;
output 	register_fifofifo_data025;
output 	register_fifofifo_data026;
output 	register_fifofifo_data027;
output 	register_fifofifo_data028;
output 	register_fifofifo_data029;
output 	register_fifofifo_data030;
output 	register_fifofifo_data031;
output 	register_fifofifo_data032;
output 	register_fifofifo_data033;
output 	register_fifofifo_data034;
output 	register_fifofifo_data035;
output 	register_fifofifo_data036;
output 	register_fifofifo_data037;
output 	register_fifofifo_data038;
output 	register_fifofifo_data039;
output 	register_fifofifo_data040;
output 	register_fifofifo_data041;
output 	register_fifofifo_data013;
input 	register_fifofifo_data0161;
output 	register_fifofifo_data012;
input 	register_fifofifo_data0171;
input 	register_fifofifo_data0181;
input 	register_fifofifo_data0191;
input 	register_fifofifo_data0201;
input 	register_fifofifo_data0211;
input 	register_fifofifo_data0221;
input 	register_fifofifo_data0231;
input 	register_fifofifo_data0241;
input 	register_fifofifo_data0251;
input 	register_fifofifo_data0261;
input 	register_fifofifo_data0271;
input 	register_fifofifo_data0281;
input 	register_fifofifo_data0291;
input 	register_fifofifo_data0301;
input 	register_fifofifo_data0311;
input 	register_fifofifo_data0321;
input 	register_fifofifo_data0331;
input 	register_fifofifo_data0341;
input 	register_fifofifo_data0351;
input 	register_fifofifo_data0361;
input 	register_fifofifo_data0371;
input 	register_fifofifo_data0381;
input 	register_fifofifo_data0391;
input 	register_fifofifo_data0401;
input 	register_fifofifo_data0411;
input 	register_fifofifo_data042;
input 	register_fifofifo_data043;
input 	register_fifofifo_data0151;
output 	register_fifofifo_data011;
input 	register_fifofifo_data0141;
output 	register_fifofifo_data010;
input 	register_fifofifo_data0131;
output 	register_fifofifo_data09;
input 	register_fifofifo_data0121;
output 	register_fifofifo_data08;
input 	register_fifofifo_data0111;
output 	register_fifofifo_data07;
input 	register_fifofifo_data0101;
output 	register_fifofifo_data06;
input 	register_fifofifo_data091;
output 	register_fifofifo_data05;
input 	register_fifofifo_data081;
output 	register_fifofifo_data04;
input 	register_fifofifo_data071;
output 	register_fifofifo_data03;
input 	register_fifofifo_data061;
output 	register_fifofifo_data02;
input 	register_fifofifo_data051;
input 	register_fifofifo_data044;
input 	register_fifofifo_data0310;
input 	register_fifofifo_data0210;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Add0~1_sumout ;
wire \Add0~2 ;
wire \Add0~5_sumout ;
wire \Add0~6 ;
wire \Add0~9_sumout ;
wire \Add0~10 ;
wire \Add0~13_sumout ;
wire \Add0~14 ;
wire \Add0~17_sumout ;
wire \Add0~18 ;
wire \Add0~21_sumout ;
wire \Add0~22 ;
wire \Add0~25_sumout ;
wire \Add0~26 ;
wire \Add0~29_sumout ;
wire \Add0~30 ;
wire \Add0~33_sumout ;
wire \Add0~34 ;
wire \Add0~37_sumout ;
wire \Add0~38 ;
wire \Add0~41_sumout ;
wire \Add0~42 ;
wire \Add0~45_sumout ;
wire \Add0~46 ;
wire \Add0~49_sumout ;
wire \Add0~50 ;
wire \Add0~53_sumout ;
wire \Add0~54 ;
wire \Add0~57_sumout ;
wire \Add0~58 ;
wire \Add0~61_sumout ;
wire \Add0~62 ;
wire \Add0~65_sumout ;
wire \Add0~66 ;
wire \Add0~69_sumout ;
wire \Add0~70 ;
wire \Add0~73_sumout ;
wire \Add0~74 ;
wire \Add0~77_sumout ;
wire \Add0~78 ;
wire \Add0~81_sumout ;
wire \Add0~82 ;
wire \Add0~85_sumout ;
wire \Add0~86 ;
wire \Add0~89_sumout ;
wire \Add0~90 ;
wire \Add0~93_sumout ;
wire \Add0~94 ;
wire \Add0~97_sumout ;
wire \Add0~98 ;
wire \Add0~101_sumout ;
wire \Add0~102 ;
wire \Add0~105_sumout ;
wire \Add0~106 ;
wire \Add0~109_sumout ;
wire \Add0~113_sumout ;
wire \Add0~114 ;
wire \Add0~117_sumout ;
wire \Add0~118 ;
wire \Add0~121_sumout ;
wire \Add0~122 ;
wire \Add0~125_sumout ;
wire \Add0~126 ;
wire \Add0~129_sumout ;
wire \Add0~130 ;
wire \Add0~133_sumout ;
wire \Add0~134 ;
wire \Add0~137_sumout ;
wire \Add0~138 ;
wire \Add0~141_sumout ;
wire \Add0~142 ;
wire \Add0~145_sumout ;
wire \Add0~146 ;
wire \Add0~149_sumout ;
wire \Add0~150 ;
wire \Add0~153_sumout ;
wire \Add0~154 ;
wire \Add0~157_sumout ;
wire \Add0~158 ;
wire \Add0~161_sumout ;
wire \Add0~162 ;
wire \Add0~165_sumout ;
wire \Add0~166 ;
wire \glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][1]~q ;
wire \glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][0]~q ;


cic_auk_dspip_delay_13 \glogic:integrator_pipeline_0_generate:u1 (
	.datain({gnd,gnd,gnd,gnd,gnd,\Add0~109_sumout ,\Add0~105_sumout ,\Add0~101_sumout ,\Add0~97_sumout ,\Add0~93_sumout ,\Add0~89_sumout ,\Add0~85_sumout ,\Add0~81_sumout ,\Add0~77_sumout ,\Add0~73_sumout ,\Add0~69_sumout ,\Add0~65_sumout ,\Add0~61_sumout ,\Add0~57_sumout ,
\Add0~53_sumout ,\Add0~49_sumout ,\Add0~45_sumout ,\Add0~41_sumout ,\Add0~37_sumout ,\Add0~33_sumout ,\Add0~29_sumout ,\Add0~25_sumout ,\Add0~21_sumout ,\Add0~17_sumout ,\Add0~13_sumout ,\Add0~9_sumout ,\Add0~5_sumout ,\Add0~1_sumout ,\Add0~113_sumout ,\Add0~117_sumout ,
\Add0~121_sumout ,\Add0~125_sumout ,\Add0~129_sumout ,\Add0~133_sumout ,\Add0~137_sumout ,\Add0~141_sumout ,\Add0~145_sumout ,\Add0~149_sumout ,\Add0~153_sumout ,\Add0~157_sumout ,\Add0~161_sumout ,\Add0~165_sumout }),
	.enable(stall_reg),
	.register_fifofifo_data014(register_fifofifo_data014),
	.register_fifofifo_data015(register_fifofifo_data015),
	.register_fifofifo_data016(register_fifofifo_data016),
	.register_fifofifo_data017(register_fifofifo_data017),
	.register_fifofifo_data018(register_fifofifo_data018),
	.register_fifofifo_data019(register_fifofifo_data019),
	.register_fifofifo_data020(register_fifofifo_data020),
	.register_fifofifo_data021(register_fifofifo_data021),
	.register_fifofifo_data022(register_fifofifo_data022),
	.register_fifofifo_data023(register_fifofifo_data023),
	.register_fifofifo_data024(register_fifofifo_data024),
	.register_fifofifo_data025(register_fifofifo_data025),
	.register_fifofifo_data026(register_fifofifo_data026),
	.register_fifofifo_data027(register_fifofifo_data027),
	.register_fifofifo_data028(register_fifofifo_data028),
	.register_fifofifo_data029(register_fifofifo_data029),
	.register_fifofifo_data030(register_fifofifo_data030),
	.register_fifofifo_data031(register_fifofifo_data031),
	.register_fifofifo_data032(register_fifofifo_data032),
	.register_fifofifo_data033(register_fifofifo_data033),
	.register_fifofifo_data034(register_fifofifo_data034),
	.register_fifofifo_data035(register_fifofifo_data035),
	.register_fifofifo_data036(register_fifofifo_data036),
	.register_fifofifo_data037(register_fifofifo_data037),
	.register_fifofifo_data038(register_fifofifo_data038),
	.register_fifofifo_data039(register_fifofifo_data039),
	.register_fifofifo_data040(register_fifofifo_data040),
	.register_fifofifo_data041(register_fifofifo_data041),
	.register_fifofifo_data013(register_fifofifo_data013),
	.register_fifofifo_data012(register_fifofifo_data012),
	.register_fifofifo_data011(register_fifofifo_data011),
	.register_fifofifo_data010(register_fifofifo_data010),
	.register_fifofifo_data09(register_fifofifo_data09),
	.register_fifofifo_data08(register_fifofifo_data08),
	.register_fifofifo_data07(register_fifofifo_data07),
	.register_fifofifo_data06(register_fifofifo_data06),
	.register_fifofifo_data05(register_fifofifo_data05),
	.register_fifofifo_data04(register_fifofifo_data04),
	.register_fifofifo_data03(register_fifofifo_data03),
	.register_fifofifo_data02(register_fifofifo_data02),
	.register_fifofifo_data01(\glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][1]~q ),
	.register_fifofifo_data00(\glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][0]~q ),
	.clk(clk),
	.reset(reset_n));

arriav_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data014),
	.datae(gnd),
	.dataf(!register_fifofifo_data0161),
	.datag(gnd),
	.cin(\Add0~114 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(\Add0~2 ),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~1 .shared_arith = "off";

arriav_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data015),
	.datae(gnd),
	.dataf(!register_fifofifo_data0171),
	.datag(gnd),
	.cin(\Add0~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~5 .shared_arith = "off";

arriav_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data016),
	.datae(gnd),
	.dataf(!register_fifofifo_data0181),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~9 .shared_arith = "off";

arriav_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data017),
	.datae(gnd),
	.dataf(!register_fifofifo_data0191),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~13 .shared_arith = "off";

arriav_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data018),
	.datae(gnd),
	.dataf(!register_fifofifo_data0201),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout());
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~17 .shared_arith = "off";

arriav_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data019),
	.datae(gnd),
	.dataf(!register_fifofifo_data0211),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout());
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~21 .shared_arith = "off";

arriav_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data020),
	.datae(gnd),
	.dataf(!register_fifofifo_data0221),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout());
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~25 .shared_arith = "off";

arriav_lcell_comb \Add0~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data021),
	.datae(gnd),
	.dataf(!register_fifofifo_data0231),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout());
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~29 .shared_arith = "off";

arriav_lcell_comb \Add0~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data022),
	.datae(gnd),
	.dataf(!register_fifofifo_data0241),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~33_sumout ),
	.cout(\Add0~34 ),
	.shareout());
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~33 .shared_arith = "off";

arriav_lcell_comb \Add0~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data023),
	.datae(gnd),
	.dataf(!register_fifofifo_data0251),
	.datag(gnd),
	.cin(\Add0~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~37_sumout ),
	.cout(\Add0~38 ),
	.shareout());
defparam \Add0~37 .extended_lut = "off";
defparam \Add0~37 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~37 .shared_arith = "off";

arriav_lcell_comb \Add0~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data024),
	.datae(gnd),
	.dataf(!register_fifofifo_data0261),
	.datag(gnd),
	.cin(\Add0~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~41_sumout ),
	.cout(\Add0~42 ),
	.shareout());
defparam \Add0~41 .extended_lut = "off";
defparam \Add0~41 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~41 .shared_arith = "off";

arriav_lcell_comb \Add0~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data025),
	.datae(gnd),
	.dataf(!register_fifofifo_data0271),
	.datag(gnd),
	.cin(\Add0~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~45_sumout ),
	.cout(\Add0~46 ),
	.shareout());
defparam \Add0~45 .extended_lut = "off";
defparam \Add0~45 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~45 .shared_arith = "off";

arriav_lcell_comb \Add0~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data026),
	.datae(gnd),
	.dataf(!register_fifofifo_data0281),
	.datag(gnd),
	.cin(\Add0~46 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~49_sumout ),
	.cout(\Add0~50 ),
	.shareout());
defparam \Add0~49 .extended_lut = "off";
defparam \Add0~49 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~49 .shared_arith = "off";

arriav_lcell_comb \Add0~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data027),
	.datae(gnd),
	.dataf(!register_fifofifo_data0291),
	.datag(gnd),
	.cin(\Add0~50 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~53_sumout ),
	.cout(\Add0~54 ),
	.shareout());
defparam \Add0~53 .extended_lut = "off";
defparam \Add0~53 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~53 .shared_arith = "off";

arriav_lcell_comb \Add0~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data028),
	.datae(gnd),
	.dataf(!register_fifofifo_data0301),
	.datag(gnd),
	.cin(\Add0~54 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~57_sumout ),
	.cout(\Add0~58 ),
	.shareout());
defparam \Add0~57 .extended_lut = "off";
defparam \Add0~57 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~57 .shared_arith = "off";

arriav_lcell_comb \Add0~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data029),
	.datae(gnd),
	.dataf(!register_fifofifo_data0311),
	.datag(gnd),
	.cin(\Add0~58 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~61_sumout ),
	.cout(\Add0~62 ),
	.shareout());
defparam \Add0~61 .extended_lut = "off";
defparam \Add0~61 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~61 .shared_arith = "off";

arriav_lcell_comb \Add0~65 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data030),
	.datae(gnd),
	.dataf(!register_fifofifo_data0321),
	.datag(gnd),
	.cin(\Add0~62 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~65_sumout ),
	.cout(\Add0~66 ),
	.shareout());
defparam \Add0~65 .extended_lut = "off";
defparam \Add0~65 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~65 .shared_arith = "off";

arriav_lcell_comb \Add0~69 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data031),
	.datae(gnd),
	.dataf(!register_fifofifo_data0331),
	.datag(gnd),
	.cin(\Add0~66 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~69_sumout ),
	.cout(\Add0~70 ),
	.shareout());
defparam \Add0~69 .extended_lut = "off";
defparam \Add0~69 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~69 .shared_arith = "off";

arriav_lcell_comb \Add0~73 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data032),
	.datae(gnd),
	.dataf(!register_fifofifo_data0341),
	.datag(gnd),
	.cin(\Add0~70 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~73_sumout ),
	.cout(\Add0~74 ),
	.shareout());
defparam \Add0~73 .extended_lut = "off";
defparam \Add0~73 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~73 .shared_arith = "off";

arriav_lcell_comb \Add0~77 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data033),
	.datae(gnd),
	.dataf(!register_fifofifo_data0351),
	.datag(gnd),
	.cin(\Add0~74 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~77_sumout ),
	.cout(\Add0~78 ),
	.shareout());
defparam \Add0~77 .extended_lut = "off";
defparam \Add0~77 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~77 .shared_arith = "off";

arriav_lcell_comb \Add0~81 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data034),
	.datae(gnd),
	.dataf(!register_fifofifo_data0361),
	.datag(gnd),
	.cin(\Add0~78 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~81_sumout ),
	.cout(\Add0~82 ),
	.shareout());
defparam \Add0~81 .extended_lut = "off";
defparam \Add0~81 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~81 .shared_arith = "off";

arriav_lcell_comb \Add0~85 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data035),
	.datae(gnd),
	.dataf(!register_fifofifo_data0371),
	.datag(gnd),
	.cin(\Add0~82 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~85_sumout ),
	.cout(\Add0~86 ),
	.shareout());
defparam \Add0~85 .extended_lut = "off";
defparam \Add0~85 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~85 .shared_arith = "off";

arriav_lcell_comb \Add0~89 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data036),
	.datae(gnd),
	.dataf(!register_fifofifo_data0381),
	.datag(gnd),
	.cin(\Add0~86 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~89_sumout ),
	.cout(\Add0~90 ),
	.shareout());
defparam \Add0~89 .extended_lut = "off";
defparam \Add0~89 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~89 .shared_arith = "off";

arriav_lcell_comb \Add0~93 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data037),
	.datae(gnd),
	.dataf(!register_fifofifo_data0391),
	.datag(gnd),
	.cin(\Add0~90 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~93_sumout ),
	.cout(\Add0~94 ),
	.shareout());
defparam \Add0~93 .extended_lut = "off";
defparam \Add0~93 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~93 .shared_arith = "off";

arriav_lcell_comb \Add0~97 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data038),
	.datae(gnd),
	.dataf(!register_fifofifo_data0401),
	.datag(gnd),
	.cin(\Add0~94 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~97_sumout ),
	.cout(\Add0~98 ),
	.shareout());
defparam \Add0~97 .extended_lut = "off";
defparam \Add0~97 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~97 .shared_arith = "off";

arriav_lcell_comb \Add0~101 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data039),
	.datae(gnd),
	.dataf(!register_fifofifo_data0411),
	.datag(gnd),
	.cin(\Add0~98 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~101_sumout ),
	.cout(\Add0~102 ),
	.shareout());
defparam \Add0~101 .extended_lut = "off";
defparam \Add0~101 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~101 .shared_arith = "off";

arriav_lcell_comb \Add0~105 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data040),
	.datae(gnd),
	.dataf(!register_fifofifo_data042),
	.datag(gnd),
	.cin(\Add0~102 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~105_sumout ),
	.cout(\Add0~106 ),
	.shareout());
defparam \Add0~105 .extended_lut = "off";
defparam \Add0~105 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~105 .shared_arith = "off";

arriav_lcell_comb \Add0~109 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data041),
	.datae(gnd),
	.dataf(!register_fifofifo_data043),
	.datag(gnd),
	.cin(\Add0~106 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~109_sumout ),
	.cout(),
	.shareout());
defparam \Add0~109 .extended_lut = "off";
defparam \Add0~109 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~109 .shared_arith = "off";

arriav_lcell_comb \Add0~113 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data013),
	.datae(gnd),
	.dataf(!register_fifofifo_data0151),
	.datag(gnd),
	.cin(\Add0~118 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~113_sumout ),
	.cout(\Add0~114 ),
	.shareout());
defparam \Add0~113 .extended_lut = "off";
defparam \Add0~113 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~113 .shared_arith = "off";

arriav_lcell_comb \Add0~117 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data012),
	.datae(gnd),
	.dataf(!register_fifofifo_data0141),
	.datag(gnd),
	.cin(\Add0~122 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~117_sumout ),
	.cout(\Add0~118 ),
	.shareout());
defparam \Add0~117 .extended_lut = "off";
defparam \Add0~117 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~117 .shared_arith = "off";

arriav_lcell_comb \Add0~121 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data011),
	.datae(gnd),
	.dataf(!register_fifofifo_data0131),
	.datag(gnd),
	.cin(\Add0~126 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~121_sumout ),
	.cout(\Add0~122 ),
	.shareout());
defparam \Add0~121 .extended_lut = "off";
defparam \Add0~121 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~121 .shared_arith = "off";

arriav_lcell_comb \Add0~125 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data010),
	.datae(gnd),
	.dataf(!register_fifofifo_data0121),
	.datag(gnd),
	.cin(\Add0~130 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~125_sumout ),
	.cout(\Add0~126 ),
	.shareout());
defparam \Add0~125 .extended_lut = "off";
defparam \Add0~125 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~125 .shared_arith = "off";

arriav_lcell_comb \Add0~129 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data09),
	.datae(gnd),
	.dataf(!register_fifofifo_data0111),
	.datag(gnd),
	.cin(\Add0~134 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~129_sumout ),
	.cout(\Add0~130 ),
	.shareout());
defparam \Add0~129 .extended_lut = "off";
defparam \Add0~129 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~129 .shared_arith = "off";

arriav_lcell_comb \Add0~133 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data08),
	.datae(gnd),
	.dataf(!register_fifofifo_data0101),
	.datag(gnd),
	.cin(\Add0~138 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~133_sumout ),
	.cout(\Add0~134 ),
	.shareout());
defparam \Add0~133 .extended_lut = "off";
defparam \Add0~133 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~133 .shared_arith = "off";

arriav_lcell_comb \Add0~137 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data07),
	.datae(gnd),
	.dataf(!register_fifofifo_data091),
	.datag(gnd),
	.cin(\Add0~142 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~137_sumout ),
	.cout(\Add0~138 ),
	.shareout());
defparam \Add0~137 .extended_lut = "off";
defparam \Add0~137 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~137 .shared_arith = "off";

arriav_lcell_comb \Add0~141 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data06),
	.datae(gnd),
	.dataf(!register_fifofifo_data081),
	.datag(gnd),
	.cin(\Add0~146 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~141_sumout ),
	.cout(\Add0~142 ),
	.shareout());
defparam \Add0~141 .extended_lut = "off";
defparam \Add0~141 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~141 .shared_arith = "off";

arriav_lcell_comb \Add0~145 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data05),
	.datae(gnd),
	.dataf(!register_fifofifo_data071),
	.datag(gnd),
	.cin(\Add0~150 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~145_sumout ),
	.cout(\Add0~146 ),
	.shareout());
defparam \Add0~145 .extended_lut = "off";
defparam \Add0~145 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~145 .shared_arith = "off";

arriav_lcell_comb \Add0~149 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data04),
	.datae(gnd),
	.dataf(!register_fifofifo_data061),
	.datag(gnd),
	.cin(\Add0~154 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~149_sumout ),
	.cout(\Add0~150 ),
	.shareout());
defparam \Add0~149 .extended_lut = "off";
defparam \Add0~149 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~149 .shared_arith = "off";

arriav_lcell_comb \Add0~153 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data03),
	.datae(gnd),
	.dataf(!register_fifofifo_data051),
	.datag(gnd),
	.cin(\Add0~158 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~153_sumout ),
	.cout(\Add0~154 ),
	.shareout());
defparam \Add0~153 .extended_lut = "off";
defparam \Add0~153 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~153 .shared_arith = "off";

arriav_lcell_comb \Add0~157 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data02),
	.datae(gnd),
	.dataf(!register_fifofifo_data044),
	.datag(gnd),
	.cin(\Add0~162 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~157_sumout ),
	.cout(\Add0~158 ),
	.shareout());
defparam \Add0~157 .extended_lut = "off";
defparam \Add0~157 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~157 .shared_arith = "off";

arriav_lcell_comb \Add0~161 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][1]~q ),
	.datae(gnd),
	.dataf(!register_fifofifo_data0310),
	.datag(gnd),
	.cin(\Add0~166 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~161_sumout ),
	.cout(\Add0~162 ),
	.shareout());
defparam \Add0~161 .extended_lut = "off";
defparam \Add0~161 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~161 .shared_arith = "off";

arriav_lcell_comb \Add0~165 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][0]~q ),
	.datae(gnd),
	.dataf(!register_fifofifo_data0210),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~165_sumout ),
	.cout(\Add0~166 ),
	.shareout());
defparam \Add0~165 .extended_lut = "off";
defparam \Add0~165 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~165 .shared_arith = "off";

endmodule

module cic_auk_dspip_delay_13 (
	datain,
	enable,
	register_fifofifo_data014,
	register_fifofifo_data015,
	register_fifofifo_data016,
	register_fifofifo_data017,
	register_fifofifo_data018,
	register_fifofifo_data019,
	register_fifofifo_data020,
	register_fifofifo_data021,
	register_fifofifo_data022,
	register_fifofifo_data023,
	register_fifofifo_data024,
	register_fifofifo_data025,
	register_fifofifo_data026,
	register_fifofifo_data027,
	register_fifofifo_data028,
	register_fifofifo_data029,
	register_fifofifo_data030,
	register_fifofifo_data031,
	register_fifofifo_data032,
	register_fifofifo_data033,
	register_fifofifo_data034,
	register_fifofifo_data035,
	register_fifofifo_data036,
	register_fifofifo_data037,
	register_fifofifo_data038,
	register_fifofifo_data039,
	register_fifofifo_data040,
	register_fifofifo_data041,
	register_fifofifo_data013,
	register_fifofifo_data012,
	register_fifofifo_data011,
	register_fifofifo_data010,
	register_fifofifo_data09,
	register_fifofifo_data08,
	register_fifofifo_data07,
	register_fifofifo_data06,
	register_fifofifo_data05,
	register_fifofifo_data04,
	register_fifofifo_data03,
	register_fifofifo_data02,
	register_fifofifo_data01,
	register_fifofifo_data00,
	clk,
	reset)/* synthesis synthesis_greybox=1 */;
input 	[46:0] datain;
input 	enable;
output 	register_fifofifo_data014;
output 	register_fifofifo_data015;
output 	register_fifofifo_data016;
output 	register_fifofifo_data017;
output 	register_fifofifo_data018;
output 	register_fifofifo_data019;
output 	register_fifofifo_data020;
output 	register_fifofifo_data021;
output 	register_fifofifo_data022;
output 	register_fifofifo_data023;
output 	register_fifofifo_data024;
output 	register_fifofifo_data025;
output 	register_fifofifo_data026;
output 	register_fifofifo_data027;
output 	register_fifofifo_data028;
output 	register_fifofifo_data029;
output 	register_fifofifo_data030;
output 	register_fifofifo_data031;
output 	register_fifofifo_data032;
output 	register_fifofifo_data033;
output 	register_fifofifo_data034;
output 	register_fifofifo_data035;
output 	register_fifofifo_data036;
output 	register_fifofifo_data037;
output 	register_fifofifo_data038;
output 	register_fifofifo_data039;
output 	register_fifofifo_data040;
output 	register_fifofifo_data041;
output 	register_fifofifo_data013;
output 	register_fifofifo_data012;
output 	register_fifofifo_data011;
output 	register_fifofifo_data010;
output 	register_fifofifo_data09;
output 	register_fifofifo_data08;
output 	register_fifofifo_data07;
output 	register_fifofifo_data06;
output 	register_fifofifo_data05;
output 	register_fifofifo_data04;
output 	register_fifofifo_data03;
output 	register_fifofifo_data02;
output 	register_fifofifo_data01;
output 	register_fifofifo_data00;
input 	clk;
input 	reset;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \register_fifo:fifo_data[0][14] (
	.clk(clk),
	.d(datain[14]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data014),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][14] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][14] .power_up = "low";

dffeas \register_fifo:fifo_data[0][15] (
	.clk(clk),
	.d(datain[15]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data015),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][15] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][15] .power_up = "low";

dffeas \register_fifo:fifo_data[0][16] (
	.clk(clk),
	.d(datain[16]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data016),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][16] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][16] .power_up = "low";

dffeas \register_fifo:fifo_data[0][17] (
	.clk(clk),
	.d(datain[17]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data017),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][17] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][17] .power_up = "low";

dffeas \register_fifo:fifo_data[0][18] (
	.clk(clk),
	.d(datain[18]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data018),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][18] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][18] .power_up = "low";

dffeas \register_fifo:fifo_data[0][19] (
	.clk(clk),
	.d(datain[19]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data019),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][19] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][19] .power_up = "low";

dffeas \register_fifo:fifo_data[0][20] (
	.clk(clk),
	.d(datain[20]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data020),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][20] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][20] .power_up = "low";

dffeas \register_fifo:fifo_data[0][21] (
	.clk(clk),
	.d(datain[21]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data021),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][21] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][21] .power_up = "low";

dffeas \register_fifo:fifo_data[0][22] (
	.clk(clk),
	.d(datain[22]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data022),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][22] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][22] .power_up = "low";

dffeas \register_fifo:fifo_data[0][23] (
	.clk(clk),
	.d(datain[23]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data023),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][23] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][23] .power_up = "low";

dffeas \register_fifo:fifo_data[0][24] (
	.clk(clk),
	.d(datain[24]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data024),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][24] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][24] .power_up = "low";

dffeas \register_fifo:fifo_data[0][25] (
	.clk(clk),
	.d(datain[25]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data025),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][25] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][25] .power_up = "low";

dffeas \register_fifo:fifo_data[0][26] (
	.clk(clk),
	.d(datain[26]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data026),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][26] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][26] .power_up = "low";

dffeas \register_fifo:fifo_data[0][27] (
	.clk(clk),
	.d(datain[27]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data027),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][27] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][27] .power_up = "low";

dffeas \register_fifo:fifo_data[0][28] (
	.clk(clk),
	.d(datain[28]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data028),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][28] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][28] .power_up = "low";

dffeas \register_fifo:fifo_data[0][29] (
	.clk(clk),
	.d(datain[29]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data029),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][29] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][29] .power_up = "low";

dffeas \register_fifo:fifo_data[0][30] (
	.clk(clk),
	.d(datain[30]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data030),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][30] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][30] .power_up = "low";

dffeas \register_fifo:fifo_data[0][31] (
	.clk(clk),
	.d(datain[31]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data031),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][31] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][31] .power_up = "low";

dffeas \register_fifo:fifo_data[0][32] (
	.clk(clk),
	.d(datain[32]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data032),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][32] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][32] .power_up = "low";

dffeas \register_fifo:fifo_data[0][33] (
	.clk(clk),
	.d(datain[33]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data033),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][33] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][33] .power_up = "low";

dffeas \register_fifo:fifo_data[0][34] (
	.clk(clk),
	.d(datain[34]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data034),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][34] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][34] .power_up = "low";

dffeas \register_fifo:fifo_data[0][35] (
	.clk(clk),
	.d(datain[35]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data035),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][35] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][35] .power_up = "low";

dffeas \register_fifo:fifo_data[0][36] (
	.clk(clk),
	.d(datain[36]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data036),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][36] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][36] .power_up = "low";

dffeas \register_fifo:fifo_data[0][37] (
	.clk(clk),
	.d(datain[37]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data037),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][37] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][37] .power_up = "low";

dffeas \register_fifo:fifo_data[0][38] (
	.clk(clk),
	.d(datain[38]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data038),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][38] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][38] .power_up = "low";

dffeas \register_fifo:fifo_data[0][39] (
	.clk(clk),
	.d(datain[39]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data039),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][39] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][39] .power_up = "low";

dffeas \register_fifo:fifo_data[0][40] (
	.clk(clk),
	.d(datain[40]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data040),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][40] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][40] .power_up = "low";

dffeas \register_fifo:fifo_data[0][41] (
	.clk(clk),
	.d(datain[41]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data041),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][41] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][41] .power_up = "low";

dffeas \register_fifo:fifo_data[0][13] (
	.clk(clk),
	.d(datain[13]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data013),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][13] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][13] .power_up = "low";

dffeas \register_fifo:fifo_data[0][12] (
	.clk(clk),
	.d(datain[12]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data012),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][12] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][12] .power_up = "low";

dffeas \register_fifo:fifo_data[0][11] (
	.clk(clk),
	.d(datain[11]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data011),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][11] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][11] .power_up = "low";

dffeas \register_fifo:fifo_data[0][10] (
	.clk(clk),
	.d(datain[10]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data010),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][10] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][10] .power_up = "low";

dffeas \register_fifo:fifo_data[0][9] (
	.clk(clk),
	.d(datain[9]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data09),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][9] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][9] .power_up = "low";

dffeas \register_fifo:fifo_data[0][8] (
	.clk(clk),
	.d(datain[8]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data08),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][8] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][8] .power_up = "low";

dffeas \register_fifo:fifo_data[0][7] (
	.clk(clk),
	.d(datain[7]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data07),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][7] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][7] .power_up = "low";

dffeas \register_fifo:fifo_data[0][6] (
	.clk(clk),
	.d(datain[6]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data06),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][6] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][6] .power_up = "low";

dffeas \register_fifo:fifo_data[0][5] (
	.clk(clk),
	.d(datain[5]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data05),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][5] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][5] .power_up = "low";

dffeas \register_fifo:fifo_data[0][4] (
	.clk(clk),
	.d(datain[4]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data04),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][4] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][4] .power_up = "low";

dffeas \register_fifo:fifo_data[0][3] (
	.clk(clk),
	.d(datain[3]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data03),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][3] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][3] .power_up = "low";

dffeas \register_fifo:fifo_data[0][2] (
	.clk(clk),
	.d(datain[2]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data02),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][2] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][2] .power_up = "low";

dffeas \register_fifo:fifo_data[0][1] (
	.clk(clk),
	.d(datain[1]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data01),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][1] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][1] .power_up = "low";

dffeas \register_fifo:fifo_data[0][0] (
	.clk(clk),
	.d(datain[0]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data00),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][0] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][0] .power_up = "low";

endmodule

module cic_auk_dspip_integrator_6 (
	stall_reg,
	register_fifofifo_data012,
	register_fifofifo_data013,
	register_fifofifo_data014,
	register_fifofifo_data015,
	register_fifofifo_data016,
	register_fifofifo_data017,
	register_fifofifo_data018,
	register_fifofifo_data019,
	register_fifofifo_data020,
	register_fifofifo_data021,
	register_fifofifo_data022,
	register_fifofifo_data023,
	register_fifofifo_data024,
	register_fifofifo_data025,
	register_fifofifo_data026,
	register_fifofifo_data027,
	register_fifofifo_data028,
	register_fifofifo_data029,
	register_fifofifo_data030,
	register_fifofifo_data031,
	register_fifofifo_data032,
	register_fifofifo_data033,
	register_fifofifo_data034,
	register_fifofifo_data035,
	register_fifofifo_data036,
	register_fifofifo_data037,
	register_fifofifo_data038,
	register_fifofifo_data039,
	register_fifofifo_data011,
	register_fifofifo_data0141,
	register_fifofifo_data010,
	register_fifofifo_data0151,
	register_fifofifo_data0161,
	register_fifofifo_data0171,
	register_fifofifo_data0181,
	register_fifofifo_data0191,
	register_fifofifo_data0201,
	register_fifofifo_data0211,
	register_fifofifo_data0221,
	register_fifofifo_data0231,
	register_fifofifo_data0241,
	register_fifofifo_data0251,
	register_fifofifo_data0261,
	register_fifofifo_data0271,
	register_fifofifo_data0281,
	register_fifofifo_data0291,
	register_fifofifo_data0301,
	register_fifofifo_data0311,
	register_fifofifo_data0321,
	register_fifofifo_data0331,
	register_fifofifo_data0341,
	register_fifofifo_data0351,
	register_fifofifo_data0361,
	register_fifofifo_data0371,
	register_fifofifo_data0381,
	register_fifofifo_data0391,
	register_fifofifo_data040,
	register_fifofifo_data041,
	register_fifofifo_data0131,
	register_fifofifo_data09,
	register_fifofifo_data0121,
	register_fifofifo_data08,
	register_fifofifo_data0111,
	register_fifofifo_data07,
	register_fifofifo_data0101,
	register_fifofifo_data06,
	register_fifofifo_data091,
	register_fifofifo_data05,
	register_fifofifo_data081,
	register_fifofifo_data04,
	register_fifofifo_data071,
	register_fifofifo_data03,
	register_fifofifo_data061,
	register_fifofifo_data02,
	register_fifofifo_data051,
	register_fifofifo_data042,
	register_fifofifo_data0310,
	register_fifofifo_data0210,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	stall_reg;
output 	register_fifofifo_data012;
output 	register_fifofifo_data013;
output 	register_fifofifo_data014;
output 	register_fifofifo_data015;
output 	register_fifofifo_data016;
output 	register_fifofifo_data017;
output 	register_fifofifo_data018;
output 	register_fifofifo_data019;
output 	register_fifofifo_data020;
output 	register_fifofifo_data021;
output 	register_fifofifo_data022;
output 	register_fifofifo_data023;
output 	register_fifofifo_data024;
output 	register_fifofifo_data025;
output 	register_fifofifo_data026;
output 	register_fifofifo_data027;
output 	register_fifofifo_data028;
output 	register_fifofifo_data029;
output 	register_fifofifo_data030;
output 	register_fifofifo_data031;
output 	register_fifofifo_data032;
output 	register_fifofifo_data033;
output 	register_fifofifo_data034;
output 	register_fifofifo_data035;
output 	register_fifofifo_data036;
output 	register_fifofifo_data037;
output 	register_fifofifo_data038;
output 	register_fifofifo_data039;
output 	register_fifofifo_data011;
input 	register_fifofifo_data0141;
output 	register_fifofifo_data010;
input 	register_fifofifo_data0151;
input 	register_fifofifo_data0161;
input 	register_fifofifo_data0171;
input 	register_fifofifo_data0181;
input 	register_fifofifo_data0191;
input 	register_fifofifo_data0201;
input 	register_fifofifo_data0211;
input 	register_fifofifo_data0221;
input 	register_fifofifo_data0231;
input 	register_fifofifo_data0241;
input 	register_fifofifo_data0251;
input 	register_fifofifo_data0261;
input 	register_fifofifo_data0271;
input 	register_fifofifo_data0281;
input 	register_fifofifo_data0291;
input 	register_fifofifo_data0301;
input 	register_fifofifo_data0311;
input 	register_fifofifo_data0321;
input 	register_fifofifo_data0331;
input 	register_fifofifo_data0341;
input 	register_fifofifo_data0351;
input 	register_fifofifo_data0361;
input 	register_fifofifo_data0371;
input 	register_fifofifo_data0381;
input 	register_fifofifo_data0391;
input 	register_fifofifo_data040;
input 	register_fifofifo_data041;
input 	register_fifofifo_data0131;
output 	register_fifofifo_data09;
input 	register_fifofifo_data0121;
output 	register_fifofifo_data08;
input 	register_fifofifo_data0111;
output 	register_fifofifo_data07;
input 	register_fifofifo_data0101;
output 	register_fifofifo_data06;
input 	register_fifofifo_data091;
output 	register_fifofifo_data05;
input 	register_fifofifo_data081;
output 	register_fifofifo_data04;
input 	register_fifofifo_data071;
output 	register_fifofifo_data03;
input 	register_fifofifo_data061;
output 	register_fifofifo_data02;
input 	register_fifofifo_data051;
input 	register_fifofifo_data042;
input 	register_fifofifo_data0310;
input 	register_fifofifo_data0210;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Add0~1_sumout ;
wire \Add0~2 ;
wire \Add0~5_sumout ;
wire \Add0~6 ;
wire \Add0~9_sumout ;
wire \Add0~10 ;
wire \Add0~13_sumout ;
wire \Add0~14 ;
wire \Add0~17_sumout ;
wire \Add0~18 ;
wire \Add0~21_sumout ;
wire \Add0~22 ;
wire \Add0~25_sumout ;
wire \Add0~26 ;
wire \Add0~29_sumout ;
wire \Add0~30 ;
wire \Add0~33_sumout ;
wire \Add0~34 ;
wire \Add0~37_sumout ;
wire \Add0~38 ;
wire \Add0~41_sumout ;
wire \Add0~42 ;
wire \Add0~45_sumout ;
wire \Add0~46 ;
wire \Add0~49_sumout ;
wire \Add0~50 ;
wire \Add0~53_sumout ;
wire \Add0~54 ;
wire \Add0~57_sumout ;
wire \Add0~58 ;
wire \Add0~61_sumout ;
wire \Add0~62 ;
wire \Add0~65_sumout ;
wire \Add0~66 ;
wire \Add0~69_sumout ;
wire \Add0~70 ;
wire \Add0~73_sumout ;
wire \Add0~74 ;
wire \Add0~77_sumout ;
wire \Add0~78 ;
wire \Add0~81_sumout ;
wire \Add0~82 ;
wire \Add0~85_sumout ;
wire \Add0~86 ;
wire \Add0~89_sumout ;
wire \Add0~90 ;
wire \Add0~93_sumout ;
wire \Add0~94 ;
wire \Add0~97_sumout ;
wire \Add0~98 ;
wire \Add0~101_sumout ;
wire \Add0~102 ;
wire \Add0~105_sumout ;
wire \Add0~106 ;
wire \Add0~109_sumout ;
wire \Add0~113_sumout ;
wire \Add0~114 ;
wire \Add0~117_sumout ;
wire \Add0~118 ;
wire \Add0~121_sumout ;
wire \Add0~122 ;
wire \Add0~125_sumout ;
wire \Add0~126 ;
wire \Add0~129_sumout ;
wire \Add0~130 ;
wire \Add0~133_sumout ;
wire \Add0~134 ;
wire \Add0~137_sumout ;
wire \Add0~138 ;
wire \Add0~141_sumout ;
wire \Add0~142 ;
wire \Add0~145_sumout ;
wire \Add0~146 ;
wire \Add0~149_sumout ;
wire \Add0~150 ;
wire \Add0~153_sumout ;
wire \Add0~154 ;
wire \Add0~157_sumout ;
wire \Add0~158 ;
wire \glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][1]~q ;
wire \glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][0]~q ;


cic_auk_dspip_delay_14 \glogic:integrator_pipeline_0_generate:u1 (
	.datain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,\Add0~109_sumout ,\Add0~105_sumout ,\Add0~101_sumout ,\Add0~97_sumout ,\Add0~93_sumout ,\Add0~89_sumout ,\Add0~85_sumout ,\Add0~81_sumout ,\Add0~77_sumout ,\Add0~73_sumout ,\Add0~69_sumout ,\Add0~65_sumout ,\Add0~61_sumout ,\Add0~57_sumout ,
\Add0~53_sumout ,\Add0~49_sumout ,\Add0~45_sumout ,\Add0~41_sumout ,\Add0~37_sumout ,\Add0~33_sumout ,\Add0~29_sumout ,\Add0~25_sumout ,\Add0~21_sumout ,\Add0~17_sumout ,\Add0~13_sumout ,\Add0~9_sumout ,\Add0~5_sumout ,\Add0~1_sumout ,\Add0~113_sumout ,\Add0~117_sumout ,
\Add0~121_sumout ,\Add0~125_sumout ,\Add0~129_sumout ,\Add0~133_sumout ,\Add0~137_sumout ,\Add0~141_sumout ,\Add0~145_sumout ,\Add0~149_sumout ,\Add0~153_sumout ,\Add0~157_sumout }),
	.enable(stall_reg),
	.register_fifofifo_data012(register_fifofifo_data012),
	.register_fifofifo_data013(register_fifofifo_data013),
	.register_fifofifo_data014(register_fifofifo_data014),
	.register_fifofifo_data015(register_fifofifo_data015),
	.register_fifofifo_data016(register_fifofifo_data016),
	.register_fifofifo_data017(register_fifofifo_data017),
	.register_fifofifo_data018(register_fifofifo_data018),
	.register_fifofifo_data019(register_fifofifo_data019),
	.register_fifofifo_data020(register_fifofifo_data020),
	.register_fifofifo_data021(register_fifofifo_data021),
	.register_fifofifo_data022(register_fifofifo_data022),
	.register_fifofifo_data023(register_fifofifo_data023),
	.register_fifofifo_data024(register_fifofifo_data024),
	.register_fifofifo_data025(register_fifofifo_data025),
	.register_fifofifo_data026(register_fifofifo_data026),
	.register_fifofifo_data027(register_fifofifo_data027),
	.register_fifofifo_data028(register_fifofifo_data028),
	.register_fifofifo_data029(register_fifofifo_data029),
	.register_fifofifo_data030(register_fifofifo_data030),
	.register_fifofifo_data031(register_fifofifo_data031),
	.register_fifofifo_data032(register_fifofifo_data032),
	.register_fifofifo_data033(register_fifofifo_data033),
	.register_fifofifo_data034(register_fifofifo_data034),
	.register_fifofifo_data035(register_fifofifo_data035),
	.register_fifofifo_data036(register_fifofifo_data036),
	.register_fifofifo_data037(register_fifofifo_data037),
	.register_fifofifo_data038(register_fifofifo_data038),
	.register_fifofifo_data039(register_fifofifo_data039),
	.register_fifofifo_data011(register_fifofifo_data011),
	.register_fifofifo_data010(register_fifofifo_data010),
	.register_fifofifo_data09(register_fifofifo_data09),
	.register_fifofifo_data08(register_fifofifo_data08),
	.register_fifofifo_data07(register_fifofifo_data07),
	.register_fifofifo_data06(register_fifofifo_data06),
	.register_fifofifo_data05(register_fifofifo_data05),
	.register_fifofifo_data04(register_fifofifo_data04),
	.register_fifofifo_data03(register_fifofifo_data03),
	.register_fifofifo_data02(register_fifofifo_data02),
	.register_fifofifo_data01(\glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][1]~q ),
	.register_fifofifo_data00(\glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][0]~q ),
	.clk(clk),
	.reset(reset_n));

arriav_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data012),
	.datae(gnd),
	.dataf(!register_fifofifo_data0141),
	.datag(gnd),
	.cin(\Add0~114 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(\Add0~2 ),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~1 .shared_arith = "off";

arriav_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data013),
	.datae(gnd),
	.dataf(!register_fifofifo_data0151),
	.datag(gnd),
	.cin(\Add0~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~5 .shared_arith = "off";

arriav_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data014),
	.datae(gnd),
	.dataf(!register_fifofifo_data0161),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~9 .shared_arith = "off";

arriav_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data015),
	.datae(gnd),
	.dataf(!register_fifofifo_data0171),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~13 .shared_arith = "off";

arriav_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data016),
	.datae(gnd),
	.dataf(!register_fifofifo_data0181),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout());
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~17 .shared_arith = "off";

arriav_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data017),
	.datae(gnd),
	.dataf(!register_fifofifo_data0191),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout());
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~21 .shared_arith = "off";

arriav_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data018),
	.datae(gnd),
	.dataf(!register_fifofifo_data0201),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout());
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~25 .shared_arith = "off";

arriav_lcell_comb \Add0~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data019),
	.datae(gnd),
	.dataf(!register_fifofifo_data0211),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout());
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~29 .shared_arith = "off";

arriav_lcell_comb \Add0~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data020),
	.datae(gnd),
	.dataf(!register_fifofifo_data0221),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~33_sumout ),
	.cout(\Add0~34 ),
	.shareout());
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~33 .shared_arith = "off";

arriav_lcell_comb \Add0~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data021),
	.datae(gnd),
	.dataf(!register_fifofifo_data0231),
	.datag(gnd),
	.cin(\Add0~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~37_sumout ),
	.cout(\Add0~38 ),
	.shareout());
defparam \Add0~37 .extended_lut = "off";
defparam \Add0~37 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~37 .shared_arith = "off";

arriav_lcell_comb \Add0~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data022),
	.datae(gnd),
	.dataf(!register_fifofifo_data0241),
	.datag(gnd),
	.cin(\Add0~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~41_sumout ),
	.cout(\Add0~42 ),
	.shareout());
defparam \Add0~41 .extended_lut = "off";
defparam \Add0~41 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~41 .shared_arith = "off";

arriav_lcell_comb \Add0~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data023),
	.datae(gnd),
	.dataf(!register_fifofifo_data0251),
	.datag(gnd),
	.cin(\Add0~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~45_sumout ),
	.cout(\Add0~46 ),
	.shareout());
defparam \Add0~45 .extended_lut = "off";
defparam \Add0~45 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~45 .shared_arith = "off";

arriav_lcell_comb \Add0~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data024),
	.datae(gnd),
	.dataf(!register_fifofifo_data0261),
	.datag(gnd),
	.cin(\Add0~46 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~49_sumout ),
	.cout(\Add0~50 ),
	.shareout());
defparam \Add0~49 .extended_lut = "off";
defparam \Add0~49 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~49 .shared_arith = "off";

arriav_lcell_comb \Add0~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data025),
	.datae(gnd),
	.dataf(!register_fifofifo_data0271),
	.datag(gnd),
	.cin(\Add0~50 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~53_sumout ),
	.cout(\Add0~54 ),
	.shareout());
defparam \Add0~53 .extended_lut = "off";
defparam \Add0~53 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~53 .shared_arith = "off";

arriav_lcell_comb \Add0~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data026),
	.datae(gnd),
	.dataf(!register_fifofifo_data0281),
	.datag(gnd),
	.cin(\Add0~54 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~57_sumout ),
	.cout(\Add0~58 ),
	.shareout());
defparam \Add0~57 .extended_lut = "off";
defparam \Add0~57 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~57 .shared_arith = "off";

arriav_lcell_comb \Add0~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data027),
	.datae(gnd),
	.dataf(!register_fifofifo_data0291),
	.datag(gnd),
	.cin(\Add0~58 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~61_sumout ),
	.cout(\Add0~62 ),
	.shareout());
defparam \Add0~61 .extended_lut = "off";
defparam \Add0~61 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~61 .shared_arith = "off";

arriav_lcell_comb \Add0~65 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data028),
	.datae(gnd),
	.dataf(!register_fifofifo_data0301),
	.datag(gnd),
	.cin(\Add0~62 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~65_sumout ),
	.cout(\Add0~66 ),
	.shareout());
defparam \Add0~65 .extended_lut = "off";
defparam \Add0~65 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~65 .shared_arith = "off";

arriav_lcell_comb \Add0~69 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data029),
	.datae(gnd),
	.dataf(!register_fifofifo_data0311),
	.datag(gnd),
	.cin(\Add0~66 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~69_sumout ),
	.cout(\Add0~70 ),
	.shareout());
defparam \Add0~69 .extended_lut = "off";
defparam \Add0~69 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~69 .shared_arith = "off";

arriav_lcell_comb \Add0~73 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data030),
	.datae(gnd),
	.dataf(!register_fifofifo_data0321),
	.datag(gnd),
	.cin(\Add0~70 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~73_sumout ),
	.cout(\Add0~74 ),
	.shareout());
defparam \Add0~73 .extended_lut = "off";
defparam \Add0~73 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~73 .shared_arith = "off";

arriav_lcell_comb \Add0~77 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data031),
	.datae(gnd),
	.dataf(!register_fifofifo_data0331),
	.datag(gnd),
	.cin(\Add0~74 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~77_sumout ),
	.cout(\Add0~78 ),
	.shareout());
defparam \Add0~77 .extended_lut = "off";
defparam \Add0~77 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~77 .shared_arith = "off";

arriav_lcell_comb \Add0~81 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data032),
	.datae(gnd),
	.dataf(!register_fifofifo_data0341),
	.datag(gnd),
	.cin(\Add0~78 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~81_sumout ),
	.cout(\Add0~82 ),
	.shareout());
defparam \Add0~81 .extended_lut = "off";
defparam \Add0~81 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~81 .shared_arith = "off";

arriav_lcell_comb \Add0~85 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data033),
	.datae(gnd),
	.dataf(!register_fifofifo_data0351),
	.datag(gnd),
	.cin(\Add0~82 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~85_sumout ),
	.cout(\Add0~86 ),
	.shareout());
defparam \Add0~85 .extended_lut = "off";
defparam \Add0~85 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~85 .shared_arith = "off";

arriav_lcell_comb \Add0~89 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data034),
	.datae(gnd),
	.dataf(!register_fifofifo_data0361),
	.datag(gnd),
	.cin(\Add0~86 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~89_sumout ),
	.cout(\Add0~90 ),
	.shareout());
defparam \Add0~89 .extended_lut = "off";
defparam \Add0~89 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~89 .shared_arith = "off";

arriav_lcell_comb \Add0~93 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data035),
	.datae(gnd),
	.dataf(!register_fifofifo_data0371),
	.datag(gnd),
	.cin(\Add0~90 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~93_sumout ),
	.cout(\Add0~94 ),
	.shareout());
defparam \Add0~93 .extended_lut = "off";
defparam \Add0~93 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~93 .shared_arith = "off";

arriav_lcell_comb \Add0~97 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data036),
	.datae(gnd),
	.dataf(!register_fifofifo_data0381),
	.datag(gnd),
	.cin(\Add0~94 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~97_sumout ),
	.cout(\Add0~98 ),
	.shareout());
defparam \Add0~97 .extended_lut = "off";
defparam \Add0~97 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~97 .shared_arith = "off";

arriav_lcell_comb \Add0~101 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data037),
	.datae(gnd),
	.dataf(!register_fifofifo_data0391),
	.datag(gnd),
	.cin(\Add0~98 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~101_sumout ),
	.cout(\Add0~102 ),
	.shareout());
defparam \Add0~101 .extended_lut = "off";
defparam \Add0~101 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~101 .shared_arith = "off";

arriav_lcell_comb \Add0~105 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data038),
	.datae(gnd),
	.dataf(!register_fifofifo_data040),
	.datag(gnd),
	.cin(\Add0~102 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~105_sumout ),
	.cout(\Add0~106 ),
	.shareout());
defparam \Add0~105 .extended_lut = "off";
defparam \Add0~105 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~105 .shared_arith = "off";

arriav_lcell_comb \Add0~109 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data039),
	.datae(gnd),
	.dataf(!register_fifofifo_data041),
	.datag(gnd),
	.cin(\Add0~106 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~109_sumout ),
	.cout(),
	.shareout());
defparam \Add0~109 .extended_lut = "off";
defparam \Add0~109 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~109 .shared_arith = "off";

arriav_lcell_comb \Add0~113 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data011),
	.datae(gnd),
	.dataf(!register_fifofifo_data0131),
	.datag(gnd),
	.cin(\Add0~118 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~113_sumout ),
	.cout(\Add0~114 ),
	.shareout());
defparam \Add0~113 .extended_lut = "off";
defparam \Add0~113 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~113 .shared_arith = "off";

arriav_lcell_comb \Add0~117 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data010),
	.datae(gnd),
	.dataf(!register_fifofifo_data0121),
	.datag(gnd),
	.cin(\Add0~122 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~117_sumout ),
	.cout(\Add0~118 ),
	.shareout());
defparam \Add0~117 .extended_lut = "off";
defparam \Add0~117 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~117 .shared_arith = "off";

arriav_lcell_comb \Add0~121 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data09),
	.datae(gnd),
	.dataf(!register_fifofifo_data0111),
	.datag(gnd),
	.cin(\Add0~126 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~121_sumout ),
	.cout(\Add0~122 ),
	.shareout());
defparam \Add0~121 .extended_lut = "off";
defparam \Add0~121 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~121 .shared_arith = "off";

arriav_lcell_comb \Add0~125 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data08),
	.datae(gnd),
	.dataf(!register_fifofifo_data0101),
	.datag(gnd),
	.cin(\Add0~130 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~125_sumout ),
	.cout(\Add0~126 ),
	.shareout());
defparam \Add0~125 .extended_lut = "off";
defparam \Add0~125 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~125 .shared_arith = "off";

arriav_lcell_comb \Add0~129 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data07),
	.datae(gnd),
	.dataf(!register_fifofifo_data091),
	.datag(gnd),
	.cin(\Add0~134 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~129_sumout ),
	.cout(\Add0~130 ),
	.shareout());
defparam \Add0~129 .extended_lut = "off";
defparam \Add0~129 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~129 .shared_arith = "off";

arriav_lcell_comb \Add0~133 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data06),
	.datae(gnd),
	.dataf(!register_fifofifo_data081),
	.datag(gnd),
	.cin(\Add0~138 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~133_sumout ),
	.cout(\Add0~134 ),
	.shareout());
defparam \Add0~133 .extended_lut = "off";
defparam \Add0~133 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~133 .shared_arith = "off";

arriav_lcell_comb \Add0~137 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data05),
	.datae(gnd),
	.dataf(!register_fifofifo_data071),
	.datag(gnd),
	.cin(\Add0~142 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~137_sumout ),
	.cout(\Add0~138 ),
	.shareout());
defparam \Add0~137 .extended_lut = "off";
defparam \Add0~137 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~137 .shared_arith = "off";

arriav_lcell_comb \Add0~141 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data04),
	.datae(gnd),
	.dataf(!register_fifofifo_data061),
	.datag(gnd),
	.cin(\Add0~146 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~141_sumout ),
	.cout(\Add0~142 ),
	.shareout());
defparam \Add0~141 .extended_lut = "off";
defparam \Add0~141 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~141 .shared_arith = "off";

arriav_lcell_comb \Add0~145 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data03),
	.datae(gnd),
	.dataf(!register_fifofifo_data051),
	.datag(gnd),
	.cin(\Add0~150 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~145_sumout ),
	.cout(\Add0~146 ),
	.shareout());
defparam \Add0~145 .extended_lut = "off";
defparam \Add0~145 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~145 .shared_arith = "off";

arriav_lcell_comb \Add0~149 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data02),
	.datae(gnd),
	.dataf(!register_fifofifo_data042),
	.datag(gnd),
	.cin(\Add0~154 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~149_sumout ),
	.cout(\Add0~150 ),
	.shareout());
defparam \Add0~149 .extended_lut = "off";
defparam \Add0~149 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~149 .shared_arith = "off";

arriav_lcell_comb \Add0~153 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][1]~q ),
	.datae(gnd),
	.dataf(!register_fifofifo_data0310),
	.datag(gnd),
	.cin(\Add0~158 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~153_sumout ),
	.cout(\Add0~154 ),
	.shareout());
defparam \Add0~153 .extended_lut = "off";
defparam \Add0~153 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~153 .shared_arith = "off";

arriav_lcell_comb \Add0~157 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][0]~q ),
	.datae(gnd),
	.dataf(!register_fifofifo_data0210),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~157_sumout ),
	.cout(\Add0~158 ),
	.shareout());
defparam \Add0~157 .extended_lut = "off";
defparam \Add0~157 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~157 .shared_arith = "off";

endmodule

module cic_auk_dspip_delay_14 (
	datain,
	enable,
	register_fifofifo_data012,
	register_fifofifo_data013,
	register_fifofifo_data014,
	register_fifofifo_data015,
	register_fifofifo_data016,
	register_fifofifo_data017,
	register_fifofifo_data018,
	register_fifofifo_data019,
	register_fifofifo_data020,
	register_fifofifo_data021,
	register_fifofifo_data022,
	register_fifofifo_data023,
	register_fifofifo_data024,
	register_fifofifo_data025,
	register_fifofifo_data026,
	register_fifofifo_data027,
	register_fifofifo_data028,
	register_fifofifo_data029,
	register_fifofifo_data030,
	register_fifofifo_data031,
	register_fifofifo_data032,
	register_fifofifo_data033,
	register_fifofifo_data034,
	register_fifofifo_data035,
	register_fifofifo_data036,
	register_fifofifo_data037,
	register_fifofifo_data038,
	register_fifofifo_data039,
	register_fifofifo_data011,
	register_fifofifo_data010,
	register_fifofifo_data09,
	register_fifofifo_data08,
	register_fifofifo_data07,
	register_fifofifo_data06,
	register_fifofifo_data05,
	register_fifofifo_data04,
	register_fifofifo_data03,
	register_fifofifo_data02,
	register_fifofifo_data01,
	register_fifofifo_data00,
	clk,
	reset)/* synthesis synthesis_greybox=1 */;
input 	[46:0] datain;
input 	enable;
output 	register_fifofifo_data012;
output 	register_fifofifo_data013;
output 	register_fifofifo_data014;
output 	register_fifofifo_data015;
output 	register_fifofifo_data016;
output 	register_fifofifo_data017;
output 	register_fifofifo_data018;
output 	register_fifofifo_data019;
output 	register_fifofifo_data020;
output 	register_fifofifo_data021;
output 	register_fifofifo_data022;
output 	register_fifofifo_data023;
output 	register_fifofifo_data024;
output 	register_fifofifo_data025;
output 	register_fifofifo_data026;
output 	register_fifofifo_data027;
output 	register_fifofifo_data028;
output 	register_fifofifo_data029;
output 	register_fifofifo_data030;
output 	register_fifofifo_data031;
output 	register_fifofifo_data032;
output 	register_fifofifo_data033;
output 	register_fifofifo_data034;
output 	register_fifofifo_data035;
output 	register_fifofifo_data036;
output 	register_fifofifo_data037;
output 	register_fifofifo_data038;
output 	register_fifofifo_data039;
output 	register_fifofifo_data011;
output 	register_fifofifo_data010;
output 	register_fifofifo_data09;
output 	register_fifofifo_data08;
output 	register_fifofifo_data07;
output 	register_fifofifo_data06;
output 	register_fifofifo_data05;
output 	register_fifofifo_data04;
output 	register_fifofifo_data03;
output 	register_fifofifo_data02;
output 	register_fifofifo_data01;
output 	register_fifofifo_data00;
input 	clk;
input 	reset;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \register_fifo:fifo_data[0][12] (
	.clk(clk),
	.d(datain[12]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data012),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][12] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][12] .power_up = "low";

dffeas \register_fifo:fifo_data[0][13] (
	.clk(clk),
	.d(datain[13]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data013),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][13] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][13] .power_up = "low";

dffeas \register_fifo:fifo_data[0][14] (
	.clk(clk),
	.d(datain[14]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data014),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][14] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][14] .power_up = "low";

dffeas \register_fifo:fifo_data[0][15] (
	.clk(clk),
	.d(datain[15]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data015),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][15] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][15] .power_up = "low";

dffeas \register_fifo:fifo_data[0][16] (
	.clk(clk),
	.d(datain[16]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data016),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][16] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][16] .power_up = "low";

dffeas \register_fifo:fifo_data[0][17] (
	.clk(clk),
	.d(datain[17]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data017),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][17] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][17] .power_up = "low";

dffeas \register_fifo:fifo_data[0][18] (
	.clk(clk),
	.d(datain[18]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data018),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][18] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][18] .power_up = "low";

dffeas \register_fifo:fifo_data[0][19] (
	.clk(clk),
	.d(datain[19]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data019),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][19] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][19] .power_up = "low";

dffeas \register_fifo:fifo_data[0][20] (
	.clk(clk),
	.d(datain[20]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data020),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][20] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][20] .power_up = "low";

dffeas \register_fifo:fifo_data[0][21] (
	.clk(clk),
	.d(datain[21]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data021),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][21] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][21] .power_up = "low";

dffeas \register_fifo:fifo_data[0][22] (
	.clk(clk),
	.d(datain[22]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data022),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][22] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][22] .power_up = "low";

dffeas \register_fifo:fifo_data[0][23] (
	.clk(clk),
	.d(datain[23]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data023),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][23] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][23] .power_up = "low";

dffeas \register_fifo:fifo_data[0][24] (
	.clk(clk),
	.d(datain[24]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data024),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][24] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][24] .power_up = "low";

dffeas \register_fifo:fifo_data[0][25] (
	.clk(clk),
	.d(datain[25]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data025),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][25] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][25] .power_up = "low";

dffeas \register_fifo:fifo_data[0][26] (
	.clk(clk),
	.d(datain[26]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data026),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][26] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][26] .power_up = "low";

dffeas \register_fifo:fifo_data[0][27] (
	.clk(clk),
	.d(datain[27]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data027),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][27] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][27] .power_up = "low";

dffeas \register_fifo:fifo_data[0][28] (
	.clk(clk),
	.d(datain[28]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data028),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][28] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][28] .power_up = "low";

dffeas \register_fifo:fifo_data[0][29] (
	.clk(clk),
	.d(datain[29]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data029),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][29] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][29] .power_up = "low";

dffeas \register_fifo:fifo_data[0][30] (
	.clk(clk),
	.d(datain[30]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data030),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][30] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][30] .power_up = "low";

dffeas \register_fifo:fifo_data[0][31] (
	.clk(clk),
	.d(datain[31]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data031),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][31] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][31] .power_up = "low";

dffeas \register_fifo:fifo_data[0][32] (
	.clk(clk),
	.d(datain[32]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data032),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][32] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][32] .power_up = "low";

dffeas \register_fifo:fifo_data[0][33] (
	.clk(clk),
	.d(datain[33]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data033),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][33] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][33] .power_up = "low";

dffeas \register_fifo:fifo_data[0][34] (
	.clk(clk),
	.d(datain[34]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data034),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][34] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][34] .power_up = "low";

dffeas \register_fifo:fifo_data[0][35] (
	.clk(clk),
	.d(datain[35]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data035),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][35] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][35] .power_up = "low";

dffeas \register_fifo:fifo_data[0][36] (
	.clk(clk),
	.d(datain[36]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data036),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][36] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][36] .power_up = "low";

dffeas \register_fifo:fifo_data[0][37] (
	.clk(clk),
	.d(datain[37]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data037),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][37] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][37] .power_up = "low";

dffeas \register_fifo:fifo_data[0][38] (
	.clk(clk),
	.d(datain[38]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data038),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][38] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][38] .power_up = "low";

dffeas \register_fifo:fifo_data[0][39] (
	.clk(clk),
	.d(datain[39]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data039),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][39] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][39] .power_up = "low";

dffeas \register_fifo:fifo_data[0][11] (
	.clk(clk),
	.d(datain[11]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data011),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][11] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][11] .power_up = "low";

dffeas \register_fifo:fifo_data[0][10] (
	.clk(clk),
	.d(datain[10]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data010),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][10] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][10] .power_up = "low";

dffeas \register_fifo:fifo_data[0][9] (
	.clk(clk),
	.d(datain[9]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data09),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][9] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][9] .power_up = "low";

dffeas \register_fifo:fifo_data[0][8] (
	.clk(clk),
	.d(datain[8]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data08),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][8] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][8] .power_up = "low";

dffeas \register_fifo:fifo_data[0][7] (
	.clk(clk),
	.d(datain[7]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data07),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][7] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][7] .power_up = "low";

dffeas \register_fifo:fifo_data[0][6] (
	.clk(clk),
	.d(datain[6]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data06),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][6] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][6] .power_up = "low";

dffeas \register_fifo:fifo_data[0][5] (
	.clk(clk),
	.d(datain[5]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data05),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][5] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][5] .power_up = "low";

dffeas \register_fifo:fifo_data[0][4] (
	.clk(clk),
	.d(datain[4]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data04),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][4] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][4] .power_up = "low";

dffeas \register_fifo:fifo_data[0][3] (
	.clk(clk),
	.d(datain[3]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data03),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][3] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][3] .power_up = "low";

dffeas \register_fifo:fifo_data[0][2] (
	.clk(clk),
	.d(datain[2]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data02),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][2] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][2] .power_up = "low";

dffeas \register_fifo:fifo_data[0][1] (
	.clk(clk),
	.d(datain[1]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data01),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][1] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][1] .power_up = "low";

dffeas \register_fifo:fifo_data[0][0] (
	.clk(clk),
	.d(datain[0]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data00),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][0] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][0] .power_up = "low";

endmodule

module cic_auk_dspip_integrator_7 (
	stall_reg,
	register_fifofifo_data010,
	register_fifofifo_data011,
	register_fifofifo_data012,
	register_fifofifo_data013,
	register_fifofifo_data014,
	register_fifofifo_data015,
	register_fifofifo_data016,
	register_fifofifo_data017,
	register_fifofifo_data018,
	register_fifofifo_data019,
	register_fifofifo_data020,
	register_fifofifo_data021,
	register_fifofifo_data022,
	register_fifofifo_data023,
	register_fifofifo_data024,
	register_fifofifo_data025,
	register_fifofifo_data026,
	register_fifofifo_data027,
	register_fifofifo_data028,
	register_fifofifo_data029,
	register_fifofifo_data030,
	register_fifofifo_data031,
	register_fifofifo_data032,
	register_fifofifo_data033,
	register_fifofifo_data034,
	register_fifofifo_data035,
	register_fifofifo_data036,
	register_fifofifo_data037,
	register_fifofifo_data09,
	register_fifofifo_data0121,
	register_fifofifo_data08,
	register_fifofifo_data0131,
	register_fifofifo_data0141,
	register_fifofifo_data0151,
	register_fifofifo_data0161,
	register_fifofifo_data0171,
	register_fifofifo_data0181,
	register_fifofifo_data0191,
	register_fifofifo_data0201,
	register_fifofifo_data0211,
	register_fifofifo_data0221,
	register_fifofifo_data0231,
	register_fifofifo_data0241,
	register_fifofifo_data0251,
	register_fifofifo_data0261,
	register_fifofifo_data0271,
	register_fifofifo_data0281,
	register_fifofifo_data0291,
	register_fifofifo_data0301,
	register_fifofifo_data0311,
	register_fifofifo_data0321,
	register_fifofifo_data0331,
	register_fifofifo_data0341,
	register_fifofifo_data0351,
	register_fifofifo_data0361,
	register_fifofifo_data0371,
	register_fifofifo_data038,
	register_fifofifo_data039,
	register_fifofifo_data0111,
	register_fifofifo_data07,
	register_fifofifo_data0101,
	register_fifofifo_data06,
	register_fifofifo_data091,
	register_fifofifo_data05,
	register_fifofifo_data081,
	register_fifofifo_data04,
	register_fifofifo_data071,
	register_fifofifo_data03,
	register_fifofifo_data061,
	register_fifofifo_data02,
	register_fifofifo_data051,
	register_fifofifo_data01,
	register_fifofifo_data041,
	register_fifofifo_data0310,
	register_fifofifo_data0210,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	stall_reg;
output 	register_fifofifo_data010;
output 	register_fifofifo_data011;
output 	register_fifofifo_data012;
output 	register_fifofifo_data013;
output 	register_fifofifo_data014;
output 	register_fifofifo_data015;
output 	register_fifofifo_data016;
output 	register_fifofifo_data017;
output 	register_fifofifo_data018;
output 	register_fifofifo_data019;
output 	register_fifofifo_data020;
output 	register_fifofifo_data021;
output 	register_fifofifo_data022;
output 	register_fifofifo_data023;
output 	register_fifofifo_data024;
output 	register_fifofifo_data025;
output 	register_fifofifo_data026;
output 	register_fifofifo_data027;
output 	register_fifofifo_data028;
output 	register_fifofifo_data029;
output 	register_fifofifo_data030;
output 	register_fifofifo_data031;
output 	register_fifofifo_data032;
output 	register_fifofifo_data033;
output 	register_fifofifo_data034;
output 	register_fifofifo_data035;
output 	register_fifofifo_data036;
output 	register_fifofifo_data037;
output 	register_fifofifo_data09;
input 	register_fifofifo_data0121;
output 	register_fifofifo_data08;
input 	register_fifofifo_data0131;
input 	register_fifofifo_data0141;
input 	register_fifofifo_data0151;
input 	register_fifofifo_data0161;
input 	register_fifofifo_data0171;
input 	register_fifofifo_data0181;
input 	register_fifofifo_data0191;
input 	register_fifofifo_data0201;
input 	register_fifofifo_data0211;
input 	register_fifofifo_data0221;
input 	register_fifofifo_data0231;
input 	register_fifofifo_data0241;
input 	register_fifofifo_data0251;
input 	register_fifofifo_data0261;
input 	register_fifofifo_data0271;
input 	register_fifofifo_data0281;
input 	register_fifofifo_data0291;
input 	register_fifofifo_data0301;
input 	register_fifofifo_data0311;
input 	register_fifofifo_data0321;
input 	register_fifofifo_data0331;
input 	register_fifofifo_data0341;
input 	register_fifofifo_data0351;
input 	register_fifofifo_data0361;
input 	register_fifofifo_data0371;
input 	register_fifofifo_data038;
input 	register_fifofifo_data039;
input 	register_fifofifo_data0111;
output 	register_fifofifo_data07;
input 	register_fifofifo_data0101;
output 	register_fifofifo_data06;
input 	register_fifofifo_data091;
output 	register_fifofifo_data05;
input 	register_fifofifo_data081;
output 	register_fifofifo_data04;
input 	register_fifofifo_data071;
output 	register_fifofifo_data03;
input 	register_fifofifo_data061;
output 	register_fifofifo_data02;
input 	register_fifofifo_data051;
output 	register_fifofifo_data01;
input 	register_fifofifo_data041;
input 	register_fifofifo_data0310;
input 	register_fifofifo_data0210;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Add0~1_sumout ;
wire \Add0~2 ;
wire \Add0~5_sumout ;
wire \Add0~6 ;
wire \Add0~9_sumout ;
wire \Add0~10 ;
wire \Add0~13_sumout ;
wire \Add0~14 ;
wire \Add0~17_sumout ;
wire \Add0~18 ;
wire \Add0~21_sumout ;
wire \Add0~22 ;
wire \Add0~25_sumout ;
wire \Add0~26 ;
wire \Add0~29_sumout ;
wire \Add0~30 ;
wire \Add0~33_sumout ;
wire \Add0~34 ;
wire \Add0~37_sumout ;
wire \Add0~38 ;
wire \Add0~41_sumout ;
wire \Add0~42 ;
wire \Add0~45_sumout ;
wire \Add0~46 ;
wire \Add0~49_sumout ;
wire \Add0~50 ;
wire \Add0~53_sumout ;
wire \Add0~54 ;
wire \Add0~57_sumout ;
wire \Add0~58 ;
wire \Add0~61_sumout ;
wire \Add0~62 ;
wire \Add0~65_sumout ;
wire \Add0~66 ;
wire \Add0~69_sumout ;
wire \Add0~70 ;
wire \Add0~73_sumout ;
wire \Add0~74 ;
wire \Add0~77_sumout ;
wire \Add0~78 ;
wire \Add0~81_sumout ;
wire \Add0~82 ;
wire \Add0~85_sumout ;
wire \Add0~86 ;
wire \Add0~89_sumout ;
wire \Add0~90 ;
wire \Add0~93_sumout ;
wire \Add0~94 ;
wire \Add0~97_sumout ;
wire \Add0~98 ;
wire \Add0~101_sumout ;
wire \Add0~102 ;
wire \Add0~105_sumout ;
wire \Add0~106 ;
wire \Add0~109_sumout ;
wire \Add0~113_sumout ;
wire \Add0~114 ;
wire \Add0~117_sumout ;
wire \Add0~118 ;
wire \Add0~121_sumout ;
wire \Add0~122 ;
wire \Add0~125_sumout ;
wire \Add0~126 ;
wire \Add0~129_sumout ;
wire \Add0~130 ;
wire \Add0~133_sumout ;
wire \Add0~134 ;
wire \Add0~137_sumout ;
wire \Add0~138 ;
wire \Add0~141_sumout ;
wire \Add0~142 ;
wire \Add0~145_sumout ;
wire \Add0~146 ;
wire \Add0~149_sumout ;
wire \Add0~150 ;
wire \glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][0]~q ;


cic_auk_dspip_delay_15 \glogic:integrator_pipeline_0_generate:u1 (
	.datain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\Add0~109_sumout ,\Add0~105_sumout ,\Add0~101_sumout ,\Add0~97_sumout ,\Add0~93_sumout ,\Add0~89_sumout ,\Add0~85_sumout ,\Add0~81_sumout ,\Add0~77_sumout ,\Add0~73_sumout ,\Add0~69_sumout ,\Add0~65_sumout ,\Add0~61_sumout ,\Add0~57_sumout ,
\Add0~53_sumout ,\Add0~49_sumout ,\Add0~45_sumout ,\Add0~41_sumout ,\Add0~37_sumout ,\Add0~33_sumout ,\Add0~29_sumout ,\Add0~25_sumout ,\Add0~21_sumout ,\Add0~17_sumout ,\Add0~13_sumout ,\Add0~9_sumout ,\Add0~5_sumout ,\Add0~1_sumout ,\Add0~113_sumout ,\Add0~117_sumout ,
\Add0~121_sumout ,\Add0~125_sumout ,\Add0~129_sumout ,\Add0~133_sumout ,\Add0~137_sumout ,\Add0~141_sumout ,\Add0~145_sumout ,\Add0~149_sumout }),
	.enable(stall_reg),
	.register_fifofifo_data010(register_fifofifo_data010),
	.register_fifofifo_data011(register_fifofifo_data011),
	.register_fifofifo_data012(register_fifofifo_data012),
	.register_fifofifo_data013(register_fifofifo_data013),
	.register_fifofifo_data014(register_fifofifo_data014),
	.register_fifofifo_data015(register_fifofifo_data015),
	.register_fifofifo_data016(register_fifofifo_data016),
	.register_fifofifo_data017(register_fifofifo_data017),
	.register_fifofifo_data018(register_fifofifo_data018),
	.register_fifofifo_data019(register_fifofifo_data019),
	.register_fifofifo_data020(register_fifofifo_data020),
	.register_fifofifo_data021(register_fifofifo_data021),
	.register_fifofifo_data022(register_fifofifo_data022),
	.register_fifofifo_data023(register_fifofifo_data023),
	.register_fifofifo_data024(register_fifofifo_data024),
	.register_fifofifo_data025(register_fifofifo_data025),
	.register_fifofifo_data026(register_fifofifo_data026),
	.register_fifofifo_data027(register_fifofifo_data027),
	.register_fifofifo_data028(register_fifofifo_data028),
	.register_fifofifo_data029(register_fifofifo_data029),
	.register_fifofifo_data030(register_fifofifo_data030),
	.register_fifofifo_data031(register_fifofifo_data031),
	.register_fifofifo_data032(register_fifofifo_data032),
	.register_fifofifo_data033(register_fifofifo_data033),
	.register_fifofifo_data034(register_fifofifo_data034),
	.register_fifofifo_data035(register_fifofifo_data035),
	.register_fifofifo_data036(register_fifofifo_data036),
	.register_fifofifo_data037(register_fifofifo_data037),
	.register_fifofifo_data09(register_fifofifo_data09),
	.register_fifofifo_data08(register_fifofifo_data08),
	.register_fifofifo_data07(register_fifofifo_data07),
	.register_fifofifo_data06(register_fifofifo_data06),
	.register_fifofifo_data05(register_fifofifo_data05),
	.register_fifofifo_data04(register_fifofifo_data04),
	.register_fifofifo_data03(register_fifofifo_data03),
	.register_fifofifo_data02(register_fifofifo_data02),
	.register_fifofifo_data01(register_fifofifo_data01),
	.register_fifofifo_data00(\glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][0]~q ),
	.clk(clk),
	.reset(reset_n));

arriav_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data010),
	.datae(gnd),
	.dataf(!register_fifofifo_data0121),
	.datag(gnd),
	.cin(\Add0~114 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(\Add0~2 ),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~1 .shared_arith = "off";

arriav_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data011),
	.datae(gnd),
	.dataf(!register_fifofifo_data0131),
	.datag(gnd),
	.cin(\Add0~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~5 .shared_arith = "off";

arriav_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data012),
	.datae(gnd),
	.dataf(!register_fifofifo_data0141),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~9 .shared_arith = "off";

arriav_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data013),
	.datae(gnd),
	.dataf(!register_fifofifo_data0151),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~13 .shared_arith = "off";

arriav_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data014),
	.datae(gnd),
	.dataf(!register_fifofifo_data0161),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout());
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~17 .shared_arith = "off";

arriav_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data015),
	.datae(gnd),
	.dataf(!register_fifofifo_data0171),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout());
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~21 .shared_arith = "off";

arriav_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data016),
	.datae(gnd),
	.dataf(!register_fifofifo_data0181),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout());
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~25 .shared_arith = "off";

arriav_lcell_comb \Add0~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data017),
	.datae(gnd),
	.dataf(!register_fifofifo_data0191),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout());
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~29 .shared_arith = "off";

arriav_lcell_comb \Add0~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data018),
	.datae(gnd),
	.dataf(!register_fifofifo_data0201),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~33_sumout ),
	.cout(\Add0~34 ),
	.shareout());
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~33 .shared_arith = "off";

arriav_lcell_comb \Add0~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data019),
	.datae(gnd),
	.dataf(!register_fifofifo_data0211),
	.datag(gnd),
	.cin(\Add0~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~37_sumout ),
	.cout(\Add0~38 ),
	.shareout());
defparam \Add0~37 .extended_lut = "off";
defparam \Add0~37 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~37 .shared_arith = "off";

arriav_lcell_comb \Add0~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data020),
	.datae(gnd),
	.dataf(!register_fifofifo_data0221),
	.datag(gnd),
	.cin(\Add0~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~41_sumout ),
	.cout(\Add0~42 ),
	.shareout());
defparam \Add0~41 .extended_lut = "off";
defparam \Add0~41 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~41 .shared_arith = "off";

arriav_lcell_comb \Add0~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data021),
	.datae(gnd),
	.dataf(!register_fifofifo_data0231),
	.datag(gnd),
	.cin(\Add0~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~45_sumout ),
	.cout(\Add0~46 ),
	.shareout());
defparam \Add0~45 .extended_lut = "off";
defparam \Add0~45 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~45 .shared_arith = "off";

arriav_lcell_comb \Add0~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data022),
	.datae(gnd),
	.dataf(!register_fifofifo_data0241),
	.datag(gnd),
	.cin(\Add0~46 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~49_sumout ),
	.cout(\Add0~50 ),
	.shareout());
defparam \Add0~49 .extended_lut = "off";
defparam \Add0~49 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~49 .shared_arith = "off";

arriav_lcell_comb \Add0~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data023),
	.datae(gnd),
	.dataf(!register_fifofifo_data0251),
	.datag(gnd),
	.cin(\Add0~50 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~53_sumout ),
	.cout(\Add0~54 ),
	.shareout());
defparam \Add0~53 .extended_lut = "off";
defparam \Add0~53 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~53 .shared_arith = "off";

arriav_lcell_comb \Add0~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data024),
	.datae(gnd),
	.dataf(!register_fifofifo_data0261),
	.datag(gnd),
	.cin(\Add0~54 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~57_sumout ),
	.cout(\Add0~58 ),
	.shareout());
defparam \Add0~57 .extended_lut = "off";
defparam \Add0~57 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~57 .shared_arith = "off";

arriav_lcell_comb \Add0~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data025),
	.datae(gnd),
	.dataf(!register_fifofifo_data0271),
	.datag(gnd),
	.cin(\Add0~58 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~61_sumout ),
	.cout(\Add0~62 ),
	.shareout());
defparam \Add0~61 .extended_lut = "off";
defparam \Add0~61 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~61 .shared_arith = "off";

arriav_lcell_comb \Add0~65 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data026),
	.datae(gnd),
	.dataf(!register_fifofifo_data0281),
	.datag(gnd),
	.cin(\Add0~62 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~65_sumout ),
	.cout(\Add0~66 ),
	.shareout());
defparam \Add0~65 .extended_lut = "off";
defparam \Add0~65 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~65 .shared_arith = "off";

arriav_lcell_comb \Add0~69 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data027),
	.datae(gnd),
	.dataf(!register_fifofifo_data0291),
	.datag(gnd),
	.cin(\Add0~66 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~69_sumout ),
	.cout(\Add0~70 ),
	.shareout());
defparam \Add0~69 .extended_lut = "off";
defparam \Add0~69 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~69 .shared_arith = "off";

arriav_lcell_comb \Add0~73 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data028),
	.datae(gnd),
	.dataf(!register_fifofifo_data0301),
	.datag(gnd),
	.cin(\Add0~70 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~73_sumout ),
	.cout(\Add0~74 ),
	.shareout());
defparam \Add0~73 .extended_lut = "off";
defparam \Add0~73 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~73 .shared_arith = "off";

arriav_lcell_comb \Add0~77 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data029),
	.datae(gnd),
	.dataf(!register_fifofifo_data0311),
	.datag(gnd),
	.cin(\Add0~74 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~77_sumout ),
	.cout(\Add0~78 ),
	.shareout());
defparam \Add0~77 .extended_lut = "off";
defparam \Add0~77 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~77 .shared_arith = "off";

arriav_lcell_comb \Add0~81 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data030),
	.datae(gnd),
	.dataf(!register_fifofifo_data0321),
	.datag(gnd),
	.cin(\Add0~78 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~81_sumout ),
	.cout(\Add0~82 ),
	.shareout());
defparam \Add0~81 .extended_lut = "off";
defparam \Add0~81 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~81 .shared_arith = "off";

arriav_lcell_comb \Add0~85 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data031),
	.datae(gnd),
	.dataf(!register_fifofifo_data0331),
	.datag(gnd),
	.cin(\Add0~82 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~85_sumout ),
	.cout(\Add0~86 ),
	.shareout());
defparam \Add0~85 .extended_lut = "off";
defparam \Add0~85 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~85 .shared_arith = "off";

arriav_lcell_comb \Add0~89 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data032),
	.datae(gnd),
	.dataf(!register_fifofifo_data0341),
	.datag(gnd),
	.cin(\Add0~86 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~89_sumout ),
	.cout(\Add0~90 ),
	.shareout());
defparam \Add0~89 .extended_lut = "off";
defparam \Add0~89 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~89 .shared_arith = "off";

arriav_lcell_comb \Add0~93 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data033),
	.datae(gnd),
	.dataf(!register_fifofifo_data0351),
	.datag(gnd),
	.cin(\Add0~90 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~93_sumout ),
	.cout(\Add0~94 ),
	.shareout());
defparam \Add0~93 .extended_lut = "off";
defparam \Add0~93 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~93 .shared_arith = "off";

arriav_lcell_comb \Add0~97 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data034),
	.datae(gnd),
	.dataf(!register_fifofifo_data0361),
	.datag(gnd),
	.cin(\Add0~94 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~97_sumout ),
	.cout(\Add0~98 ),
	.shareout());
defparam \Add0~97 .extended_lut = "off";
defparam \Add0~97 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~97 .shared_arith = "off";

arriav_lcell_comb \Add0~101 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data035),
	.datae(gnd),
	.dataf(!register_fifofifo_data0371),
	.datag(gnd),
	.cin(\Add0~98 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~101_sumout ),
	.cout(\Add0~102 ),
	.shareout());
defparam \Add0~101 .extended_lut = "off";
defparam \Add0~101 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~101 .shared_arith = "off";

arriav_lcell_comb \Add0~105 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data036),
	.datae(gnd),
	.dataf(!register_fifofifo_data038),
	.datag(gnd),
	.cin(\Add0~102 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~105_sumout ),
	.cout(\Add0~106 ),
	.shareout());
defparam \Add0~105 .extended_lut = "off";
defparam \Add0~105 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~105 .shared_arith = "off";

arriav_lcell_comb \Add0~109 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data037),
	.datae(gnd),
	.dataf(!register_fifofifo_data039),
	.datag(gnd),
	.cin(\Add0~106 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~109_sumout ),
	.cout(),
	.shareout());
defparam \Add0~109 .extended_lut = "off";
defparam \Add0~109 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~109 .shared_arith = "off";

arriav_lcell_comb \Add0~113 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data09),
	.datae(gnd),
	.dataf(!register_fifofifo_data0111),
	.datag(gnd),
	.cin(\Add0~118 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~113_sumout ),
	.cout(\Add0~114 ),
	.shareout());
defparam \Add0~113 .extended_lut = "off";
defparam \Add0~113 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~113 .shared_arith = "off";

arriav_lcell_comb \Add0~117 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data08),
	.datae(gnd),
	.dataf(!register_fifofifo_data0101),
	.datag(gnd),
	.cin(\Add0~122 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~117_sumout ),
	.cout(\Add0~118 ),
	.shareout());
defparam \Add0~117 .extended_lut = "off";
defparam \Add0~117 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~117 .shared_arith = "off";

arriav_lcell_comb \Add0~121 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data07),
	.datae(gnd),
	.dataf(!register_fifofifo_data091),
	.datag(gnd),
	.cin(\Add0~126 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~121_sumout ),
	.cout(\Add0~122 ),
	.shareout());
defparam \Add0~121 .extended_lut = "off";
defparam \Add0~121 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~121 .shared_arith = "off";

arriav_lcell_comb \Add0~125 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data06),
	.datae(gnd),
	.dataf(!register_fifofifo_data081),
	.datag(gnd),
	.cin(\Add0~130 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~125_sumout ),
	.cout(\Add0~126 ),
	.shareout());
defparam \Add0~125 .extended_lut = "off";
defparam \Add0~125 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~125 .shared_arith = "off";

arriav_lcell_comb \Add0~129 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data05),
	.datae(gnd),
	.dataf(!register_fifofifo_data071),
	.datag(gnd),
	.cin(\Add0~134 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~129_sumout ),
	.cout(\Add0~130 ),
	.shareout());
defparam \Add0~129 .extended_lut = "off";
defparam \Add0~129 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~129 .shared_arith = "off";

arriav_lcell_comb \Add0~133 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data04),
	.datae(gnd),
	.dataf(!register_fifofifo_data061),
	.datag(gnd),
	.cin(\Add0~138 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~133_sumout ),
	.cout(\Add0~134 ),
	.shareout());
defparam \Add0~133 .extended_lut = "off";
defparam \Add0~133 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~133 .shared_arith = "off";

arriav_lcell_comb \Add0~137 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data03),
	.datae(gnd),
	.dataf(!register_fifofifo_data051),
	.datag(gnd),
	.cin(\Add0~142 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~137_sumout ),
	.cout(\Add0~138 ),
	.shareout());
defparam \Add0~137 .extended_lut = "off";
defparam \Add0~137 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~137 .shared_arith = "off";

arriav_lcell_comb \Add0~141 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data02),
	.datae(gnd),
	.dataf(!register_fifofifo_data041),
	.datag(gnd),
	.cin(\Add0~146 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~141_sumout ),
	.cout(\Add0~142 ),
	.shareout());
defparam \Add0~141 .extended_lut = "off";
defparam \Add0~141 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~141 .shared_arith = "off";

arriav_lcell_comb \Add0~145 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!register_fifofifo_data01),
	.datae(gnd),
	.dataf(!register_fifofifo_data0310),
	.datag(gnd),
	.cin(\Add0~150 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~145_sumout ),
	.cout(\Add0~146 ),
	.shareout());
defparam \Add0~145 .extended_lut = "off";
defparam \Add0~145 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~145 .shared_arith = "off";

arriav_lcell_comb \Add0~149 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][0]~q ),
	.datae(gnd),
	.dataf(!register_fifofifo_data0210),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~149_sumout ),
	.cout(\Add0~150 ),
	.shareout());
defparam \Add0~149 .extended_lut = "off";
defparam \Add0~149 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~149 .shared_arith = "off";

endmodule

module cic_auk_dspip_delay_15 (
	datain,
	enable,
	register_fifofifo_data010,
	register_fifofifo_data011,
	register_fifofifo_data012,
	register_fifofifo_data013,
	register_fifofifo_data014,
	register_fifofifo_data015,
	register_fifofifo_data016,
	register_fifofifo_data017,
	register_fifofifo_data018,
	register_fifofifo_data019,
	register_fifofifo_data020,
	register_fifofifo_data021,
	register_fifofifo_data022,
	register_fifofifo_data023,
	register_fifofifo_data024,
	register_fifofifo_data025,
	register_fifofifo_data026,
	register_fifofifo_data027,
	register_fifofifo_data028,
	register_fifofifo_data029,
	register_fifofifo_data030,
	register_fifofifo_data031,
	register_fifofifo_data032,
	register_fifofifo_data033,
	register_fifofifo_data034,
	register_fifofifo_data035,
	register_fifofifo_data036,
	register_fifofifo_data037,
	register_fifofifo_data09,
	register_fifofifo_data08,
	register_fifofifo_data07,
	register_fifofifo_data06,
	register_fifofifo_data05,
	register_fifofifo_data04,
	register_fifofifo_data03,
	register_fifofifo_data02,
	register_fifofifo_data01,
	register_fifofifo_data00,
	clk,
	reset)/* synthesis synthesis_greybox=1 */;
input 	[46:0] datain;
input 	enable;
output 	register_fifofifo_data010;
output 	register_fifofifo_data011;
output 	register_fifofifo_data012;
output 	register_fifofifo_data013;
output 	register_fifofifo_data014;
output 	register_fifofifo_data015;
output 	register_fifofifo_data016;
output 	register_fifofifo_data017;
output 	register_fifofifo_data018;
output 	register_fifofifo_data019;
output 	register_fifofifo_data020;
output 	register_fifofifo_data021;
output 	register_fifofifo_data022;
output 	register_fifofifo_data023;
output 	register_fifofifo_data024;
output 	register_fifofifo_data025;
output 	register_fifofifo_data026;
output 	register_fifofifo_data027;
output 	register_fifofifo_data028;
output 	register_fifofifo_data029;
output 	register_fifofifo_data030;
output 	register_fifofifo_data031;
output 	register_fifofifo_data032;
output 	register_fifofifo_data033;
output 	register_fifofifo_data034;
output 	register_fifofifo_data035;
output 	register_fifofifo_data036;
output 	register_fifofifo_data037;
output 	register_fifofifo_data09;
output 	register_fifofifo_data08;
output 	register_fifofifo_data07;
output 	register_fifofifo_data06;
output 	register_fifofifo_data05;
output 	register_fifofifo_data04;
output 	register_fifofifo_data03;
output 	register_fifofifo_data02;
output 	register_fifofifo_data01;
output 	register_fifofifo_data00;
input 	clk;
input 	reset;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \register_fifo:fifo_data[0][10] (
	.clk(clk),
	.d(datain[10]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data010),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][10] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][10] .power_up = "low";

dffeas \register_fifo:fifo_data[0][11] (
	.clk(clk),
	.d(datain[11]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data011),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][11] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][11] .power_up = "low";

dffeas \register_fifo:fifo_data[0][12] (
	.clk(clk),
	.d(datain[12]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data012),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][12] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][12] .power_up = "low";

dffeas \register_fifo:fifo_data[0][13] (
	.clk(clk),
	.d(datain[13]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data013),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][13] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][13] .power_up = "low";

dffeas \register_fifo:fifo_data[0][14] (
	.clk(clk),
	.d(datain[14]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data014),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][14] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][14] .power_up = "low";

dffeas \register_fifo:fifo_data[0][15] (
	.clk(clk),
	.d(datain[15]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data015),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][15] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][15] .power_up = "low";

dffeas \register_fifo:fifo_data[0][16] (
	.clk(clk),
	.d(datain[16]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data016),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][16] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][16] .power_up = "low";

dffeas \register_fifo:fifo_data[0][17] (
	.clk(clk),
	.d(datain[17]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data017),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][17] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][17] .power_up = "low";

dffeas \register_fifo:fifo_data[0][18] (
	.clk(clk),
	.d(datain[18]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data018),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][18] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][18] .power_up = "low";

dffeas \register_fifo:fifo_data[0][19] (
	.clk(clk),
	.d(datain[19]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data019),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][19] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][19] .power_up = "low";

dffeas \register_fifo:fifo_data[0][20] (
	.clk(clk),
	.d(datain[20]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data020),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][20] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][20] .power_up = "low";

dffeas \register_fifo:fifo_data[0][21] (
	.clk(clk),
	.d(datain[21]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data021),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][21] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][21] .power_up = "low";

dffeas \register_fifo:fifo_data[0][22] (
	.clk(clk),
	.d(datain[22]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data022),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][22] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][22] .power_up = "low";

dffeas \register_fifo:fifo_data[0][23] (
	.clk(clk),
	.d(datain[23]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data023),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][23] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][23] .power_up = "low";

dffeas \register_fifo:fifo_data[0][24] (
	.clk(clk),
	.d(datain[24]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data024),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][24] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][24] .power_up = "low";

dffeas \register_fifo:fifo_data[0][25] (
	.clk(clk),
	.d(datain[25]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data025),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][25] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][25] .power_up = "low";

dffeas \register_fifo:fifo_data[0][26] (
	.clk(clk),
	.d(datain[26]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data026),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][26] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][26] .power_up = "low";

dffeas \register_fifo:fifo_data[0][27] (
	.clk(clk),
	.d(datain[27]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data027),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][27] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][27] .power_up = "low";

dffeas \register_fifo:fifo_data[0][28] (
	.clk(clk),
	.d(datain[28]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data028),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][28] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][28] .power_up = "low";

dffeas \register_fifo:fifo_data[0][29] (
	.clk(clk),
	.d(datain[29]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data029),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][29] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][29] .power_up = "low";

dffeas \register_fifo:fifo_data[0][30] (
	.clk(clk),
	.d(datain[30]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data030),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][30] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][30] .power_up = "low";

dffeas \register_fifo:fifo_data[0][31] (
	.clk(clk),
	.d(datain[31]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data031),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][31] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][31] .power_up = "low";

dffeas \register_fifo:fifo_data[0][32] (
	.clk(clk),
	.d(datain[32]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data032),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][32] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][32] .power_up = "low";

dffeas \register_fifo:fifo_data[0][33] (
	.clk(clk),
	.d(datain[33]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data033),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][33] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][33] .power_up = "low";

dffeas \register_fifo:fifo_data[0][34] (
	.clk(clk),
	.d(datain[34]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data034),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][34] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][34] .power_up = "low";

dffeas \register_fifo:fifo_data[0][35] (
	.clk(clk),
	.d(datain[35]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data035),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][35] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][35] .power_up = "low";

dffeas \register_fifo:fifo_data[0][36] (
	.clk(clk),
	.d(datain[36]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data036),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][36] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][36] .power_up = "low";

dffeas \register_fifo:fifo_data[0][37] (
	.clk(clk),
	.d(datain[37]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data037),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][37] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][37] .power_up = "low";

dffeas \register_fifo:fifo_data[0][9] (
	.clk(clk),
	.d(datain[9]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data09),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][9] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][9] .power_up = "low";

dffeas \register_fifo:fifo_data[0][8] (
	.clk(clk),
	.d(datain[8]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data08),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][8] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][8] .power_up = "low";

dffeas \register_fifo:fifo_data[0][7] (
	.clk(clk),
	.d(datain[7]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data07),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][7] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][7] .power_up = "low";

dffeas \register_fifo:fifo_data[0][6] (
	.clk(clk),
	.d(datain[6]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data06),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][6] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][6] .power_up = "low";

dffeas \register_fifo:fifo_data[0][5] (
	.clk(clk),
	.d(datain[5]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data05),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][5] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][5] .power_up = "low";

dffeas \register_fifo:fifo_data[0][4] (
	.clk(clk),
	.d(datain[4]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data04),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][4] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][4] .power_up = "low";

dffeas \register_fifo:fifo_data[0][3] (
	.clk(clk),
	.d(datain[3]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data03),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][3] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][3] .power_up = "low";

dffeas \register_fifo:fifo_data[0][2] (
	.clk(clk),
	.d(datain[2]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data02),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][2] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][2] .power_up = "low";

dffeas \register_fifo:fifo_data[0][1] (
	.clk(clk),
	.d(datain[1]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data01),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][1] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][1] .power_up = "low";

dffeas \register_fifo:fifo_data[0][0] (
	.clk(clk),
	.d(datain[0]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data00),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][0] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][0] .power_up = "low";

endmodule

module cic_counter_module_3 (
	stall_reg,
	count_0,
	count_1,
	count_2,
	count_3,
	count_4,
	Equal0,
	sample_state,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	stall_reg;
output 	count_0;
output 	count_1;
output 	count_2;
output 	count_3;
output 	count_4;
output 	Equal0;
input 	sample_state;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \count[0]~0_combout ;
wire \count[1]~1_combout ;
wire \count[2]~4_combout ;
wire \count[3]~2_combout ;
wire \Add0~0_combout ;
wire \count[4]~3_combout ;


dffeas \count[0] (
	.clk(clk),
	.d(\count[0]~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(count_0),
	.prn(vcc));
defparam \count[0] .is_wysiwyg = "true";
defparam \count[0] .power_up = "low";

dffeas \count[1] (
	.clk(clk),
	.d(\count[1]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(count_1),
	.prn(vcc));
defparam \count[1] .is_wysiwyg = "true";
defparam \count[1] .power_up = "low";

dffeas \count[2] (
	.clk(clk),
	.d(\count[2]~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(count_2),
	.prn(vcc));
defparam \count[2] .is_wysiwyg = "true";
defparam \count[2] .power_up = "low";

dffeas \count[3] (
	.clk(clk),
	.d(\count[3]~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(count_3),
	.prn(vcc));
defparam \count[3] .is_wysiwyg = "true";
defparam \count[3] .power_up = "low";

dffeas \count[4] (
	.clk(clk),
	.d(\count[4]~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(count_4),
	.prn(vcc));
defparam \count[4] .is_wysiwyg = "true";
defparam \count[4] .power_up = "low";

arriav_lcell_comb \Equal0~0 (
	.dataa(!count_1),
	.datab(!count_2),
	.datac(!count_3),
	.datad(!count_4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Equal0),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~0 .extended_lut = "off";
defparam \Equal0~0 .lut_mask = 64'hFEFFFEFFFEFFFEFF;
defparam \Equal0~0 .shared_arith = "off";

arriav_lcell_comb \count[0]~0 (
	.dataa(!reset_n),
	.datab(!stall_reg),
	.datac(!count_0),
	.datad(!Equal0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\count[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \count[0]~0 .extended_lut = "off";
defparam \count[0]~0 .lut_mask = 64'hFF7DFF7DFF7DFF7D;
defparam \count[0]~0 .shared_arith = "off";

arriav_lcell_comb \count[1]~1 (
	.dataa(!reset_n),
	.datab(!stall_reg),
	.datac(!count_0),
	.datad(!count_1),
	.datae(!Equal0),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\count[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \count[1]~1 .extended_lut = "off";
defparam \count[1]~1 .lut_mask = 64'hFFFFD77DFFFFD77D;
defparam \count[1]~1 .shared_arith = "off";

arriav_lcell_comb \count[2]~4 (
	.dataa(!count_2),
	.datab(!count_1),
	.datac(!count_0),
	.datad(!stall_reg),
	.datae(!reset_n),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\count[2]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \count[2]~4 .extended_lut = "off";
defparam \count[2]~4 .lut_mask = 64'h6996FFFF6996FFFF;
defparam \count[2]~4 .shared_arith = "off";

arriav_lcell_comb \count[3]~2 (
	.dataa(!reset_n),
	.datab(!stall_reg),
	.datac(!count_0),
	.datad(!count_3),
	.datae(!Equal0),
	.dataf(!sample_state),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\count[3]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \count[3]~2 .extended_lut = "off";
defparam \count[3]~2 .lut_mask = 64'hF7FDFDF7FDF7F7FD;
defparam \count[3]~2 .shared_arith = "off";

arriav_lcell_comb \Add0~0 (
	.dataa(!count_3),
	.datab(!sample_state),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~0 .extended_lut = "off";
defparam \Add0~0 .lut_mask = 64'h7777777777777777;
defparam \Add0~0 .shared_arith = "off";

arriav_lcell_comb \count[4]~3 (
	.dataa(!reset_n),
	.datab(!stall_reg),
	.datac(!count_0),
	.datad(!count_4),
	.datae(!Equal0),
	.dataf(!\Add0~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\count[4]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \count[4]~3 .extended_lut = "off";
defparam \count[4]~3 .lut_mask = 64'hF7FDFDF7FDF7F7FD;
defparam \count[4]~3 .shared_arith = "off";

endmodule

module cic_auk_dspip_avalon_streaming_controller (
	rd_addr_ptr_2,
	dffe_nae,
	dffe_af,
	Equal2,
	Mux0,
	sink_ready_ctrl,
	usedw_process,
	stall_reg1,
	sink_ready_ctrl1,
	sink_ready_ctrl2,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	rd_addr_ptr_2;
input 	dffe_nae;
input 	dffe_af;
output 	Equal2;
output 	Mux0;
output 	sink_ready_ctrl;
output 	usedw_process;
output 	stall_reg1;
output 	sink_ready_ctrl1;
output 	sink_ready_ctrl2;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \ready_FIFO|fifo_array[4][0]~q ;
wire \ready_FIFO|fifo_array[5][0]~q ;
wire \ready_FIFO|rd_addr_ptr[0]~q ;
wire \ready_FIFO|rd_addr_ptr[1]~q ;
wire \stall_reg~0_combout ;


cic_auk_dspip_avalon_streaming_small_fifo ready_FIFO(
	.rd_addr_ptr_2(rd_addr_ptr_2),
	.fifo_array_0_4(\ready_FIFO|fifo_array[4][0]~q ),
	.fifo_array_0_5(\ready_FIFO|fifo_array[5][0]~q ),
	.dffe_nae(dffe_nae),
	.dffe_af(dffe_af),
	.Equal2(Equal2),
	.rd_addr_ptr_0(\ready_FIFO|rd_addr_ptr[0]~q ),
	.rd_addr_ptr_1(\ready_FIFO|rd_addr_ptr[1]~q ),
	.Mux0(Mux0),
	.usedw_process(usedw_process),
	.stall_reg(stall_reg1),
	.clock(clk),
	.reset_n(reset_n));

arriav_lcell_comb \sink_ready_ctrl~0 (
	.dataa(!\ready_FIFO|rd_addr_ptr[0]~q ),
	.datab(!\ready_FIFO|rd_addr_ptr[1]~q ),
	.datac(!rd_addr_ptr_2),
	.datad(!\ready_FIFO|fifo_array[4][0]~q ),
	.datae(!\ready_FIFO|fifo_array[5][0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(sink_ready_ctrl),
	.sumout(),
	.cout(),
	.shareout());
defparam \sink_ready_ctrl~0 .extended_lut = "off";
defparam \sink_ready_ctrl~0 .lut_mask = 64'h8DFFFFFF8DFFFFFF;
defparam \sink_ready_ctrl~0 .shared_arith = "off";

dffeas stall_reg(
	.clk(clk),
	.d(\stall_reg~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(stall_reg1),
	.prn(vcc));
defparam stall_reg.is_wysiwyg = "true";
defparam stall_reg.power_up = "low";

arriav_lcell_comb \sink_ready_ctrl~1 (
	.dataa(!Equal2),
	.datab(!Mux0),
	.datac(!rd_addr_ptr_2),
	.datad(!sink_ready_ctrl),
	.datae(!usedw_process),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(sink_ready_ctrl1),
	.sumout(),
	.cout(),
	.shareout());
defparam \sink_ready_ctrl~1 .extended_lut = "off";
defparam \sink_ready_ctrl~1 .lut_mask = 64'hF7FFFFFFF7FFFFFF;
defparam \sink_ready_ctrl~1 .shared_arith = "off";

arriav_lcell_comb \sink_ready_ctrl~2 (
	.dataa(!Equal2),
	.datab(!\ready_FIFO|rd_addr_ptr[0]~q ),
	.datac(!\ready_FIFO|rd_addr_ptr[1]~q ),
	.datad(!rd_addr_ptr_2),
	.datae(!\ready_FIFO|fifo_array[4][0]~q ),
	.dataf(!\ready_FIFO|fifo_array[5][0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(sink_ready_ctrl2),
	.sumout(),
	.cout(),
	.shareout());
defparam \sink_ready_ctrl~2 .extended_lut = "off";
defparam \sink_ready_ctrl~2 .lut_mask = 64'hFFFFFFFFFFFFBF8F;
defparam \sink_ready_ctrl~2 .shared_arith = "off";

arriav_lcell_comb \stall_reg~0 (
	.dataa(!dffe_nae),
	.datab(!dffe_af),
	.datac(!reset_n),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\stall_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \stall_reg~0 .extended_lut = "off";
defparam \stall_reg~0 .lut_mask = 64'hFBFBFBFBFBFBFBFB;
defparam \stall_reg~0 .shared_arith = "off";

endmodule

module cic_auk_dspip_avalon_streaming_small_fifo (
	rd_addr_ptr_2,
	fifo_array_0_4,
	fifo_array_0_5,
	dffe_nae,
	dffe_af,
	Equal2,
	rd_addr_ptr_0,
	rd_addr_ptr_1,
	Mux0,
	usedw_process,
	stall_reg,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	rd_addr_ptr_2;
output 	fifo_array_0_4;
output 	fifo_array_0_5;
input 	dffe_nae;
input 	dffe_af;
output 	Equal2;
output 	rd_addr_ptr_0;
output 	rd_addr_ptr_1;
output 	Mux0;
output 	usedw_process;
input 	stall_reg;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \rd_addr_ptr~3_combout ;
wire \fifo_usedw[1]~2_combout ;
wire \fifo_usedw[1]~q ;
wire \usedw_process~1_combout ;
wire \fifo_usedw[0]~1_combout ;
wire \fifo_usedw[0]~q ;
wire \fifo_usedw[2]~0_combout ;
wire \fifo_usedw[2]~q ;
wire \rd_addr_ptr[2]~1_combout ;
wire \usedw_process~2_combout ;
wire \wr_addr_ptr~2_combout ;
wire \wr_addr_ptr[2]~1_combout ;
wire \wr_addr_ptr[0]~q ;
wire \wr_addr_ptr~3_combout ;
wire \wr_addr_ptr[1]~q ;
wire \wr_addr_ptr~0_combout ;
wire \wr_addr_ptr[2]~q ;
wire \fifo_array~4_combout ;
wire \fifo_array~5_combout ;
wire \rd_addr_ptr~0_combout ;
wire \rd_addr_ptr~2_combout ;
wire \fifo_array~0_combout ;
wire \fifo_array[0][0]~q ;
wire \fifo_array~1_combout ;
wire \fifo_array[1][0]~q ;
wire \fifo_array~2_combout ;
wire \fifo_array[2][0]~q ;
wire \fifo_array~3_combout ;
wire \fifo_array[3][0]~q ;


dffeas \rd_addr_ptr[2] (
	.clk(clock),
	.d(\rd_addr_ptr~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\rd_addr_ptr[2]~1_combout ),
	.q(rd_addr_ptr_2),
	.prn(vcc));
defparam \rd_addr_ptr[2] .is_wysiwyg = "true";
defparam \rd_addr_ptr[2] .power_up = "low";

dffeas \fifo_array[4][0] (
	.clk(clock),
	.d(\fifo_array~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(vcc),
	.q(fifo_array_0_4),
	.prn(vcc));
defparam \fifo_array[4][0] .is_wysiwyg = "true";
defparam \fifo_array[4][0] .power_up = "low";

dffeas \fifo_array[5][0] (
	.clk(clock),
	.d(\fifo_array~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(vcc),
	.q(fifo_array_0_5),
	.prn(vcc));
defparam \fifo_array[5][0] .is_wysiwyg = "true";
defparam \fifo_array[5][0] .power_up = "low";

arriav_lcell_comb \Equal2~0 (
	.dataa(!\fifo_usedw[2]~q ),
	.datab(!\fifo_usedw[0]~q ),
	.datac(!\fifo_usedw[1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Equal2),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal2~0 .extended_lut = "off";
defparam \Equal2~0 .lut_mask = 64'hFEFEFEFEFEFEFEFE;
defparam \Equal2~0 .shared_arith = "off";

dffeas \rd_addr_ptr[0] (
	.clk(clock),
	.d(\rd_addr_ptr~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\rd_addr_ptr[2]~1_combout ),
	.q(rd_addr_ptr_0),
	.prn(vcc));
defparam \rd_addr_ptr[0] .is_wysiwyg = "true";
defparam \rd_addr_ptr[0] .power_up = "low";

dffeas \rd_addr_ptr[1] (
	.clk(clock),
	.d(\rd_addr_ptr~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\rd_addr_ptr[2]~1_combout ),
	.q(rd_addr_ptr_1),
	.prn(vcc));
defparam \rd_addr_ptr[1] .is_wysiwyg = "true";
defparam \rd_addr_ptr[1] .power_up = "low";

arriav_lcell_comb \Mux0~0 (
	.dataa(!\fifo_array[0][0]~q ),
	.datab(!\fifo_array[1][0]~q ),
	.datac(!\fifo_array[2][0]~q ),
	.datad(!\fifo_array[3][0]~q ),
	.datae(!rd_addr_ptr_0),
	.dataf(!rd_addr_ptr_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Mux0),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux0~0 .extended_lut = "off";
defparam \Mux0~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux0~0 .shared_arith = "off";

arriav_lcell_comb \usedw_process~0 (
	.dataa(!dffe_nae),
	.datab(!dffe_af),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(usedw_process),
	.sumout(),
	.cout(),
	.shareout());
defparam \usedw_process~0 .extended_lut = "off";
defparam \usedw_process~0 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \usedw_process~0 .shared_arith = "off";

arriav_lcell_comb \rd_addr_ptr~3 (
	.dataa(!rd_addr_ptr_0),
	.datab(!rd_addr_ptr_1),
	.datac(!rd_addr_ptr_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rd_addr_ptr~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rd_addr_ptr~3 .extended_lut = "off";
defparam \rd_addr_ptr~3 .lut_mask = 64'h7B7B7B7B7B7B7B7B;
defparam \rd_addr_ptr~3 .shared_arith = "off";

arriav_lcell_comb \fifo_usedw[1]~2 (
	.dataa(!\fifo_usedw[2]~q ),
	.datab(!\fifo_usedw[0]~q ),
	.datac(!\fifo_usedw[1]~q ),
	.datad(!usedw_process),
	.datae(!reset_n),
	.dataf(!stall_reg),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fifo_usedw[1]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fifo_usedw[1]~2 .extended_lut = "off";
defparam \fifo_usedw[1]~2 .lut_mask = 64'h9669FFFF6996FFFF;
defparam \fifo_usedw[1]~2 .shared_arith = "off";

dffeas \fifo_usedw[1] (
	.clk(clock),
	.d(\fifo_usedw[1]~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\fifo_usedw[1]~q ),
	.prn(vcc));
defparam \fifo_usedw[1] .is_wysiwyg = "true";
defparam \fifo_usedw[1] .power_up = "low";

arriav_lcell_comb \usedw_process~1 (
	.dataa(!\fifo_usedw[2]~q ),
	.datab(!\fifo_usedw[0]~q ),
	.datac(!\fifo_usedw[1]~q ),
	.datad(!stall_reg),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\usedw_process~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \usedw_process~1 .extended_lut = "off";
defparam \usedw_process~1 .lut_mask = 64'hFFFBFFFBFFFBFFFB;
defparam \usedw_process~1 .shared_arith = "off";

arriav_lcell_comb \fifo_usedw[0]~1 (
	.dataa(!\fifo_usedw[0]~q ),
	.datab(!Equal2),
	.datac(!dffe_nae),
	.datad(!dffe_af),
	.datae(!reset_n),
	.dataf(!\usedw_process~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fifo_usedw[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fifo_usedw[0]~1 .extended_lut = "off";
defparam \fifo_usedw[0]~1 .lut_mask = 64'h9669FFFF6996FFFF;
defparam \fifo_usedw[0]~1 .shared_arith = "off";

dffeas \fifo_usedw[0] (
	.clk(clock),
	.d(\fifo_usedw[0]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\fifo_usedw[0]~q ),
	.prn(vcc));
defparam \fifo_usedw[0] .is_wysiwyg = "true";
defparam \fifo_usedw[0] .power_up = "low";

arriav_lcell_comb \fifo_usedw[2]~0 (
	.dataa(!\fifo_usedw[2]~q ),
	.datab(!\fifo_usedw[0]~q ),
	.datac(!\fifo_usedw[1]~q ),
	.datad(!usedw_process),
	.datae(!reset_n),
	.dataf(!stall_reg),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fifo_usedw[2]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fifo_usedw[2]~0 .extended_lut = "off";
defparam \fifo_usedw[2]~0 .lut_mask = 64'h9669FFFF6996FFFF;
defparam \fifo_usedw[2]~0 .shared_arith = "off";

dffeas \fifo_usedw[2] (
	.clk(clock),
	.d(\fifo_usedw[2]~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\fifo_usedw[2]~q ),
	.prn(vcc));
defparam \fifo_usedw[2] .is_wysiwyg = "true";
defparam \fifo_usedw[2] .power_up = "low";

arriav_lcell_comb \rd_addr_ptr[2]~1 (
	.dataa(!\fifo_usedw[2]~q ),
	.datab(!\fifo_usedw[0]~q ),
	.datac(!\fifo_usedw[1]~q ),
	.datad(!dffe_nae),
	.datae(!dffe_af),
	.dataf(!reset_n),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rd_addr_ptr[2]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rd_addr_ptr[2]~1 .extended_lut = "off";
defparam \rd_addr_ptr[2]~1 .lut_mask = 64'hFFFFFFFFFFFF7FFF;
defparam \rd_addr_ptr[2]~1 .shared_arith = "off";

arriav_lcell_comb \usedw_process~2 (
	.dataa(!\fifo_usedw[2]~q ),
	.datab(!\fifo_usedw[0]~q ),
	.datac(!\fifo_usedw[1]~q ),
	.datad(!dffe_nae),
	.datae(!dffe_af),
	.dataf(!stall_reg),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\usedw_process~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \usedw_process~2 .extended_lut = "off";
defparam \usedw_process~2 .lut_mask = 64'hFFFFFFFFFF7BFFFF;
defparam \usedw_process~2 .shared_arith = "off";

arriav_lcell_comb \wr_addr_ptr~2 (
	.dataa(!reset_n),
	.datab(!\wr_addr_ptr[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wr_addr_ptr~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wr_addr_ptr~2 .extended_lut = "off";
defparam \wr_addr_ptr~2 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \wr_addr_ptr~2 .shared_arith = "off";

arriav_lcell_comb \wr_addr_ptr[2]~1 (
	.dataa(!Equal2),
	.datab(!dffe_nae),
	.datac(!dffe_af),
	.datad(!reset_n),
	.datae(!\usedw_process~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wr_addr_ptr[2]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wr_addr_ptr[2]~1 .extended_lut = "off";
defparam \wr_addr_ptr[2]~1 .lut_mask = 64'hFFEFFFFFFFEFFFFF;
defparam \wr_addr_ptr[2]~1 .shared_arith = "off";

dffeas \wr_addr_ptr[0] (
	.clk(clock),
	.d(\wr_addr_ptr~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_addr_ptr[2]~1_combout ),
	.q(\wr_addr_ptr[0]~q ),
	.prn(vcc));
defparam \wr_addr_ptr[0] .is_wysiwyg = "true";
defparam \wr_addr_ptr[0] .power_up = "low";

arriav_lcell_comb \wr_addr_ptr~3 (
	.dataa(!reset_n),
	.datab(!\wr_addr_ptr[2]~q ),
	.datac(!\wr_addr_ptr[0]~q ),
	.datad(!\wr_addr_ptr[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wr_addr_ptr~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wr_addr_ptr~3 .extended_lut = "off";
defparam \wr_addr_ptr~3 .lut_mask = 64'hDFFDDFFDDFFDDFFD;
defparam \wr_addr_ptr~3 .shared_arith = "off";

dffeas \wr_addr_ptr[1] (
	.clk(clock),
	.d(\wr_addr_ptr~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_addr_ptr[2]~1_combout ),
	.q(\wr_addr_ptr[1]~q ),
	.prn(vcc));
defparam \wr_addr_ptr[1] .is_wysiwyg = "true";
defparam \wr_addr_ptr[1] .power_up = "low";

arriav_lcell_comb \wr_addr_ptr~0 (
	.dataa(!\wr_addr_ptr[2]~q ),
	.datab(!\wr_addr_ptr[0]~q ),
	.datac(!\wr_addr_ptr[1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wr_addr_ptr~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wr_addr_ptr~0 .extended_lut = "off";
defparam \wr_addr_ptr~0 .lut_mask = 64'h6F6F6F6F6F6F6F6F;
defparam \wr_addr_ptr~0 .shared_arith = "off";

dffeas \wr_addr_ptr[2] (
	.clk(clock),
	.d(\wr_addr_ptr~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\wr_addr_ptr[2]~1_combout ),
	.q(\wr_addr_ptr[2]~q ),
	.prn(vcc));
defparam \wr_addr_ptr[2] .is_wysiwyg = "true";
defparam \wr_addr_ptr[2] .power_up = "low";

arriav_lcell_comb \fifo_array~4 (
	.dataa(!fifo_array_0_4),
	.datab(!\usedw_process~2_combout ),
	.datac(!\wr_addr_ptr[2]~q ),
	.datad(!\wr_addr_ptr[0]~q ),
	.datae(!\wr_addr_ptr[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fifo_array~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fifo_array~4 .extended_lut = "off";
defparam \fifo_array~4 .lut_mask = 64'hFFFFFF7FFFFFFF7F;
defparam \fifo_array~4 .shared_arith = "off";

arriav_lcell_comb \fifo_array~5 (
	.dataa(!fifo_array_0_5),
	.datab(!\usedw_process~2_combout ),
	.datac(!\wr_addr_ptr[2]~q ),
	.datad(!\wr_addr_ptr[0]~q ),
	.datae(!\wr_addr_ptr[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fifo_array~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fifo_array~5 .extended_lut = "off";
defparam \fifo_array~5 .lut_mask = 64'hFFFF7FFFFFFF7FFF;
defparam \fifo_array~5 .shared_arith = "off";

arriav_lcell_comb \rd_addr_ptr~0 (
	.dataa(!rd_addr_ptr_0),
	.datab(!reset_n),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rd_addr_ptr~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rd_addr_ptr~0 .extended_lut = "off";
defparam \rd_addr_ptr~0 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \rd_addr_ptr~0 .shared_arith = "off";

arriav_lcell_comb \rd_addr_ptr~2 (
	.dataa(!rd_addr_ptr_0),
	.datab(!rd_addr_ptr_1),
	.datac(!rd_addr_ptr_2),
	.datad(!reset_n),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rd_addr_ptr~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rd_addr_ptr~2 .extended_lut = "off";
defparam \rd_addr_ptr~2 .lut_mask = 64'hF6FFF6FFF6FFF6FF;
defparam \rd_addr_ptr~2 .shared_arith = "off";

arriav_lcell_comb \fifo_array~0 (
	.dataa(!\fifo_array[0][0]~q ),
	.datab(!\usedw_process~2_combout ),
	.datac(!\wr_addr_ptr[2]~q ),
	.datad(!\wr_addr_ptr[0]~q ),
	.datae(!\wr_addr_ptr[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fifo_array~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fifo_array~0 .extended_lut = "off";
defparam \fifo_array~0 .lut_mask = 64'hFFFFFFF7FFFFFFF7;
defparam \fifo_array~0 .shared_arith = "off";

dffeas \fifo_array[0][0] (
	.clk(clock),
	.d(\fifo_array~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(vcc),
	.q(\fifo_array[0][0]~q ),
	.prn(vcc));
defparam \fifo_array[0][0] .is_wysiwyg = "true";
defparam \fifo_array[0][0] .power_up = "low";

arriav_lcell_comb \fifo_array~1 (
	.dataa(!\fifo_array[1][0]~q ),
	.datab(!\usedw_process~2_combout ),
	.datac(!\wr_addr_ptr[2]~q ),
	.datad(!\wr_addr_ptr[0]~q ),
	.datae(!\wr_addr_ptr[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fifo_array~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fifo_array~1 .extended_lut = "off";
defparam \fifo_array~1 .lut_mask = 64'hFFFFF7FFFFFFF7FF;
defparam \fifo_array~1 .shared_arith = "off";

dffeas \fifo_array[1][0] (
	.clk(clock),
	.d(\fifo_array~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(vcc),
	.q(\fifo_array[1][0]~q ),
	.prn(vcc));
defparam \fifo_array[1][0] .is_wysiwyg = "true";
defparam \fifo_array[1][0] .power_up = "low";

arriav_lcell_comb \fifo_array~2 (
	.dataa(!\fifo_array[2][0]~q ),
	.datab(!\usedw_process~2_combout ),
	.datac(!\wr_addr_ptr[2]~q ),
	.datad(!\wr_addr_ptr[0]~q ),
	.datae(!\wr_addr_ptr[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fifo_array~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fifo_array~2 .extended_lut = "off";
defparam \fifo_array~2 .lut_mask = 64'hFFF7FFFFFFF7FFFF;
defparam \fifo_array~2 .shared_arith = "off";

dffeas \fifo_array[2][0] (
	.clk(clock),
	.d(\fifo_array~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(vcc),
	.q(\fifo_array[2][0]~q ),
	.prn(vcc));
defparam \fifo_array[2][0] .is_wysiwyg = "true";
defparam \fifo_array[2][0] .power_up = "low";

arriav_lcell_comb \fifo_array~3 (
	.dataa(!\fifo_array[3][0]~q ),
	.datab(!\usedw_process~2_combout ),
	.datac(!\wr_addr_ptr[2]~q ),
	.datad(!\wr_addr_ptr[0]~q ),
	.datae(!\wr_addr_ptr[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fifo_array~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fifo_array~3 .extended_lut = "off";
defparam \fifo_array~3 .lut_mask = 64'hF7FFFFFFF7FFFFFF;
defparam \fifo_array~3 .shared_arith = "off";

dffeas \fifo_array[3][0] (
	.clk(clock),
	.d(\fifo_array~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(vcc),
	.q(\fifo_array[3][0]~q ),
	.prn(vcc));
defparam \fifo_array[3][0] .is_wysiwyg = "true";
defparam \fifo_array[3][0] .power_up = "low";

endmodule

module cic_auk_dspip_avalon_streaming_sink (
	full_dff,
	rd_addr_ptr_2,
	dffe_nae,
	data,
	Equal2,
	Mux0,
	sink_ready_ctrl,
	usedw_process,
	sink_ready_ctrl1,
	sink_ready_ctrl2,
	clk,
	in_valid,
	reset_n,
	at_sink_data)/* synthesis synthesis_greybox=1 */;
output 	full_dff;
input 	rd_addr_ptr_2;
output 	dffe_nae;
output 	[19:0] data;
input 	Equal2;
input 	Mux0;
input 	sink_ready_ctrl;
input 	usedw_process;
input 	sink_ready_ctrl1;
input 	sink_ready_ctrl2;
input 	clk;
input 	in_valid;
input 	reset_n;
input 	[19:0] at_sink_data;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cic_scfifo_2 sink_FIFO(
	.full_dff(full_dff),
	.rd_addr_ptr_2(rd_addr_ptr_2),
	.dffe_nae(dffe_nae),
	.q({q_unconnected_wire_37,q_unconnected_wire_36,q_unconnected_wire_35,q_unconnected_wire_34,q_unconnected_wire_33,q_unconnected_wire_32,q_unconnected_wire_31,q_unconnected_wire_30,q_unconnected_wire_29,q_unconnected_wire_28,q_unconnected_wire_27,q_unconnected_wire_26,
q_unconnected_wire_25,q_unconnected_wire_24,q_unconnected_wire_23,q_unconnected_wire_22,q_unconnected_wire_21,q_unconnected_wire_20,data[19],data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.Equal2(Equal2),
	.Mux0(Mux0),
	.sink_ready_ctrl(sink_ready_ctrl),
	.usedw_process(usedw_process),
	.sink_ready_ctrl1(sink_ready_ctrl1),
	.sink_ready_ctrl2(sink_ready_ctrl2),
	.clock(clk),
	.in_valid(in_valid),
	.sclr(reset_n),
	.data({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,at_sink_data[19],at_sink_data[18],at_sink_data[17],at_sink_data[16],at_sink_data[15],at_sink_data[14],at_sink_data[13],at_sink_data[12],at_sink_data[11],at_sink_data[10],at_sink_data[9],at_sink_data[8],at_sink_data[7],at_sink_data[6],at_sink_data[5],at_sink_data[4],
at_sink_data[3],at_sink_data[2],at_sink_data[1],at_sink_data[0]}));

endmodule

module cic_scfifo_2 (
	full_dff,
	rd_addr_ptr_2,
	dffe_nae,
	q,
	Equal2,
	Mux0,
	sink_ready_ctrl,
	usedw_process,
	sink_ready_ctrl1,
	sink_ready_ctrl2,
	clock,
	in_valid,
	sclr,
	data)/* synthesis synthesis_greybox=1 */;
output 	full_dff;
input 	rd_addr_ptr_2;
output 	dffe_nae;
output 	[37:0] q;
input 	Equal2;
input 	Mux0;
input 	sink_ready_ctrl;
input 	usedw_process;
input 	sink_ready_ctrl1;
input 	sink_ready_ctrl2;
input 	clock;
input 	in_valid;
input 	sclr;
input 	[37:0] data;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cic_scfifo_ted1 auto_generated(
	.full_dff(full_dff),
	.rd_addr_ptr_2(rd_addr_ptr_2),
	.dffe_nae1(dffe_nae),
	.q({q_unconnected_wire_21,q_unconnected_wire_20,q[19],q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.Equal2(Equal2),
	.Mux0(Mux0),
	.sink_ready_ctrl(sink_ready_ctrl),
	.usedw_process(usedw_process),
	.sink_ready_ctrl1(sink_ready_ctrl1),
	.sink_ready_ctrl2(sink_ready_ctrl2),
	.clock(clock),
	.in_valid(in_valid),
	.sclr(sclr),
	.data({gnd,gnd,data[19],data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}));

endmodule

module cic_scfifo_ted1 (
	full_dff,
	rd_addr_ptr_2,
	dffe_nae1,
	q,
	Equal2,
	Mux0,
	sink_ready_ctrl,
	usedw_process,
	sink_ready_ctrl1,
	sink_ready_ctrl2,
	clock,
	in_valid,
	sclr,
	data)/* synthesis synthesis_greybox=1 */;
output 	full_dff;
input 	rd_addr_ptr_2;
output 	dffe_nae1;
output 	[21:0] q;
input 	Equal2;
input 	Mux0;
input 	sink_ready_ctrl;
input 	usedw_process;
input 	sink_ready_ctrl1;
input 	sink_ready_ctrl2;
input 	clock;
input 	in_valid;
input 	sclr;
input 	[21:0] data;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \dpfifo|usedw_counter|counter_reg_bit[2]~q ;
wire \dpfifo|usedw_counter|counter_reg_bit[1]~q ;
wire \dpfifo|usedw_counter|counter_reg_bit[0]~q ;
wire \dffe_nae~0_combout ;


cic_a_dpfifo_ek51 dpfifo(
	.full_dff1(full_dff),
	.rd_addr_ptr_2(rd_addr_ptr_2),
	.counter_reg_bit_2(\dpfifo|usedw_counter|counter_reg_bit[2]~q ),
	.counter_reg_bit_1(\dpfifo|usedw_counter|counter_reg_bit[1]~q ),
	.counter_reg_bit_0(\dpfifo|usedw_counter|counter_reg_bit[0]~q ),
	.q({q_unconnected_wire_21,q_unconnected_wire_20,q[19],q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.Equal2(Equal2),
	.Mux0(Mux0),
	.sink_ready_ctrl(sink_ready_ctrl),
	.usedw_process(usedw_process),
	.sink_ready_ctrl1(sink_ready_ctrl2),
	.clock(clock),
	.in_valid(in_valid),
	.sclr(sclr),
	.data({gnd,gnd,data[19],data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}));

dffeas dffe_nae(
	.clk(clock),
	.d(\dffe_nae~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!sclr),
	.sload(gnd),
	.ena(vcc),
	.q(dffe_nae1),
	.prn(vcc));
defparam dffe_nae.is_wysiwyg = "true";
defparam dffe_nae.power_up = "low";

arriav_lcell_comb \dffe_nae~0 (
	.dataa(!dffe_nae1),
	.datab(!sink_ready_ctrl1),
	.datac(!\dpfifo|usedw_counter|counter_reg_bit[2]~q ),
	.datad(!in_valid),
	.datae(!\dpfifo|usedw_counter|counter_reg_bit[1]~q ),
	.dataf(!\dpfifo|usedw_counter|counter_reg_bit[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dffe_nae~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dffe_nae~0 .extended_lut = "off";
defparam \dffe_nae~0 .lut_mask = 64'hFDFFFFFFFFFFFFFF;
defparam \dffe_nae~0 .shared_arith = "off";

endmodule

module cic_a_dpfifo_ek51 (
	full_dff1,
	rd_addr_ptr_2,
	counter_reg_bit_2,
	counter_reg_bit_1,
	counter_reg_bit_0,
	q,
	Equal2,
	Mux0,
	sink_ready_ctrl,
	usedw_process,
	sink_ready_ctrl1,
	clock,
	in_valid,
	sclr,
	data)/* synthesis synthesis_greybox=1 */;
output 	full_dff1;
input 	rd_addr_ptr_2;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
output 	counter_reg_bit_0;
output 	[21:0] q;
input 	Equal2;
input 	Mux0;
input 	sink_ready_ctrl;
input 	usedw_process;
input 	sink_ready_ctrl1;
input 	clock;
input 	in_valid;
input 	sclr;
input 	[21:0] data;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \wr_ptr|counter_reg_bit[0]~q ;
wire \wr_ptr|counter_reg_bit[1]~q ;
wire \wr_ptr|counter_reg_bit[2]~q ;
wire \rd_ptr_msb|counter_reg_bit[0]~q ;
wire \rd_ptr_msb|counter_reg_bit[1]~q ;
wire \low_addressa[0]~q ;
wire \rd_ptr_lsb~q ;
wire \ram_read_address[0]~0_combout ;
wire \low_addressa[1]~q ;
wire \ram_read_address[1]~1_combout ;
wire \low_addressa[2]~q ;
wire \ram_read_address[2]~2_combout ;
wire \low_addressa[0]~0_combout ;
wire \rd_ptr_lsb~0_combout ;
wire \rd_ptr_lsb~1_combout ;
wire \low_addressa[1]~1_combout ;
wire \low_addressa[2]~2_combout ;
wire \valid_wreq~combout ;
wire \empty_dff~1_combout ;
wire \usedw_is_0_dff~q ;
wire \usedw_will_be_1~0_combout ;
wire \usedw_will_be_1~1_combout ;
wire \usedw_is_1_dff~q ;
wire \empty_dff~0_combout ;
wire \empty_dff~q ;
wire \valid_rreq~combout ;
wire \_~0_combout ;


cic_cntr_gra wr_ptr(
	.full_dff(full_dff1),
	.counter_reg_bit_0(\wr_ptr|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\wr_ptr|counter_reg_bit[1]~q ),
	.counter_reg_bit_2(\wr_ptr|counter_reg_bit[2]~q ),
	.clock(clock),
	.in_valid(in_valid),
	.sclr(sclr));

cic_cntr_sr6 usedw_counter(
	.full_dff(full_dff1),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_1(counter_reg_bit_1),
	.counter_reg_bit_0(counter_reg_bit_0),
	.valid_rreq(\valid_rreq~combout ),
	.valid_wreq(\valid_wreq~combout ),
	.clock(clock),
	.in_valid(in_valid),
	.sclr(sclr));

cic_cntr_fra_1 rd_ptr_msb(
	.counter_reg_bit_0(\rd_ptr_msb|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\rd_ptr_msb|counter_reg_bit[1]~q ),
	.valid_rreq(\valid_rreq~combout ),
	.rd_ptr_lsb(\rd_ptr_lsb~q ),
	.clock(clock),
	.sclr(sclr));

cic_altsyncram_t6n1 FIFOram(
	.q_b({q_b_unconnected_wire_21,q_b_unconnected_wire_20,q[19],q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.address_a({\wr_ptr|counter_reg_bit[2]~q ,\wr_ptr|counter_reg_bit[1]~q ,\wr_ptr|counter_reg_bit[0]~q }),
	.clocken1(\valid_rreq~combout ),
	.wren_a(\valid_wreq~combout ),
	.address_b({\ram_read_address[2]~2_combout ,\ram_read_address[1]~1_combout ,\ram_read_address[0]~0_combout }),
	.clock1(clock),
	.clock0(clock),
	.data_a({gnd,gnd,data[19],data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}));

dffeas \low_addressa[0] (
	.clk(clock),
	.d(\low_addressa[0]~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[0]~q ),
	.prn(vcc));
defparam \low_addressa[0] .is_wysiwyg = "true";
defparam \low_addressa[0] .power_up = "low";

dffeas rd_ptr_lsb(
	.clk(clock),
	.d(\rd_ptr_lsb~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\rd_ptr_lsb~1_combout ),
	.q(\rd_ptr_lsb~q ),
	.prn(vcc));
defparam rd_ptr_lsb.is_wysiwyg = "true";
defparam rd_ptr_lsb.power_up = "low";

arriav_lcell_comb \ram_read_address[0]~0 (
	.dataa(!\valid_rreq~combout ),
	.datab(!\low_addressa[0]~q ),
	.datac(!\rd_ptr_lsb~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ram_read_address[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ram_read_address[0]~0 .extended_lut = "off";
defparam \ram_read_address[0]~0 .lut_mask = 64'hB1B1B1B1B1B1B1B1;
defparam \ram_read_address[0]~0 .shared_arith = "off";

dffeas \low_addressa[1] (
	.clk(clock),
	.d(\low_addressa[1]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[1]~q ),
	.prn(vcc));
defparam \low_addressa[1] .is_wysiwyg = "true";
defparam \low_addressa[1] .power_up = "low";

arriav_lcell_comb \ram_read_address[1]~1 (
	.dataa(!\valid_rreq~combout ),
	.datab(!\rd_ptr_msb|counter_reg_bit[0]~q ),
	.datac(!\low_addressa[1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ram_read_address[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ram_read_address[1]~1 .extended_lut = "off";
defparam \ram_read_address[1]~1 .lut_mask = 64'h2727272727272727;
defparam \ram_read_address[1]~1 .shared_arith = "off";

dffeas \low_addressa[2] (
	.clk(clock),
	.d(\low_addressa[2]~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[2]~q ),
	.prn(vcc));
defparam \low_addressa[2] .is_wysiwyg = "true";
defparam \low_addressa[2] .power_up = "low";

arriav_lcell_comb \ram_read_address[2]~2 (
	.dataa(!\valid_rreq~combout ),
	.datab(!\rd_ptr_msb|counter_reg_bit[1]~q ),
	.datac(!\low_addressa[2]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ram_read_address[2]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ram_read_address[2]~2 .extended_lut = "off";
defparam \ram_read_address[2]~2 .lut_mask = 64'h2727272727272727;
defparam \ram_read_address[2]~2 .shared_arith = "off";

arriav_lcell_comb \low_addressa[0]~0 (
	.dataa(!\valid_rreq~combout ),
	.datab(!sclr),
	.datac(!\low_addressa[0]~q ),
	.datad(!\rd_ptr_lsb~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\low_addressa[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \low_addressa[0]~0 .extended_lut = "off";
defparam \low_addressa[0]~0 .lut_mask = 64'hBF1FBF1FBF1FBF1F;
defparam \low_addressa[0]~0 .shared_arith = "off";

arriav_lcell_comb \rd_ptr_lsb~0 (
	.dataa(!sclr),
	.datab(!\rd_ptr_lsb~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rd_ptr_lsb~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rd_ptr_lsb~0 .extended_lut = "off";
defparam \rd_ptr_lsb~0 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \rd_ptr_lsb~0 .shared_arith = "off";

arriav_lcell_comb \rd_ptr_lsb~1 (
	.dataa(!\empty_dff~q ),
	.datab(!Mux0),
	.datac(!rd_addr_ptr_2),
	.datad(!usedw_process),
	.datae(!sink_ready_ctrl1),
	.dataf(!sclr),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rd_ptr_lsb~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rd_ptr_lsb~1 .extended_lut = "off";
defparam \rd_ptr_lsb~1 .lut_mask = 64'hFFFFFFFFFFFFF7FF;
defparam \rd_ptr_lsb~1 .shared_arith = "off";

arriav_lcell_comb \low_addressa[1]~1 (
	.dataa(!\valid_rreq~combout ),
	.datab(!sclr),
	.datac(!\rd_ptr_msb|counter_reg_bit[0]~q ),
	.datad(!\low_addressa[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\low_addressa[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \low_addressa[1]~1 .extended_lut = "off";
defparam \low_addressa[1]~1 .lut_mask = 64'h27FF27FF27FF27FF;
defparam \low_addressa[1]~1 .shared_arith = "off";

arriav_lcell_comb \low_addressa[2]~2 (
	.dataa(!\valid_rreq~combout ),
	.datab(!sclr),
	.datac(!\rd_ptr_msb|counter_reg_bit[1]~q ),
	.datad(!\low_addressa[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\low_addressa[2]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \low_addressa[2]~2 .extended_lut = "off";
defparam \low_addressa[2]~2 .lut_mask = 64'h27FF27FF27FF27FF;
defparam \low_addressa[2]~2 .shared_arith = "off";

dffeas full_dff(
	.clk(clock),
	.d(\_~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!sclr),
	.sload(gnd),
	.ena(vcc),
	.q(full_dff1),
	.prn(vcc));
defparam full_dff.is_wysiwyg = "true";
defparam full_dff.power_up = "low";

arriav_lcell_comb valid_wreq(
	.dataa(!full_dff1),
	.datab(!in_valid),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\valid_wreq~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam valid_wreq.extended_lut = "off";
defparam valid_wreq.lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam valid_wreq.shared_arith = "off";

arriav_lcell_comb \empty_dff~1 (
	.dataa(!full_dff1),
	.datab(!\valid_rreq~combout ),
	.datac(!in_valid),
	.datad(!sclr),
	.datae(!\usedw_is_1_dff~q ),
	.dataf(!\usedw_is_0_dff~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\empty_dff~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \empty_dff~1 .extended_lut = "off";
defparam \empty_dff~1 .lut_mask = 64'hFFFF96FFFFFFFFFF;
defparam \empty_dff~1 .shared_arith = "off";

dffeas usedw_is_0_dff(
	.clk(clock),
	.d(\empty_dff~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\usedw_is_0_dff~q ),
	.prn(vcc));
defparam usedw_is_0_dff.is_wysiwyg = "true";
defparam usedw_is_0_dff.power_up = "low";

arriav_lcell_comb \usedw_will_be_1~0 (
	.dataa(!counter_reg_bit_2),
	.datab(!counter_reg_bit_1),
	.datac(!counter_reg_bit_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\usedw_will_be_1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \usedw_will_be_1~0 .extended_lut = "off";
defparam \usedw_will_be_1~0 .lut_mask = 64'hFBFBFBFBFBFBFBFB;
defparam \usedw_will_be_1~0 .shared_arith = "off";

arriav_lcell_comb \usedw_will_be_1~1 (
	.dataa(!\valid_rreq~combout ),
	.datab(!sclr),
	.datac(!\valid_wreq~combout ),
	.datad(!\usedw_is_1_dff~q ),
	.datae(!\usedw_is_0_dff~q ),
	.dataf(!\usedw_will_be_1~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\usedw_will_be_1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \usedw_will_be_1~1 .extended_lut = "off";
defparam \usedw_will_be_1~1 .lut_mask = 64'hFFFF7BFFFFFFFFFF;
defparam \usedw_will_be_1~1 .shared_arith = "off";

dffeas usedw_is_1_dff(
	.clk(clock),
	.d(\usedw_will_be_1~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\usedw_is_1_dff~q ),
	.prn(vcc));
defparam usedw_is_1_dff.is_wysiwyg = "true";
defparam usedw_is_1_dff.power_up = "low";

arriav_lcell_comb \empty_dff~0 (
	.dataa(!\valid_rreq~combout ),
	.datab(!sclr),
	.datac(!\valid_wreq~combout ),
	.datad(!\usedw_is_1_dff~q ),
	.datae(!\usedw_is_0_dff~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\empty_dff~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \empty_dff~0 .extended_lut = "off";
defparam \empty_dff~0 .lut_mask = 64'hF7B3FFFFF7B3FFFF;
defparam \empty_dff~0 .shared_arith = "off";

dffeas empty_dff(
	.clk(clock),
	.d(\empty_dff~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\empty_dff~q ),
	.prn(vcc));
defparam empty_dff.is_wysiwyg = "true";
defparam empty_dff.power_up = "low";

arriav_lcell_comb valid_rreq(
	.dataa(!\empty_dff~q ),
	.datab(!Equal2),
	.datac(!Mux0),
	.datad(!rd_addr_ptr_2),
	.datae(!sink_ready_ctrl),
	.dataf(!usedw_process),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\valid_rreq~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam valid_rreq.extended_lut = "off";
defparam valid_rreq.lut_mask = 64'hFF7FFFFFFFFFFFFF;
defparam valid_rreq.shared_arith = "off";

arriav_lcell_comb \_~0 (
	.dataa(!full_dff1),
	.datab(!\valid_rreq~combout ),
	.datac(!counter_reg_bit_2),
	.datad(!in_valid),
	.datae(!counter_reg_bit_1),
	.dataf(!counter_reg_bit_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\_~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \_~0 .extended_lut = "off";
defparam \_~0 .lut_mask = 64'hDFFFFFFFFFFFFFFF;
defparam \_~0 .shared_arith = "off";

endmodule

module cic_altsyncram_t6n1 (
	q_b,
	address_a,
	clocken1,
	wren_a,
	address_b,
	clock1,
	clock0,
	data_a)/* synthesis synthesis_greybox=1 */;
output 	[21:0] q_b;
input 	[2:0] address_a;
input 	clocken1;
input 	wren_a;
input 	[2:0] address_b;
input 	clock1;
input 	clock0;
input 	[21:0] data_a;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a19_PORTBDATAOUT_bus;
wire [143:0] ram_block1a18_PORTBDATAOUT_bus;
wire [143:0] ram_block1a17_PORTBDATAOUT_bus;
wire [143:0] ram_block1a16_PORTBDATAOUT_bus;
wire [143:0] ram_block1a15_PORTBDATAOUT_bus;
wire [143:0] ram_block1a14_PORTBDATAOUT_bus;
wire [143:0] ram_block1a13_PORTBDATAOUT_bus;
wire [143:0] ram_block1a12_PORTBDATAOUT_bus;
wire [143:0] ram_block1a11_PORTBDATAOUT_bus;
wire [143:0] ram_block1a10_PORTBDATAOUT_bus;
wire [143:0] ram_block1a9_PORTBDATAOUT_bus;
wire [143:0] ram_block1a8_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a1_PORTBDATAOUT_bus;
wire [143:0] ram_block1a0_PORTBDATAOUT_bus;

assign q_b[19] = ram_block1a19_PORTBDATAOUT_bus[0];

assign q_b[18] = ram_block1a18_PORTBDATAOUT_bus[0];

assign q_b[17] = ram_block1a17_PORTBDATAOUT_bus[0];

assign q_b[16] = ram_block1a16_PORTBDATAOUT_bus[0];

assign q_b[15] = ram_block1a15_PORTBDATAOUT_bus[0];

assign q_b[14] = ram_block1a14_PORTBDATAOUT_bus[0];

assign q_b[13] = ram_block1a13_PORTBDATAOUT_bus[0];

assign q_b[12] = ram_block1a12_PORTBDATAOUT_bus[0];

assign q_b[11] = ram_block1a11_PORTBDATAOUT_bus[0];

assign q_b[10] = ram_block1a10_PORTBDATAOUT_bus[0];

assign q_b[9] = ram_block1a9_PORTBDATAOUT_bus[0];

assign q_b[8] = ram_block1a8_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

arriav_ram_block ram_block1a19(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[19]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a19_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a19.clk1_output_clock_enable = "ena1";
defparam ram_block1a19.data_interleave_offset_in_bits = 1;
defparam ram_block1a19.data_interleave_width_in_bits = 1;
defparam ram_block1a19.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_ted1:auto_generated|a_dpfifo_ek51:dpfifo|altsyncram_t6n1:FIFOram|ALTSYNCRAM";
defparam ram_block1a19.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a19.operation_mode = "dual_port";
defparam ram_block1a19.port_a_address_clear = "none";
defparam ram_block1a19.port_a_address_width = 3;
defparam ram_block1a19.port_a_data_out_clear = "none";
defparam ram_block1a19.port_a_data_out_clock = "none";
defparam ram_block1a19.port_a_data_width = 1;
defparam ram_block1a19.port_a_first_address = 0;
defparam ram_block1a19.port_a_first_bit_number = 19;
defparam ram_block1a19.port_a_last_address = 7;
defparam ram_block1a19.port_a_logical_ram_depth = 8;
defparam ram_block1a19.port_a_logical_ram_width = 22;
defparam ram_block1a19.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a19.port_b_address_clear = "none";
defparam ram_block1a19.port_b_address_clock = "clock1";
defparam ram_block1a19.port_b_address_width = 3;
defparam ram_block1a19.port_b_data_out_clear = "none";
defparam ram_block1a19.port_b_data_out_clock = "clock1";
defparam ram_block1a19.port_b_data_width = 1;
defparam ram_block1a19.port_b_first_address = 0;
defparam ram_block1a19.port_b_first_bit_number = 19;
defparam ram_block1a19.port_b_last_address = 7;
defparam ram_block1a19.port_b_logical_ram_depth = 8;
defparam ram_block1a19.port_b_logical_ram_width = 22;
defparam ram_block1a19.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a19.port_b_read_enable_clock = "clock1";
defparam ram_block1a19.ram_block_type = "auto";

arriav_ram_block ram_block1a18(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[18]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a18_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a18.clk1_output_clock_enable = "ena1";
defparam ram_block1a18.data_interleave_offset_in_bits = 1;
defparam ram_block1a18.data_interleave_width_in_bits = 1;
defparam ram_block1a18.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_ted1:auto_generated|a_dpfifo_ek51:dpfifo|altsyncram_t6n1:FIFOram|ALTSYNCRAM";
defparam ram_block1a18.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a18.operation_mode = "dual_port";
defparam ram_block1a18.port_a_address_clear = "none";
defparam ram_block1a18.port_a_address_width = 3;
defparam ram_block1a18.port_a_data_out_clear = "none";
defparam ram_block1a18.port_a_data_out_clock = "none";
defparam ram_block1a18.port_a_data_width = 1;
defparam ram_block1a18.port_a_first_address = 0;
defparam ram_block1a18.port_a_first_bit_number = 18;
defparam ram_block1a18.port_a_last_address = 7;
defparam ram_block1a18.port_a_logical_ram_depth = 8;
defparam ram_block1a18.port_a_logical_ram_width = 22;
defparam ram_block1a18.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a18.port_b_address_clear = "none";
defparam ram_block1a18.port_b_address_clock = "clock1";
defparam ram_block1a18.port_b_address_width = 3;
defparam ram_block1a18.port_b_data_out_clear = "none";
defparam ram_block1a18.port_b_data_out_clock = "clock1";
defparam ram_block1a18.port_b_data_width = 1;
defparam ram_block1a18.port_b_first_address = 0;
defparam ram_block1a18.port_b_first_bit_number = 18;
defparam ram_block1a18.port_b_last_address = 7;
defparam ram_block1a18.port_b_logical_ram_depth = 8;
defparam ram_block1a18.port_b_logical_ram_width = 22;
defparam ram_block1a18.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a18.port_b_read_enable_clock = "clock1";
defparam ram_block1a18.ram_block_type = "auto";

arriav_ram_block ram_block1a17(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[17]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a17_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a17.clk1_output_clock_enable = "ena1";
defparam ram_block1a17.data_interleave_offset_in_bits = 1;
defparam ram_block1a17.data_interleave_width_in_bits = 1;
defparam ram_block1a17.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_ted1:auto_generated|a_dpfifo_ek51:dpfifo|altsyncram_t6n1:FIFOram|ALTSYNCRAM";
defparam ram_block1a17.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a17.operation_mode = "dual_port";
defparam ram_block1a17.port_a_address_clear = "none";
defparam ram_block1a17.port_a_address_width = 3;
defparam ram_block1a17.port_a_data_out_clear = "none";
defparam ram_block1a17.port_a_data_out_clock = "none";
defparam ram_block1a17.port_a_data_width = 1;
defparam ram_block1a17.port_a_first_address = 0;
defparam ram_block1a17.port_a_first_bit_number = 17;
defparam ram_block1a17.port_a_last_address = 7;
defparam ram_block1a17.port_a_logical_ram_depth = 8;
defparam ram_block1a17.port_a_logical_ram_width = 22;
defparam ram_block1a17.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a17.port_b_address_clear = "none";
defparam ram_block1a17.port_b_address_clock = "clock1";
defparam ram_block1a17.port_b_address_width = 3;
defparam ram_block1a17.port_b_data_out_clear = "none";
defparam ram_block1a17.port_b_data_out_clock = "clock1";
defparam ram_block1a17.port_b_data_width = 1;
defparam ram_block1a17.port_b_first_address = 0;
defparam ram_block1a17.port_b_first_bit_number = 17;
defparam ram_block1a17.port_b_last_address = 7;
defparam ram_block1a17.port_b_logical_ram_depth = 8;
defparam ram_block1a17.port_b_logical_ram_width = 22;
defparam ram_block1a17.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a17.port_b_read_enable_clock = "clock1";
defparam ram_block1a17.ram_block_type = "auto";

arriav_ram_block ram_block1a16(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a16_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a16.clk1_output_clock_enable = "ena1";
defparam ram_block1a16.data_interleave_offset_in_bits = 1;
defparam ram_block1a16.data_interleave_width_in_bits = 1;
defparam ram_block1a16.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_ted1:auto_generated|a_dpfifo_ek51:dpfifo|altsyncram_t6n1:FIFOram|ALTSYNCRAM";
defparam ram_block1a16.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a16.operation_mode = "dual_port";
defparam ram_block1a16.port_a_address_clear = "none";
defparam ram_block1a16.port_a_address_width = 3;
defparam ram_block1a16.port_a_data_out_clear = "none";
defparam ram_block1a16.port_a_data_out_clock = "none";
defparam ram_block1a16.port_a_data_width = 1;
defparam ram_block1a16.port_a_first_address = 0;
defparam ram_block1a16.port_a_first_bit_number = 16;
defparam ram_block1a16.port_a_last_address = 7;
defparam ram_block1a16.port_a_logical_ram_depth = 8;
defparam ram_block1a16.port_a_logical_ram_width = 22;
defparam ram_block1a16.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a16.port_b_address_clear = "none";
defparam ram_block1a16.port_b_address_clock = "clock1";
defparam ram_block1a16.port_b_address_width = 3;
defparam ram_block1a16.port_b_data_out_clear = "none";
defparam ram_block1a16.port_b_data_out_clock = "clock1";
defparam ram_block1a16.port_b_data_width = 1;
defparam ram_block1a16.port_b_first_address = 0;
defparam ram_block1a16.port_b_first_bit_number = 16;
defparam ram_block1a16.port_b_last_address = 7;
defparam ram_block1a16.port_b_logical_ram_depth = 8;
defparam ram_block1a16.port_b_logical_ram_width = 22;
defparam ram_block1a16.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a16.port_b_read_enable_clock = "clock1";
defparam ram_block1a16.ram_block_type = "auto";

arriav_ram_block ram_block1a15(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a15_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a15.clk1_output_clock_enable = "ena1";
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_ted1:auto_generated|a_dpfifo_ek51:dpfifo|altsyncram_t6n1:FIFOram|ALTSYNCRAM";
defparam ram_block1a15.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a15.operation_mode = "dual_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 3;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 7;
defparam ram_block1a15.port_a_logical_ram_depth = 8;
defparam ram_block1a15.port_a_logical_ram_width = 22;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a15.port_b_address_clear = "none";
defparam ram_block1a15.port_b_address_clock = "clock1";
defparam ram_block1a15.port_b_address_width = 3;
defparam ram_block1a15.port_b_data_out_clear = "none";
defparam ram_block1a15.port_b_data_out_clock = "clock1";
defparam ram_block1a15.port_b_data_width = 1;
defparam ram_block1a15.port_b_first_address = 0;
defparam ram_block1a15.port_b_first_bit_number = 15;
defparam ram_block1a15.port_b_last_address = 7;
defparam ram_block1a15.port_b_logical_ram_depth = 8;
defparam ram_block1a15.port_b_logical_ram_width = 22;
defparam ram_block1a15.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a15.port_b_read_enable_clock = "clock1";
defparam ram_block1a15.ram_block_type = "auto";

arriav_ram_block ram_block1a14(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a14_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a14.clk1_output_clock_enable = "ena1";
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_ted1:auto_generated|a_dpfifo_ek51:dpfifo|altsyncram_t6n1:FIFOram|ALTSYNCRAM";
defparam ram_block1a14.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a14.operation_mode = "dual_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 3;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 7;
defparam ram_block1a14.port_a_logical_ram_depth = 8;
defparam ram_block1a14.port_a_logical_ram_width = 22;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a14.port_b_address_clear = "none";
defparam ram_block1a14.port_b_address_clock = "clock1";
defparam ram_block1a14.port_b_address_width = 3;
defparam ram_block1a14.port_b_data_out_clear = "none";
defparam ram_block1a14.port_b_data_out_clock = "clock1";
defparam ram_block1a14.port_b_data_width = 1;
defparam ram_block1a14.port_b_first_address = 0;
defparam ram_block1a14.port_b_first_bit_number = 14;
defparam ram_block1a14.port_b_last_address = 7;
defparam ram_block1a14.port_b_logical_ram_depth = 8;
defparam ram_block1a14.port_b_logical_ram_width = 22;
defparam ram_block1a14.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a14.port_b_read_enable_clock = "clock1";
defparam ram_block1a14.ram_block_type = "auto";

arriav_ram_block ram_block1a13(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a13_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a13.clk1_output_clock_enable = "ena1";
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_ted1:auto_generated|a_dpfifo_ek51:dpfifo|altsyncram_t6n1:FIFOram|ALTSYNCRAM";
defparam ram_block1a13.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a13.operation_mode = "dual_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 3;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 7;
defparam ram_block1a13.port_a_logical_ram_depth = 8;
defparam ram_block1a13.port_a_logical_ram_width = 22;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a13.port_b_address_clear = "none";
defparam ram_block1a13.port_b_address_clock = "clock1";
defparam ram_block1a13.port_b_address_width = 3;
defparam ram_block1a13.port_b_data_out_clear = "none";
defparam ram_block1a13.port_b_data_out_clock = "clock1";
defparam ram_block1a13.port_b_data_width = 1;
defparam ram_block1a13.port_b_first_address = 0;
defparam ram_block1a13.port_b_first_bit_number = 13;
defparam ram_block1a13.port_b_last_address = 7;
defparam ram_block1a13.port_b_logical_ram_depth = 8;
defparam ram_block1a13.port_b_logical_ram_width = 22;
defparam ram_block1a13.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a13.port_b_read_enable_clock = "clock1";
defparam ram_block1a13.ram_block_type = "auto";

arriav_ram_block ram_block1a12(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a12_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a12.clk1_output_clock_enable = "ena1";
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_ted1:auto_generated|a_dpfifo_ek51:dpfifo|altsyncram_t6n1:FIFOram|ALTSYNCRAM";
defparam ram_block1a12.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a12.operation_mode = "dual_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 3;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 7;
defparam ram_block1a12.port_a_logical_ram_depth = 8;
defparam ram_block1a12.port_a_logical_ram_width = 22;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a12.port_b_address_clear = "none";
defparam ram_block1a12.port_b_address_clock = "clock1";
defparam ram_block1a12.port_b_address_width = 3;
defparam ram_block1a12.port_b_data_out_clear = "none";
defparam ram_block1a12.port_b_data_out_clock = "clock1";
defparam ram_block1a12.port_b_data_width = 1;
defparam ram_block1a12.port_b_first_address = 0;
defparam ram_block1a12.port_b_first_bit_number = 12;
defparam ram_block1a12.port_b_last_address = 7;
defparam ram_block1a12.port_b_logical_ram_depth = 8;
defparam ram_block1a12.port_b_logical_ram_width = 22;
defparam ram_block1a12.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a12.port_b_read_enable_clock = "clock1";
defparam ram_block1a12.ram_block_type = "auto";

arriav_ram_block ram_block1a11(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a11_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a11.clk1_output_clock_enable = "ena1";
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_ted1:auto_generated|a_dpfifo_ek51:dpfifo|altsyncram_t6n1:FIFOram|ALTSYNCRAM";
defparam ram_block1a11.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a11.operation_mode = "dual_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 3;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 7;
defparam ram_block1a11.port_a_logical_ram_depth = 8;
defparam ram_block1a11.port_a_logical_ram_width = 22;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a11.port_b_address_clear = "none";
defparam ram_block1a11.port_b_address_clock = "clock1";
defparam ram_block1a11.port_b_address_width = 3;
defparam ram_block1a11.port_b_data_out_clear = "none";
defparam ram_block1a11.port_b_data_out_clock = "clock1";
defparam ram_block1a11.port_b_data_width = 1;
defparam ram_block1a11.port_b_first_address = 0;
defparam ram_block1a11.port_b_first_bit_number = 11;
defparam ram_block1a11.port_b_last_address = 7;
defparam ram_block1a11.port_b_logical_ram_depth = 8;
defparam ram_block1a11.port_b_logical_ram_width = 22;
defparam ram_block1a11.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a11.port_b_read_enable_clock = "clock1";
defparam ram_block1a11.ram_block_type = "auto";

arriav_ram_block ram_block1a10(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a10_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a10.clk1_output_clock_enable = "ena1";
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_ted1:auto_generated|a_dpfifo_ek51:dpfifo|altsyncram_t6n1:FIFOram|ALTSYNCRAM";
defparam ram_block1a10.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a10.operation_mode = "dual_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 3;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 7;
defparam ram_block1a10.port_a_logical_ram_depth = 8;
defparam ram_block1a10.port_a_logical_ram_width = 22;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a10.port_b_address_clear = "none";
defparam ram_block1a10.port_b_address_clock = "clock1";
defparam ram_block1a10.port_b_address_width = 3;
defparam ram_block1a10.port_b_data_out_clear = "none";
defparam ram_block1a10.port_b_data_out_clock = "clock1";
defparam ram_block1a10.port_b_data_width = 1;
defparam ram_block1a10.port_b_first_address = 0;
defparam ram_block1a10.port_b_first_bit_number = 10;
defparam ram_block1a10.port_b_last_address = 7;
defparam ram_block1a10.port_b_logical_ram_depth = 8;
defparam ram_block1a10.port_b_logical_ram_width = 22;
defparam ram_block1a10.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a10.port_b_read_enable_clock = "clock1";
defparam ram_block1a10.ram_block_type = "auto";

arriav_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a9.clk1_output_clock_enable = "ena1";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_ted1:auto_generated|a_dpfifo_ek51:dpfifo|altsyncram_t6n1:FIFOram|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a9.operation_mode = "dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 3;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 7;
defparam ram_block1a9.port_a_logical_ram_depth = 8;
defparam ram_block1a9.port_a_logical_ram_width = 22;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a9.port_b_address_clear = "none";
defparam ram_block1a9.port_b_address_clock = "clock1";
defparam ram_block1a9.port_b_address_width = 3;
defparam ram_block1a9.port_b_data_out_clear = "none";
defparam ram_block1a9.port_b_data_out_clock = "clock1";
defparam ram_block1a9.port_b_data_width = 1;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 7;
defparam ram_block1a9.port_b_logical_ram_depth = 8;
defparam ram_block1a9.port_b_logical_ram_width = 22;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock1";
defparam ram_block1a9.ram_block_type = "auto";

arriav_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a8.clk1_output_clock_enable = "ena1";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_ted1:auto_generated|a_dpfifo_ek51:dpfifo|altsyncram_t6n1:FIFOram|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a8.operation_mode = "dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 3;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 7;
defparam ram_block1a8.port_a_logical_ram_depth = 8;
defparam ram_block1a8.port_a_logical_ram_width = 22;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a8.port_b_address_clear = "none";
defparam ram_block1a8.port_b_address_clock = "clock1";
defparam ram_block1a8.port_b_address_width = 3;
defparam ram_block1a8.port_b_data_out_clear = "none";
defparam ram_block1a8.port_b_data_out_clock = "clock1";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 7;
defparam ram_block1a8.port_b_logical_ram_depth = 8;
defparam ram_block1a8.port_b_logical_ram_width = 22;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock1";
defparam ram_block1a8.ram_block_type = "auto";

arriav_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a7.clk1_output_clock_enable = "ena1";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_ted1:auto_generated|a_dpfifo_ek51:dpfifo|altsyncram_t6n1:FIFOram|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 3;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 7;
defparam ram_block1a7.port_a_logical_ram_depth = 8;
defparam ram_block1a7.port_a_logical_ram_width = 22;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock1";
defparam ram_block1a7.port_b_address_width = 3;
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "clock1";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 7;
defparam ram_block1a7.port_b_logical_ram_depth = 8;
defparam ram_block1a7.port_b_logical_ram_width = 22;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock1";
defparam ram_block1a7.ram_block_type = "auto";

arriav_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a6.clk1_output_clock_enable = "ena1";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_ted1:auto_generated|a_dpfifo_ek51:dpfifo|altsyncram_t6n1:FIFOram|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 3;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 7;
defparam ram_block1a6.port_a_logical_ram_depth = 8;
defparam ram_block1a6.port_a_logical_ram_width = 22;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock1";
defparam ram_block1a6.port_b_address_width = 3;
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "clock1";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 7;
defparam ram_block1a6.port_b_logical_ram_depth = 8;
defparam ram_block1a6.port_b_logical_ram_width = 22;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock1";
defparam ram_block1a6.ram_block_type = "auto";

arriav_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a5.clk1_output_clock_enable = "ena1";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_ted1:auto_generated|a_dpfifo_ek51:dpfifo|altsyncram_t6n1:FIFOram|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 3;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 7;
defparam ram_block1a5.port_a_logical_ram_depth = 8;
defparam ram_block1a5.port_a_logical_ram_width = 22;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock1";
defparam ram_block1a5.port_b_address_width = 3;
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "clock1";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 7;
defparam ram_block1a5.port_b_logical_ram_depth = 8;
defparam ram_block1a5.port_b_logical_ram_width = 22;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock1";
defparam ram_block1a5.ram_block_type = "auto";

arriav_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a4.clk1_output_clock_enable = "ena1";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_ted1:auto_generated|a_dpfifo_ek51:dpfifo|altsyncram_t6n1:FIFOram|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a4.operation_mode = "dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 3;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 7;
defparam ram_block1a4.port_a_logical_ram_depth = 8;
defparam ram_block1a4.port_a_logical_ram_width = 22;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_address_clear = "none";
defparam ram_block1a4.port_b_address_clock = "clock1";
defparam ram_block1a4.port_b_address_width = 3;
defparam ram_block1a4.port_b_data_out_clear = "none";
defparam ram_block1a4.port_b_data_out_clock = "clock1";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 7;
defparam ram_block1a4.port_b_logical_ram_depth = 8;
defparam ram_block1a4.port_b_logical_ram_width = 22;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock1";
defparam ram_block1a4.ram_block_type = "auto";

arriav_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a3.clk1_output_clock_enable = "ena1";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_ted1:auto_generated|a_dpfifo_ek51:dpfifo|altsyncram_t6n1:FIFOram|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a3.operation_mode = "dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 3;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 7;
defparam ram_block1a3.port_a_logical_ram_depth = 8;
defparam ram_block1a3.port_a_logical_ram_width = 22;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_address_clear = "none";
defparam ram_block1a3.port_b_address_clock = "clock1";
defparam ram_block1a3.port_b_address_width = 3;
defparam ram_block1a3.port_b_data_out_clear = "none";
defparam ram_block1a3.port_b_data_out_clock = "clock1";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 7;
defparam ram_block1a3.port_b_logical_ram_depth = 8;
defparam ram_block1a3.port_b_logical_ram_width = 22;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock1";
defparam ram_block1a3.ram_block_type = "auto";

arriav_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a2.clk1_output_clock_enable = "ena1";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_ted1:auto_generated|a_dpfifo_ek51:dpfifo|altsyncram_t6n1:FIFOram|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a2.operation_mode = "dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 3;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 7;
defparam ram_block1a2.port_a_logical_ram_depth = 8;
defparam ram_block1a2.port_a_logical_ram_width = 22;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_address_clear = "none";
defparam ram_block1a2.port_b_address_clock = "clock1";
defparam ram_block1a2.port_b_address_width = 3;
defparam ram_block1a2.port_b_data_out_clear = "none";
defparam ram_block1a2.port_b_data_out_clock = "clock1";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 7;
defparam ram_block1a2.port_b_logical_ram_depth = 8;
defparam ram_block1a2.port_b_logical_ram_width = 22;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock1";
defparam ram_block1a2.ram_block_type = "auto";

arriav_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a1.clk1_output_clock_enable = "ena1";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_ted1:auto_generated|a_dpfifo_ek51:dpfifo|altsyncram_t6n1:FIFOram|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 3;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 7;
defparam ram_block1a1.port_a_logical_ram_depth = 8;
defparam ram_block1a1.port_a_logical_ram_width = 22;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_address_clear = "none";
defparam ram_block1a1.port_b_address_clock = "clock1";
defparam ram_block1a1.port_b_address_width = 3;
defparam ram_block1a1.port_b_data_out_clear = "none";
defparam ram_block1a1.port_b_data_out_clock = "clock1";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 7;
defparam ram_block1a1.port_b_logical_ram_depth = 8;
defparam ram_block1a1.port_b_logical_ram_width = 22;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock1";
defparam ram_block1a1.ram_block_type = "auto";

arriav_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a0.clk1_output_clock_enable = "ena1";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_ted1:auto_generated|a_dpfifo_ek51:dpfifo|altsyncram_t6n1:FIFOram|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 3;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 7;
defparam ram_block1a0.port_a_logical_ram_depth = 8;
defparam ram_block1a0.port_a_logical_ram_width = 22;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_address_clear = "none";
defparam ram_block1a0.port_b_address_clock = "clock1";
defparam ram_block1a0.port_b_address_width = 3;
defparam ram_block1a0.port_b_data_out_clear = "none";
defparam ram_block1a0.port_b_data_out_clock = "clock1";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 7;
defparam ram_block1a0.port_b_logical_ram_depth = 8;
defparam ram_block1a0.port_b_logical_ram_width = 22;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock1";
defparam ram_block1a0.ram_block_type = "auto";

endmodule

module cic_cntr_fra_1 (
	counter_reg_bit_0,
	counter_reg_bit_1,
	valid_rreq,
	rd_ptr_lsb,
	clock,
	sclr)/* synthesis synthesis_greybox=1 */;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
input 	valid_rreq;
input 	rd_ptr_lsb;
input 	clock;
input 	sclr;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~sumout ;
wire \_~0_combout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~sumout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!sclr),
	.sload(gnd),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!sclr),
	.sload(gnd),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

arriav_lcell_comb counter_comb_bita0(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita0~sumout ),
	.cout(\counter_comb_bita0~COUT ),
	.shareout());
defparam counter_comb_bita0.extended_lut = "off";
defparam counter_comb_bita0.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita0.shared_arith = "off";

arriav_lcell_comb \_~0 (
	.dataa(!valid_rreq),
	.datab(!sclr),
	.datac(!rd_ptr_lsb),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\_~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \_~0 .extended_lut = "off";
defparam \_~0 .lut_mask = 64'hFDFDFDFDFDFDFDFD;
defparam \_~0 .shared_arith = "off";

arriav_lcell_comb counter_comb_bita1(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita0~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita1~sumout ),
	.cout(),
	.shareout());
defparam counter_comb_bita1.extended_lut = "off";
defparam counter_comb_bita1.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita1.shared_arith = "off";

endmodule

module cic_cntr_gra (
	full_dff,
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_2,
	clock,
	in_valid,
	sclr)/* synthesis synthesis_greybox=1 */;
input 	full_dff;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
input 	clock;
input 	in_valid;
input 	sclr;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~sumout ;
wire \_~0_combout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~sumout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~sumout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!sclr),
	.sload(gnd),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!sclr),
	.sload(gnd),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!sclr),
	.sload(gnd),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

arriav_lcell_comb counter_comb_bita0(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita0~sumout ),
	.cout(\counter_comb_bita0~COUT ),
	.shareout());
defparam counter_comb_bita0.extended_lut = "off";
defparam counter_comb_bita0.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita0.shared_arith = "off";

arriav_lcell_comb \_~0 (
	.dataa(!full_dff),
	.datab(!in_valid),
	.datac(!sclr),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\_~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \_~0 .extended_lut = "off";
defparam \_~0 .lut_mask = 64'hFBFBFBFBFBFBFBFB;
defparam \_~0 .shared_arith = "off";

arriav_lcell_comb counter_comb_bita1(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita0~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita1~sumout ),
	.cout(\counter_comb_bita1~COUT ),
	.shareout());
defparam counter_comb_bita1.extended_lut = "off";
defparam counter_comb_bita1.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita1.shared_arith = "off";

arriav_lcell_comb counter_comb_bita2(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita1~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita2~sumout ),
	.cout(),
	.shareout());
defparam counter_comb_bita2.extended_lut = "off";
defparam counter_comb_bita2.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita2.shared_arith = "off";

endmodule

module cic_cntr_sr6 (
	full_dff,
	counter_reg_bit_2,
	counter_reg_bit_1,
	counter_reg_bit_0,
	valid_rreq,
	valid_wreq,
	clock,
	in_valid,
	sclr)/* synthesis synthesis_greybox=1 */;
input 	full_dff;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
output 	counter_reg_bit_0;
input 	valid_rreq;
input 	valid_wreq;
input 	clock;
input 	in_valid;
input 	sclr;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~sumout ;
wire \_~0_combout ;
wire \counter_comb_bita1~sumout ;
wire \counter_comb_bita0~sumout ;


dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!sclr),
	.sload(gnd),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!sclr),
	.sload(gnd),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!sclr),
	.sload(gnd),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

arriav_lcell_comb counter_comb_bita0(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita0~sumout ),
	.cout(\counter_comb_bita0~COUT ),
	.shareout());
defparam counter_comb_bita0.extended_lut = "off";
defparam counter_comb_bita0.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita0.shared_arith = "off";

arriav_lcell_comb counter_comb_bita1(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_1),
	.datae(gnd),
	.dataf(!valid_wreq),
	.datag(gnd),
	.cin(\counter_comb_bita0~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita1~sumout ),
	.cout(\counter_comb_bita1~COUT ),
	.shareout());
defparam counter_comb_bita1.extended_lut = "off";
defparam counter_comb_bita1.lut_mask = 64'h000000FF000000FF;
defparam counter_comb_bita1.shared_arith = "off";

arriav_lcell_comb counter_comb_bita2(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_2),
	.datae(gnd),
	.dataf(!valid_wreq),
	.datag(gnd),
	.cin(\counter_comb_bita1~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita2~sumout ),
	.cout(),
	.shareout());
defparam counter_comb_bita2.extended_lut = "off";
defparam counter_comb_bita2.lut_mask = 64'h000000FF000000FF;
defparam counter_comb_bita2.shared_arith = "off";

arriav_lcell_comb \_~0 (
	.dataa(!full_dff),
	.datab(!valid_rreq),
	.datac(!in_valid),
	.datad(!sclr),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\_~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \_~0 .extended_lut = "off";
defparam \_~0 .lut_mask = 64'hFF96FF96FF96FF96;
defparam \_~0 .shared_arith = "off";

endmodule

module cic_auk_dspip_avalon_streaming_source (
	at_source_data,
	source_valid_s1,
	dffe_af,
	dout_valid,
	state_0,
	data,
	stall_reg,
	clk,
	reset_n,
	out_ready)/* synthesis synthesis_greybox=1 */;
output 	[27:0] at_source_data;
output 	source_valid_s1;
output 	dffe_af;
input 	dout_valid;
input 	state_0;
input 	[27:0] data;
input 	stall_reg;
input 	clk;
input 	reset_n;
input 	out_ready;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \source_FIFO|auto_generated|dpfifo|empty_dff~q ;
wire \source_valid_s_process~0_combout ;
wire \source_valid_s~0_combout ;


cic_scfifo_3 source_FIFO(
	.q({q_unconnected_wire_37,q_unconnected_wire_36,q_unconnected_wire_35,q_unconnected_wire_34,q_unconnected_wire_33,q_unconnected_wire_32,q_unconnected_wire_31,q_unconnected_wire_30,q_unconnected_wire_29,q_unconnected_wire_28,at_source_data[27],at_source_data[26],at_source_data[25],
at_source_data[24],at_source_data[23],at_source_data[22],at_source_data[21],at_source_data[20],at_source_data[19],at_source_data[18],at_source_data[17],at_source_data[16],at_source_data[15],at_source_data[14],at_source_data[13],at_source_data[12],at_source_data[11],at_source_data[10],at_source_data[9],at_source_data[8],at_source_data[7],
at_source_data[6],at_source_data[5],at_source_data[4],at_source_data[3],at_source_data[2],at_source_data[1],at_source_data[0]}),
	.source_valid_s(source_valid_s1),
	.dffe_af(dffe_af),
	.dout_valid(dout_valid),
	.state_0(state_0),
	.data({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data[27],data[26],data[25],data[24],data[23],data[22],data[21],data[20],data[19],data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.stall_reg(stall_reg),
	.empty_dff(\source_FIFO|auto_generated|dpfifo|empty_dff~q ),
	.source_valid_s_process(\source_valid_s_process~0_combout ),
	.clock(clk),
	.sclr(reset_n),
	.out_ready(out_ready));

arriav_lcell_comb \source_valid_s_process~0 (
	.dataa(!source_valid_s1),
	.datab(!\source_FIFO|auto_generated|dpfifo|empty_dff~q ),
	.datac(!out_ready),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\source_valid_s_process~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \source_valid_s_process~0 .extended_lut = "off";
defparam \source_valid_s_process~0 .lut_mask = 64'hBFBFBFBFBFBFBFBF;
defparam \source_valid_s_process~0 .shared_arith = "off";

dffeas source_valid_s(
	.clk(clk),
	.d(\source_valid_s~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(vcc),
	.q(source_valid_s1),
	.prn(vcc));
defparam source_valid_s.is_wysiwyg = "true";
defparam source_valid_s.power_up = "low";

arriav_lcell_comb \source_valid_s~0 (
	.dataa(!source_valid_s1),
	.datab(!\source_FIFO|auto_generated|dpfifo|empty_dff~q ),
	.datac(!out_ready),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\source_valid_s~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \source_valid_s~0 .extended_lut = "off";
defparam \source_valid_s~0 .lut_mask = 64'hF7F7F7F7F7F7F7F7;
defparam \source_valid_s~0 .shared_arith = "off";

endmodule

module cic_scfifo_3 (
	q,
	source_valid_s,
	dffe_af,
	dout_valid,
	state_0,
	data,
	stall_reg,
	empty_dff,
	source_valid_s_process,
	clock,
	sclr,
	out_ready)/* synthesis synthesis_greybox=1 */;
output 	[37:0] q;
input 	source_valid_s;
output 	dffe_af;
input 	dout_valid;
input 	state_0;
input 	[37:0] data;
input 	stall_reg;
output 	empty_dff;
input 	source_valid_s_process;
input 	clock;
input 	sclr;
input 	out_ready;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cic_scfifo_1id1 auto_generated(
	.q({q_unconnected_wire_28,q[27],q[26],q[25],q[24],q[23],q[22],q[21],q[20],q[19],q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.source_valid_s(source_valid_s),
	.dffe_af1(dffe_af),
	.dout_valid(dout_valid),
	.state_0(state_0),
	.data({gnd,data[27],data[26],data[25],data[24],data[23],data[22],data[21],data[20],data[19],data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.stall_reg(stall_reg),
	.empty_dff(empty_dff),
	.source_valid_s_process(source_valid_s_process),
	.clock(clock),
	.sclr(sclr),
	.out_ready(out_ready));

endmodule

module cic_scfifo_1id1 (
	q,
	source_valid_s,
	dffe_af1,
	dout_valid,
	state_0,
	data,
	stall_reg,
	empty_dff,
	source_valid_s_process,
	clock,
	sclr,
	out_ready)/* synthesis synthesis_greybox=1 */;
output 	[28:0] q;
input 	source_valid_s;
output 	dffe_af1;
input 	dout_valid;
input 	state_0;
input 	[28:0] data;
input 	stall_reg;
output 	empty_dff;
input 	source_valid_s_process;
input 	clock;
input 	sclr;
input 	out_ready;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \dpfifo|usedw_counter|counter_reg_bit[0]~q ;
wire \dpfifo|usedw_counter|counter_reg_bit[4]~q ;
wire \dpfifo|usedw_counter|counter_reg_bit[3]~q ;
wire \dpfifo|usedw_counter|counter_reg_bit[2]~q ;
wire \dpfifo|usedw_counter|counter_reg_bit[1]~q ;
wire \dpfifo|valid_wreq~1_combout ;
wire \dffe_af~0_combout ;
wire \dffe_af~1_combout ;


cic_a_dpfifo_up51 dpfifo(
	.q({q_unconnected_wire_28,q[27],q[26],q[25],q[24],q[23],q[22],q[21],q[20],q[19],q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.source_valid_s(source_valid_s),
	.dout_valid(dout_valid),
	.state_0(state_0),
	.data({gnd,data[27],data[26],data[25],data[24],data[23],data[22],data[21],data[20],data[19],data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.counter_reg_bit_0(\dpfifo|usedw_counter|counter_reg_bit[0]~q ),
	.counter_reg_bit_4(\dpfifo|usedw_counter|counter_reg_bit[4]~q ),
	.counter_reg_bit_3(\dpfifo|usedw_counter|counter_reg_bit[3]~q ),
	.counter_reg_bit_2(\dpfifo|usedw_counter|counter_reg_bit[2]~q ),
	.counter_reg_bit_1(\dpfifo|usedw_counter|counter_reg_bit[1]~q ),
	.stall_reg(stall_reg),
	.empty_dff1(empty_dff),
	.source_valid_s_process(source_valid_s_process),
	.valid_wreq(\dpfifo|valid_wreq~1_combout ),
	.clock(clock),
	.sclr(sclr),
	.out_ready(out_ready));

dffeas dffe_af(
	.clk(clock),
	.d(\dffe_af~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!sclr),
	.sload(gnd),
	.ena(vcc),
	.q(dffe_af1),
	.prn(vcc));
defparam dffe_af.is_wysiwyg = "true";
defparam dffe_af.power_up = "low";

arriav_lcell_comb \dffe_af~0 (
	.dataa(!\dpfifo|usedw_counter|counter_reg_bit[4]~q ),
	.datab(!\dpfifo|usedw_counter|counter_reg_bit[3]~q ),
	.datac(!\dpfifo|usedw_counter|counter_reg_bit[2]~q ),
	.datad(!\dpfifo|usedw_counter|counter_reg_bit[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dffe_af~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dffe_af~0 .extended_lut = "off";
defparam \dffe_af~0 .lut_mask = 64'hFFBFFFBFFFBFFFBF;
defparam \dffe_af~0 .shared_arith = "off";

arriav_lcell_comb \dffe_af~1 (
	.dataa(!source_valid_s),
	.datab(!dffe_af1),
	.datac(!\dpfifo|valid_wreq~1_combout ),
	.datad(!out_ready),
	.datae(!\dpfifo|usedw_counter|counter_reg_bit[0]~q ),
	.dataf(!\dffe_af~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dffe_af~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dffe_af~1 .extended_lut = "off";
defparam \dffe_af~1 .lut_mask = 64'hFF7FFF7FFFFF7F7F;
defparam \dffe_af~1 .shared_arith = "off";

endmodule

module cic_a_dpfifo_up51 (
	q,
	source_valid_s,
	dout_valid,
	state_0,
	data,
	counter_reg_bit_0,
	counter_reg_bit_4,
	counter_reg_bit_3,
	counter_reg_bit_2,
	counter_reg_bit_1,
	stall_reg,
	empty_dff1,
	source_valid_s_process,
	valid_wreq,
	clock,
	sclr,
	out_ready)/* synthesis synthesis_greybox=1 */;
output 	[28:0] q;
input 	source_valid_s;
input 	dout_valid;
input 	state_0;
input 	[28:0] data;
output 	counter_reg_bit_0;
output 	counter_reg_bit_4;
output 	counter_reg_bit_3;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
input 	stall_reg;
output 	empty_dff1;
input 	source_valid_s_process;
output 	valid_wreq;
input 	clock;
input 	sclr;
input 	out_ready;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \wr_ptr|counter_reg_bit[0]~q ;
wire \wr_ptr|counter_reg_bit[1]~q ;
wire \wr_ptr|counter_reg_bit[2]~q ;
wire \wr_ptr|counter_reg_bit[3]~q ;
wire \wr_ptr|counter_reg_bit[4]~q ;
wire \rd_ptr_msb|counter_reg_bit[0]~q ;
wire \rd_ptr_msb|counter_reg_bit[1]~q ;
wire \rd_ptr_msb|counter_reg_bit[2]~q ;
wire \rd_ptr_msb|counter_reg_bit[3]~q ;
wire \low_addressa[0]~q ;
wire \rd_ptr_lsb~q ;
wire \ram_read_address[0]~0_combout ;
wire \low_addressa[1]~q ;
wire \ram_read_address[1]~1_combout ;
wire \low_addressa[2]~q ;
wire \ram_read_address[2]~2_combout ;
wire \low_addressa[3]~q ;
wire \ram_read_address[3]~3_combout ;
wire \low_addressa[4]~q ;
wire \ram_read_address[4]~4_combout ;
wire \low_addressa[0]~0_combout ;
wire \rd_ptr_lsb~0_combout ;
wire \rd_ptr_lsb~1_combout ;
wire \low_addressa[1]~1_combout ;
wire \low_addressa[2]~2_combout ;
wire \low_addressa[3]~3_combout ;
wire \low_addressa[4]~4_combout ;
wire \_~0_combout ;
wire \_~1_combout ;
wire \full_dff~q ;
wire \valid_wreq~0_combout ;
wire \empty_dff~1_combout ;
wire \usedw_is_0_dff~q ;
wire \usedw_will_be_1~0_combout ;
wire \usedw_will_be_1~1_combout ;
wire \usedw_is_1_dff~q ;
wire \empty_dff~0_combout ;


cic_cntr_hra rd_ptr_msb(
	.source_valid_s(source_valid_s),
	.counter_reg_bit_0(\rd_ptr_msb|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\rd_ptr_msb|counter_reg_bit[1]~q ),
	.counter_reg_bit_2(\rd_ptr_msb|counter_reg_bit[2]~q ),
	.counter_reg_bit_3(\rd_ptr_msb|counter_reg_bit[3]~q ),
	.empty_dff(empty_dff1),
	.rd_ptr_lsb(\rd_ptr_lsb~q ),
	.clock(clock),
	.sclr(sclr),
	.out_ready(out_ready));

cic_altsyncram_9an1 FIFOram(
	.q_b({q_b_unconnected_wire_28,q[27],q[26],q[25],q[24],q[23],q[22],q[21],q[20],q[19],q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.data_a({gnd,data[27],data[26],data[25],data[24],data[23],data[22],data[21],data[20],data[19],data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.address_a({\wr_ptr|counter_reg_bit[4]~q ,\wr_ptr|counter_reg_bit[3]~q ,\wr_ptr|counter_reg_bit[2]~q ,\wr_ptr|counter_reg_bit[1]~q ,\wr_ptr|counter_reg_bit[0]~q }),
	.wren_a(\valid_wreq~0_combout ),
	.clocken1(source_valid_s_process),
	.address_b({\ram_read_address[4]~4_combout ,\ram_read_address[3]~3_combout ,\ram_read_address[2]~2_combout ,\ram_read_address[1]~1_combout ,\ram_read_address[0]~0_combout }),
	.clock1(clock),
	.clock0(clock));

cic_cntr_ira wr_ptr(
	.full_dff(\full_dff~q ),
	.dout_valid(dout_valid),
	.state_0(state_0),
	.counter_reg_bit_0(\wr_ptr|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\wr_ptr|counter_reg_bit[1]~q ),
	.counter_reg_bit_2(\wr_ptr|counter_reg_bit[2]~q ),
	.counter_reg_bit_3(\wr_ptr|counter_reg_bit[3]~q ),
	.counter_reg_bit_4(\wr_ptr|counter_reg_bit[4]~q ),
	.stall_reg(stall_reg),
	.clock(clock),
	.sclr(sclr));

cic_cntr_ur6 usedw_counter(
	.source_valid_s(source_valid_s),
	.counter_reg_bit_0(counter_reg_bit_0),
	.counter_reg_bit_4(counter_reg_bit_4),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_1(counter_reg_bit_1),
	.valid_wreq(\valid_wreq~0_combout ),
	.empty_dff(empty_dff1),
	.clock(clock),
	.sclr(sclr),
	.out_ready(out_ready));

dffeas \low_addressa[0] (
	.clk(clock),
	.d(\low_addressa[0]~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[0]~q ),
	.prn(vcc));
defparam \low_addressa[0] .is_wysiwyg = "true";
defparam \low_addressa[0] .power_up = "low";

dffeas rd_ptr_lsb(
	.clk(clock),
	.d(\rd_ptr_lsb~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\rd_ptr_lsb~1_combout ),
	.q(\rd_ptr_lsb~q ),
	.prn(vcc));
defparam rd_ptr_lsb.is_wysiwyg = "true";
defparam rd_ptr_lsb.power_up = "low";

arriav_lcell_comb \ram_read_address[0]~0 (
	.dataa(!source_valid_s),
	.datab(!empty_dff1),
	.datac(!out_ready),
	.datad(!\low_addressa[0]~q ),
	.datae(!\rd_ptr_lsb~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ram_read_address[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ram_read_address[0]~0 .extended_lut = "off";
defparam \ram_read_address[0]~0 .lut_mask = 64'hFFFF96FFFFFF96FF;
defparam \ram_read_address[0]~0 .shared_arith = "off";

dffeas \low_addressa[1] (
	.clk(clock),
	.d(\low_addressa[1]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[1]~q ),
	.prn(vcc));
defparam \low_addressa[1] .is_wysiwyg = "true";
defparam \low_addressa[1] .power_up = "low";

arriav_lcell_comb \ram_read_address[1]~1 (
	.dataa(!source_valid_s),
	.datab(!empty_dff1),
	.datac(!out_ready),
	.datad(!\rd_ptr_msb|counter_reg_bit[0]~q ),
	.datae(!\low_addressa[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ram_read_address[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ram_read_address[1]~1 .extended_lut = "off";
defparam \ram_read_address[1]~1 .lut_mask = 64'h96FFFFFF96FFFFFF;
defparam \ram_read_address[1]~1 .shared_arith = "off";

dffeas \low_addressa[2] (
	.clk(clock),
	.d(\low_addressa[2]~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[2]~q ),
	.prn(vcc));
defparam \low_addressa[2] .is_wysiwyg = "true";
defparam \low_addressa[2] .power_up = "low";

arriav_lcell_comb \ram_read_address[2]~2 (
	.dataa(!source_valid_s),
	.datab(!empty_dff1),
	.datac(!out_ready),
	.datad(!\rd_ptr_msb|counter_reg_bit[1]~q ),
	.datae(!\low_addressa[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ram_read_address[2]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ram_read_address[2]~2 .extended_lut = "off";
defparam \ram_read_address[2]~2 .lut_mask = 64'h96FFFFFF96FFFFFF;
defparam \ram_read_address[2]~2 .shared_arith = "off";

dffeas \low_addressa[3] (
	.clk(clock),
	.d(\low_addressa[3]~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[3]~q ),
	.prn(vcc));
defparam \low_addressa[3] .is_wysiwyg = "true";
defparam \low_addressa[3] .power_up = "low";

arriav_lcell_comb \ram_read_address[3]~3 (
	.dataa(!source_valid_s),
	.datab(!empty_dff1),
	.datac(!out_ready),
	.datad(!\rd_ptr_msb|counter_reg_bit[2]~q ),
	.datae(!\low_addressa[3]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ram_read_address[3]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ram_read_address[3]~3 .extended_lut = "off";
defparam \ram_read_address[3]~3 .lut_mask = 64'h96FFFFFF96FFFFFF;
defparam \ram_read_address[3]~3 .shared_arith = "off";

dffeas \low_addressa[4] (
	.clk(clock),
	.d(\low_addressa[4]~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[4]~q ),
	.prn(vcc));
defparam \low_addressa[4] .is_wysiwyg = "true";
defparam \low_addressa[4] .power_up = "low";

arriav_lcell_comb \ram_read_address[4]~4 (
	.dataa(!source_valid_s),
	.datab(!empty_dff1),
	.datac(!out_ready),
	.datad(!\rd_ptr_msb|counter_reg_bit[3]~q ),
	.datae(!\low_addressa[4]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ram_read_address[4]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ram_read_address[4]~4 .extended_lut = "off";
defparam \ram_read_address[4]~4 .lut_mask = 64'h96FFFFFF96FFFFFF;
defparam \ram_read_address[4]~4 .shared_arith = "off";

arriav_lcell_comb \low_addressa[0]~0 (
	.dataa(!source_valid_s),
	.datab(!sclr),
	.datac(!empty_dff1),
	.datad(!out_ready),
	.datae(!\low_addressa[0]~q ),
	.dataf(!\rd_ptr_lsb~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\low_addressa[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \low_addressa[0]~0 .extended_lut = "off";
defparam \low_addressa[0]~0 .lut_mask = 64'hFFFFFFFFB77BFFFF;
defparam \low_addressa[0]~0 .shared_arith = "off";

arriav_lcell_comb \rd_ptr_lsb~0 (
	.dataa(!sclr),
	.datab(!\rd_ptr_lsb~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rd_ptr_lsb~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rd_ptr_lsb~0 .extended_lut = "off";
defparam \rd_ptr_lsb~0 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \rd_ptr_lsb~0 .shared_arith = "off";

arriav_lcell_comb \rd_ptr_lsb~1 (
	.dataa(!source_valid_s),
	.datab(!sclr),
	.datac(!empty_dff1),
	.datad(!out_ready),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rd_ptr_lsb~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rd_ptr_lsb~1 .extended_lut = "off";
defparam \rd_ptr_lsb~1 .lut_mask = 64'hEFFFEFFFEFFFEFFF;
defparam \rd_ptr_lsb~1 .shared_arith = "off";

arriav_lcell_comb \low_addressa[1]~1 (
	.dataa(!source_valid_s),
	.datab(!sclr),
	.datac(!empty_dff1),
	.datad(!out_ready),
	.datae(!\rd_ptr_msb|counter_reg_bit[0]~q ),
	.dataf(!\low_addressa[1]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\low_addressa[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \low_addressa[1]~1 .extended_lut = "off";
defparam \low_addressa[1]~1 .lut_mask = 64'hB77BFFFFFFFFFFFF;
defparam \low_addressa[1]~1 .shared_arith = "off";

arriav_lcell_comb \low_addressa[2]~2 (
	.dataa(!source_valid_s),
	.datab(!sclr),
	.datac(!empty_dff1),
	.datad(!out_ready),
	.datae(!\rd_ptr_msb|counter_reg_bit[1]~q ),
	.dataf(!\low_addressa[2]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\low_addressa[2]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \low_addressa[2]~2 .extended_lut = "off";
defparam \low_addressa[2]~2 .lut_mask = 64'hB77BFFFFFFFFFFFF;
defparam \low_addressa[2]~2 .shared_arith = "off";

arriav_lcell_comb \low_addressa[3]~3 (
	.dataa(!source_valid_s),
	.datab(!sclr),
	.datac(!empty_dff1),
	.datad(!out_ready),
	.datae(!\rd_ptr_msb|counter_reg_bit[2]~q ),
	.dataf(!\low_addressa[3]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\low_addressa[3]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \low_addressa[3]~3 .extended_lut = "off";
defparam \low_addressa[3]~3 .lut_mask = 64'hB77BFFFFFFFFFFFF;
defparam \low_addressa[3]~3 .shared_arith = "off";

arriav_lcell_comb \low_addressa[4]~4 (
	.dataa(!source_valid_s),
	.datab(!sclr),
	.datac(!empty_dff1),
	.datad(!out_ready),
	.datae(!\rd_ptr_msb|counter_reg_bit[3]~q ),
	.dataf(!\low_addressa[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\low_addressa[4]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \low_addressa[4]~4 .extended_lut = "off";
defparam \low_addressa[4]~4 .lut_mask = 64'hB77BFFFFFFFFFFFF;
defparam \low_addressa[4]~4 .shared_arith = "off";

dffeas empty_dff(
	.clk(clock),
	.d(\empty_dff~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(empty_dff1),
	.prn(vcc));
defparam empty_dff.is_wysiwyg = "true";
defparam empty_dff.power_up = "low";

arriav_lcell_comb \valid_wreq~1 (
	.dataa(!stall_reg),
	.datab(!dout_valid),
	.datac(!state_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(valid_wreq),
	.sumout(),
	.cout(),
	.shareout());
defparam \valid_wreq~1 .extended_lut = "off";
defparam \valid_wreq~1 .lut_mask = 64'hBFBFBFBFBFBFBFBF;
defparam \valid_wreq~1 .shared_arith = "off";

arriav_lcell_comb \_~0 (
	.dataa(!counter_reg_bit_0),
	.datab(!counter_reg_bit_4),
	.datac(!counter_reg_bit_3),
	.datad(!counter_reg_bit_2),
	.datae(!counter_reg_bit_1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\_~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \_~0 .extended_lut = "off";
defparam \_~0 .lut_mask = 64'hFFFFFBFFFFFFFBFF;
defparam \_~0 .shared_arith = "off";

arriav_lcell_comb \_~1 (
	.dataa(!source_valid_s),
	.datab(!\full_dff~q ),
	.datac(!\valid_wreq~0_combout ),
	.datad(!empty_dff1),
	.datae(!out_ready),
	.dataf(!\_~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\_~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \_~1 .extended_lut = "off";
defparam \_~1 .lut_mask = 64'hFFFFFF7FFFFFFFFF;
defparam \_~1 .shared_arith = "off";

dffeas full_dff(
	.clk(clock),
	.d(\_~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!sclr),
	.sload(gnd),
	.ena(vcc),
	.q(\full_dff~q ),
	.prn(vcc));
defparam full_dff.is_wysiwyg = "true";
defparam full_dff.power_up = "low";

arriav_lcell_comb \valid_wreq~0 (
	.dataa(!\full_dff~q ),
	.datab(!stall_reg),
	.datac(!dout_valid),
	.datad(!state_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\valid_wreq~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \valid_wreq~0 .extended_lut = "off";
defparam \valid_wreq~0 .lut_mask = 64'hEFFFEFFFEFFFEFFF;
defparam \valid_wreq~0 .shared_arith = "off";

arriav_lcell_comb \empty_dff~1 (
	.dataa(!sclr),
	.datab(!\valid_wreq~0_combout ),
	.datac(!source_valid_s_process),
	.datad(!\usedw_is_1_dff~q ),
	.datae(!\usedw_is_0_dff~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\empty_dff~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \empty_dff~1 .extended_lut = "off";
defparam \empty_dff~1 .lut_mask = 64'hFF7DFFFFFF7DFFFF;
defparam \empty_dff~1 .shared_arith = "off";

dffeas usedw_is_0_dff(
	.clk(clock),
	.d(\empty_dff~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\usedw_is_0_dff~q ),
	.prn(vcc));
defparam usedw_is_0_dff.is_wysiwyg = "true";
defparam usedw_is_0_dff.power_up = "low";

arriav_lcell_comb \usedw_will_be_1~0 (
	.dataa(!counter_reg_bit_0),
	.datab(!counter_reg_bit_4),
	.datac(!counter_reg_bit_3),
	.datad(!counter_reg_bit_2),
	.datae(!counter_reg_bit_1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\usedw_will_be_1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \usedw_will_be_1~0 .extended_lut = "off";
defparam \usedw_will_be_1~0 .lut_mask = 64'hFFFEFFFFFFFEFFFF;
defparam \usedw_will_be_1~0 .shared_arith = "off";

arriav_lcell_comb \usedw_will_be_1~1 (
	.dataa(!sclr),
	.datab(!\valid_wreq~0_combout ),
	.datac(!source_valid_s_process),
	.datad(!\usedw_is_1_dff~q ),
	.datae(!\usedw_is_0_dff~q ),
	.dataf(!\usedw_will_be_1~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\usedw_will_be_1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \usedw_will_be_1~1 .extended_lut = "off";
defparam \usedw_will_be_1~1 .lut_mask = 64'hFFFF7DFFFFFFFFFF;
defparam \usedw_will_be_1~1 .shared_arith = "off";

dffeas usedw_is_1_dff(
	.clk(clock),
	.d(\usedw_will_be_1~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\usedw_is_1_dff~q ),
	.prn(vcc));
defparam usedw_is_1_dff.is_wysiwyg = "true";
defparam usedw_is_1_dff.power_up = "low";

arriav_lcell_comb \empty_dff~0 (
	.dataa(!sclr),
	.datab(!\valid_wreq~0_combout ),
	.datac(!source_valid_s_process),
	.datad(!\usedw_is_1_dff~q ),
	.datae(!\usedw_is_0_dff~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\empty_dff~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \empty_dff~0 .extended_lut = "off";
defparam \empty_dff~0 .lut_mask = 64'hDFD5FFFFDFD5FFFF;
defparam \empty_dff~0 .shared_arith = "off";

endmodule

module cic_altsyncram_9an1 (
	q_b,
	data_a,
	address_a,
	wren_a,
	clocken1,
	address_b,
	clock1,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[28:0] q_b;
input 	[28:0] data_a;
input 	[4:0] address_a;
input 	wren_a;
input 	clocken1;
input 	[4:0] address_b;
input 	clock1;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a0_PORTBDATAOUT_bus;
wire [143:0] ram_block1a1_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a8_PORTBDATAOUT_bus;
wire [143:0] ram_block1a9_PORTBDATAOUT_bus;
wire [143:0] ram_block1a10_PORTBDATAOUT_bus;
wire [143:0] ram_block1a11_PORTBDATAOUT_bus;
wire [143:0] ram_block1a12_PORTBDATAOUT_bus;
wire [143:0] ram_block1a13_PORTBDATAOUT_bus;
wire [143:0] ram_block1a14_PORTBDATAOUT_bus;
wire [143:0] ram_block1a15_PORTBDATAOUT_bus;
wire [143:0] ram_block1a16_PORTBDATAOUT_bus;
wire [143:0] ram_block1a17_PORTBDATAOUT_bus;
wire [143:0] ram_block1a18_PORTBDATAOUT_bus;
wire [143:0] ram_block1a19_PORTBDATAOUT_bus;
wire [143:0] ram_block1a20_PORTBDATAOUT_bus;
wire [143:0] ram_block1a21_PORTBDATAOUT_bus;
wire [143:0] ram_block1a22_PORTBDATAOUT_bus;
wire [143:0] ram_block1a23_PORTBDATAOUT_bus;
wire [143:0] ram_block1a24_PORTBDATAOUT_bus;
wire [143:0] ram_block1a25_PORTBDATAOUT_bus;
wire [143:0] ram_block1a26_PORTBDATAOUT_bus;
wire [143:0] ram_block1a27_PORTBDATAOUT_bus;

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[8] = ram_block1a8_PORTBDATAOUT_bus[0];

assign q_b[9] = ram_block1a9_PORTBDATAOUT_bus[0];

assign q_b[10] = ram_block1a10_PORTBDATAOUT_bus[0];

assign q_b[11] = ram_block1a11_PORTBDATAOUT_bus[0];

assign q_b[12] = ram_block1a12_PORTBDATAOUT_bus[0];

assign q_b[13] = ram_block1a13_PORTBDATAOUT_bus[0];

assign q_b[14] = ram_block1a14_PORTBDATAOUT_bus[0];

assign q_b[15] = ram_block1a15_PORTBDATAOUT_bus[0];

assign q_b[16] = ram_block1a16_PORTBDATAOUT_bus[0];

assign q_b[17] = ram_block1a17_PORTBDATAOUT_bus[0];

assign q_b[18] = ram_block1a18_PORTBDATAOUT_bus[0];

assign q_b[19] = ram_block1a19_PORTBDATAOUT_bus[0];

assign q_b[20] = ram_block1a20_PORTBDATAOUT_bus[0];

assign q_b[21] = ram_block1a21_PORTBDATAOUT_bus[0];

assign q_b[22] = ram_block1a22_PORTBDATAOUT_bus[0];

assign q_b[23] = ram_block1a23_PORTBDATAOUT_bus[0];

assign q_b[24] = ram_block1a24_PORTBDATAOUT_bus[0];

assign q_b[25] = ram_block1a25_PORTBDATAOUT_bus[0];

assign q_b[26] = ram_block1a26_PORTBDATAOUT_bus[0];

assign q_b[27] = ram_block1a27_PORTBDATAOUT_bus[0];

arriav_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.clk1_output_clock_enable = "ena1";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_source:output_source_0|scfifo:source_FIFO|scfifo_1id1:auto_generated|a_dpfifo_up51:dpfifo|altsyncram_9an1:FIFOram|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 5;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 31;
defparam ram_block1a0.port_a_logical_ram_depth = 32;
defparam ram_block1a0.port_a_logical_ram_width = 29;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_address_clear = "none";
defparam ram_block1a0.port_b_address_clock = "clock1";
defparam ram_block1a0.port_b_address_width = 5;
defparam ram_block1a0.port_b_data_out_clear = "none";
defparam ram_block1a0.port_b_data_out_clock = "clock1";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 31;
defparam ram_block1a0.port_b_logical_ram_depth = 32;
defparam ram_block1a0.port_b_logical_ram_width = 29;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock1";
defparam ram_block1a0.ram_block_type = "auto";

arriav_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.clk1_output_clock_enable = "ena1";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_source:output_source_0|scfifo:source_FIFO|scfifo_1id1:auto_generated|a_dpfifo_up51:dpfifo|altsyncram_9an1:FIFOram|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 5;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 31;
defparam ram_block1a1.port_a_logical_ram_depth = 32;
defparam ram_block1a1.port_a_logical_ram_width = 29;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_address_clear = "none";
defparam ram_block1a1.port_b_address_clock = "clock1";
defparam ram_block1a1.port_b_address_width = 5;
defparam ram_block1a1.port_b_data_out_clear = "none";
defparam ram_block1a1.port_b_data_out_clock = "clock1";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 31;
defparam ram_block1a1.port_b_logical_ram_depth = 32;
defparam ram_block1a1.port_b_logical_ram_width = 29;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock1";
defparam ram_block1a1.ram_block_type = "auto";

arriav_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.clk1_output_clock_enable = "ena1";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_source:output_source_0|scfifo:source_FIFO|scfifo_1id1:auto_generated|a_dpfifo_up51:dpfifo|altsyncram_9an1:FIFOram|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a2.operation_mode = "dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 5;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 31;
defparam ram_block1a2.port_a_logical_ram_depth = 32;
defparam ram_block1a2.port_a_logical_ram_width = 29;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_address_clear = "none";
defparam ram_block1a2.port_b_address_clock = "clock1";
defparam ram_block1a2.port_b_address_width = 5;
defparam ram_block1a2.port_b_data_out_clear = "none";
defparam ram_block1a2.port_b_data_out_clock = "clock1";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 31;
defparam ram_block1a2.port_b_logical_ram_depth = 32;
defparam ram_block1a2.port_b_logical_ram_width = 29;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock1";
defparam ram_block1a2.ram_block_type = "auto";

arriav_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.clk1_output_clock_enable = "ena1";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_source:output_source_0|scfifo:source_FIFO|scfifo_1id1:auto_generated|a_dpfifo_up51:dpfifo|altsyncram_9an1:FIFOram|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a3.operation_mode = "dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 5;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 31;
defparam ram_block1a3.port_a_logical_ram_depth = 32;
defparam ram_block1a3.port_a_logical_ram_width = 29;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_address_clear = "none";
defparam ram_block1a3.port_b_address_clock = "clock1";
defparam ram_block1a3.port_b_address_width = 5;
defparam ram_block1a3.port_b_data_out_clear = "none";
defparam ram_block1a3.port_b_data_out_clock = "clock1";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 31;
defparam ram_block1a3.port_b_logical_ram_depth = 32;
defparam ram_block1a3.port_b_logical_ram_width = 29;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock1";
defparam ram_block1a3.ram_block_type = "auto";

arriav_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.clk1_output_clock_enable = "ena1";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_source:output_source_0|scfifo:source_FIFO|scfifo_1id1:auto_generated|a_dpfifo_up51:dpfifo|altsyncram_9an1:FIFOram|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a4.operation_mode = "dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 5;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 31;
defparam ram_block1a4.port_a_logical_ram_depth = 32;
defparam ram_block1a4.port_a_logical_ram_width = 29;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_address_clear = "none";
defparam ram_block1a4.port_b_address_clock = "clock1";
defparam ram_block1a4.port_b_address_width = 5;
defparam ram_block1a4.port_b_data_out_clear = "none";
defparam ram_block1a4.port_b_data_out_clock = "clock1";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 31;
defparam ram_block1a4.port_b_logical_ram_depth = 32;
defparam ram_block1a4.port_b_logical_ram_width = 29;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock1";
defparam ram_block1a4.ram_block_type = "auto";

arriav_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.clk1_output_clock_enable = "ena1";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_source:output_source_0|scfifo:source_FIFO|scfifo_1id1:auto_generated|a_dpfifo_up51:dpfifo|altsyncram_9an1:FIFOram|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 5;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 31;
defparam ram_block1a5.port_a_logical_ram_depth = 32;
defparam ram_block1a5.port_a_logical_ram_width = 29;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock1";
defparam ram_block1a5.port_b_address_width = 5;
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "clock1";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 31;
defparam ram_block1a5.port_b_logical_ram_depth = 32;
defparam ram_block1a5.port_b_logical_ram_width = 29;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock1";
defparam ram_block1a5.ram_block_type = "auto";

arriav_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.clk1_output_clock_enable = "ena1";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_source:output_source_0|scfifo:source_FIFO|scfifo_1id1:auto_generated|a_dpfifo_up51:dpfifo|altsyncram_9an1:FIFOram|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 5;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 31;
defparam ram_block1a6.port_a_logical_ram_depth = 32;
defparam ram_block1a6.port_a_logical_ram_width = 29;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock1";
defparam ram_block1a6.port_b_address_width = 5;
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "clock1";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 31;
defparam ram_block1a6.port_b_logical_ram_depth = 32;
defparam ram_block1a6.port_b_logical_ram_width = 29;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock1";
defparam ram_block1a6.ram_block_type = "auto";

arriav_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.clk1_output_clock_enable = "ena1";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_source:output_source_0|scfifo:source_FIFO|scfifo_1id1:auto_generated|a_dpfifo_up51:dpfifo|altsyncram_9an1:FIFOram|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 5;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 31;
defparam ram_block1a7.port_a_logical_ram_depth = 32;
defparam ram_block1a7.port_a_logical_ram_width = 29;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock1";
defparam ram_block1a7.port_b_address_width = 5;
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "clock1";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 31;
defparam ram_block1a7.port_b_logical_ram_depth = 32;
defparam ram_block1a7.port_b_logical_ram_width = 29;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock1";
defparam ram_block1a7.ram_block_type = "auto";

arriav_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a8.clk0_core_clock_enable = "ena0";
defparam ram_block1a8.clk1_output_clock_enable = "ena1";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_source:output_source_0|scfifo:source_FIFO|scfifo_1id1:auto_generated|a_dpfifo_up51:dpfifo|altsyncram_9an1:FIFOram|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a8.operation_mode = "dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 5;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 31;
defparam ram_block1a8.port_a_logical_ram_depth = 32;
defparam ram_block1a8.port_a_logical_ram_width = 29;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a8.port_b_address_clear = "none";
defparam ram_block1a8.port_b_address_clock = "clock1";
defparam ram_block1a8.port_b_address_width = 5;
defparam ram_block1a8.port_b_data_out_clear = "none";
defparam ram_block1a8.port_b_data_out_clock = "clock1";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 31;
defparam ram_block1a8.port_b_logical_ram_depth = 32;
defparam ram_block1a8.port_b_logical_ram_width = 29;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock1";
defparam ram_block1a8.ram_block_type = "auto";

arriav_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a9.clk0_core_clock_enable = "ena0";
defparam ram_block1a9.clk1_output_clock_enable = "ena1";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_source:output_source_0|scfifo:source_FIFO|scfifo_1id1:auto_generated|a_dpfifo_up51:dpfifo|altsyncram_9an1:FIFOram|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a9.operation_mode = "dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 5;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 31;
defparam ram_block1a9.port_a_logical_ram_depth = 32;
defparam ram_block1a9.port_a_logical_ram_width = 29;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a9.port_b_address_clear = "none";
defparam ram_block1a9.port_b_address_clock = "clock1";
defparam ram_block1a9.port_b_address_width = 5;
defparam ram_block1a9.port_b_data_out_clear = "none";
defparam ram_block1a9.port_b_data_out_clock = "clock1";
defparam ram_block1a9.port_b_data_width = 1;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 31;
defparam ram_block1a9.port_b_logical_ram_depth = 32;
defparam ram_block1a9.port_b_logical_ram_width = 29;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock1";
defparam ram_block1a9.ram_block_type = "auto";

arriav_ram_block ram_block1a10(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a10_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a10.clk0_core_clock_enable = "ena0";
defparam ram_block1a10.clk1_output_clock_enable = "ena1";
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_source:output_source_0|scfifo:source_FIFO|scfifo_1id1:auto_generated|a_dpfifo_up51:dpfifo|altsyncram_9an1:FIFOram|ALTSYNCRAM";
defparam ram_block1a10.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a10.operation_mode = "dual_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 5;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 31;
defparam ram_block1a10.port_a_logical_ram_depth = 32;
defparam ram_block1a10.port_a_logical_ram_width = 29;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a10.port_b_address_clear = "none";
defparam ram_block1a10.port_b_address_clock = "clock1";
defparam ram_block1a10.port_b_address_width = 5;
defparam ram_block1a10.port_b_data_out_clear = "none";
defparam ram_block1a10.port_b_data_out_clock = "clock1";
defparam ram_block1a10.port_b_data_width = 1;
defparam ram_block1a10.port_b_first_address = 0;
defparam ram_block1a10.port_b_first_bit_number = 10;
defparam ram_block1a10.port_b_last_address = 31;
defparam ram_block1a10.port_b_logical_ram_depth = 32;
defparam ram_block1a10.port_b_logical_ram_width = 29;
defparam ram_block1a10.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a10.port_b_read_enable_clock = "clock1";
defparam ram_block1a10.ram_block_type = "auto";

arriav_ram_block ram_block1a11(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a11_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a11.clk0_core_clock_enable = "ena0";
defparam ram_block1a11.clk1_output_clock_enable = "ena1";
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_source:output_source_0|scfifo:source_FIFO|scfifo_1id1:auto_generated|a_dpfifo_up51:dpfifo|altsyncram_9an1:FIFOram|ALTSYNCRAM";
defparam ram_block1a11.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a11.operation_mode = "dual_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 5;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 31;
defparam ram_block1a11.port_a_logical_ram_depth = 32;
defparam ram_block1a11.port_a_logical_ram_width = 29;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a11.port_b_address_clear = "none";
defparam ram_block1a11.port_b_address_clock = "clock1";
defparam ram_block1a11.port_b_address_width = 5;
defparam ram_block1a11.port_b_data_out_clear = "none";
defparam ram_block1a11.port_b_data_out_clock = "clock1";
defparam ram_block1a11.port_b_data_width = 1;
defparam ram_block1a11.port_b_first_address = 0;
defparam ram_block1a11.port_b_first_bit_number = 11;
defparam ram_block1a11.port_b_last_address = 31;
defparam ram_block1a11.port_b_logical_ram_depth = 32;
defparam ram_block1a11.port_b_logical_ram_width = 29;
defparam ram_block1a11.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a11.port_b_read_enable_clock = "clock1";
defparam ram_block1a11.ram_block_type = "auto";

arriav_ram_block ram_block1a12(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a12_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a12.clk0_core_clock_enable = "ena0";
defparam ram_block1a12.clk1_output_clock_enable = "ena1";
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_source:output_source_0|scfifo:source_FIFO|scfifo_1id1:auto_generated|a_dpfifo_up51:dpfifo|altsyncram_9an1:FIFOram|ALTSYNCRAM";
defparam ram_block1a12.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a12.operation_mode = "dual_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 5;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 31;
defparam ram_block1a12.port_a_logical_ram_depth = 32;
defparam ram_block1a12.port_a_logical_ram_width = 29;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a12.port_b_address_clear = "none";
defparam ram_block1a12.port_b_address_clock = "clock1";
defparam ram_block1a12.port_b_address_width = 5;
defparam ram_block1a12.port_b_data_out_clear = "none";
defparam ram_block1a12.port_b_data_out_clock = "clock1";
defparam ram_block1a12.port_b_data_width = 1;
defparam ram_block1a12.port_b_first_address = 0;
defparam ram_block1a12.port_b_first_bit_number = 12;
defparam ram_block1a12.port_b_last_address = 31;
defparam ram_block1a12.port_b_logical_ram_depth = 32;
defparam ram_block1a12.port_b_logical_ram_width = 29;
defparam ram_block1a12.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a12.port_b_read_enable_clock = "clock1";
defparam ram_block1a12.ram_block_type = "auto";

arriav_ram_block ram_block1a13(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a13_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a13.clk0_core_clock_enable = "ena0";
defparam ram_block1a13.clk1_output_clock_enable = "ena1";
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_source:output_source_0|scfifo:source_FIFO|scfifo_1id1:auto_generated|a_dpfifo_up51:dpfifo|altsyncram_9an1:FIFOram|ALTSYNCRAM";
defparam ram_block1a13.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a13.operation_mode = "dual_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 5;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 31;
defparam ram_block1a13.port_a_logical_ram_depth = 32;
defparam ram_block1a13.port_a_logical_ram_width = 29;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a13.port_b_address_clear = "none";
defparam ram_block1a13.port_b_address_clock = "clock1";
defparam ram_block1a13.port_b_address_width = 5;
defparam ram_block1a13.port_b_data_out_clear = "none";
defparam ram_block1a13.port_b_data_out_clock = "clock1";
defparam ram_block1a13.port_b_data_width = 1;
defparam ram_block1a13.port_b_first_address = 0;
defparam ram_block1a13.port_b_first_bit_number = 13;
defparam ram_block1a13.port_b_last_address = 31;
defparam ram_block1a13.port_b_logical_ram_depth = 32;
defparam ram_block1a13.port_b_logical_ram_width = 29;
defparam ram_block1a13.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a13.port_b_read_enable_clock = "clock1";
defparam ram_block1a13.ram_block_type = "auto";

arriav_ram_block ram_block1a14(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a14_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a14.clk0_core_clock_enable = "ena0";
defparam ram_block1a14.clk1_output_clock_enable = "ena1";
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_source:output_source_0|scfifo:source_FIFO|scfifo_1id1:auto_generated|a_dpfifo_up51:dpfifo|altsyncram_9an1:FIFOram|ALTSYNCRAM";
defparam ram_block1a14.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a14.operation_mode = "dual_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 5;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 31;
defparam ram_block1a14.port_a_logical_ram_depth = 32;
defparam ram_block1a14.port_a_logical_ram_width = 29;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a14.port_b_address_clear = "none";
defparam ram_block1a14.port_b_address_clock = "clock1";
defparam ram_block1a14.port_b_address_width = 5;
defparam ram_block1a14.port_b_data_out_clear = "none";
defparam ram_block1a14.port_b_data_out_clock = "clock1";
defparam ram_block1a14.port_b_data_width = 1;
defparam ram_block1a14.port_b_first_address = 0;
defparam ram_block1a14.port_b_first_bit_number = 14;
defparam ram_block1a14.port_b_last_address = 31;
defparam ram_block1a14.port_b_logical_ram_depth = 32;
defparam ram_block1a14.port_b_logical_ram_width = 29;
defparam ram_block1a14.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a14.port_b_read_enable_clock = "clock1";
defparam ram_block1a14.ram_block_type = "auto";

arriav_ram_block ram_block1a15(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a15_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a15.clk0_core_clock_enable = "ena0";
defparam ram_block1a15.clk1_output_clock_enable = "ena1";
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_source:output_source_0|scfifo:source_FIFO|scfifo_1id1:auto_generated|a_dpfifo_up51:dpfifo|altsyncram_9an1:FIFOram|ALTSYNCRAM";
defparam ram_block1a15.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a15.operation_mode = "dual_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 5;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 31;
defparam ram_block1a15.port_a_logical_ram_depth = 32;
defparam ram_block1a15.port_a_logical_ram_width = 29;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a15.port_b_address_clear = "none";
defparam ram_block1a15.port_b_address_clock = "clock1";
defparam ram_block1a15.port_b_address_width = 5;
defparam ram_block1a15.port_b_data_out_clear = "none";
defparam ram_block1a15.port_b_data_out_clock = "clock1";
defparam ram_block1a15.port_b_data_width = 1;
defparam ram_block1a15.port_b_first_address = 0;
defparam ram_block1a15.port_b_first_bit_number = 15;
defparam ram_block1a15.port_b_last_address = 31;
defparam ram_block1a15.port_b_logical_ram_depth = 32;
defparam ram_block1a15.port_b_logical_ram_width = 29;
defparam ram_block1a15.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a15.port_b_read_enable_clock = "clock1";
defparam ram_block1a15.ram_block_type = "auto";

arriav_ram_block ram_block1a16(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a16_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a16.clk0_core_clock_enable = "ena0";
defparam ram_block1a16.clk1_output_clock_enable = "ena1";
defparam ram_block1a16.data_interleave_offset_in_bits = 1;
defparam ram_block1a16.data_interleave_width_in_bits = 1;
defparam ram_block1a16.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_source:output_source_0|scfifo:source_FIFO|scfifo_1id1:auto_generated|a_dpfifo_up51:dpfifo|altsyncram_9an1:FIFOram|ALTSYNCRAM";
defparam ram_block1a16.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a16.operation_mode = "dual_port";
defparam ram_block1a16.port_a_address_clear = "none";
defparam ram_block1a16.port_a_address_width = 5;
defparam ram_block1a16.port_a_data_out_clear = "none";
defparam ram_block1a16.port_a_data_out_clock = "none";
defparam ram_block1a16.port_a_data_width = 1;
defparam ram_block1a16.port_a_first_address = 0;
defparam ram_block1a16.port_a_first_bit_number = 16;
defparam ram_block1a16.port_a_last_address = 31;
defparam ram_block1a16.port_a_logical_ram_depth = 32;
defparam ram_block1a16.port_a_logical_ram_width = 29;
defparam ram_block1a16.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a16.port_b_address_clear = "none";
defparam ram_block1a16.port_b_address_clock = "clock1";
defparam ram_block1a16.port_b_address_width = 5;
defparam ram_block1a16.port_b_data_out_clear = "none";
defparam ram_block1a16.port_b_data_out_clock = "clock1";
defparam ram_block1a16.port_b_data_width = 1;
defparam ram_block1a16.port_b_first_address = 0;
defparam ram_block1a16.port_b_first_bit_number = 16;
defparam ram_block1a16.port_b_last_address = 31;
defparam ram_block1a16.port_b_logical_ram_depth = 32;
defparam ram_block1a16.port_b_logical_ram_width = 29;
defparam ram_block1a16.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a16.port_b_read_enable_clock = "clock1";
defparam ram_block1a16.ram_block_type = "auto";

arriav_ram_block ram_block1a17(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[17]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a17_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a17.clk0_core_clock_enable = "ena0";
defparam ram_block1a17.clk1_output_clock_enable = "ena1";
defparam ram_block1a17.data_interleave_offset_in_bits = 1;
defparam ram_block1a17.data_interleave_width_in_bits = 1;
defparam ram_block1a17.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_source:output_source_0|scfifo:source_FIFO|scfifo_1id1:auto_generated|a_dpfifo_up51:dpfifo|altsyncram_9an1:FIFOram|ALTSYNCRAM";
defparam ram_block1a17.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a17.operation_mode = "dual_port";
defparam ram_block1a17.port_a_address_clear = "none";
defparam ram_block1a17.port_a_address_width = 5;
defparam ram_block1a17.port_a_data_out_clear = "none";
defparam ram_block1a17.port_a_data_out_clock = "none";
defparam ram_block1a17.port_a_data_width = 1;
defparam ram_block1a17.port_a_first_address = 0;
defparam ram_block1a17.port_a_first_bit_number = 17;
defparam ram_block1a17.port_a_last_address = 31;
defparam ram_block1a17.port_a_logical_ram_depth = 32;
defparam ram_block1a17.port_a_logical_ram_width = 29;
defparam ram_block1a17.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a17.port_b_address_clear = "none";
defparam ram_block1a17.port_b_address_clock = "clock1";
defparam ram_block1a17.port_b_address_width = 5;
defparam ram_block1a17.port_b_data_out_clear = "none";
defparam ram_block1a17.port_b_data_out_clock = "clock1";
defparam ram_block1a17.port_b_data_width = 1;
defparam ram_block1a17.port_b_first_address = 0;
defparam ram_block1a17.port_b_first_bit_number = 17;
defparam ram_block1a17.port_b_last_address = 31;
defparam ram_block1a17.port_b_logical_ram_depth = 32;
defparam ram_block1a17.port_b_logical_ram_width = 29;
defparam ram_block1a17.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a17.port_b_read_enable_clock = "clock1";
defparam ram_block1a17.ram_block_type = "auto";

arriav_ram_block ram_block1a18(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[18]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a18_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a18.clk0_core_clock_enable = "ena0";
defparam ram_block1a18.clk1_output_clock_enable = "ena1";
defparam ram_block1a18.data_interleave_offset_in_bits = 1;
defparam ram_block1a18.data_interleave_width_in_bits = 1;
defparam ram_block1a18.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_source:output_source_0|scfifo:source_FIFO|scfifo_1id1:auto_generated|a_dpfifo_up51:dpfifo|altsyncram_9an1:FIFOram|ALTSYNCRAM";
defparam ram_block1a18.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a18.operation_mode = "dual_port";
defparam ram_block1a18.port_a_address_clear = "none";
defparam ram_block1a18.port_a_address_width = 5;
defparam ram_block1a18.port_a_data_out_clear = "none";
defparam ram_block1a18.port_a_data_out_clock = "none";
defparam ram_block1a18.port_a_data_width = 1;
defparam ram_block1a18.port_a_first_address = 0;
defparam ram_block1a18.port_a_first_bit_number = 18;
defparam ram_block1a18.port_a_last_address = 31;
defparam ram_block1a18.port_a_logical_ram_depth = 32;
defparam ram_block1a18.port_a_logical_ram_width = 29;
defparam ram_block1a18.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a18.port_b_address_clear = "none";
defparam ram_block1a18.port_b_address_clock = "clock1";
defparam ram_block1a18.port_b_address_width = 5;
defparam ram_block1a18.port_b_data_out_clear = "none";
defparam ram_block1a18.port_b_data_out_clock = "clock1";
defparam ram_block1a18.port_b_data_width = 1;
defparam ram_block1a18.port_b_first_address = 0;
defparam ram_block1a18.port_b_first_bit_number = 18;
defparam ram_block1a18.port_b_last_address = 31;
defparam ram_block1a18.port_b_logical_ram_depth = 32;
defparam ram_block1a18.port_b_logical_ram_width = 29;
defparam ram_block1a18.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a18.port_b_read_enable_clock = "clock1";
defparam ram_block1a18.ram_block_type = "auto";

arriav_ram_block ram_block1a19(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[19]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a19_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a19.clk0_core_clock_enable = "ena0";
defparam ram_block1a19.clk1_output_clock_enable = "ena1";
defparam ram_block1a19.data_interleave_offset_in_bits = 1;
defparam ram_block1a19.data_interleave_width_in_bits = 1;
defparam ram_block1a19.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_source:output_source_0|scfifo:source_FIFO|scfifo_1id1:auto_generated|a_dpfifo_up51:dpfifo|altsyncram_9an1:FIFOram|ALTSYNCRAM";
defparam ram_block1a19.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a19.operation_mode = "dual_port";
defparam ram_block1a19.port_a_address_clear = "none";
defparam ram_block1a19.port_a_address_width = 5;
defparam ram_block1a19.port_a_data_out_clear = "none";
defparam ram_block1a19.port_a_data_out_clock = "none";
defparam ram_block1a19.port_a_data_width = 1;
defparam ram_block1a19.port_a_first_address = 0;
defparam ram_block1a19.port_a_first_bit_number = 19;
defparam ram_block1a19.port_a_last_address = 31;
defparam ram_block1a19.port_a_logical_ram_depth = 32;
defparam ram_block1a19.port_a_logical_ram_width = 29;
defparam ram_block1a19.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a19.port_b_address_clear = "none";
defparam ram_block1a19.port_b_address_clock = "clock1";
defparam ram_block1a19.port_b_address_width = 5;
defparam ram_block1a19.port_b_data_out_clear = "none";
defparam ram_block1a19.port_b_data_out_clock = "clock1";
defparam ram_block1a19.port_b_data_width = 1;
defparam ram_block1a19.port_b_first_address = 0;
defparam ram_block1a19.port_b_first_bit_number = 19;
defparam ram_block1a19.port_b_last_address = 31;
defparam ram_block1a19.port_b_logical_ram_depth = 32;
defparam ram_block1a19.port_b_logical_ram_width = 29;
defparam ram_block1a19.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a19.port_b_read_enable_clock = "clock1";
defparam ram_block1a19.ram_block_type = "auto";

arriav_ram_block ram_block1a20(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[20]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a20_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a20.clk0_core_clock_enable = "ena0";
defparam ram_block1a20.clk1_output_clock_enable = "ena1";
defparam ram_block1a20.data_interleave_offset_in_bits = 1;
defparam ram_block1a20.data_interleave_width_in_bits = 1;
defparam ram_block1a20.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_source:output_source_0|scfifo:source_FIFO|scfifo_1id1:auto_generated|a_dpfifo_up51:dpfifo|altsyncram_9an1:FIFOram|ALTSYNCRAM";
defparam ram_block1a20.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a20.operation_mode = "dual_port";
defparam ram_block1a20.port_a_address_clear = "none";
defparam ram_block1a20.port_a_address_width = 5;
defparam ram_block1a20.port_a_data_out_clear = "none";
defparam ram_block1a20.port_a_data_out_clock = "none";
defparam ram_block1a20.port_a_data_width = 1;
defparam ram_block1a20.port_a_first_address = 0;
defparam ram_block1a20.port_a_first_bit_number = 20;
defparam ram_block1a20.port_a_last_address = 31;
defparam ram_block1a20.port_a_logical_ram_depth = 32;
defparam ram_block1a20.port_a_logical_ram_width = 29;
defparam ram_block1a20.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a20.port_b_address_clear = "none";
defparam ram_block1a20.port_b_address_clock = "clock1";
defparam ram_block1a20.port_b_address_width = 5;
defparam ram_block1a20.port_b_data_out_clear = "none";
defparam ram_block1a20.port_b_data_out_clock = "clock1";
defparam ram_block1a20.port_b_data_width = 1;
defparam ram_block1a20.port_b_first_address = 0;
defparam ram_block1a20.port_b_first_bit_number = 20;
defparam ram_block1a20.port_b_last_address = 31;
defparam ram_block1a20.port_b_logical_ram_depth = 32;
defparam ram_block1a20.port_b_logical_ram_width = 29;
defparam ram_block1a20.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a20.port_b_read_enable_clock = "clock1";
defparam ram_block1a20.ram_block_type = "auto";

arriav_ram_block ram_block1a21(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[21]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a21_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a21.clk0_core_clock_enable = "ena0";
defparam ram_block1a21.clk1_output_clock_enable = "ena1";
defparam ram_block1a21.data_interleave_offset_in_bits = 1;
defparam ram_block1a21.data_interleave_width_in_bits = 1;
defparam ram_block1a21.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_source:output_source_0|scfifo:source_FIFO|scfifo_1id1:auto_generated|a_dpfifo_up51:dpfifo|altsyncram_9an1:FIFOram|ALTSYNCRAM";
defparam ram_block1a21.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a21.operation_mode = "dual_port";
defparam ram_block1a21.port_a_address_clear = "none";
defparam ram_block1a21.port_a_address_width = 5;
defparam ram_block1a21.port_a_data_out_clear = "none";
defparam ram_block1a21.port_a_data_out_clock = "none";
defparam ram_block1a21.port_a_data_width = 1;
defparam ram_block1a21.port_a_first_address = 0;
defparam ram_block1a21.port_a_first_bit_number = 21;
defparam ram_block1a21.port_a_last_address = 31;
defparam ram_block1a21.port_a_logical_ram_depth = 32;
defparam ram_block1a21.port_a_logical_ram_width = 29;
defparam ram_block1a21.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a21.port_b_address_clear = "none";
defparam ram_block1a21.port_b_address_clock = "clock1";
defparam ram_block1a21.port_b_address_width = 5;
defparam ram_block1a21.port_b_data_out_clear = "none";
defparam ram_block1a21.port_b_data_out_clock = "clock1";
defparam ram_block1a21.port_b_data_width = 1;
defparam ram_block1a21.port_b_first_address = 0;
defparam ram_block1a21.port_b_first_bit_number = 21;
defparam ram_block1a21.port_b_last_address = 31;
defparam ram_block1a21.port_b_logical_ram_depth = 32;
defparam ram_block1a21.port_b_logical_ram_width = 29;
defparam ram_block1a21.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a21.port_b_read_enable_clock = "clock1";
defparam ram_block1a21.ram_block_type = "auto";

arriav_ram_block ram_block1a22(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[22]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a22_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a22.clk0_core_clock_enable = "ena0";
defparam ram_block1a22.clk1_output_clock_enable = "ena1";
defparam ram_block1a22.data_interleave_offset_in_bits = 1;
defparam ram_block1a22.data_interleave_width_in_bits = 1;
defparam ram_block1a22.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_source:output_source_0|scfifo:source_FIFO|scfifo_1id1:auto_generated|a_dpfifo_up51:dpfifo|altsyncram_9an1:FIFOram|ALTSYNCRAM";
defparam ram_block1a22.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a22.operation_mode = "dual_port";
defparam ram_block1a22.port_a_address_clear = "none";
defparam ram_block1a22.port_a_address_width = 5;
defparam ram_block1a22.port_a_data_out_clear = "none";
defparam ram_block1a22.port_a_data_out_clock = "none";
defparam ram_block1a22.port_a_data_width = 1;
defparam ram_block1a22.port_a_first_address = 0;
defparam ram_block1a22.port_a_first_bit_number = 22;
defparam ram_block1a22.port_a_last_address = 31;
defparam ram_block1a22.port_a_logical_ram_depth = 32;
defparam ram_block1a22.port_a_logical_ram_width = 29;
defparam ram_block1a22.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a22.port_b_address_clear = "none";
defparam ram_block1a22.port_b_address_clock = "clock1";
defparam ram_block1a22.port_b_address_width = 5;
defparam ram_block1a22.port_b_data_out_clear = "none";
defparam ram_block1a22.port_b_data_out_clock = "clock1";
defparam ram_block1a22.port_b_data_width = 1;
defparam ram_block1a22.port_b_first_address = 0;
defparam ram_block1a22.port_b_first_bit_number = 22;
defparam ram_block1a22.port_b_last_address = 31;
defparam ram_block1a22.port_b_logical_ram_depth = 32;
defparam ram_block1a22.port_b_logical_ram_width = 29;
defparam ram_block1a22.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a22.port_b_read_enable_clock = "clock1";
defparam ram_block1a22.ram_block_type = "auto";

arriav_ram_block ram_block1a23(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[23]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a23_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a23.clk0_core_clock_enable = "ena0";
defparam ram_block1a23.clk1_output_clock_enable = "ena1";
defparam ram_block1a23.data_interleave_offset_in_bits = 1;
defparam ram_block1a23.data_interleave_width_in_bits = 1;
defparam ram_block1a23.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_source:output_source_0|scfifo:source_FIFO|scfifo_1id1:auto_generated|a_dpfifo_up51:dpfifo|altsyncram_9an1:FIFOram|ALTSYNCRAM";
defparam ram_block1a23.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a23.operation_mode = "dual_port";
defparam ram_block1a23.port_a_address_clear = "none";
defparam ram_block1a23.port_a_address_width = 5;
defparam ram_block1a23.port_a_data_out_clear = "none";
defparam ram_block1a23.port_a_data_out_clock = "none";
defparam ram_block1a23.port_a_data_width = 1;
defparam ram_block1a23.port_a_first_address = 0;
defparam ram_block1a23.port_a_first_bit_number = 23;
defparam ram_block1a23.port_a_last_address = 31;
defparam ram_block1a23.port_a_logical_ram_depth = 32;
defparam ram_block1a23.port_a_logical_ram_width = 29;
defparam ram_block1a23.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a23.port_b_address_clear = "none";
defparam ram_block1a23.port_b_address_clock = "clock1";
defparam ram_block1a23.port_b_address_width = 5;
defparam ram_block1a23.port_b_data_out_clear = "none";
defparam ram_block1a23.port_b_data_out_clock = "clock1";
defparam ram_block1a23.port_b_data_width = 1;
defparam ram_block1a23.port_b_first_address = 0;
defparam ram_block1a23.port_b_first_bit_number = 23;
defparam ram_block1a23.port_b_last_address = 31;
defparam ram_block1a23.port_b_logical_ram_depth = 32;
defparam ram_block1a23.port_b_logical_ram_width = 29;
defparam ram_block1a23.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a23.port_b_read_enable_clock = "clock1";
defparam ram_block1a23.ram_block_type = "auto";

arriav_ram_block ram_block1a24(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[24]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a24_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a24.clk0_core_clock_enable = "ena0";
defparam ram_block1a24.clk1_output_clock_enable = "ena1";
defparam ram_block1a24.data_interleave_offset_in_bits = 1;
defparam ram_block1a24.data_interleave_width_in_bits = 1;
defparam ram_block1a24.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_source:output_source_0|scfifo:source_FIFO|scfifo_1id1:auto_generated|a_dpfifo_up51:dpfifo|altsyncram_9an1:FIFOram|ALTSYNCRAM";
defparam ram_block1a24.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a24.operation_mode = "dual_port";
defparam ram_block1a24.port_a_address_clear = "none";
defparam ram_block1a24.port_a_address_width = 5;
defparam ram_block1a24.port_a_data_out_clear = "none";
defparam ram_block1a24.port_a_data_out_clock = "none";
defparam ram_block1a24.port_a_data_width = 1;
defparam ram_block1a24.port_a_first_address = 0;
defparam ram_block1a24.port_a_first_bit_number = 24;
defparam ram_block1a24.port_a_last_address = 31;
defparam ram_block1a24.port_a_logical_ram_depth = 32;
defparam ram_block1a24.port_a_logical_ram_width = 29;
defparam ram_block1a24.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a24.port_b_address_clear = "none";
defparam ram_block1a24.port_b_address_clock = "clock1";
defparam ram_block1a24.port_b_address_width = 5;
defparam ram_block1a24.port_b_data_out_clear = "none";
defparam ram_block1a24.port_b_data_out_clock = "clock1";
defparam ram_block1a24.port_b_data_width = 1;
defparam ram_block1a24.port_b_first_address = 0;
defparam ram_block1a24.port_b_first_bit_number = 24;
defparam ram_block1a24.port_b_last_address = 31;
defparam ram_block1a24.port_b_logical_ram_depth = 32;
defparam ram_block1a24.port_b_logical_ram_width = 29;
defparam ram_block1a24.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a24.port_b_read_enable_clock = "clock1";
defparam ram_block1a24.ram_block_type = "auto";

arriav_ram_block ram_block1a25(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[25]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a25_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a25.clk0_core_clock_enable = "ena0";
defparam ram_block1a25.clk1_output_clock_enable = "ena1";
defparam ram_block1a25.data_interleave_offset_in_bits = 1;
defparam ram_block1a25.data_interleave_width_in_bits = 1;
defparam ram_block1a25.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_source:output_source_0|scfifo:source_FIFO|scfifo_1id1:auto_generated|a_dpfifo_up51:dpfifo|altsyncram_9an1:FIFOram|ALTSYNCRAM";
defparam ram_block1a25.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a25.operation_mode = "dual_port";
defparam ram_block1a25.port_a_address_clear = "none";
defparam ram_block1a25.port_a_address_width = 5;
defparam ram_block1a25.port_a_data_out_clear = "none";
defparam ram_block1a25.port_a_data_out_clock = "none";
defparam ram_block1a25.port_a_data_width = 1;
defparam ram_block1a25.port_a_first_address = 0;
defparam ram_block1a25.port_a_first_bit_number = 25;
defparam ram_block1a25.port_a_last_address = 31;
defparam ram_block1a25.port_a_logical_ram_depth = 32;
defparam ram_block1a25.port_a_logical_ram_width = 29;
defparam ram_block1a25.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a25.port_b_address_clear = "none";
defparam ram_block1a25.port_b_address_clock = "clock1";
defparam ram_block1a25.port_b_address_width = 5;
defparam ram_block1a25.port_b_data_out_clear = "none";
defparam ram_block1a25.port_b_data_out_clock = "clock1";
defparam ram_block1a25.port_b_data_width = 1;
defparam ram_block1a25.port_b_first_address = 0;
defparam ram_block1a25.port_b_first_bit_number = 25;
defparam ram_block1a25.port_b_last_address = 31;
defparam ram_block1a25.port_b_logical_ram_depth = 32;
defparam ram_block1a25.port_b_logical_ram_width = 29;
defparam ram_block1a25.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a25.port_b_read_enable_clock = "clock1";
defparam ram_block1a25.ram_block_type = "auto";

arriav_ram_block ram_block1a26(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[26]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a26_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a26.clk0_core_clock_enable = "ena0";
defparam ram_block1a26.clk1_output_clock_enable = "ena1";
defparam ram_block1a26.data_interleave_offset_in_bits = 1;
defparam ram_block1a26.data_interleave_width_in_bits = 1;
defparam ram_block1a26.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_source:output_source_0|scfifo:source_FIFO|scfifo_1id1:auto_generated|a_dpfifo_up51:dpfifo|altsyncram_9an1:FIFOram|ALTSYNCRAM";
defparam ram_block1a26.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a26.operation_mode = "dual_port";
defparam ram_block1a26.port_a_address_clear = "none";
defparam ram_block1a26.port_a_address_width = 5;
defparam ram_block1a26.port_a_data_out_clear = "none";
defparam ram_block1a26.port_a_data_out_clock = "none";
defparam ram_block1a26.port_a_data_width = 1;
defparam ram_block1a26.port_a_first_address = 0;
defparam ram_block1a26.port_a_first_bit_number = 26;
defparam ram_block1a26.port_a_last_address = 31;
defparam ram_block1a26.port_a_logical_ram_depth = 32;
defparam ram_block1a26.port_a_logical_ram_width = 29;
defparam ram_block1a26.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a26.port_b_address_clear = "none";
defparam ram_block1a26.port_b_address_clock = "clock1";
defparam ram_block1a26.port_b_address_width = 5;
defparam ram_block1a26.port_b_data_out_clear = "none";
defparam ram_block1a26.port_b_data_out_clock = "clock1";
defparam ram_block1a26.port_b_data_width = 1;
defparam ram_block1a26.port_b_first_address = 0;
defparam ram_block1a26.port_b_first_bit_number = 26;
defparam ram_block1a26.port_b_last_address = 31;
defparam ram_block1a26.port_b_logical_ram_depth = 32;
defparam ram_block1a26.port_b_logical_ram_width = 29;
defparam ram_block1a26.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a26.port_b_read_enable_clock = "clock1";
defparam ram_block1a26.ram_block_type = "auto";

arriav_ram_block ram_block1a27(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[27]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a27_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a27.clk0_core_clock_enable = "ena0";
defparam ram_block1a27.clk1_output_clock_enable = "ena1";
defparam ram_block1a27.data_interleave_offset_in_bits = 1;
defparam ram_block1a27.data_interleave_width_in_bits = 1;
defparam ram_block1a27.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_source:output_source_0|scfifo:source_FIFO|scfifo_1id1:auto_generated|a_dpfifo_up51:dpfifo|altsyncram_9an1:FIFOram|ALTSYNCRAM";
defparam ram_block1a27.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a27.operation_mode = "dual_port";
defparam ram_block1a27.port_a_address_clear = "none";
defparam ram_block1a27.port_a_address_width = 5;
defparam ram_block1a27.port_a_data_out_clear = "none";
defparam ram_block1a27.port_a_data_out_clock = "none";
defparam ram_block1a27.port_a_data_width = 1;
defparam ram_block1a27.port_a_first_address = 0;
defparam ram_block1a27.port_a_first_bit_number = 27;
defparam ram_block1a27.port_a_last_address = 31;
defparam ram_block1a27.port_a_logical_ram_depth = 32;
defparam ram_block1a27.port_a_logical_ram_width = 29;
defparam ram_block1a27.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a27.port_b_address_clear = "none";
defparam ram_block1a27.port_b_address_clock = "clock1";
defparam ram_block1a27.port_b_address_width = 5;
defparam ram_block1a27.port_b_data_out_clear = "none";
defparam ram_block1a27.port_b_data_out_clock = "clock1";
defparam ram_block1a27.port_b_data_width = 1;
defparam ram_block1a27.port_b_first_address = 0;
defparam ram_block1a27.port_b_first_bit_number = 27;
defparam ram_block1a27.port_b_last_address = 31;
defparam ram_block1a27.port_b_logical_ram_depth = 32;
defparam ram_block1a27.port_b_logical_ram_width = 29;
defparam ram_block1a27.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a27.port_b_read_enable_clock = "clock1";
defparam ram_block1a27.ram_block_type = "auto";

endmodule

module cic_cntr_hra (
	source_valid_s,
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_2,
	counter_reg_bit_3,
	empty_dff,
	rd_ptr_lsb,
	clock,
	sclr,
	out_ready)/* synthesis synthesis_greybox=1 */;
input 	source_valid_s;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
output 	counter_reg_bit_3;
input 	empty_dff;
input 	rd_ptr_lsb;
input 	clock;
input 	sclr;
input 	out_ready;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~sumout ;
wire \_~0_combout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~sumout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~sumout ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~sumout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!sclr),
	.sload(gnd),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!sclr),
	.sload(gnd),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!sclr),
	.sload(gnd),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!sclr),
	.sload(gnd),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

arriav_lcell_comb counter_comb_bita0(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita0~sumout ),
	.cout(\counter_comb_bita0~COUT ),
	.shareout());
defparam counter_comb_bita0.extended_lut = "off";
defparam counter_comb_bita0.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita0.shared_arith = "off";

arriav_lcell_comb \_~0 (
	.dataa(!source_valid_s),
	.datab(!sclr),
	.datac(!empty_dff),
	.datad(!out_ready),
	.datae(!rd_ptr_lsb),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\_~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \_~0 .extended_lut = "off";
defparam \_~0 .lut_mask = 64'hFFFFEFFFFFFFEFFF;
defparam \_~0 .shared_arith = "off";

arriav_lcell_comb counter_comb_bita1(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita0~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita1~sumout ),
	.cout(\counter_comb_bita1~COUT ),
	.shareout());
defparam counter_comb_bita1.extended_lut = "off";
defparam counter_comb_bita1.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita1.shared_arith = "off";

arriav_lcell_comb counter_comb_bita2(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita1~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita2~sumout ),
	.cout(\counter_comb_bita2~COUT ),
	.shareout());
defparam counter_comb_bita2.extended_lut = "off";
defparam counter_comb_bita2.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita2.shared_arith = "off";

arriav_lcell_comb counter_comb_bita3(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita2~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita3~sumout ),
	.cout(),
	.shareout());
defparam counter_comb_bita3.extended_lut = "off";
defparam counter_comb_bita3.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita3.shared_arith = "off";

endmodule

module cic_cntr_ira (
	full_dff,
	dout_valid,
	state_0,
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_2,
	counter_reg_bit_3,
	counter_reg_bit_4,
	stall_reg,
	clock,
	sclr)/* synthesis synthesis_greybox=1 */;
input 	full_dff;
input 	dout_valid;
input 	state_0;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
output 	counter_reg_bit_3;
output 	counter_reg_bit_4;
input 	stall_reg;
input 	clock;
input 	sclr;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~sumout ;
wire \_~0_combout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~sumout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~sumout ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~sumout ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~sumout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!sclr),
	.sload(gnd),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!sclr),
	.sload(gnd),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!sclr),
	.sload(gnd),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!sclr),
	.sload(gnd),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!sclr),
	.sload(gnd),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

arriav_lcell_comb counter_comb_bita0(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita0~sumout ),
	.cout(\counter_comb_bita0~COUT ),
	.shareout());
defparam counter_comb_bita0.extended_lut = "off";
defparam counter_comb_bita0.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita0.shared_arith = "off";

arriav_lcell_comb \_~0 (
	.dataa(!sclr),
	.datab(!full_dff),
	.datac(!stall_reg),
	.datad(!dout_valid),
	.datae(!state_0),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\_~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \_~0 .extended_lut = "off";
defparam \_~0 .lut_mask = 64'hFEFFFFFFFEFFFFFF;
defparam \_~0 .shared_arith = "off";

arriav_lcell_comb counter_comb_bita1(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita0~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita1~sumout ),
	.cout(\counter_comb_bita1~COUT ),
	.shareout());
defparam counter_comb_bita1.extended_lut = "off";
defparam counter_comb_bita1.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita1.shared_arith = "off";

arriav_lcell_comb counter_comb_bita2(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita1~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita2~sumout ),
	.cout(\counter_comb_bita2~COUT ),
	.shareout());
defparam counter_comb_bita2.extended_lut = "off";
defparam counter_comb_bita2.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita2.shared_arith = "off";

arriav_lcell_comb counter_comb_bita3(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita2~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita3~sumout ),
	.cout(\counter_comb_bita3~COUT ),
	.shareout());
defparam counter_comb_bita3.extended_lut = "off";
defparam counter_comb_bita3.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita3.shared_arith = "off";

arriav_lcell_comb counter_comb_bita4(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita3~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita4~sumout ),
	.cout(),
	.shareout());
defparam counter_comb_bita4.extended_lut = "off";
defparam counter_comb_bita4.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita4.shared_arith = "off";

endmodule

module cic_cntr_ur6 (
	source_valid_s,
	counter_reg_bit_0,
	counter_reg_bit_4,
	counter_reg_bit_3,
	counter_reg_bit_2,
	counter_reg_bit_1,
	valid_wreq,
	empty_dff,
	clock,
	sclr,
	out_ready)/* synthesis synthesis_greybox=1 */;
input 	source_valid_s;
output 	counter_reg_bit_0;
output 	counter_reg_bit_4;
output 	counter_reg_bit_3;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
input 	valid_wreq;
input 	empty_dff;
input 	clock;
input 	sclr;
input 	out_ready;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~sumout ;
wire \_~0_combout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~sumout ;
wire \counter_comb_bita3~sumout ;
wire \counter_comb_bita2~sumout ;
wire \counter_comb_bita1~sumout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!sclr),
	.sload(gnd),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!sclr),
	.sload(gnd),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!sclr),
	.sload(gnd),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!sclr),
	.sload(gnd),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!sclr),
	.sload(gnd),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

arriav_lcell_comb counter_comb_bita0(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita0~sumout ),
	.cout(\counter_comb_bita0~COUT ),
	.shareout());
defparam counter_comb_bita0.extended_lut = "off";
defparam counter_comb_bita0.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita0.shared_arith = "off";

arriav_lcell_comb \_~0 (
	.dataa(!source_valid_s),
	.datab(!sclr),
	.datac(!valid_wreq),
	.datad(!empty_dff),
	.datae(!out_ready),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\_~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \_~0 .extended_lut = "off";
defparam \_~0 .lut_mask = 64'hDEEDEDDEDEEDEDDE;
defparam \_~0 .shared_arith = "off";

arriav_lcell_comb counter_comb_bita1(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_1),
	.datae(gnd),
	.dataf(!valid_wreq),
	.datag(gnd),
	.cin(\counter_comb_bita0~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita1~sumout ),
	.cout(\counter_comb_bita1~COUT ),
	.shareout());
defparam counter_comb_bita1.extended_lut = "off";
defparam counter_comb_bita1.lut_mask = 64'h000000FF000000FF;
defparam counter_comb_bita1.shared_arith = "off";

arriav_lcell_comb counter_comb_bita2(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_2),
	.datae(gnd),
	.dataf(!valid_wreq),
	.datag(gnd),
	.cin(\counter_comb_bita1~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita2~sumout ),
	.cout(\counter_comb_bita2~COUT ),
	.shareout());
defparam counter_comb_bita2.extended_lut = "off";
defparam counter_comb_bita2.lut_mask = 64'h000000FF000000FF;
defparam counter_comb_bita2.shared_arith = "off";

arriav_lcell_comb counter_comb_bita3(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_3),
	.datae(gnd),
	.dataf(!valid_wreq),
	.datag(gnd),
	.cin(\counter_comb_bita2~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita3~sumout ),
	.cout(\counter_comb_bita3~COUT ),
	.shareout());
defparam counter_comb_bita3.extended_lut = "off";
defparam counter_comb_bita3.lut_mask = 64'h000000FF000000FF;
defparam counter_comb_bita3.shared_arith = "off";

arriav_lcell_comb counter_comb_bita4(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_4),
	.datae(gnd),
	.dataf(!valid_wreq),
	.datag(gnd),
	.cin(\counter_comb_bita3~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita4~sumout ),
	.cout(),
	.shareout());
defparam counter_comb_bita4.extended_lut = "off";
defparam counter_comb_bita4.lut_mask = 64'h000000FF000000FF;
defparam counter_comb_bita4.shared_arith = "off";

endmodule
