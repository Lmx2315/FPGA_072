// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.0std
// ALTERA_TIMESTAMP:Wed Apr 26 13:33:39 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
fy1Y6+d7PbnCXWpBVuyIoXcNSuU8esUUcfJQbuUF5KReLnyXzNZ1EXYUFQqM4mOf
/WhaJiNl8FyCVaSZbMztG1CM1/tp1d1fvgfX5kS+Skt4RdI44s1twWXVpP7aipbN
96zhCcMX8YTcoiuNuCNRJ3jSyt3VNlCwdqBWgndpMs0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7696)
DvfBmtTIZQf2mdkSVgLBgo/S5RWIjixLxXS92UD7MXfNb7FqeJvfd+oDWbV/maEE
yQBn4Bb1oi8eKTlIY2/y1rGy9leDkz46s87+LvMS9VsUEwiYfXy0JSZDBLaYvWcb
92XB/U1EZhrfO8Ht86nvHk4ryjci1VlA18DW9Z4tM0ZmUJguTU0ocqelk9+dKsdi
+zkAMo8UlyyU5zo4toxevTTvC9sjLTxIUVlIoCisz07I8vdmkv9Wgw8iNStw9dAr
dpfyNjOcZGeLysdiRm1+1Pr2fRettm69mtOjXNnRmXbnhtyDfK+mSuKInjKjuJ9L
W2hM+gHL4LB6Bb3dkTjctmMP1ysJvjon3cvVPinqIDzT+317EezECBmOgFpGSwZh
tiT3va1UXma2UYo6rP6ibqIEAqD8/oG4rfnSJH0yd3J2MDZBCpozSFwysRyWnbPN
2p7RVQQrFQOsTIvCji03yRkBo1GO6ckWXM+fD9x2N+UOls+UULpgPtd0x7jJ+MTe
0nWMd0gruSEErUdcsqKY6r1jXI7DF5vqL2Oid9b6qpslYL8CF6aqetK7xXGakXGk
koPWLj5IxRDcsaW5+zkxKBUq/7uLjdZZD/wY7I54PfOglIdHj22PhycrEUf3YzQG
8dgSrktGAGn/qqSCo6nBJsxrh6luMFCz0pIvi2odU487TJCV56SGJi3wS3NKLtV8
XG/B+/DdFmw+W7d9da8ctlv6hOz0Wt9+zoFatU6P6+2Llsbyi8nLzF6aAYLHf4DK
nRUapRDwgZdpzAhGjA3PFzsEtlnqe0AFWbcoUqSncFZJZHJDxQrtqD5oXUViosf8
c2kZRJPhRaProeQStSB/D8lVP/wHJkb/aTF7mMIBPNVmjONP7p0I5isgeKIPYxq+
5MIo8mC6/81WtD20fTENAbWjc3ci/OPjXOy4xNRn2PEb/LX6qWVck31v6N1bEy9j
LF4BnWDX3v6yiVIqNiBjFhwnhNAThZxArgq29GyOZQLMevzBa0r+flG15tLXeFl1
bxmh69tASe/stjPKsTDZAwT8w7WhqesG0wK/lVscOHaA+HoRhImtgOiljt5uC1qu
xw9DM13T0LCORUwYUYSpIRa2Ra4rZfjTa4bkhD4R7MS8Fvs1dyBwV0Y4BZqrYRqp
GxlUBTUVTAeo3+uiHHBXX1OLW+fWupU3j3APcmheecYpGDQG8+LXaHngT/lBHHln
nKVNNDbd87NglWPXPxyo6J1H1DlKkePF8iFd1RwkNkl5U83DIEInFLq0K2sJON45
r/sxtDq3Xqj4fcCYCw9k3V8hbmfwuEpeup1y+8i+BOokZLJeyjfq4qebGpdQcnJ7
EBe+/FZm/izExTbTySBHUaRsb2Yuvw16myFe+FPAuwzTI9Oqed/Qolv33p1m2tlT
4tliDcngPEvPLzLz6HrNSCTsZpeYufFZqhkH7ku0ExKbeDpdnEQOSqRK6Ybytnwe
gGqzDONeyMijdsOzTic9Gj0i5T9ebC55fMsaq3bHbPDglUHYUTYGwpgyFtb1asRU
uYX6VL+MKGAKjfGhsWDeshsgyEEASZgfLTs554kP3qGMnVBcLFprfa4ekqwW5JZp
XjmMeHxkGX2wrpkPsIg8lL9sbNIuEmfoTOOPh7rCek0oo5vxIsprvMshFNuQpWBd
V62v1dySNq9p4x911bym0ENFz8x1gSFohqJjvk78fLiiEtRSYCHSpb2HbtxZCj/K
nyucE5rywhe9DQTf7QDqvrTOwqBzNYLnJ3bUWWyG+d1CFajLX1KQFOlKbcxrwoG5
1BhPezvifiwzIcBjArL6OpdbY33KwfxiJf3UZKF6gdNDJL2cfXYPjQlL86SlK1GD
Nt79Dvt60OCtWYpbT6Xy48Cb79hPs5B3xFzCg3UBZp+XGt2m3kwuXO1XVTQRmDyW
fzLHvVTuV4KX97oeDdmALCBz25ul7x1yo5q+AMLvTgjsTbD4Kudh3NCXWhzudGzW
Z3sCYANn0kJEL+2acCjgapVGVdG1XNlKLEHVVIrRQa+w2OCw7Hh35jNAAAaPGMqY
OzyWeykRODPbbSs1kUMl5hoIMQqhMr1CxGWHCa6DG+lpMAQOMpfpXyl86BXD5uby
XAP5dlSnFvmE0woul5h8ETYXFZeI9gXYmrX7sLIItKiOeuggn24fSpH13qrEJFuq
+/ZjPZNj9yGDh3T4Xn8eKipNpvVbUV24lR52QBXu4TUxlSoMdvfyCnIvmvxZ3Omb
YUU3nA9or28WaghAfWzwr3saGF87pCOeV4yYBWgzPXJemlKFA4XzUrp1u4b5L1IB
YWljKLL1OvRF68G6A+6e5pvGdin6XewuRTmLcRsmxApYkNw4dTW21GBoeluJrSGi
9MmJAfQU55HTLJCik+xEGjoydmX7m+Ilm9rWbRumQtKMkTvFfHpt5fOHoN1MpW8f
rcADuZR33t8b56J/aLWvApWZ6TIXNpxoca2MmBo6csr7GTK1GbTxlmyVN+0dl45Q
1C1zAtA9RAtUwqFZzes/SHVSqHH8mBUNKendxurzPwM1yWmUe0mtAYKriSDTVA15
pohWD1P3O8GiQTU4UsfvkZkCJyHDz/0Wg9bXquy792Y93kPAqvAV4d1V+5C6/60i
PWYfm2ywqoKBuNQ6amA/colvJRQ978CZixERss0wJqStdqP5Ru/ceRxGKrYE59zj
mW6Mo/QM0xUdq/UiLNffwNJxLdNAbHzkxHpazqJ7HhytCuSZNjCCIJ/sq5hluB52
B3OAQi4OKi0WE9m7PV9yICYdGjxwCfBYQmdCI7OGo6T4kO9RLUMEXvPj2M2v56ID
KbeP+eOlzEKNM9+4lsf2BXVGmzAvWQlonN/YaCUZJ5v2w25HJExrA57TO8ZOb9/v
ylY+ghKF4bYfk2E8mM48vG3h9DhtoDOXzlQSzxrawSQ0UaC2BlybiTisc/C1cSbb
KDuCwSDgqf7vJbhjX/YY2ewCgh4XH/gpvvjPaGATLgMSeWzYJvAU1YKI2M555FSL
jU8EJIyG52WQSGHURzVyqEYMbkpebd/U+YyEe3sJ0AoFlvcdaaTfNJbwx/tXrGUW
w1ImtT5NHqKbnSqkVa3KVjHCNk9jdokSlW/uyxmJWH3JdIbHPvqRK0tjmlUGhPjm
zEVvxckThs8mWB/rpZeC/syUKnXLKZqfFhvDCwJOlYodZBtuDvQ4M9XGaOMaLcD0
cM7o2eIQO/QbVPj8YH33L1NzYu+Yj+o8SLydzx7dOg/ReQJ28ofKL5ZOgR7h4kni
zhg1lt+ungbmLqoAV10CXPvffD7oMHA4ZxcWO78GJmfmjDItg0X+TTZCCBBvHuCC
jitKSyuZAGnNmn3l+tvJWnLWuulfldzMEvRImEXl6e8DNxni9eNkx4mHKQDweKOl
RIz/MncfGYRNSj+HQUqvplH4ptUz/C11teUzJ8T9+ZNokCiihaTxRr9sAzF7Cds6
ohmHaufoICfMNflIbNrtEDKGx5TkHpbu1ZIt6xus5gsuANi8R0ZW4w1TXcjivROD
9Nf6y57BLjYJqPGYv+njBiqWUGxgkgrzjlezjlTyFv+l3WUDqZCr4hHYMuVm+V9V
cOqc69wFE9vPRaa5cS/P3IXDxexOl5KN5i5XttmzN2RSHRVEA3UTxXztx/m+pf4e
S/vQNyeYZxF0SB/tMU1V9nQJNuTvP3MXJYJ5VXkjBTGSAghUxpmAdyMCxSxv0OxC
UWf0ECEp04j8GgHpfSdZWcmmAm15BamZkpUPzvtUkkfCecAo+Ts9MXGnOHeCXm4D
X6iyboSVmDUElXATusEjBna98AREOho/GH3hX0VuPbRaIZa0/dN3FPTIozVdyNBI
5TW2pGSIHfTflt67xTriwZKA9T4l2zMtLdKFbdvS3zE0Oj1PuhHcjH3eL5uhwJ+B
jigfxI+7AMnEeRxNExY9gXXWErvUQwHMua/GcJMreAj6dyocfkRfli/SG/of06Kd
kH5aIqZ8QEwo6QCgNq57fjkgiXyteiJ8N9rAs7goJ+ymb+9/aoSudYeHMLGXJrgr
maGmjvQvf/q3oxdeqFLXkwqqPBpHrvhEKeyi+Mp9RQT57B5trxgC9OTcXi/lTrWF
d+ofpr72UwGNT7Qy1xjImAhyVpaKYbbsH5at4Bvp3mvUPpr7DVeVWb84W7/3A1l5
F/Sfi3+3SJJ2Wi0WJYxQdsBl7Q8wvY1NIDEdXTWDADBggju4PUKtMnRhJdCj+wc2
hnkpMAFMVLuAaFmzZFDQRPiSFbIQ/LFSnd2R58nQ77ITBV89OSh44xzhMzdZXZX0
1DqVJ/M/xPhPorZv9uhislobTQLd51jcBOt3eT51KrxKKcTfBS//tC0CWxQ5Xi7s
DD8cMsH1M9RM49TsLn5PuAIq55l1IQrsL5rfDNf0lMytqp1MrDSpbJY5w7rASMHN
O0gYChrDPZo9gu71VCahcjsIdFDjAQBC8ioXf47tWfIQOFBC4bvMKGBjoTYY2HlS
sLaKJlFmQy7Me/lPcMWkGPXcnLTLbzB8kRLD/894+vX4Do8n1qCZiY3aJrK4u94E
8SKj2HS6Nl4u5MXsQ5R8ZSyYw/Kr79V64CdFLU7BoZuAnVelQW8W/pbP8u3v8h/l
8Z0sT4S0nGbcnt8K8xdU/07S+VQQO0D0XgcxdW+qg6CuLxjBJptczSNNbOJkmzl0
p6MfbM2oD7D2wHUrzIUz8Ers6AHb69nGJqrF51k2405/bsIuRhoUkGwiqn5FYASl
cBQyaAF7bREECY1yguVKI6IANbsWG4A6xkbsnAOH351+8PoHyGO2yPTNek/QCAQZ
szb6H+xlj1au/ASeAgg/V/HBT1ZvA3KcPGi6/wNc47HYONynQGVTiQUzoEc55PuV
TcDD3u51pOib+fR9oktMgnh8Hjwzt3emdUyJ1ZwStMmJJjtljuLVLn6+GgszgJI6
ZUGE3GQYqjUOgTT3Eytb9hQjlk4LwsVzdE1hKxfqFQmTqE8fJ+Gy29pk0B5cbB3q
Gtefa3gLr5Wa4U+X3ayZ0dmb62niEihz6HOb4cUXdC76A1UdOU4o/RsLAdvrA6vw
+uRAOTpGkeGNL4lR41pi5l/Lfala+4YvYNfNkSblZvQjJ+tbjx/OoiggKE8cQBIc
AjgzcV4zXbp7MLA8uR16729VZy+rNRC0z2QA5peeUWkG2dmoPbfWJs+qiara1A4/
7n9MaAyjgl9UELzcbVbySiXqrnjC5yVdaB19UBTiK8C4tqxtcuaMMLbBP2nEs0ZQ
ccahwidLagNMPmuK4tu8hCR3yVXbHkOMNNT6nFI+cGnpxxB/y1QC2xJ2WM5Ll0fY
SvH5xicVxbSXT+Mhut40oOxbmwLoRuqBhDeHtauCwGlZP8cX+dZeMZe3uZzJsKus
cAp6pAaXLHTMpTfyEEckGRYeKp8ZZSvvZWFhIe9SVoYsJPlpPxxlx0YfdSQfCFlY
cUrN7pgTTJQ4oZIpRj/CEWbdipq5w3A5xCF/iSe3GdpVTY8g7OWqOFSLXLVM2Jbo
TKbWsL8keBio8sks1amS36tgQZJAFzwnTlxhXyj1hRF8EmySeGjpph+OKItOcbAd
f/Lis5c7UGSZ08rRXEVbTLymgAuCeEpBIQQEeyXukV4shEjgIw/2I4K8K83RZXqt
F2ejXaTbF6dnw0utRgRu/OfKzoWrDb5cDKMoCkdS8LJ90Y7NecM2rlHPJze0NghO
w8983Oj2EQFNOgj383In+TUCdMwFs4eokvJZzMAumN58n491+E5B+RXMrTggYMrl
5lAe3OjiKJ1Om6UJubpB4mL3wh9BuLEuV8+rpS0uyyJSsaYYx2dEYOqSVzqRjTlo
x6NWgppaqnTOWAqVXapoSfmXMstOtElxh1j3IRsBKXulwB15+woMi8dGp6v1JBgG
4vIPJWpgfXZGtVUdNnGEHcedzDeqbvT4Zumunob46QMkIKmdahvWuraYni1eoPO6
fbfThXKffZuG7Ayt+dbUheNgjkPiouhXOiQCaE5Wiv1slNefEEeGyJcAqAYdtOjf
AaRI+xs2MagsVg7iSxU/CJszcWZ3r8d8nVmXsQ8k0VXUkPoLBPDrot3uJ5B/QJY7
Zq4OIEkRtyagjvOh46Lnq9tbPAwwSR/2xR1/Yr242tdEhyPFwMxS4QkjKdX0sbN7
U8V1H+f010Rft7eEY5JIG70oFKfAXa4/Xxbi30H4CoGy4XlRbQEHn6zgPzLhx66h
r3+NQSJwlb6EBSUwfFA+5VLYpgHrFKx7SOw3N+1R4PFSl+egp91KIELzOTf6MtAi
NCiqU+H9ITecTI8gloZhV75DLxPh9BGjZ4Db/Z8axcKk+SaQFJtACs+dW59zyvl7
xMuii+yZWAgExFpr1r/ICcaxBEFQAFj3MOB0LYaSvEHa61TR0x8Ik/k5nXnJRCTL
NuFbPN83wm293l3p3dmvWhFRphJQwt2G9n3CCtdKAlqVUGUR6i2ZJxXAwL1ZSW4Y
8+ivMhgEP/eooajTC3F29wa+a90i95nmXPnauz2KwD8DCHHFLjHBhgLbY8FYI8Bo
yT3Ym2og7WSFRHsRBgk0GoePVY9x5WMpyX6LLfAvdp22PRLrcv3Xdd13fQy5dNB4
8y7zGnx5MUlG/Za9SpFliRE4lFbhz6SrJ8m9pHESuEK24CEtnfEWOf/6EG55cat8
U6YiR48QQAPL4h+elkfZQNl/rwSHng/ka6RxHJK91re19DSR27clxpQx+AuGodYO
Jz5gDdWyNQAlc2UB3tumF8VuJIOV2f4hi+Pcj0m5ey1lEaQ7skBZYDKo9BuqZ6ZH
xXlLaFbJ7fIp5HCFXMPRYKknzcuh//WQkXaSDpeKL66Wegn9buzxp7I8px7MwBdh
LgcL5AMTIPd3SOhJWJwbg9LyUq5Oj+V2mmszg/zX2ghQFN+843FZN333rtG1Lw6t
oncCXpn5cdPLQdfq5ikAV07E8nhQHpIoWc54wNlRgrELbslTbKGaBRzHTxYZrhsb
KhM/+5SaI0gPujtTEgSEcJ0y/uNYNlRQmiQfJN5rJWgHX+ViU4G+MwFRl4VRblaj
yp/Xh3Z7UatM+vg0IyXP5gUGcZ3eVEQA36VNMCuOkxA6EcFgnLTnI/2zyfs5eJOx
set87BNYB5k2uzVEs9a8f60MQu5rpv2faBQIaHlioIBvqMvo47fvB502dWIjfvfk
165jK++1v7kATVYVLwk+EZOSsZBG3v2A6YGRmeX/aoy/JHDtl7WN3XIXAkxCdv6S
lGLp44JNqBAJ75PgXxzcuX64RbLqeZ91i2Cefws9zV1pNczAnZ+Mqqk9hPtars1H
VxZFvlju0LdZUq1H3jlrGOfvJExc8bufJHsNLYK+/lWyqcbu4RT5ETU91+QZ+5qb
8/7dfixuCvmL9L/o16GMIXcCwhqMA2q5hMt8lSbzRQqM8GfiqApBKQDgQiepcYtU
N20RBVJkXftAxOrwdHBiGYJPPQwfcmzmVVqVWaW0/BxY2dqHQwcZdEKXt3ZYm2KY
lmQUDRgyYjBeta/c6sT5RC3W7uwy5w0LLjyYniQy7gyf+X7PdEx45sCJuITGQaAG
B6dpCEGV9A7ckhxz9VnG46PmnSigQNBrn4vt715LFVz78tOlIIwZKYokQ3pZ88z4
4dHrLNb62OfgD3mXcynd4ruO7X1WiuSp8ZjEcMq0Bc47Ogr4jZ52Cuh+KEXh+XZT
yP7gOxvWzX63bHnwM091OXgZ1zyQs60LZof5+FxsGK+bTDZqr+n3/MIfKLbrY8SP
7K5smV8cuW7B7TG1ZH3fewS4V+s0PRnwWO9pHqnyuwzUUGOlzomC6pAwibFrn70G
E7oQb9w4Kc8xoJy4byXutVhAvErKPXsDlT4gB3Zj25zBAXRKSelFrN2ZY4KdfFHb
nygXTk7c7JnmlELkGf5slU/hP4kRwMsOdVhQUUmvviLqmGiQt4gxpvYRNR8H6+Ql
kLCWM0+uNfJfjCGVqOU6fvhqOCKt+nO8lgBAY1OOY1+IkSWL5LwKAdb9k8NjBuDJ
9rQlbfzekG4s3AZl3CaIL6ouFv6uJx5F36wgfPR1AoemNPncXG/TpI2htzrbzY1l
2QP4YkJ9L5AonQI9zyHCM/3dN468GeKDnJjHR9CT/PdoRYTZXRAjKytUIvRW8J8u
w1BLvNm99YHCneKGK2NBbhbggBSGCASLATA5cJXJiwWXAwum+aLYtP5p6AbiRjls
Z7g/OGEnqwSe52sITArARos3mUEeS1yZAa+/rLa3N1B8ZUIe2LJrLyM0rzdXqCXG
gnVRKNibbPyyLj1dLPbVTfBCZVgPWpXHDKCKDRDKsKysH3qhzHLoyNlJvEaaP6B5
8waui7diyREGohU91dtcvc3c6bdE1qyinUVxsAG+oIXvFCCQuH/JckVEmh5hkRBf
lwzBZdAqgGCvnRs+BS1BBfKhNaMSwJFxJtHtZGZWwOKe0yfw6PU0PshfPPMyWQzP
scEF6RFK8pbAcXN3rUpSxD2AhrcsQc5Eb0k/kle4DmJb7WCGbCG2evxI7dH634LQ
hfjxpQdkdZ8ceIAq+obQu9eTr3ONGo3WsB3MrFkvBGwHBMg0/1qzFzpI5JrfWrRg
9AKWeaIdciy+3/uUjIiH2W67f6GlJs+gq+Efa762DpcQK5/JYsPw5BHjOnPlrZ4I
EAIU7or1cWtQVc02xF0GXqq2YFQj1cO/ykzOFeVBoep9wCF8exN2MmiKF0mTY9ca
MUeXI2LKNFhIxhJiwlDrTK2RaWfeCXhcmrfBQjXrL8n2B8pDg+Mw1OK9vqOw2dx6
jRfa/mf7UvlTNcXY3cARcsYlnv88g+wRfQsONvzrRa7qnbxdmoq8BHu2nX+YavRS
WSJw4NDW23xM0HMZAl4hzuSfrAwLLkO64Q1dO1ce73OQM6QDbLQ9rER1t6Z7nlMR
KdcmTZfp2PIlsPna4/73bJv3v10IGjvX3wmFQEXDJydN8UlCbT0iYELxJzzMPEyw
Yb8btm/58x5HHoygiHPlhY6Uyb6A/anLe1+Zqq3WodVC/qmzAzZeuOn1qxlm+0Aa
YtFGqCLnQt8jGKB39zzjbXAQ/00YV5Nc0CgsgB43KaDfu3Z/WBy0diDDkfzGDrSF
zxiee2CysEDslj8yIraT3RvgKMMQ8YFq4VLI9txO1TndViod5SMC8AXNwL/7FuQK
Cf3g2p44/ZQgCfXa0ZSGS8HhnOv8BxURrFCxLxPgRBfiew2kdas8wsoPpGxvUFeh
0w2i5FgLD5qsDhLQoev1ed295ZIav2tmGjgykMTfrMHPhn/7nbLkXOl1RzA8AD+C
9aWEY0WrRRvOevF9kM/oRsh9qLWM0aO5I4OwGq4qVJnsxAxJXtTcY4Le5tnglGQZ
fQMlm/X7vYQ1jZ9n2KDjimfcl2bcW920ncavV/++Y1V9PTUrOfQKvvt1rZYpi5C/
gjQYTb8Q/kL4eHKdKIxYk7jVeKXLOLtqQZaEFpQHN50pgOxPjwEFAUGKN8kXsNZD
kffdYy0EFmo7NR0/9dvWncDB0fR36nPyauvLKjmdxUANNtH8kL8ifNgA9oYXXA+Z
ajRrcFuFUyWMY7hTdBlHBGg/cUZH4l34I/zFcm8DTjK8QfSGJ2N9iPIHyuTa08Jy
+abjyYe+SPSZcFYFitslWscGwdZxl54rmWWqfm28thpFdEx1/sfnpZqipaJ+Ihcu
Tphf6C34kV0m6OFEu6kzZMVnlvbv2SM6AojI08KbzQicTGPMDiq77fI/gVloQW6c
6kVPB2b5oG6M1pntnR131nKA+OoINuvwLPrTCQHF3tb2H4Hv7flGApVrJ/kfjGjn
1S3LVpjCPCDdcmQ7NiZbk9nrd6dWcKZrosEctbHUGchpHxz2L25g0L7+g9EYHctv
9CswtA6zmunyu/WkMKpERD3Q3Pg9rlEq4iq6ErADjNx+uwY7lha3H97mDXX0a4HG
tjM1XKeWBFQYcPGWVmUZ5qznPFNcoq1qrAi3eTuWl1qSI1JY2EnrvwxbNxhb1SXK
89FrYR5ds/Zeoioa8eoQvigUeiEfDFbginUg/B5ymqu7cv4t/A8gQ/6Uj/fo+EnZ
ASeA4xHPXv0wAbpqHvqpSWCep6zoOZIPTkIUohAV2ebzEtzMjvBd/xJ9J3JXMGQl
vbGuARG6qHnaPH6ZDTwOZlvkEwcxnooV2G0tA3Cjckwufyy6rlApAuUhO7JEOGHE
m+wdHzA4tKrouQjgOwRhFx3zS0Wuju94LIAAaHkTqQGL5DqR4vjwGT1ijhEkJnWb
mA1sCnxZbeSHB6fPYPyY9Q==
`pragma protect end_protected
