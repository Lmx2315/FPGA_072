// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:36:58 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
OTYlOth7yQaPe6IxU08tdCYxD8UxiYuboncPckbXcXHb0UXMSklIZLGY4Fz1koJB
izZI/NVQJaLwwIWbHNsbrV5qANGkg/yRyzzJgrTOIJNvMN1Ln33P7Gl6fZb/3f9g
utne3EPp5oy9axAC33arXfoTdwme3DHZv4wflV0r0Zc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 20976)
aCDjBDAgamX1DgJHNa6Pk5J+VBY/aDZfeLtmVvURD5GQuUQwYtghJDZ8Hc98S1OG
cJb7w+EkNzOkjZAy+vLy7XZOiGYLrWECyxMMZxbwpgAjmSb6scJf3mozAIjJqDO9
XPEdTYncFzZxgeCNftudmbyDN3wn+KR9wvPrhrT+WlbzDDaJnZlEq9utS7RAvpjD
NOmGcxrl+lgWI/XovwlzhcfiQtbq1OX1yfVfhZm0HyA0350ogeKvzKiLSGHZoRv5
+IsTo/+lU3Xd6WZUkMf54d6rfhtKFWDdVaKn5jrHn+BFwFXG8QTLD5tOGlK0euhM
r0H6lGebyV/ZejL0IGgY/VeT0OGYnA5sdEnMA4dhL0Z6s/StPDhjmvf5jrX0t4E8
WSnPptLDDAvdtP2w70RtwgursCba3KO7cXRK5hFDcETVgYxtMUNpEgT/m9uaK/2a
JH07kFc5GXMPo+3+7scJEaxY5c8uiywUfK03K15Xb5A0uJSKd5Lud4w68ORfv/7e
60YYyMPS2perE6PM5wpcnL9YKub3EMyKXjpGzzf9nTN+xw0SQjaKWnjF0k4HE8rh
awj7vGZfgg5ILH78pyHk5wiejYa/uFBuzFCyW/bPSIU/WFfKiwluEpfbUirgncdV
zIV6/R0v50Aga+khmTOx8UTyBaGf65YntakSwYTqz9HD8ewN2tBBGXcZat2LaAhJ
Cvai03JD4oWzWSnk3QA8FTAkTdvdnctTqqYwCV1ErgDWiSD26gm58a1ftpiLyo0N
LOHGLoN7zCbVIi+ZkxU71fWWwkHQ/olRGKWTevwI705OrelvjqciB0PaCbKUEeTz
ULz98cBGlbFbDO5gyIlxoGAnURZCkVjaQTXZwdmwhC8NgtDhvOpBIafJm2rONEhp
fNYwhufkwbK1W6OrfduuBv4yoGCs2adzYfcDFFacu3hUhj3KZjY3TNcKkI4NHbcy
SnjDP4jYW0C2s8dqOOuiGViRSDFodd3LDcrMCZETE3pBFHlkwDSKv3MLTf4iLw6X
xj0Nc+uflDLxRD9bagkHjAHcceAOMrJcq5ywkspgQqEYQFVB35hGLdyDXwBNHvc/
7My7N02MFbIJ/ii9kEzpNpYOW1SMFvvK+VG708EDFZQ9vbjK1HPYn2AoHWh6gf8J
W1KTnWESKgS3VLGq/pbaTTsBvorYzeHJ9tYz9DpZ3Xn5VG7tlYKnnNisVHJrcRhD
jsG/7tRwEcshXBEjCgwtgVZ2JB1ifV04sZ36UrQIf6HSot6nhVOoslltQLSbnryJ
gsnYHz9P81C6R5jQIyMuGQZ7Ltve/BkfMGefJ2tHILqKLcsHJDCepfPiNzd+KDM9
ehFxYnorceA8ItDHgQAUejwkHTAQ7xgtuW70n6vejkEOQQJHr238+xIC8myVF88p
eseYa7bqE6dtHhF1OxnLf+cAfFbTQ1EQEKAMgXz8WW37A8gMpleNCjzUTSh3aZvZ
RB67EPvBtCvkccrrDwBETDDW8l8Zv1Q5YlfysmCC/shwIMIIKziswQrwGulOdaa3
Uyx5OyVJ3P5NUSYgZELqm8vitJBD8ZeH9pD/PzKQx8dU3ZYFTNp/BZuY6ZevCkVh
AVKO1lquTi6NvOgcXHkxD7mOH3gYrLUgB4oinKgBFfbqtX7O+dxCx4UINE6KkVyr
v9Ihu6Vm/LUERD3oPcVXmLmscB0FHM1dfHr6wNhroPP/393aqMzwGFXn+uReJO/M
KAEPH48Hz3wjnWxf9i04iXNVtJlhg2gupLNRNGhqghcMDM/n2RZGhpMFpqfw3mi9
eABdF9QD+dAPOQzDdtoGj+iNHfSq/n7r9SxyfVaXGMMCh5Nom3iOTLhHJ+/T/3fg
1f6W9w/9t6ZH+ZmwUQPELM9rTNkvisIJ55HTL9vuhyveL3W4wCnHi2ZZW1NOYMOZ
cuYIbzgofNTrLZgxNFoyAkc59Bg+zxyUE/tj2jehgIG7l3DLFkIlGVOJEqEAOMdZ
4IThUovKYoN3Yj51yTEkBcRKP5NNnwJfMCkR7Twz7rbLxik3a1okBiZDtybzMh69
XVKlCejTvIt9+lMI2O/wxis+/4d0yr2o4sg3xqHuKsAT0mk+0IBH35ErCXiPkzHS
apak5cSUPvhm7FcQi+Vzs2sQfdu/0M7lWFFDEGKJq26dBz6DBlmlOCowVeUbfQzX
fM7igVxrZFw0a50B7qBVSWHJ2+RyuekMiX6Ws5R/hQ1buX4gUFaSdfYPY7QAg+Dz
T62LbZqJTiTbAxq7omxVIaG6XOGG8EH3mbCrENyLpOQnyfG9JlR5voY80K0S5Gy6
h8p3+RR4CfsBMc0yAttLpNw1C+IHfJ2FRE49smBUvsGAh65EkHTwP5LE6XwD1QYW
ToDXeit0uWlyYhw3Y3FmF1S2k83ZE3nTaDQgSoBFT0XSBuhNjG+kTL/HuP2It/0W
EaWjahPYgkGciM5p12Y+WGz29V6YcDxQHTodpiE4GEZRNQPLtDV7Kl6kV6+D+FQF
ywX1t0dubsIRgv5kair/vBQd/6j3OMIHWdspaWJwtUwJYR20LCXO2HM2TToIWlBg
nfNk76P4xUoBjUBu5t9M+LpxWulR5d/r4OHuAp8icoxgqv60CwZRuKublTTB1EyE
or4dxklzjW1NW6kQGsg07wUdZ8ruwIpfFQIJZ+73lqxp3mq+UmRvIt+xWET6uPzT
EG6qkjTUgsP7kOkYgv7W+VB8WIa/b7IOwvoWmlx2URFt9c61XYwVOKEPYm1Hnr7b
mEwWmCkj99dTnFus403TvxZceeD6T5HbyAzUobW0/y36h6y1dVPcdkJXf3ZGBA6a
IvUlTYTOEY9Ye3lo7u5i188zdwDl68vcVipkjqayryG4VodXafQtr/DLx5Unnt87
W+PL+bAjwXBef+t88n/E5JrDLASYbZfxUeIDzhozx4BHUM4AA1F7XTjdWn5WjOTN
LD08V/JYojm1DpUabe/riCppj6DBBft6+O00O93gfVhG9DH/BK90EFtaONZSmhVy
ozOAuSAxuYd0akmvhGUoOwBgeintTZNMBOqJlPvSOzCP5YcFAUcUcESPN5AUPQX7
yr/Iw1mCbNTiFT/hcNxxERP6JEtdnfHyxIrOR+M1/OJSfAyG2DVwN+W0c0gKE0/y
xjCVS7lSlY92/rNyFUu7KxLruu5ip8wcWYTps9GzYI40ZTejDuim14DN7cUsqLJE
mFiS8E7sqWBJZRK4gvU5nqSclY67NBhZFfOjSw8395LlI4jU16kNcUqn6kJkjZW5
T/Wjc+fsTmonCBExgVoJRSQ4uCJCcmwDFQGjlV/LgKH3dAvQAZP4WOr0y6gqDCTU
hrWEd6O9LHaXw5fxcMruhuwuvDqPkPOa6EtDiPjDfHeO+ciyOeH7VHsz2RmqzqwB
3pPKjELsaeGx5WWQdA91Qf90ZPZAxT4JhOTurrBXnLYWA0kMQ5qCxSUH6u6uJKz5
ypkoAOHxZE5ZFaqn3OS/AJume0dw+5aC3onpagzY8rEK3abbK+gvgLv7fG229M8q
YqK2l+FBQPbMkJoaeQDxlv/4MwE1XpFCpOJo0XS1HczvrSfp63l+P/o/aOldwEV1
XYFMLDCAqHZkUsvgh24+aAYaMWrQPSOBKUr9ft0pEffX0MI5wbih7caSAxbUSwD9
FIwFiACAVrSvnEYYldS2NhttTzo6ZVlM11e+WD58D6+CFDcLCo72pvSn8leOeP9S
9gkS8DYjpMcD84ACTcrWl62ouXVNBlLjvzxtciZmSHA1kUBcs1TyiFUA/2TgJSqo
clU0OXg/taFgSFKzppjdl2FLkk4ozFwXfYeqy5R47YRKXAheHNKjC8q0cYdqamCV
y2CC+BGe5mLdGePh8rTYe1tNLyvAym0/B3qRmGPx039La9wjRQfYi2rEAnKvQEh5
+V5mw7Vvdg7yTRgqzDuhKrubFvjDIywpprANbl1cZH4M9BmyHdaGyXlLaOBBPdjB
Dds7YlFNXnUXSFPluzeJ1hr4JCNTpXSaveN7gtXlMYVwPmJLXA6+RzdKLx9XgImQ
JUpQYyPspkqEByMmxnDrmkfdlJ9GUP+pscCN7xo8YB8EPGm8JnjPNoNHtTszv1H2
RlwuB3BesraQbq2iAKrVroC2qShSr9OgOsxphCS3tI4+DqJR1Biova0ydxMEw4pe
RxehE4Z2jLc+I1jkMRosnO+ra3UHFHsevcHEv4J3G2rDib9ahUHQCvHF1ED1bred
gRRY9YfHqkCciOW4PYkvOvaxl3+Rz5kNrvABmWugPtuvjlxcjwGzcy5oKqUkqx7i
zmnoHd63rPLZAcTAVtmJq8KdOBLWTJFBlTz97ufow1Mqk+9HafRynLDRTMWG1+HZ
3hAP4X9FsBakg77j8ULSjh/X6ncUvk/vOhW2nhZT0kQhL/FhUHQi8vgjKRQa8Mw/
Ee8A4jQFzqLI+dFa7lvcDWnTTd6k0zVwu5I3REUgkyrXV03HBT2UruIeubvqK0ty
xIGnNn6raTwhnSzAw9muyyh/55HdeSvSP5dA3qXS4vWV0BuzTvCZbszs6PJrylUJ
uabtAUkvuHIfwixSy/a22SbVIBw3EE2ur+HuTpx6DbvpkbhHV1ur/lI+FRAcwIjd
AdnbZueEjIaKq9jFwbfANuq7oi1AwYnZkXVEhdbHu7Oglp7L4hJtySEN6VSTk8FG
/W2hmJ1KELx4p//Cnk3Evyp9YL1T9QMGTuLdQQ/9jpQYjbGDSYI7IXJu7ose4n9Y
EA0wp/i6qptpHFuizD9igBVBhI+5lYQPHehmgO/PUu63NUzNMI23oh3bz7G8YK64
xjn4yyONh5W6ZpXny77Jyb2ZnFI+Uxspohg1L3YErKIhkoejhJoTPj3Lr5Y1ygZB
rBnZFzltLVwKz7dmuLDox0ZeT0P/Tybu3p0rJuMainDGAj2OmucXePQvALqjFjbn
zBOAStQy6sc8ckqBlmdRv++ZFOfbNHeUnV4HVM9VSKqH4vvJLxJQtsWtQJUemuzP
gPbzJpWWVwgdyOl7qQHrTnmXFR0HDP2uP//kWyEPbZ6ejLRVTa7yQiZU2LNgTgG/
JP1tfQ+C+95waUQ+phbYvXAJmysjPtjmI99qi1UIvW0hE2sp+NbAPmwG4Xu2Z4i+
vD5OL648a+zCTWksLIMglGBHg0abtNLNA5Lu2KhBYU79N8Hp37gbHzlNrXzvhL8A
85v8+aQl1uY8fkKB+qTtq0HzgITXFdiAWuMqSVssOE2qJdybrCqStnO7C2TvbqgA
geJ93uEMohX3FKSnt1Gpoghq8dnHpgofMcIWS9Gm4N2RQAHIiIwx2ea2RMTE1jN4
Q56vRlwBde24VoaxtJBLKSEMQl3Su64H+StUB70yYB5/GwznSLHTzMFo+WOwKMe7
DnFyz1sLT8c4h2avuz1Hx2tAwMA4wNp4bUVqg8XfjX7d1eVqL3ygEjLc/XP9BzQ3
f9gGAImHir6TeKX0e3Vq73GwGbeNfCQX/tc52bUX9V2pWCV6UW03no2cYiud3a2a
4LelUb/zBqKNGJpjVi0HITAbFIiiyBM/xfjTg3MIOHV+QTHFt2t2E7nKADbpmFCh
q9cJp8HZc3tc49kZt5k9YVu+4wooDoT5Y/rsFPpWXND32NdZ6DT4sncecuQ5o9e3
+lZ3uNjcv/mN/CF7jzQXjEf2NdA6n5gA+hPaykdWklt42k6feWXhJAe3xJ7ofJ0D
vf2KvzNagLcpYUVSoY/S7qombPtrDQ27af9Yq4+q7PIdzOnKgYQYkgDEMkjo93bR
qdWs7nrALoKPbr7QJsKk1LJg4xe64vBDGZHGodGR0H6iQWBuj/F93jrf/JPqILMp
kyIpPxZ/MdE+1YSwWtO4FHk3xKaRnSCOBLM1N6wNQwVJGIp9cit95N0prsx/a2y+
zKJEwPigvXoqq6OT+sPmc3larLoIii8Z01/LrcZdNw96UsntGsZYPOirmmkVQq5V
HC3JgTaVSg4fyHndDKYiQpY063WSGoi19qUg9gCjsHFIFFAUbQRb30L1kW6mkyA0
CX+YQtBKHhjW6LMC+JlLo3kKeVidTTRdp4H9oO4NL5pChKAQ4t3nAppTwSkx94C5
hh4Gqg54Y3NGA3+4eK79e+7Wk+ItEi8ui7tg4MqZufj+dCAR+7FQpqDVOUDvquGa
+gg/oBRr60+A0TVwuTgx3SroEOg/8sNBGb5I8Iidym36d3z3I3hMrM1w7SmnOGQs
tVy+9xeu7gU5A049wnR2vGNeyPrxplx+voIXNyR9eikd+YeYRfyk14Bf/A52a1Ng
M1E4Lyv7U5f4WcSU0KDpKlR3BSJCHkSio8WrJRAuTyAdoL/h/pdiA9KkG1zWTrIl
pU4bcpOXXyXxUm8Rpxtv6x/5hMO1qJNIb3jBe9Bpt9HivpjIyvbjKOaI8blZMpNo
4s9mc9z2Uar+8yYR9yOB32uECuZTsDJTN+7ckOiYxeP5KxPghd8KCcJnslEpOVAQ
aXYqq5yyfyrBzPta0J1MCMJeKqdcOCzZNqylZMoGSKL7y3eL2qDTod1bz70OQxMA
Ys7lwt/Ha7J2iZb9n+8jZBByvDVQnOoEAsmhVMsCHrMNM62qcBvWKL1qOM7mJo34
Kv73JcviH2E1RET8ZOwGXd2FwKLT9pjd8slqOEYb/twYXhKEiX+NSyFUZUnI2ADC
XiVn5qlDZADyet7awbwamqfzrk7aYBJm8U57owVgLcPC0RcNcKMoF8cMvWq284bP
8OXLQYJyVVnk0PURQmuElrcsy09yyDSvw6xXSm4S81yUXOt1XGr5I5SUmTaOYL2Q
JBUeY0vF/zHO5EER7OEQPxGqL9x+sz5hGIPlQkyfgQCM+1biVFnq1bXwU7r2nkPS
Lshj7MydyNPVfi3Sz6AF4EASlDyr1PZN6luMpMcIAfZZWnMvVg7igbiRLa5yWToy
Vgyav+/j6r6EM2tz9D8jhXE8QWnjgO4MEMJ3pi7MGz3/IneUNT7aZ6Cr0kj0Ygyz
SMgyxmTzICaBcLD4nGPfBR/m8IIwD6emNwe1IbXWKfmN1dhCSl3oe6qm3WMFXjfv
Vh2l+vKxmZNUGdwm1OOtw88+C9EthAhckeMHEcHu0ESyTHFdcbcSeVurw0ZGchfI
3q1e6UJECfQW3nBaNhhwyquF1k2f+dQJazoYdkm4eDysHdW0eDHHWttNZ51ArmLO
iMUuNtYHnkft/xwxgLyEgU6yapZF2Qw0HmRV5cWOq+6MLj6RQN6AkMiip4y4q2Pa
UK5H46yn8i6nofQg+Gblrwqmj1e2iOGOvubLZwqa5O+7gMdJQdz0fd+ta4AVyQYL
6GYHFAgebIoVndkcXOIurNwUJ/VYCdTk/j9a7qETYyVfZ1BdwCBjf40ePTLb0n1N
8x84/PpN5WiU1Fmg+s5ghb0kynRuVKoMkrlruauhUBX6HWG50OlKXGDYq36rMuhV
ya4Uda1MzSyik5u6ReA6f7PI7HecB+/00KV+LkeFrUNXPqx79YsLWq76XyUWQ0um
x/z+i4sm6Xbk/8zg1P0FqDSky2btpq3q8q1nDOS3Bnf/YZo0Sg87v1r7FdUvWmef
1/NAjqEZRryfOOxlQLBqnHaGYRGjWac5zI5eNWbEdocf/nXQbYtLxpxHNqW1MHQs
HL4exp/ZRoDUsFkH2SSjEEhegduK0cOtYH0bcgNZL24EwTG23nhlec4Z4jArsgff
np219wLnsYsw5L6eTwNx1GkrifwsRvSFtiGpGoh4sXleFgryzcYoB5m65gzyIoc5
HPVvhcGSZYsjf0H/ilhgMoLarzpMKUEBjfefWtFRvw//wWZmOetCHzcKe057IoLo
0V0O9bfQwzrVDVQrEp+L5KtASZBpp0/QqRhPbx5uv/TlcqEq3nydZysWKU7g9oI3
K74ye4UcKHtVkR7L7fFCq/9S9wwAEf1PKD8MQayCyVrHAJUZ1QCDgsDCh6idKYMr
BzZY9chheIlXO+wCeiE5hHmVEQ9Yr6go4+AvUWGvGStq0viepDRxX4avFD8PwHHy
o0ejcCFijC+mEL3I/aa+0sYfhN33RLyLJwNv2nuT2i5GD2pSEkvyVbGyfI6Zp8rB
/C8EM2XgkFFtB+5OjNNBR57CU65GXbn2cipKbsiEyL33uTSoMlA/WPs7Vxl+VKKi
gSVNUYiFwg6Kw4NnWwJeeBbkzZKCpXeSfqq1FWKpDWXCvANceMR9auhQdLV7V2LZ
hxYTz3dH0VXbVDkPrmOOK4h2XO0qCx9iBfQQuuHWoMbQtw3bJE7/jyhQDO9x0Yla
GtIMYio7AIdRlH7mSp/floDKtxJJGCJf2+yo6zVzhmxKUceMGdW6eQvEDocfNTpD
tyMBRiQ/KITzpq/iLbvEo9Qh/xgM4UwQi6pH7P7MMb5Ji0yDi9/aVV289XrNkIdy
47kdcHiQI6Li1XKb0N9uUaVDEcC6Mt0H9uGddn356AVZtAN7zlVeRE79kbT1jghn
LJNKBE3cTtB/GAxgpcgejsqOvlaCB9iwWxylXpVw7FW3JlOK0YokF8IxmmF2RJ7Q
aQdV30af8NzPKkYpbWsy84KV91vdffPhahS1IJcyk+DKFupgky2YciCQRavyLPrT
22cp+LKJoP9NFh8d3t/YEhfcSiSS67eCvYwfeNovdxqXWhSanTHTX7BuP9VRDzPc
wIsBkP7Yc3JHkXm4vmG/cYkjeSSjY8TFyb/6tO3hdWijAqa9ssQsUE9drBEGuJCB
fxt9weEynsXXNpgPgO1g3EeLHUYsugnwsKwtGFrv7RVmya8byw4vzoUG7Kt+eCD8
Iej/C1XMcuFtTpxPOQQEIn+5XS2OrCj9/4oEYYQsqURMtgAgt7ZsKIPy1x1CdfhC
6SqqvrNWXlS80JpVLB+6i/M+oyQrDfIFt4nXtTd42BbzdACnbBDa72up9/knzeyN
gjo5JfsKKgztcAWaiC2+IBhb4SZUACzQ6HvIhR8daLVU1NQuvoFLCUk1vMbae1TE
bL9L9D04J3IxcwNMKGc2W0HBtsLYKOlafi50ymdbq1+EcMFmM8bbPinnh91/33BB
uEWZkWAzjAsSc4yZWHCnbMU6onjSkMyJeoYtpV+BH3jlVESvhFot3bObkRCLh8wQ
bXUM8zM4Jvy+QABmp2WeCbYFaC8X/foFAT7q6euovKL6fy1TOkhe0mAAv8irJBgT
s/VjGDk3xwpxogqNym8FLthyWkXUcDMiawM2GBH/1pvhIK7grt1tlzbdiQG8tDc9
Kjwx7UIh7O9gbrezepMocjTd/4FEEtWAFY6T31uMgwzTa5m2vsZYfzgsQwGK0sIW
UVLBNDbhXWX/uryZQGZsQorEZSWNa8zjAwrYvyTKNsAWH41sHvATKGuhODfUZk5p
MXjksYO7vnnlVPKzTSTfuCX8Mgf6ExgABfL3RvHdbxHBJH8BP0ottcqJYNBSp9oK
LaXAQaIfPvUXiirIsNrh73/2auuAI7a2hPgyjvF6oOvJ7NMjcnetE036ALHrH/h6
LOgHxLbuMUJCi7L1+yN2cl+iFAETMXGPA2f2wEQCd7g22PfB3uSp/NvsHHFn1AaB
3QVwu+WRx9ZWp/nJGoABwwPA0pJMff1MPijUiXDTZ4tMBzZJgVW6meVlNF1NTcKV
pvTWreTTgL5SpoQvHty2SdSQ157JlWCohtMQFpinvUtg2cKrA/Qx2e9m8mWRUcc3
k+rvnsj4yNKWZxJ7c5dF5bTrjiaecQ66OmixLb7/DRsmWpLzaDKaFunUtozp1gLA
E2Tl/lwN+z9ILf6pqBlupp3ysmCFBqwxSVfsXepSbY9qpJbY44TxfsXMlI5DB/Ct
EtUFXdSQdW3LA8rSW/qRTPBQqWpqBeF4nV81TOs0OuBMeeHAzu0fGWFYlU1SzrQA
vrnsu0aq/aqSZThV5WN6OZJcDPkk827WNDfI+RtY80JDtwNSaukAOrLIySF0nnBH
umqdNz9vwPCnrcZhnrflCxNr+ZPCOijjR87Pv3fdaDBdN5siOCTScQi/fwkRxNhi
ZazpRO9LRox3OhcnzfxRYEaI8AwkLJkD5kpM7l2JD+TMzgRa39KOSjW6xDbfY9wG
hvw3TT5l+UUSHMRX68hQyMJ9S9zra85xp0JBuHq8u+3J6mrhKtk1BAxsdXsJ0TK7
WyXqwhO2DPgzfBqy2d5i0t5tQHMPJEhET2e5mmBl3dAnbDi35IZ/sTkiShrI2f0M
K7JQ0C7OgOUAyxMb78yriafxWIEvDvQGVhC88yiQwrXUQebWd/e7WmU4fWhJWFYi
Xrpj3oCYXJhbeH5w+YyAg4e5S0rWq66+AT4V0H/wbpMrIuUBTgYJIKd2n/0n7+tp
ynWMNz7sBik8fWGYJat9XgyzRI9FfT52ixs0D601EYSITny4AiXcZfDGdLQjV5vE
Og6jZ/kIQIwc4ZnXSOVWZeRi0fHh5CorqFUXiZq6AL//wbCWNTecVmo+r7AXjRjY
/4wdWlytpN8mkhM13kW4a7d9EehrTV+ypqsKboDFJiEA1JMlebNjzvYxT3EhNVaS
NK7XED3GyvK9N3+yP9W3LlqRhUKBuhBaUukrRcYCh+I3CccgFqvVsXJIEBA04ZNM
0e/uRn4BTWFRHK3PxGOlAZBNjmcoUkK3WNWGFSyc1gizxB86Jlnb9bk9m5AgONyd
vVqSJxEovljZyVkxFR5dlYmWHZtvzltoCc3OalnQ9GHtEe0v49bse9F2CU35K4p/
ODFy213kjzIFTiFxbHaBHtukK4D1OQfo7bzcG6VAnowaQwHguv+egu0M6Qzz7g7b
Eaf0Lvd3WTamkmDBcCIIX8Fx7WHbfhcyxF0AGpX4Pomubik7HvDf90SjhNsCONGF
TrvnTEQFmiIip8bOG6nR6nJYD8Ktw7OSh+xTZnzxh5ep9wLnIVHx+vkKDLTfwX/c
zJdw0PwxF8i298BG42Qlg48UiF+dPNrazSguUibWmIVvfl/yjHWY8JU6qW9+kOFT
K/XWH286HOGsTku9THnI8sF2Oztl4f8xY5cs7lRpfEGiVKhF+FIpiKtPGpe68Vov
DbEByBKvAuIH/1SPgufAkLPD32npR9neWk26KitXGpWkRom1USj4Up59hxx7fuGp
9ZdLsUppOWyT6RFrVvOL4KZW2+Py96xvMFunfcGdUAOZZaqAHLlf9/TvyDT353ZE
io0nqvyuSb7htyxuOq2MCPJ9EX690hFQKa7lDbka0RyMfW+uE6Jh0PobqnCcyY3x
ZEALYrakUih2gTSsAVmZ4dP42Zpr6F2/HVwsRY1YQjt3S+l0CQGspS9gDUGU7wo+
+Mhdf6/dB3X3qC0mgO1JZJ9ndw/YxpRANjUMZ6P8v8I2HkK41UNOwMcJEbqCXQ44
pNaULxV3IMoHUceVZY2cJthWUyo9WD73OUL4t/KVQEmOqcqb1yF7ztVQVaT9NnCk
oS3vFr7E+szSBCZ8cNSa+2d0pqD5zrItGwDCXY1+gwcXmIUxCJilUIa7ol0bwRZt
MqBuf2wXaEmeEDpYvAUxwYILkqBDT1i7Mmwzya6TPLc54+1GHh8wuBejS68gBXTw
KNgQ2mdOp/2OGQH5CGwOUVteCaxDO+fwtqhoiqTjAdbsNAi96FpnGgtkn1Ix/f0X
qmEj38+Ft5auSj9MtQxtdlNFbEJAyJplvy70QTLEYEYcUKG0WsBVHVjxoq9wpNJf
NIhYj5oZb0eDxhDUODoeRraUzVz12eFk3YCUb76kqu1YGe8yLAMdmc0Fb8Pxs32f
0pIVIU63UTmpIfvpLDgQyGX8T8g/vn8/ROQEcf60qqU9/IMaSRrdkC8X7fpcm5sc
/k3tFVjLZJPI3Wo4rsrMQTPWxwdUP4DfVwXnsyYxZLDqSKKWIyvWGEl7wHb076bG
ZEnfRs0YlmNMW305Lxllv118/UGLERHG+mgPVWFReqKtRMl5//rPtCkb+YKAQbui
/vWvqqOFGU/8AYikoO7Jcc4JnXwL4FG2sl7YXG07lIXd/C6Bu5kBy/9jtk5Bt18k
+sUvjjYgWtXmQMnCVKTAHIUaoPhliG9C8ZqARQlV58V8W7N/UKAVz6eY1Ibs0GBM
oQ2geFceVY2keHJnYDIH0hvusUY9wvE0mnecrYTs+0VeTme5XWKs186zv0qIj1fS
FvLITVqd35gm/Ht3GQVyRJf2zedmBpUSwY/lyTEL6dLk40/wW1WJKhXUJ5FP79G6
30Vecir6FQi4hXMOeXM6C14PHv+EaOpYW5UYAo3GUchUPN/8YGsfTlhZrvrYLGO0
vSPDBqIjUBhP4Q81A4jrJcB/tPB4ZPOadkWsa+rTp8iXu8smRurE1uMl9DrjkMI/
R1hGXCYd03cXDHY4DhJuJ/O+WMDjuzFGGzHwkjG4qXNbQVrmDgaa2KfRvuS/Y9PX
Aq83c2RZY8RUcKOZwJnp6DaBeccjjKR8PR0i+KaV/wdP2dFvYGW6NQTHznsFYCkG
ruvNeh5EeL2HT1tKoS5AQh4qZ2Fhnvn7GwRmU7MW6+yhzQhlkcGQJ+VQunMfj7L/
ncwZTLoZ0mEqgrWkQr0EhaoMSduqAFv8VEmDgYHhMDgr5SkI/kcXjymvIWTnUJsl
O4uJ8ujKpCXw1o6wP5MXbxyrU1e1OQwh8ploIXUn1BzkzKeuU82EgujCtwwFX5eB
xMKs1UyLO7DIL4zwdmAxjysoMHTTzMTJ/XiLmgF+Nw3G5kx6PV4b2FMxTEnwSIvZ
bvN7EnkyO4Q7etd2rylUsNmY8SQeG151WvtHnMdsN8Sbose4xfK8c7BOVtKGFaa/
RyLYQd76kaQd40pVahdF/pau0+4WJeifdcMfB7Tkf3h5YdWM+gDRnJrKx/XRmwF0
fMqeGfvbQVnd2KLwaP+717kpS7nABXaqT1OAAtLMT/+0TxYdoKijaRbHkP1CCclU
kITbykiUxfE6ot3saSZu6GcAiOSbyWNnrmm75rgAem5++zN5Yv3aTAanVArZ7EHR
VBm5IbfRmPFjP+M7D8vLue+MYcwvkArruDd8+5/Mgm2n9rxD3updoS9jjrLNAAXP
zytd74qJT3KgirjD6jAIh+JGeaij+s29q7gatf196+hYYt2l+FRuhi23c9fdWL2S
U1WQz8i+c/wPtSNRNiZBpQmdVBsg/dPlc1cXWogXj0JRROaiQm3I/oz0hC9U/qmU
vScMZAlrBjhgDeEswxR72+UdwuMZt7tq1p6JaBjZxXHXk/ttK7SQtZg2lLUvVbaZ
Xm0Uyn2mkt9PkMlQER7g2OcSGyKYjJQ/Ravjop2PKSQ66oF5OASemM6J/Qlrj0t/
VWVnZX0ILvorudv8oMe2wn2r80J3IsjCFW4w+3KCEjKnlked1D3f2Zn+unZlYl9z
L1AC0HaMRfE4xjhjP6TVEfc1hvbuVk1qVexdqR8oN8vhXb9etP0dBrsJAjGElxxf
mIaR+OXU5z4HzNdR2YRuJR9eV2QzpYFu3H6tKH2PAm4RLyLArpBPD3Z+ctYb3j4H
nr2zmdNTNPH1wOnPkQc8Q/9PqMdsQllVwx6Qx4BYZHMIEzV54RP9U5Bmm2JB6nAC
iXpEV+5x+3ZutPvTXZtLD9eUAo8mPXSmJk1nwb7VY7OfGe3Y+3CvuQLXIAMFaw44
OvQ+0rj+c89klVUwCVt6jk6RZOuvK4cKv5OwD86SIqrCaSAHOCnAxI9JCsdVgetN
swny/3QmeBmY7AFl5ftXPd/Z/V1x+LNaUfVMGqUEel68F/B4qY7ugSfIo4sgzZzV
gKePJK8KkLEJfNvqtIxLJVQrcDZTnxZSCtobkhBEjzJWhiIhTtKniKW+kNo9WUBQ
zIsIPL5IWDMJdE9Qem1AIbawcQasF5AGzOmGU76LzNmShABQFRbhn5YC5RYLv/wc
Dp9Rp3fH2u3Ee4N1poKxlrBbJXWeYeWIPe2QAmXEIfx0dbVJbebcUxFbsBTWb1cS
1SsfRPraDMBYPn4zvWLdVZZIPQg1DVNX5WdWDB3sS+TWq6u0o5HMctQ/6QfPY/Fk
/HrN4LYUBiStJqwsGJ0o95RVatOMbNVrVCriGwxi4rg3HsLu2RJv+tjj7eT3VFo2
fjAiQ+k/I5iGIQY4a5xHieOl15Cr5eWhNtNIyO9IyKLbTsNIXbN4oFgADQb6RMt2
RdM2DydZeqfkEgxRnQp4PMK1SchnMFWFU4+3xxch3SoSDYbbB9fKk5DyqkFKqMyd
a0tJ3v5MLQhNiJWws3X4BmNJmnDIrTtvx0LZR6QmpKfe+mgeESpzQpq1TH+PnAkc
46ZyA7y3doArPo5q6hbZNJoPPzumlw+Fxdm4CtKfpxD4X73PQRy18hWj3aYWYLgX
/3+L7uPDV8M7LPw6tfO292JzQPVtaWtjAd1B3wVPf/07pdhlLA0Idtb8am61fYYz
OtwnZc1QHLZ9+Gfk0fjXzv4rfb4it5t+gUDw0ZItFhtvj3YQjSj7O6EVfuuFtWWz
Cn7T2n+PzCn35liF2Nlmx9eX/YoJSGtDMJ0FvPEWF2/DM9ShosN1CRb8MNhWs5St
k8ifZ0b5rcppZXYbY7GfNJeXyH2aVg8PhvmpGmdHcErHLpEmMmuI15yCtFe0JMUz
ofeY4Yg4E/nkt0hUru9kBJCh/OyglM2QvslAV2PQCBcvE6IzLAeGHhPelZouqxJP
k8hZ0xyv+Jsn7W1AMC309BnlsJZg6n1va5ujRcL3/iuk/iEfdC5UnNEa0l+JRGb1
7nM3o3rwyq0Qn9eXrNt5RHIwQ/nDR7ZjDUVBY24Jypy/XiEMlbYYc+yFQ9txTp/L
XW4qS4F3zYUIMq8PEr1+cHqbqHTuRc+m7sm3ixgNeq1UUe5ORuxk0LEbvjgqvq76
MRXDfesNNNUMZG+8B0n/7OcgveFPAwOJaKyOw8k15Zv2ESNbk8bbh8D5X1Sm/HFU
3D7i3wuOtF7ztK7FPS/MXx4voDBg6vqzdNPcuTx4J1MCxe/eiP9oIL7WHReXsRLB
mbJFLC/uc0LXWpBeRwxfALmMUch6pogKecq/c/a1hLaYSq9+U6plSOLn8W/0gBpo
8/QiNb+bOcXzXhiUW4suvMIzlJ3ICtSedEJTXpO0VG+x9KYtyeSI0vYgC529puzp
xGF/IaIndFIIDBVSk+DZaG6oeg6M/R8od59KDlk0nx4iQdc2AAuHoI4uEqPFVi64
yngHS3b+9E45zavmzPY4d+GCWGDWCCP353ouKs8t/vKpbRCN8mMGILwyVVwltE7x
soeoK0JiNIW8osNqkWnFYrwGrNJ3ctWHWm7/mlGRkp0QzOW0vFwvL+UTal/EB2w4
TVphz6JowKd6sxteiLm2EWqTGfSrpTKnOMR8cSYr+CK2iDRx0W5kJwCaDkOrQ0h3
ni6w5S50iMta/Psti4ud63CIVR3l2cBhdimLwXtBy0Zi14ajvOZr8uAYP1ANswgn
BjwSx1rYcnncygkESwxpCQf2Wd6mcEkjtRBvq+B/82t6/RXarYlWxPMDr+iQgsay
+hBIhw4BQIbk20n1c92xbxrJ1pkwI0yWQdTEq3dHYl+G6s0tYXp4uIndfliCVtqT
DAsyHYONPPtkcfVBHxazCLdBgv/XpEe4yjc8p3I56AAsMcX078hc/ODfldQsFFXy
dFTSsC+JUUvpAnDf/x070OFWbdRgQnTrogLgjb8wYJDV/gba1OkVp2M6E5oblkgv
EWM94QkkVwapbfrz2nRtpbNN+g4G6l+JSIly3uSHswMYesYHUbTXGqidIacAuucZ
jQHFZp3BdfLpCCfJWGSFqtVyv+pvHHS4e69DmlW2A7at44YJ68zlyvNyKlzBrN1Q
G7sW2bFHKsW2Ia9mS+/mjcp4VIs1GN2Q2J1N9Y6be63jD7/bZDIaxUY102+2P4rR
18RLrYnCFbVbZLR6bwkYBCB4r7eRa425O8okoKP06BUO6MXZseKoO1K+jbxFn4lg
QZ9NW2Cgxe3m/O3uDCOacaD6K1bySLJqtnrdnqBSKftmcETVzjMMZ5HXl2Qbuvmn
z4KNIc9jycjVnoXfmsNXLC6DKtrIg+EiHv98YRIMOdzptFrurdBwdvAdGmp+ymMN
OPS8jnH4XJIaF5uyNBLeem5GePCo0nefnQhEChapiVjewp8k92XcC7YtKfVud81W
r3IL+CVEMwal4Cpj1wIIPF3at8lADBn+BSkXTYw5jgRKOY3K+Nzmnj25qy+L4PZd
ie+NDKAFaSXgeFgiMu/OAz3CsCt0kdSU8Vcb+UaNvcX1/lJogMC5cLjt03wNiaCw
oJCC6lyfs4Dmac5njAXIsXmkvZ499m3CZNoLQGUykwaIgKVAnCMLdr8nCjLHT+Ld
sXc3lhfUNhcwWxfhdCBniiSq2S8JkahFE12j6nPMzd8FzkxOKh+0q86+SJoKi7qx
VHLeadr403Rc5QLGGUrLrqMIY5gdeyFc9RoHid3BZLK0d2OyWYXOebdNXQse2Yk/
Mr+2g4z2t7zjrtxPXe8A+6P0frwPsef/8za/SJQFVYk624g0tfUb2UVfMIhQufDD
KJ4RH2YLMHK8ozb8k6boo9+6h6eRas+HeGBllPnE3BQPXxhfT1El5sXDnlj7tuRD
pLr516TpRpQ7naRDLK682uH+nW18whOoJ9mVFUyHTvMkqHfgOcqSa4oqghFR9L4S
vJWnTdd10XKUk9cmT0UlaDFZOwj7uvfXY5wKlsaFWKqOACw/nWP9PhNGHmY54tEj
xRMzLNjAq0TPEOzvhRfmnEB8H4iCxB/N9PDeoujc+dpiDcghQzMano2JOPICgl68
Q9cZWOIo3Z6W+KqDCz4g29dylt3mo+7tNbMmg5uQbrZb/2oQgXoS98ezcz7VLsmj
o9FQ6VVJytM+CnVp/7wV1iIAaLgv4q+Iba2etTAi5GrlNqBtZiB3E2BpmkNRxhQv
Cb8cc+LlfFRJHT14FVwADDsJI4ubeXW7XlFTuN03ogo8gI1o1Fca8nl/8AKjWTy+
nnKub5g7ZDNxkmoI6/T/L3s6uYkXgegnpLYfGqyeQkCpL2gLmh2PwZ9rXpu2bElh
oR5VbugCq4hBIovk0GxSl40viI1+lz1NGEpw4menxpR6Ss2AUTH7ux/cTZ+Fcb/i
JSy0vTtsRAwaaRx/3xyig/4R2oHGz+gDsX4LyIy9kAN3vJSC4HogP9VdfYAiAcuv
qqYJ85jRBh2JGt/Dwp5G1eZV29G59WoshSsDbqknWwts5FCGBdcnmNOYdJQl9utZ
PJz0L3shqOgR9Wr1LKdmDPLZGvjx4NeKZQMqIyZh39A0BQhiPMUtzCaYhbNA8Q3R
0QFvdUNI87QvcdUtjmLJMkTaRUT5EEz2VNMalU/NfOATuTWvxO2aGKO0bLz/6M4e
NCM3drLvxKNfcEhZnrMtTltsLAv+k61SiVsai+uWBOyYxVS1z6+3ePJ9e1cUVxoD
xLKiAr/xgzDbWIxKMV48dLoiZ4wBuJXKSWFcvAMy6fPWXXkdJ3SkSKn42Lu2iOE2
fkQ6E9H8QfsK0aLG8ilL4qg9sdF6VqhsbJ5HCNLOfC9zdUMi+ROu8kLBnReUtuyn
vBQ7tDUAqy+kXOyjr3agwb6bMTOFhJWeMDZS+7p2vAuc13yrezpNtgyQj3iQLkoV
sGumhDc3AtBHBL23eHt87FSNFnU7HWZv4Xl6Fv5sEhHasawA40cieBzSvDENltys
G3VpGn92vUFlQkiwLscqVpI3Qh3v+nhVkjT4oZ515lr0NErmDqBm5FUy43wx7Ik4
jhM5Kvj/VadzKAujRSe/jTVjlTMAwqjNLBT/yTDCT3DlBvQ5QmLlbk7atwmfuE3H
eCAu/Lf7akriLW31ykxA37uRV7OBjjgSLZPocNXoeTacYPzKSeMkZUcSp1HI7Kgo
OTJxk8x1Nhw3XfgZXxyJsZLK/522SfGPzRQyzI+h29O6n+SHt90AUcCBE7Kp2MHh
+iL1AKdavIxpsk+UWZ2SRPMxFwM0KtBvuPmR8kkw/U6lQGf0yVBnZ2IZyeO19hRs
IIvT4KGQWRYuO7IDSv/7pEMkt4YGiHx/7riAbyO7xay3aGLsfycl+wF1k4zAmolk
GzD4fxKeePvDgzRAZwWIeonMQO2PHAMn9MOtx1AgIgrZSTHBc2Xpf7dqPDud6GcQ
/+yKxpNo5n/9/aZovIQ2+pWLGl8ZOzk8HJm1Ayrg3aDytMWPgP6nTBD48T0nXfWy
p1sjIAGQl8k4cxiWfvibkm3lWSi5sk5RnD2my2AOP4d+785EvGYpXPmRvjNrHm+Z
mGLcaB8bJ5jHKaSN3w/zvpVs3dG+Wegepwl9GzTOHhUsjTQoW4lD4vBdyIGmjCIX
X89f5OqM7fZpgXXTRSbsfxZnJ/ZlsKA7eMl48XRaUjnVPqXNOFgLwPLOdsZbfniq
Nma2KUy/yOTY3BpCVyJPqLYoFBDUaPtYg2ve5mHgBpxCDtfiuzYn+ynWEHdVUaZE
ACZVRC3scBR1ya9TF7ITxO9tMgt+xAyDmPhrhFfqI/NsSR2+BDwle1X3g33hy51j
iZqAg9e+Y5E86/ErDzRRWPzDCgSOrmtxkODO6qPkiwkV2POqXeISmn2JJkdKJDFY
mRkfC5uZvXZot4y2K2EMWQhUnGN/bghIAgEGwls5G2V2JTm2kmHcpt1NZF0XHxhz
1f8hwxaSFjVGLcXgQvtCvN6jFeyaDQAIP3/3zFr806ifoxaWbQZPTtcIH0nZFRHD
5fxrcHZPD/XoljhflAcnFztkSNnJllQM96aNJNBM6qzLYOHZLadvWfwlpK7++XC4
QnmLq++BoSXaSr44SUV94Fd/djKd1q3Y2jnB5szgHd4UU6/T+LcfX5CQT/3YEnnL
3hZSPBzaiQnRbdHXtC0CNOD7SpDkTeEF/77f0jtHxkFvMDjVg0iYsXPeI5nZ18gb
WWhRTxsV5ZzOqd0QgVriPrNJ9VCZye8a8k8IiVVen3Kp083jmvRhyBslGNpiMPPi
+fZtgM0TX2Wwt9t/HrHmkCAwGLPQ6NDZoXywFEC5H8cF8y6lh4swimow8kHAXYBK
q7c12S5qVMsUxqigIXhlyhCEZKICtlbvREZ8zNmEMWu2eU/I1iiqZTqayawf6MY6
21e5zshdeE7etUJ1YJLsMvI+mt8BAJT9B8yrXJpHUtHOYOTD4rEeBnvuHeKlHA7i
CQ88U/9u2z3xhoytGkhp1lSSz4mtJuxWeLPN2q3D7C09PhTZUrHK7G3HJPlXa/tw
Uguevbr8wX8Rmz/qtQzoJm5qF38hJZ3RJl+HH7VEbymtnks4AiXu5DCmIAwwHCAe
BrzUFiOohQuEA4+xWBgZsxbdoc5HMROWNYeWm7o77AGplC+IWVbZPlUPueIXo9dB
DCvOVJmwcwLK4a48a4JkdQ/+610CaU1VWyC4LGc64dYstDvGgb9QznGuGlVR8xOZ
jvSMabscyV74UXwSll9Rty2z2imzkN910j4JrWsDoo8g6yKDIWb5gvHlA2kt8SoL
9Wqq81cHSw6y9t/upcGQ/jXMjtJrNXdUCLonjLLZibKj5Kij0SO8G4vItLaNTHyy
ksvvhbH+ZfqHPc7eHGFPtqL2RaXGVYfHbDjI57/Eqjg1h4Eteukwq1DkfZMmZHYA
kf7Er67CP2hE0DyOmkANe1wj0LCtCCDdwIz5lFCJEX4waylnEmprRjT2HJYhYzT8
VaY7lXfxyar/IqO5jAfXYhSwxwqF2BSMTvPPxVUdpl1a7U3r+Q3xtQUS83o5h0zM
GRl9k0cuq+7NAk60/5YUvaX9DAvMb/U+5A+IiIlsp6crMyqCne+UJrnebvHtyZN8
DXy1tqo0RCV3g9DH+R1YXN5ToAvhmBXyL1TWkWznYN4pfwVOOgEQePnG1orcqBwC
8LC2Ethzl5QiuiKKmx1W+xz2HQM8J/VAg9BaOl0Sl8QF1/7eRBhos1X0zToBO5pd
Gruj4XqK+tbCAUcOz8SgI+yHmKSLYtGcTbjRFPXQ/kdBcLzPyOUz/MwZC2r+DMDJ
q5r1e+YW8fkaR2bnyCEtra7IseKMdBwRQiJU8PhkFVHNQZ7B0oBt30UvYA6Jnlbc
KnjXdvXk/7FI7A3zmjVVWqktLwrNG/MuHzGhLU2OmszHQ7jKDKxH8bx9AD8eZ9tD
pJcPG059mIOmX1W0HeulnUNgrbQhUHXwSaCjBv5bmJkfUiucVBQTi+hlVfrtfeej
j7Cmj7hW3BHsYk1pZKPE56vjX61JciTRpFXUDy8fmkt1nI35xJgjGPUhLkuk5jVw
x7gOgsb+ruNXfp+R2vydyvIpRPQI/38L7voaOXO4tcqSy7GSU+ehZBraJXgZ16CS
IFV2XsJwxtPXIuK1lmbMF/RaaMHmaHE1YjKcv3nqfKlKeA/M7+lou+x3kjJ5LRh9
fw7PlTM8aFh3JDSvNDLUcPVkuRWxnhG9DNqXpmo9cZik23stq+Qh5kCCC4PPbUsX
RNqdoBt5inOVoqMR4cXVtuccah6yhIHPk2IjPniMsEy0kWKlgYPQaCeAnmA1bQ6U
zOcYehLl5XbKg4oUdOt4v8I3cvQJIyzc/rqATkJumoRJye9Vjsd5IZ9YETPB7jAj
XOeU+yn2xjyM8noTMQlDaia+dPBwEdU3C8dK/ltyQCkbSx8iRbOLfG/3YZGS7FRA
fgEVa4KW0IQhue4hsCRcNn9SbCAfK2lEsJUTf7Bl5hLtWeUGyNKiPF1PkWNpwsWx
jybTLR80zO3PXg0yzho82BQR49PqZIgLLqtfQ4epb4gr4zFL/HTb8Lkh9MalZc5d
+B/htjLmYF3k/T33D5V2ZsTwzEXYoQIos7X6Le8M0LIY4NnkvqqH+xoJFaZ0MUab
IwMMguqSTYRVspKrDxaWk3Pp/7sovy09lL5iwajgzZkX73QpWFc5/hsNTWvSDQpz
9Dhrqx8W4W/81ECCrWj1bz6WLmHKRoIg4DYCqxWtsrY9nq6TFsa0yxVGJwcGIlrG
0PVFoXdO8nGoFM7lxUMksoaXZ6wZSCDOFXzsHqx4P/DY/MthTkLVl4VdSCZ8LlNa
7QIBu4Nhb9+f8b9cyLBr78LYh1QY+3ToYAGh7x0OKmyduQ1Pk9xmIgd8OLYf172t
Tpf5xcCCxRU2KMrxMDGnsyUALH3r2wop46CIL0UtKfXn6oujxWsJ4HNqsBfE02JG
929J1snwwGT76hJr+8JHIh11+wh+cjQZcn1g+5Hxgnd1AJyBrgAlOpV8zVgTh2kX
xkfBbdihQsva517sRo1ZA8ielMsGE58TgcGhGDfVZ92BRaWF7U8/0u7L/3Mjg/gn
m9H4hVatDuj2z3oi8ideU5aj5u8ywTZhq5ujUCyPL7iSPIprjjO7n3QJ8mlBO5z0
yGxJW05iqd9xvJjXfarqu3KfL15hnoCJ3nNLNFCTzeJiS1EDcWCgz+caRVSPK+8R
Glh7JlZ/DmcFKqNUpo2ShcGvHIP0QgtEqKjvy6AzJPwh786eRLywnqP7q8zay/Z/
ymS/+xPolvcAVOfBrN2BgeGCnXieeMsNy4QYGaqpE68hdgUBKkxh45ZCo3r2iLNP
Tz+oqvZSjMt9bGIZhe2z5tXjCU1GWi/2zcftOR58zxbyXRfX2qnaXPAVFbJh5okC
D4vnu7GO+2JbLqIZkS7uWmiSCEjDfrPPnjXB7x1JfiuT2AlnRCAY+XqdWmFOlkoF
QYj3/JaP78PjDNqpBFLqWBGHQHSps6kKdGFOMFyFRF7NppmwMtPSlE4+Truxn3Qp
qCKYDsWehsZvdzsyHv9YLK26tIEY3BpcCmjRlPRz53rSr+zkaMatkXP0SGSykhFU
mk0ddGgQ94K7vRFrDTyMz+uaBaztjQiunrX0KJYDEDtZff4LuV/u2YcAMEDhqnWQ
4MvKs8xoZInrxvIKuCwJ28HuUaEI3yvRQc63ijx0bAXJaxEm62Rv9L+MNu3+DUsd
+lxjBimm8wC19OwUFLVeD4dkY5zeMV6Rq97ZUt1R60lh3BtfD8hwMjZyByo6wqa2
h4bIHhqameXpFTDP8QqjC2d2T4cOOaEFJicx6X9mg0/H2QpjLNkZhNhcw+HhmVM7
iOX94F2ce3qRfQY+zTTv8JK4bF+BbxDwVp+G5AYzU7kzQPrb6MMv+XiL4SU9O8LZ
AbRl+l2O1NajiIdV6t+P+lWEOw4mli5Tgw1UIUyRMf/vs55CBt4/TQkgNsch55+x
QxCIMAUtQ/+o4jnH83yclVZy/fC0cEtTF5NITBDx4lATua3BlPumHTs/HOYk8rRk
+kGi/Jsu50sAQflBykFhVviwlM0f6QZFjmM+E3jxCXTnOe/uagYv4L4BmTO+pvnE
xKwD2pP6A9slrlHZeGSKhS8tBWDYXE6FwBZNV0cEzQDVwyO70v1NMqz2/SBIrQaX
3yQ1WmFFtewEYeOmIBB1LKzwIGjb4EW35hrdl9tgD3fCR1yVkF18icCHsAr3TSED
9iQit1i2Q6tETDLHhZUGxMEoIHytKUL7Q2GjK+rSfY7tCHA5H7HysxzJcn4jQq/B
k1AOFiJH+a1y0XoknKx5L1ebaIUT/fl40UuJa0q9KOH9QonCdwVNeqK6HLZx1Jna
yXrDyhWBROlYbiDCiWaPnwWhgotW1/0PG8KQ9+FtJ0fjTVSP1RTEtyqKoNCebzmx
zfCO/nd1e9RKu1XW7L4c+A7drSAS0R+/XRxMPT+SLM3aipZ0oIjWGX1HvEY85N0W
WkQKBOVLAQ+dFlHRLZWpjCPbUSA0Q7mVx3rgYzfb8BJDJ8gFHv97FiREk6D7uXYL
9Du9YxMNcJHc4G9ncvCeZzYjGgppXlNmJ+YuYBXlu2TZGu2qjUwBCHr8by2wBeoO
PquKhLu512qAus0F6uzpLYcpY4q3pNsXhC02z2gk6vZ9Om6ZNXjzkPSTZpnw3pkF
gkUWt/SZQj7gZAxIlvJEcVv+/iJx6KC8IC6Mrj7tLifTUsFvcevLYRamNJodyH88
u/pYJsbDyTaS+n3E0/IrLO/1Zm+SRtH3/2MHtmrZedOH+6GPYqNhd8rJ/cvG6S/l
5Dh8SSq8rUyWT7DFpCScI9fwCz6vqZNe55Mb+ZA0YcNsX0VMxewtsni48bRDPvLD
0KdD7LGZRk0yzoxAYAudf1c0y4c1by/ZFSe78ABcdOSyn+1XyP+RiYb47rMAiC0O
kpABCtGxJ26aTRVX/RGYw1i8OcnbqRP/0GlVeoOSRk7CC+Vy7jEVvZQK57RPP/YK
RyzJxq5f2arlVIorcP7zXP3TIs21tvaNky68MArUu8cZEC1GHrXXdfPWFJ9GuXOz
qnMaV78uxkt0enbOAlof7EDS7iRoSyRjcZsyDhI70J0SY/HQFHlzEP/58jnSmImi
JN+/CQsQrPUiAtsR5z9uct4V4ItzMlVzuQpgWEo9hg4SHSUEABA8KbTYsEwQo3kb
uP1spiDYUZHP5nbWoI6wgbLEGneyoeOKBgt1X2zdSpsqUVrTe6b0DFh0m90TpOH2
0Wblg/3oiUq97f10izX2OiiED6FT0M97tY0IJmOZQvLdNp8WmPg0/TC+1xLNTuFV
CKJTtW1G+0z7BcPxICw0FZH1szVjl+a7bbfdOcpGgp4SVAApuN+nEP/igR3dm3vY
BdOz333JAcuPdstL5aAVPTweNVHmOs0T7aNKSbuYpMfpXNAw6iCF9AzumNC28JyW
HkItTRm62/so4v/1Q2QakvIB8UfppidZyeo1Us3bXrZP1+NV6DhH1xONzNXC3ubk
EYSzd8Td6yrXZvtLFazNtDlJN0vF3Xjqn8X7ZDpclr31sfIsgAdvZCNU+XjoWLCV
aO+zU8vGbxjb3jpgcZxTyWQOY8kNMdXrQ2yDbcit0ODHXBYIkGgYWzXgRgvocfOB
HiI9EfkaHyAub59Kgn2RoSclGhhqULSDn9LjqBcn1v/s6dp6hluEZ2/jnGwG2c3q
HNY6+XwtuFa8qe9bIXOEcCovPUjCFSmzbU6wV4EkyguioWaZTEJxgMFDTTO/5imK
AUvQblXrlgr+hbwb+4B7fxMsrSd+zDKjtmer0gX+0WaWIzJVV5AtI2gnDxFqGNCH
IgbSpwt4heXhvhf8mp5C5WvUjUkBv0gWy9dkY2YENkTXUeRfCLbN4URTsCaRfZqR
tCLe+6PwEhqybN6n8wJkIsGFqsd0+RDDPjlFYFBAKRPnQTHN9+2+ybto0sCfvI+n
XyJnZTgm1u3Jh0gvh9aFSTxltBAQshWkHj7hXsIS+EiztwS2U8BfrqzidxDpQDEJ
/hm2uEJ6wxdTg9i1It0uFo5KStvRagMIfBZtWTXNtnTDPG5IiIZO0sWK9Uk1h5N+
lcRF3UyirQshGgotQda8XMCo+KcKMoVxeor8GFdrMahrkSAyNuFkhAOBoqtA6cUu
uY/CqFedD31BYfJumoG0O0y9DnwCapmH7tOy9OhurYsLPSYg/eZpjL/sRmL7iSq/
50EW/pDkhEkfXxA8Y1wGSYNWngwZOT/K4mXOpzaIwWM/QZMLcfvTqcgN1lysKuf0
uFZ9nmlpGmDGeEGPj82PWMFQbxjyyESEwbfLiCS9cG63SU6dt+9NcJ1tN2P1aSzA
YWcrK/oNaCT2bgnq+phY7RzWq+++RMwFFfKK62ss7uCViYtxWvtUusI5kqAZiSrm
QcvloxyCfLH+FsdR9MGEVftbFIOTtVMQIFnjoRxha/T1aITAvusoDXMY9AKOwziS
Io9S3o5bKAcgt7h3fSXlO8OcPmddCkbxkKMgtc4BBOZcUYI891IGNGC7/1wc3uY+
mVOL4972j9sh/v/IdLcW0eWPkhuazwRjwwqa5DchAKCKclGlWB5cYio6Bw0kYKqF
kbcvziiHNXB132MhiHKLFdPxuhKRP9DTVoTW+2ZdJUK7Y0FdkNe6yv/wgUj1n1Rq
lcvcS7vvX9exZxF9Dn8ZTJPTEPq+h3eSub+KJyL31zCd52THBZ1leRl6YLPR63F8
zl2aQUxgWbxQd1WOZ6nLJYlF8foIGtIfDjjF9D9VSEmIgCzcB7PmaAPvyLr9+F3h
c1le8vcZ6GWj2BaBWax89zctEdPrINpFm8s8+trzKQUa1sY2XRGrF/x0a+Ns10fG
0XcA2wg+cwrlnbQFPFNfNZ96ZXgU3uRhCLuOnclmlIhGV5xP6uERxPwBYgzcgRHB
BLLC+upfeVPez1tetLd7hvn0f2tvFYnfWhOW1zADGlhr80joJeekNvVjZvToZ1zi
8LW7lg/WpFZx1cC4ZsZh54NjxO2gqoM0xZlbDKHl/ha6edejEOHOtZM0ZUjTar2l
q+mXF/ozkOFu3040NlHsdPgoZ9ghf2nEOy5steye42DOkRaaNPzmGhj3nSNPBX1o
0bkHhl2/TfZ49l4Yg1hB7VF1+MUKczq5VC08SigGDxPA7nBuUDfzpHJbIrwdOrB9
6b7zdLhGnIVRBJg1RsNcXilyti0B8eDYeCRunYbRX6kbngLepv7uzCo0tXeMMGfl
ZLG/cgdhZUQHD2Pcpq6qWWapHbYD+eV76pKaYUo3q6ey+W7hRrKPOIcl941IIPYv
8k8weZpP7YgM3QWK76Yaen0ERJqGnzcuTKQBZqAq9qKakH/xosIdOJ+SYIoSWzVC
Py86kbCLuNRXfPXEEUwu+5Mmh9p6F52G4nlskXV0Gy2EgU1XdhAjA7eRprCBEKvq
uIIA/uk13MBdt99ARsBE5jXpWYbiF6D4/2619111qJRDQsAlUDCXY7/YslxvzvMs
IYTWPHCIB+sCbziEi9ehwyGl9Cq77i0LuNHQhOwLHaUqUV14T4bmWM7Yn5STioEH
Eq1qj1wGH5Tqu5pwuEdTcEpUb5J447IekpgEe5lDFVsKs3M/TIdjmh2/C9y8OUgS
s/vz9Av5eTaDhHIKHBpJx3UxekNY78kRKaIvJxwkmuhIh6Tq0ygHFQANI3s6cN+t
2FbsaoBlQjJ1NBxjdDgiqP0nCggIkG29TW8QYlkZg32OAh4gBfyv+M/FU1gUCKTz
nvAsnG4K2O68fXxyxW6styzWNpaFVzjOrK6UitYa4/zUWjsifvKZyaP7xAo13rTV
mJ6UJ4jkgcgEo0UWGsxl5A1nigbNCEpm21Tqc8yFqt45KEAxe3IyjJr0e1bn3OAt
bfeRCT8JAol6c+g3f1zSgijFLChBgMzE7sVfWPzW+B7os4qZ6gPoe8maDZKInHgs
NKGa5HlEsOLfqDC5pPl9tt9XDnntU/VVQhv9+0twzHk1xf9UsyAhcCPJDe5yJEwx
Qn2HPge1byXpLRFmJVihIlAhXoX8eRPbs6aFRLbgx4JIivF/toD0yPTEy/CZ1adi
zpMeoxygFxqaB7SAKMkaf6eY47KaUEtHYACAZc72ajNGVaveN9YfrVnjjD2l5dPy
n1xm6bdYcJ3QIIZ4hpTvtFejZqsKcT4wEjTfoOZSChIKpDfpRbovWn0Ju9W8dnbQ
CtquVV5Y672068sRx38EVujQuR3nsTqEHwlyPR3na+OANNX1RIOI6WhLTkvo8cq9
Wmb44N+J7+iURgoWKg7/bMeWCRs8mHOUzxxUsyMiaQyM3cx/Q10K8c4Y91KQnjNk
3hskTDp7ZT7LnB+8XEIT4IeKKgR18FpKoObEJVekQOw4/ruItLOwop1LmQ6rV5n9
TXuDdRrLXECqrnfRTtviiAs1pF6sVlBTSEyVounPlDVX+9qZyIfvDzCUX1q3gtsx
O4rQFxl/sRUdYwRr2QJ2Ln4xsinMzT9tDCy9+B+ZAD43LzURCVwF+dHXfy40ppIa
EojSMWEEJysGqViVCwhpMqRGb29qoMEhMK28rylWR/K7RO8iChIg8J575uO7eNVD
lOMHTrG16fL1PSYliEky4biFKanE13DlYar4QVcdRnrjUXv2rE7Z6rWD3vWO3hnq
lXWOI46Kh+pqNuXzaZ7YvHi/GgQDxAkFKyABQn/Rm90UX+0JsBD2MNR1EXTWKz22
mspbRr9jV742Cdwolkua8mtIxEtOq239BW0XtqOoZEAJ4n0OD14Z54RC6OtqeFoG
bbW4c2Qaher/uvQb51Zd0B9kREzWDrkkNR3et5J9c9uadSEmpttR3yOoO4SYGafv
DalFBdCLS0iYqlY4emMejdlWCcD6mqhaS2CvUe1192KIJ9hq79wk6s/9f+ZnkBag
/8JMua34BCsI3yQBqL6eJskDVwdR+/gPB8ThZKIApUW0YVc5MYMz+MNmSyeqbOCT
dSl9lkC77P2qXqtg7bKNeZm7mk+YQ0HMJJg3p6DgLfuZi/0tgWeY/VDYuIYJ0Xel
Q4N4nwDeg40FZM3dPLzZ+ZYi5SDyaK6rMyDBtul9Ub9bxMzd+aJ/hJgm7boIz9Eo
i275QIyFTgfOR1dxQH6AmhUZ/LQC62zQTI/S6WvvEPWsFkrDbAmk2qBSDrVQPUBT
LQmH49uFzBBnSnbeyOuR8oauyeS/Ghcs+ZZkAmi6Qlxa7Rxq2b8FVGeABuzKRBJd
EmFa8bVLrQeIJsEbszcdoDSJeP/yHaAJvJMJBAzlV5LEq+VjQ3HCkMugybr7ylLw
4KCCSKCQjUqE9EKznekoNspgVG18nLyirPiPGkAeeZ5NSdHbPEVKu58BKv5DbVjD
nhMglI037rfVNWAdMFovXgeJg6guIWLNONgPlOK8grN04cdBh7esjJr3xpxFiR9y
EhLNe906OWa+G/O7z7WgJX7FsjRI1KlUdF3J3Zb7nLPK73v6abCrfV36bQDASw0p
zdBfr+66m2toqFzG9S+CvfZwhzLMzbuLOEqIkykkyKWeI0aAdU6s0+/WEgrJgyuW
HLYp3qrmx2bXuKej23+U7HXH5jkLKJ2096em6K8aekxzQIGdE9oUEcZx1MOwCgfg
MB0ml4eE75qRPJvXWoRyrEUCqZDr2CMlGyD9jXiItsjmeseXhB0rniiThKzJxBkW
ahKspeDwKRdojVAR/aLKIPmcE+gB//T1pXcwvPWLvbsWlFkHnosvlEvBaX94OXzO
+7gW5iBBRMGyEVdsjo9rIvjN7KgAFRSZCdEMJPQ5/WvHpUin6d2IoutlnMvVYG5w
Ks9P0/njXlOQRk72Wr7JK2xE7J5EgdgUeh/ZL02hZxJ0HepTANUFKB07A3f5ocbO
`pragma protect end_protected
