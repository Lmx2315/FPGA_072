// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.0std
// ALTERA_TIMESTAMP:Wed Apr 26 13:36:54 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
JwvEUeuE7d4xxWpuZdS355aYBxRWR0O0O/h2gmBttc/AOZ8PT03Wef/JnSMBHpr1
a2ijPlL3fyQnlPvEjQXVbiYYsLQv9muYGl0r1qb9o/Ru7haoW2TN+LsYB6p5UNCv
fFOxZguKGARIYqp4cM0243Sml5RoLTUiyEJeTX0qil0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5792)
wV0wHwwXTpbqgWWYxKyepAzS0BgP4a3DGi6yRFnSE7+bstqxcbYKa3ML1PgyxUrE
5kI7RYQT46JDUAPiSd1/4kcly79RWW4NI4i4QfLG8TN1VjgfbR31nKe1r67dqguK
Fjs3NRNOLtAmqWMA52B7v7B5VPCy1cyHqTwvoZFEirs2pbUoifjXlenmvtoeTvma
g/3L7DQgGVqlSxRfib9ZPSSukdXNeUYMj2pvLGOFAExwyQYMfFBdLMYDHSKM7bAU
S4wsKO6loNjFzjT4Do47SACks50OeMxLqqsyNsuuFxOmpk123YZSVNosWN7pXip8
zQyKPhfd2dEqFmLMSLs3pB/jG7K6+Z7lvLsZ1CPezfJr5t9yw9dJhGWAV4Ft9gXH
z05VaGlSBCqexNYv/KQHKNaVs4gH2qV/e7FMlj3hwYmP0D7fvAg9GlozBnfZvkQU
UIyQjsE3o6gAUd64N09c+NO8KRDy2CQAOrNmD9K2CbKRuq/X7BV9KNIk6aN83/PU
bKhzHfeCT3gS/mDp1z8JsI8+3wN1asMFntvMp+yY9v2tvZq7NdWkX0kZco0xIRUZ
OnoPZbxzqJFLu3n4Ky/IQn4i6Ldla58eVI/XK4s6+AU+ypaB24N01f/M5vSt/9Dt
ynpFA9poE1AA36Fv7sAJJmDZqqF1FXCuqOCsMie59+iuVq6yhivKeOSSDVFd30Rr
JcxgLnOqkItbX7z0/9JSJ0/mb6uomCfbkxFhg1FCsRjNTXQVujA6bCUgLIyEaBxg
4RjGMaarwtC0XrDggNvUQhGpmWSnwsJI4miJcxHpqSqbmXlbMEDt6Ng0qIaFW7lg
dMNyTXE8lYsfygey9cUq/5999LFGi0ovXYg+1tu5L2TXgrWkPPWt26kPEg56xdZP
KKpSDeUDilM7fIP8mnReli+bQa7ISIdJtb5iXPCeM6Pe5iQdr90OlX9t/vMQ3CLj
3Pgwvis8BbZ+PNNF43NqyHHaoH3VY/ofyZFMW5aw0Dg/ePR9bEQYJlFOrrrjLQC0
TbaMgTfkcMqnaCYI69EbLZqlsEuLT2dqrUheblJdJ+78Egc/NNxSKSlp6P2JPcQl
WDEMt8NPmWaxQnYXgYLtCt/Q0hGG3U/eYJsfG3xYoR7sNVpWpdjg1aaugAqTBj8H
zluUZSgczs05PkWDLbmyxcZFuOaJfsDjIy90LmPFdI1ulHMnWyt1V2ALBIrgJRjD
xi3TbcJEs0im/5KU3nDY2nt8PM0omTRCnr/1l52bOhYmZ6EKCAmZHUF+6dIywt+A
uPVNujcnSeoK/ZN/KYlC8ztzr4FyH6hYR4yQtw2gbmNSQrYzScHhxLjEMAoQ+HCy
BGUt3DWAcG70GlbwK1//qG17j7VVCAbhfSKWW1qvvDP1FgMol3OxgNdtMdFBS8rY
e5j72yVWTL4xEKN/Qy59g3xle0x1jEqxCdg/L/xRUG6A9C/i5HP1QxT5A7r9UEE/
fBA0YQ6v6tyckePfv/Gd8NEILsup0kCN/8HbNAPXcTfDCybB9iTp3UOiBmCBR99L
L9/0zEspepp7XSU+hBHKafQdqe0dEadNFX8XqjSxaG4hx5LrdQBRC5B3YNQz3+dL
arHqqkFojaJimJ6+Sr4SsxpMoCYDV6PzGXKYtE8IWLJnmOZyx2AWinxwiXcCA91f
DbNMpyagFp26Da1IHRIM7WC8SoQ9VAYaCWBYGc6/P5UMdZdl8h0vRG7ZwcfDx859
5ccVPavnpfqffDjgvRc1sQGkICd48PkZDcu2hFiLx9soskTBk8YUCldZFkIOGsDY
uelJZFEwa/w3nKEpCLihruswA1VvikCU0m1l9HSkZ981xtEvpEuB9g3pAOI3VP7+
KuahJjd1GP6M8HXSzCh/g1dtkC7EfmAh7Jdk1NGsCeMAvtKU99CybdLBuYkWVa4V
uPpeDKymOwxU0+cG2MpBfopzcIi83Dr8PqMO76mBHyJLOqHmoHS575zV3VGHKN3L
FF4ail1iT8q2aJ405agO1YjGEOObgd2pWQB266rAQbJbotXMKKx1tTD8hrhv1sEC
8IAp1OeW76ouYFYO7iFrEGdc0f1M+q3UYagEy4G+fl7anuvzxQqk87HBS1HNeHFK
0WQVN7vR2RMN04jLC0Y+0NfIq0+ThhmGgLfJkxikw5mJtx5woJ0Ui0KCP5/NvG8a
TA1dy0ZwsJFzMC8JSkU6rg+pa21e8wA9Q42XQwEDW/EjF29pwld+yuTDQ9wfmvK5
0yzsF9BZu+Y3croEkcDrzhEDVnU+MldlmYtoktSDDXOXlXPeqja61nndyeYN5i4f
QKjYBpJqrvGjWTv2eBxQyTRLAtj558GU5llFSlzhaa6M9bcOS8RT8bn+H+P1IxtD
q8UiMMjkmszE5HA1MX6NT1ZgvQ40X2Vl7oXx4x9IJCQNk5v0d7blo1Ku4Ks6DQVT
CPxDPxPPIlKvPpPJf6QTZKoXY9Gj0jo4cisG7UWjbm9D/uP6gt2nFq2WdcTJJOjF
Tdg4J0UTbZZcDNNwS4oXd+KmcaMqgELdCQ9pHMcvGqZ0mgDKOv+wbBr8dt2qS82K
+n+nwWzx2SgHE4Xig0kj7D9opK4L+284b3/Q50mNyEMcLTAuO9cEJHgP5CAV89oR
W66WVvUwswLXGHNlmV84AF6MZa0jS7Ml2/2oTdC3PY7ZibNb7k85G4O+RTQaByKw
rP8PLGWJJYnevmDj0+bG2h3io2Pw/otmd5HOakJYEpVQUOozczh5SulTHXDoI0nF
/6rEhO7eTfFlAhzchWekoGUvU9Npa6/RayR0yqNCYOslVEofJ3+o35n4xq4k/glB
D4L8cCzIUAkcqivBa7Rc8olriFJ7wUUHz57Jw6cxqJBbSRppy2b+D5Txh0zn0XzC
Ziw4eb2Oqqa8+MgX7JeYYa/DA+/5ewAaxnvwSlVj+vxr2ZajbTN2Ao4G+q1SNijX
2/2wSVBohuaVLcunOz6Xodn0Ai/2g3W1mDHLvZacIyZb5UNFIgrRuoMVG22D8WxY
JQxxutnGwnR0bpy+RYu+oz5A/pdi5f+qzQkMrvNhUu+gqzcHZzsDrbw5cNKMjFEh
s+9bof5QBbFBodiArK12vCF+OvYgdQx29JlAET+nTAvxcv/6J0xKYLIhBEs6zw/9
Y69Tm8D6Lbqkcm1m+OJJFAWJIWYMFymJNARUuRqXrBg1KVTdocxSWSaKmAuVKoDL
OGRnleAQwNwEuYBDWwQaJN84b1EAbYjK8nj2ZsMrurOxu4vuadHN11QhOgY/Rdvi
tU2gUab2azNiion4YPTHC+FEWxvQt77G7N40OFUITxw9shu1S61YFL/hmJMUvpQH
oVzegEtXYTSVmIZGEsGggRdeU3vAobvVXygRMK4qxUGXpEuSUBeAKbRJQXUIiulS
OZPjUCIFAWwDJYnBi3UqnRgU3epKZNfPiTZXLBwaxa/lvelKaJ+pk6Ys26SZ3VWC
BoY/NBtlkA2KcGjVgN79UFZedMHzpA8PZMLWr2y6vrRKfzfW0A4QHdpmWduwov4Y
VO/udtN05DOuCEmuxSvVzd+ftkUK6OJreJlc5ljCdZZn3h3ZkYaB+KUmEzBvV6VT
smsvqOdAGvHCezB1s8eaZW7msz7FrREReW0BljSATYHpSEWWOuAb0CgQG/xa/mhb
F01tuRA1+uF6b+p6hwGBtmbyuKOxzbhzRQIKxjeIUTg5zD2A+z0IUdneTqwcszxw
SptW73oEby8uKB7cy7NL6kto8DKrTlznpScBCruze3uqWTUmSG7O+6mqxSPVj1YE
zHZ9HIGibndOtPvKGJYjDHCRd85/Rf7LfNmKLzI3aVTajfGAsoWzf3E/xkHlQDAK
ncCaI8pb/ePlmeFbVsDeaOJG/9GMUWSKxtsuqwsrGYB283+SJnHczfUOkODQozJa
t30FpogtCBRU2J9ad3qs4RwrmFluzxnHV9OnufTxs8bCYcqqQbFO06Z5zBa0gpJj
KYU6qBoP/uT4e6dfvY2wvHkIKcsBu1R2phcy64fkImE6W9x5GrkMlJynOWx8ocV9
wfpyx/wJw8qE+SasMLaF70TYUf2B6AXzyCVFwrawHnRcFstslz727W+Lo3D1yU0E
fEE7nlIbfBRzEOA1a3TJNIAh4IeFtGR8Nzk9fV+FM+/Zk/b84Ve0GdybmSWda1Ud
C4fTLXGbDBkK305mv49uswN7ZIS748JZOtirx7b4ZyGgQynsttGhOLMZo+67k0o5
6QPU69/tvDIcykaPAMhAnVvLyBP76brfB20zVB6+Lq2AbWEkEzIQ0PPcCzDd3bur
94M+x3YzUQYUykLuYr10YZ92GiVxegziuv3u7Wp8m/n0hig//RvWvJyZ4XW0Sj8w
hl2seiw/0dsJ3bbc4f0deSsQ9K+atPj8APvNBEKuZCFIZZryBDUsH7ZDE2OgEb4l
fRtYMLbIcETnazqLJxwx7dJWCnevE1OTLUE++a0GGI3uiTm7Cuqs+rF1LAt8q/j9
tRN9BX2QDM4DZ40Cj3VsCXh/hJTWvEIcFqCbgO93uMfUQxwEq63PRSq8YHlrnMwg
8YzbGHdgLMrAXgSFmTjYOkFdid561NSPHX9vPQX7C+kUOMZi6Izr+jRJKWAoFVdH
chWORndFVB2Ms0XvaWtA9FjF/C6VphDYKRuOAOVAH50IDIV6qjV3STqwUCLEFHyG
++lkEXaJs007XE66t/MDwkoAvq4sqrFU8rmkY7Qe/eGhbqu22wl4xXn+KcCrAdpr
FpSmbBtU6ytIiiNgjS7ZSw79+2JNAN/wmuk6ckSRtoN++U1lewmH/YKEDBWvrY49
X+qVrKFDBAkeGCt7TMrFGYn8IMd7/Aaan1j7Yjrcbgunl7CZ+LY96zHPrKJFXv0V
nOYntDlCGFSDsiJp75WxIskQc2TgPJ3A2DswblpPScDtCkq/P9Zc45VbZJ9YOuc8
mggAVU1iGuT4yMq3PKVnv3eCqVEy3iO8QziG5P43YnO43OyE6IAisoNfaoku9pez
dt5QbOgOT9Eh+UMQZLbzIMoSqC137rm3hC3lmqoeGLlLeOPrKoRyP3SC4hkB6Lxf
UsRPo8z7FmTBViHhmPW2CHvY+6vrJwgasC6AUS47qceuTC2ZpjKqIAnsZ34Vw4zp
EAJd4Ai7pgo38RjuCbg755XsynqZdGHcPI47EJ3AjQGgWkEhqUd/bM4DwqxG6dFf
9coGAkBxJ3lxbewy/jGvnypaIscuQ3ZxjIZtfR+D7CTplNagZXfPlkQLp3j+ubSx
+ZZ2BG6TqiPpMPrgEBO1PtrtFzVQOdGnlfhxwdqUGFoZXLYk0Rre5cMuHFwPy1R4
f1ShDo57f0DPopl3NALrtf5YYtC8Dcu2MLOr6GLr3yaM3slBUaUjAoUj+xFhxOkl
CSMdBrg5rjFQiGp2qPPWinGTYeGHPbjiCTxpKWgkHZikouWvFift0Ta20XnSxEcY
H6kyO/LU3B9ijJKQi8dQRyQo8pv37AkGVx+bzH87+UzrYqq/EjDUAY94vIAZobia
Za7tLZyo0LPyN/sDDfQivZJ+wzpJJ39SzTwxVHZGN0BXNI9ARPCBsY4+oZhi7AKW
2hjvPYgRBiByWtiObjVvvelijFtJyWQNpJsXOdZgaNiHJn2Qg3lAWUkacrIzJB4r
o3s88UOYasWTiWGeoZjtpTKO3JOhvOD8+1DbnLlboH/cyhVHFxvo8x4goxY/DW70
6EyDbfRtoZ9BlQVWRfvA3sbNsSx+hvqo8cZMzYld98pgidhYq9TVZY7lbbK8wltL
60CsSssGbqIjqiW2nMKfxp/L7VHuET66hbRZ/9cC6HeyBUB/LNkugmXt4imqAvFZ
+cs6ZNYdiP1/+hwt7paJ6Ed7g4pUDdKDtqUhZkxm2ASMQMfxeOWvP0+fU3hwVeQ3
U1icoK8Sl9j9ABMmLWsrqsPQYNReix+fRkR6CndtoLLIBCHe0nmVv/E608q56Xn+
hHNbLIePc4BgSPTNt3Tj7XxKjLBShSnb/6SntJ6+TuRIl2PIiYi600/cO8O5jLqx
Hwl1odMiidQxrk21cJRU0MaQjCWi6JzzMvUysU31FC2TZ5zZtN14V2ZGdD0pLu5X
t9NCNGjLA5/0y/I+I/0a9EMJr80Q387mT5bPmT8vS8TVVp4OVQq3Iv7KYR7Pdtc6
REN6mldzWomM8tuRaByVnEvZ8jqQpNX/WFMwSNT7cel319mMWZaMq4HWJqiX0Oky
mXv+2DVbUwWJnmCWeXcssxeR5tYizZWos5hgqJLSql2dQ5SFNFzybCTps+7tLpV1
f9p+vpsJQVumb6BvZzthhxm5UhJ/vHfcf+7hN46pVlkrm6YZDK7F11fq7qqq+Cfv
x7nrGdZVmiE6N2HjPkHJ27mSopVWpg1Wexs2V8GeG7tiqAy/N8fQWSwW88AD3KbA
0ENXEp2U3tbKV6Uj8PPwLKXrqwCFnCNr+kgumIh3xKzK4BOQyduA+WrsZeWjmsTw
fPwZLXJc50j1CvpqyjpeRAIUjS1vxY0M868XDJ3aXmcFryRCTpiVPbcHr1cU8fsP
908jgWmCnExOzuDD0xMvI6hEiNVPLXpab1RXAm2BJXRCZ7zF4qDUXNKfC/+qadOD
Dz+RAYKSub+mTGPEqcedBpOk+SvqmdTJxv3WgledkgAUtmHYdeBh9JbNhPnw0TSE
5xBqma5YkAOcZafyYxnlYw4k42asZ2HKuZwR+vniI5m/NgfukdkZyCkYS94UC+Qm
iOsycIOP154F23Buw6ICIBWR+YatdpB6NhfPHjcMkTzjTpDSK1Z4QSMf9gB7Zsix
7b7DdGG0lcqM3ri4/8Pafd/oKnSqYwUEhFgvrDCCf00yQk5NWljrL9a8DxlNhhb4
45ReEph6rwhKG0F3d/KPKPO7X3zvJ61FwR7LBiyEiVrx63OGQncaD4NYNTfimvz4
w8rRYFBOfUeRnuB49/q9DBvkynCSHHtYloh6KKjaCGaZ7unCHX/RRFl2tK7R/Mse
y0lvpvh0RrVrfv9r1YTR3cOb2nkG63qcf6PhmJInc507+PhxMSWCU0mQbUplLxMr
kpx58xZ61zZZZpRyKshxd9DUIaJkzY6Gm9lkn+dyhVk/JSLwAJNue6mygLIpq7Bi
sojVqLu0voE0mhTgcsEP+8Ij14WUxbPYpOea1v5jnQ2r0idlZnArcNsJgv+KMBep
7I0WuCJE37sqdLELTn25XexxjZBlKhFfajI6S0l07yn3f2y2ozOHDnWFFWlFAV+g
hj4W2AIfNMjbeUfwxmuZ2qCVzBBhXsnyjeV1fEMZP+1pERd2lx+2ZtMTQzpUZJ28
Ksvbw7VuXSqPSqy33OlBi2rRIVSxVz5QZp4k3UwlDuU7OiTCBLG1xYwOcfghgcRZ
qGF7KpBfCSLJxniWuSNjXRy5k176nX3/OH0LwJ7XyFQol70dJ4QX4Vo71MCTgcOn
ovnEenySiqwJrYY0eSib6EIntWwl3UQuI6W6ttmTgK7naDsyfhK6kfuFWwwjQNAz
Bxw1Y1ZbdSB9buTluIUHy4Db0K9r6BSnyKRweAzSdb18Xc2wSa/wII9Z8i4fQPQA
Y7+1QPx7ypJkJz9GFFczgr8YZ0CpEwcE4OWlW/z4LgRnINXKc09/4rvdL3CwPDrh
Jq1jD6idrcmvlF97cFE2Na/pHGmrtSxbd9gARjfab5mYRa/ly7MLJvjvp2TtJucW
1amnb9TZN5Ffq5rSAHPPnMcQ2P0Txl6+N9eqtCY5W5s=
`pragma protect end_protected
