// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.0std
// ALTERA_TIMESTAMP:Wed Apr 26 13:33:38 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ENARmbOB3AY1b+WLAJkYrE62BDsLgy9VcTk5vd+WG6VNSbpLssLXCJYVcJYV9QeU
GjBOgRgNZhptOQ5z51j6/Cf2DGdQN0TuhGhv5y0S6yUDsY2K2p2uk2sOHpT3vmEk
8UsngGLeYWe4y+Kx/TC1q3nJ0ScC0UtwedB++IfP7I4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8400)
JVuUsx5G6zEd1l0+hCgKOpD4Uuf2J4J9fEOeud50R2zSNMlgZiT3X33sSJEepAr7
aUW1A0hWu7Ov9H2jhMx3vvjfzzxExiefi3ePj8/e4NP76WgflXdfbSV3UfnxRNRt
B2iaMMVKPTnDHL9PRDSyzJQbVfOM4x2QOCNqw0M2EEgDn5JhCyuv2FE8puPZzCyi
/CMlZ20kSfvkeapgqKaPEUjv4/pzhq0i+JXSvG78gnwWCsAYgORyPrnAsGrmvAVA
LQJmYbKMlUHxyPVCBxAXMWCgwYXw5tixnz9OOMv4gvl9DhEWmNHColZLpJYeW6lg
xw+zejZGX78CHeDZcLn0l6QxeqTSZoqpmHjlbV6fbI95m2z8M87pwk9WFks+5c4w
h2l31THMMXLhkk1ev2U2GnwOr0XiYI/8BohwKwmMznW1xAfA8oxXcCHZARGJmgGp
1ZC0xdt+oDN7oWPu6Sfa9Zg1AeSaxbtG+gMsg7Sau9w8SJerGDhWNqYcSuqPiKr3
T3MrjpkXBy5c8b8wb+a4Lnya7OjXqFzQLdbWDBYdx/d9b0vPlizxmSHEK7145R4O
wP8zAabEKWKV0MDo7B2k6Euff39f1cygcJho5hZXBqHdsaE7xdc3vYs1mhMfXzPz
Bw89LnNemEuxAyykR58+7ToSk8MWxQF8H4bx1JjhflLVLVL/ugq6C7HT9dNVaGGr
TId4/i3RRPNzo7OXf93/PKEcg4jBhIweZDYTMpDgmkSu69d6P+lEb1WP1Df9uE8Z
XKTAxLFiGDya9S4oUbeNKuNOk1Cc+bRgwi1FzFEN+1vMXTQNzlLQ6w/tLKbv9sqd
U4ylj0vTwzvibLMpCmAd+RXpLpgTtvkT5L9rXSfOqmud/jbGoItZZYkUsFkHvAuv
o3pHAJ+hDD4iReybvujqtBV+pQ22oO1UmFSwsUZnPHS6ix14LbGDcjh6zsbM1qox
wJ7JAReFnBuylWsLhRYVsA01oZOoBVMfslMve4iIojzE60UKyJm5+csOa7Wnf5uw
GIWHjXWQQd65uH8oalBzMwHNN1yFvxLoIbFxmDuwNNxuCh/pEHre9Wpf0DN5GhDx
wVdNMX730kG8we8v4htIdooenRg1KV4eXFZcyCYhc4/sPpIwoJ1a7coLn8ofly/O
ZmMw04RqH19npnzIPfKYOwqwxvBOZSJSwJq/8i4iVTRqKCus9SfHN6ythA+WwhTK
0GYUjqa9PRgy2qjBf6oHVltDNlf+yIB8q31FyBFYcLbPJe7XaDOsPebK3QjGsvfF
DKqLlRaXQz2GMo6fEbWkrQ0wYdCfsAqUMjCG6Mv0fMHtDLWyxydNmYgSwJJMMzY7
xuL8/Tf83EoOlP1SmQ/LkNNGyPCDL0j89sdW1HYEovOO6UO3DW2pDKjafzL8e4P+
EADVy/eOp7bDHtA3qTvCsbWfrJWBPAtJL1dA2UXtimg257vTFXyh39K8qu0WqwdT
BcoTH9g7DS/2qNSzDYXn/KK/MeGCC4BGfBh8U2AaND8ZrOw2dota71tqJ00v2Fmm
oGZ8cul8vbcswjksPdchcWDqxmnNoJPxVa3TTd/qWL7jvkDkMuJOf5h8ZL3nwzZ5
ie1E9j1LQPiuUKV4TKUwwa9iI+yy6HkLgn+sxu50TqLy0y9Fh+AgxYQJCnrLShUa
OHTo4AFJN6dB0kInFD0qS7rBWk9ztIepj+n9/zvQ0+jBghvQlUjVzoHZMr0phiqh
4SYQ23jy4QuRPx68CwqFeBfjf62btwI7E0uJbvSiwn06cn+Tsoqyf5FcoIFp0fLI
4aIXmlqPvJT8eirCgs68M4YwOnvpUu+O1s5DkpZOxcQX/swuZDKhaQmJ9YuJp/el
E6T2SVrxsr40dXzWRMRlgA4VMYFF4fsq9kyhoYEfBPO+tSvAzirYQJnQamijDMF2
AjSltY8sf6iBQsTCK4HabhlHW/DiXvsA/cUWOfTmiUI058TFxj4vHDeir0MLEOBY
6gIC+H1MiJDVyYo4d/Dx83hirnLS9yZEqJ+J0nLMtQVkutvDrVUXM9cghtVHNnCZ
XITOaRyG9rj+ULNK1q3CAbw1s2m9brkXbcgdVQGz2m9Gfoilw0mbKZSi1QRbxLoz
eZ3g0uOVTYR/GU1J4VkOvMnjXhtUW0tbVojANoAG6NM6cBqLpH7WjLnUb5CKOohJ
lPMg3ZEx+pG+DaZmIFsTJMmRFMM1TI7sOsmeVoMtaqBugj0RLNsbtSUvPBCV4vZI
SJfgI3S9+QCd8YEdc8LJgG67yaiL7iPUo1CeZzQHoDtyKZw2aVDvSkPiYIIDDZd9
jCAFcpo61bFwCuMCHRQCcO15G/qXNG1Y/IZ6VxiB9+KgdbqMUxwzMTE0r3AJ3prF
HAK00sPakbE6L2D7S3IebmcYCT/VO6Urf/ERo2EPt4zQtW76yZi2fJcIIdtsR++C
N13iKlUl9a6aJzrRwk9CAWy9FdDesUVB0pjVuMqYIISm23OkfsCKxSRURFebOC/v
ByXcZUF95egIYXwkXH/tB1N3AyFPPzA4M+jdSIjv2lNjpkzA0Tw8gB7Cl4Au2UYv
/Ze8nPniTERULFrzIXXOMP99aYcUwJb7EyQklL/zYb+Ex2auxmqfkMg736GIrKCR
rcUu/Zm8sFjRYsvaEAE0b1MWwOHoqylUVFsy93gd35DOpoTwcQi4bijvmzEHGWDk
XqcYXuHRtFWSUJY424G12exDl6s64kokt6YAlKL1ahP0tepZkw6QacR8P/b3rkLe
Tx6fsVcFdgGzR/sKVD610xTEhl7mlOlcSEOy2a4vfrxsQUmcfw+4YGLSheLtU9dp
7VS/t8oqFn+TGuFNqCmE7wy0atnEjw26dm7COriHwVh/pozR1L0ujBYwMnUVfDQ6
5ssP6P59AWVFhvVLC3AFigMuuOnPmOb1TvJDNYwpIXVP3KuN/yL/O7uqtaco/Mhc
b+RfDusojvkuAfb2/L/T9I+fUX6TUxIwCyrOzswrwnS4gtzyhyu4rOM499cet8pt
qx5Td5CFvmqY0AZNc1CHaE2jt+CQs5+OC4ttulJuEjLFngltVhlqPrloPLWrLxsN
m2rInLiS17Lt5lmd2R3Nr3mBGkgz8rxn96UYX3X79aWzaNTbJoJndaz6yo9qzU6n
NghFtn5rbjKjmONSuEWcwmmV5jlZpLJCezgSwOUfub/bHth1/Zc8qB1wu6e4x/HF
95QHRFfA0PjRhzWD5mDo85xR32YE3Uynec3NjjbbLnVeck6IgJSh+pnkJQxfy0Ul
LLFFekdigDP6UfHOAQrWK0AOOuzQ4Sm5aWVqBz3E4Ip60FV1NLX7Z/RZtKEoY3BY
bw6gYlBmqtad7Ytgor0y0KAJyhZqTkDRq9fiTZZnAMQpzqC1gyKLd+QrjFSgx7ng
z4WNGPVE+m3oKjuZzFBOxVmIVVPIZDoWGwSZ1lXdd2AdeHifqgaxHSX2oc4HqIiM
TY5xPtmY/P4uJ+FFNvMhWXO0YA3cWJHFtsDSI/o9Q5fTxZdlBTQUBee4hR9T0u+G
q4GT7Fywbk4PHYaRD/FWL1Q7yMRqPWbIDaD6KfE/IgLr48JQ4zzx7XSaTXvS5NCH
fdhmbvTWEGnzy0eABRUNeqmnbGJOAv1yGMFjK4TUcaLDkVeTzN8K6f4irZ7PrlKw
TGz2y8UB9nw5HAMFpIV9wS6kJLnES/rkvakpfvsaLXESSW2KXbTWN/AN8E+ALFrf
/f3+BpZqfOXLBNGeMn/CrYYZdWjk/vhAhC850XhlkXvSfQstySem+wQbfN66Qgom
tWSk2RLxRV/cI4LZs7mAxD464y7o/ZEVU9yLyrsELvGP6CkcvTCgOv+a2nB6iz/j
/dtr/16pvbCKbbaJZECbYofpPLmmkV58HjavkU5Ew0mhekFvOGB3Uco/EYZS9QFs
v6eTbPCn1REiSQb8IQ91FK2U9co+lIBdwavXBwKcW+2zA5ei41HuIdfgzZXof/Jm
6uPqqM0tVsd6wLFnJuCVe+3Cf59xkAnfb6mOcF3xwoa1RHMJw/Io1b80qMfvvvHY
N3tytQwHaTJ5ZGazXH4niE8y6gKh7pkLgRKlyvIujR5XvgVDF93OVGNWStKTV3Kf
/rK1ScCwVTaMSt0n98RGnCaWEiFiFKK/aoPm09Pqn9gyIEu21YOFaShM+KDMZ6Ql
vP3roKC9ESZmmwehgBTyAaEFhQoBr9iTbKpX/gA27ALDtCGAowk9CM3HUDrYTRqZ
GXULGXFAulF2+GvX1wlFdldXH4UTQSCEFQxJYB+lZ/svCCGXOtvY4Due2AkausGk
+LqU24w32OTTObC9hUQ+uisk+UphfqgSLzpd0sh4xbWlvTVSLsucqr+rw7UporM7
e+w5ThBmqtbQ3XmyKJ7orsvnRqHf95NOeY84fUoH4cMHUKWOxNSxWSO4ykpAgrxT
9LJy/IhV3P2VlU+Fod/OltRPe/nyDirEz8k9vx5BddotEPgREhMGmIvrRA2IRzn9
uSQ9LRmkdrY8kilgRHBsXo1NBu+b+8GkdWLleNwUm908zcahsFyM5GDEbyfvU2cN
5n5Wp0daqm9s48PBF0LCf11B2Kg2LgVy6vE+aos6zvkuBTCwetxjSRDQHrMAeTU0
uwRM78plt7F/XWZfg+NKKcxpYbek+zZIFs2ze4MoVrcZmxMHknzCrZnIb1OtcL26
VAons8obcTXrYP/NATTgmAyrz2UY9KStmxufbMqjbqPqWoaBwH2b1TJT/MaMAnBO
YM2ks1NkDt24c9bQaThGCv57etnvMOjZJhouewrOSsv/rf5oDxY4YZTl32OPDRIa
sj92A3CORAtqp8Jg9imDw1DdNtm1T1S0SHieEud9SseerVP2civFPM7X0yt0fHRW
BmFvZs4YukKc65lFV35e9ckFC7FkV5nunXhxz5tL2lLWeotmoTb0tU45WXdJjYkv
Zl04oKthY+9YqTRBl8fxXVtUuG9bFEkyhMZDUeyID4Onjsyn6q0XY8pi7LMQTYIx
TLxmhCekhYRCB0W3EHNZdrQqd8MKqQP0sBSLyDn/J4bkZzyJOk2SCaXLi8BurI2Z
HhRgsA+bwYOtYEb2T0aa0BLiEj+0CIx2nTvEUm1q1J6HeN4kWn9HelCtPB1ayJMz
Oxza7dLuemJ/gApxC3oR39ZokkR/qdBnNNpWGcuLBN43H53B9idSvCsm5yx1Krb9
9A3HN7n6dkHPY+TKHOJr/gC6RVL63Y2JklkOPp1bvWAQUmC0mJ0ggNqLgCvVPR3T
KtLtpxE4tgXEUgZ36VOVjzB+IK18bflPy7w/2IzsL53h1e+qvZqZ12uKyB0iGqS8
gcCErOuD3Vx6Kf2ei9weSf4AnWub+NLnhOyCdCSHVzBEBBGMhmqHQcliGAxha8Q3
7E1UJD9CmdRBb97Gb+PO3egYoYNGFcyM8ThtCQPjyUmlQ5yWRq5F2Ommd/OK8O8o
pcijm1u6qr0pxpbAtwDvwNpAvGZ/DdewCFCp39otUPcdjhpqt08AlfehHE9ckMbR
OoaJlkd0wdaZHi5SUM1jlHI48sVs4klBDnoiNFtJGB2+UoZj1+6/obGgB6yu//Va
XpLvFyLIIBmhrLCl03cJlSwePKvEubmJuhcn4nbSjYe+Iu4XqvxEs7wFbLPZn3Bs
4igK2i+gE4vrqpfKP5Z+dsZkATpZx+TLPtSa3dpkZhp1JobMmeK/Qozx26QKzxgp
wcUAJT52jgJJPjchNh/BsuGHbrE8ssPuieuj2aWF9lNY9MycQ/Kn6s/uP80thsF8
gILmjXrMcTRuM2eXRLRm1UVA2sLPjuXhY7dHWNyfg2RPMldZr0Oe+4Z0rLaVg8jZ
0HkA7iuJSMbyRHctfSa9KubJFttTQliQTc5iawitIAIIV8HoyFO8YiVmVSZHrjW+
HNeUw1IBpO80Sz+YjEW+KGnTNMCekI8WFzu4StPGO1K9SjfrYoly69V6jQ3w82p5
Fu5iYqTZsM3uGmDKJY43Y5rPOkjHEf6OpomLDyzsDkIOo15mxPaF9FCxYV0lP3kD
hBAYnDBqE7n3p9YqqXC2amopUaBddx9tZHqWGqRfRWmdoh7CuTeG0hwWLCeisxrJ
xg/jc3rlX7qzgykEsi8ZNdj2YI49Le/USGGdUlsFgyto4i5ShSDpk9jNYVPkVgBg
quY9LMRd2KKlMzwbO4FwPS7sr6f4HOVqLnQ498+pzg+/Ss/BSeokzA4pqBc/yyh+
NXdSdrr7bVQx3/owZwg5s9JH1bMoS5IWEl0POxNluB9GRI/tEZ/JFrSB4UqbBFVJ
LZzfsslUmGOLfBtJrvphCk4/RadJL0CnnEIK2xLWHR/ThW9ObbScWIDPT9v6Qi+1
kI80pGyeLSsvVg9NTgYgM6IwvFpF/2SU2C/gstn4zL2vZw7n9phSBXDsTXjrUydJ
/V6g9zNzn0jD+QtcWh1gsRhqHT3Xe7/yA/W6LKZdbCkzj7CSbdU/NJ5lqYvowePP
a53taxyl+nmppb7UgfF4xzx1P2V6PvCo4mkIRe7/eXFM/vu6TrFLkIx264CyrAPB
uy+ImzeKCF5ejMLgxmKIlPhYTdNDhaw3AmQaK06I8teW5fhXaMfhhyndQhQ212gG
l6DXe/pjm9cTDgWIZMiyTItm6WmgSkE7mMmenFHD1nuHUzSG/FUJ44Jn7RViG8f4
sTJ6u5BXChKcyhyx7K0kDS4AQDFWZfxKbXilLwdUH3jeTSiAlPBYz2/6/o4HC/Og
vAx4ekSKvvF8QxeOtNpaCIeq1qWGxBTH0Xb1BOEFNO+0MG03tqjXBQaw7Z8Cg1Hl
N9Pgrg79h4qFy+E0hScQ0Au65zsnVxaXFBtGSFmPDnRiPhk1aAyKGLZLa/VBWM/L
Z8gi7k/sUCPI9dVHqjBT71MPbnpZJi50xKwppOFGdRnlU7Dl24bztR4Jm6TcTV/C
xAKLX4Ya0f+9tSwyxzfoTer3JrXOWwbBtBiDzd4+0HWUqZLegoytQ3Hj6h6GjdBM
lhZdMM9Wh3IgqRlnub+mj92TdosElgjsmduKwBR/zu96upUud9A5fkk5hcMSy1WH
nSHi+jp2QkWBlmT0ej2LUToIaNRznEsqNp6T4R0h7KovehTFMbIa1SD0wJTGUCc6
IAZzId2C8BkkOSly/bGMyQEGblTJg3ob5T/Ge9mn4nIhx+my6lXsoqPPE41HiSZc
NbcQaUKDrW5f9weYefE9oqeZhVl5/DBxO+wF44v8z8kA3h+QJtIm2vD4lfkQ2JtU
jHxSzd5h4+dnoPTr4VqLRhI6CrBAOdZ9R3bJsZo31Ugs9X66hlwfI6bZSp3t3BYB
TwIS9Oz+8mskUGq5kajjLgdxg21BsCHjGtyehcujFyEYgxE+xljC489voOXS1EH7
2l3qQXkR7YFQqvkBVD45d8ey6ZpqYSno4YLsRQvl8Nx/SJocD7O2imZGPqrFZgkk
E/4SiIwxyc2m8nll7KUwrybPY9hIQph5Z/aXfGp4zXIxQCQVc8RY+ALUn0pA5rCm
iBrAK/Wi5kx+y6gelGhIWd3Y0tDw26XIBmX2ulS/Q1axOIM0lYlc9N7x30vjJA4M
zHSPq5DoM+EpZTJhdElCTWdchgHUHAj1jeKDxPkpd9VZsjHr7XYgzB3fuJFg485Q
BILclA4WziRUz/fbXhjZHc8CwO/qOWKRsKswOEz7St6ECRSCbyOS3aH9qlnANwJq
zyLDXC/WXg/jKuVtCxOMBLH+zdPB41aM1A44VJZzgUK+cHcoM3KwuLbCwNFZe/mj
CUqb8sOEaopO8Jj5NfafB5Mc9RP9Lcpy++Tz58FZBmivHAEW8fKWSIWj6lRJQFez
QntIq8J0KTcq42lmPrJVFI6oE7U6eZsriMMdRFtRfwubjxLyRiavoGvt/drKShaz
76LKAlfaKoHDjwenGG3dr53sF6aYmSJPzS1iFewFCu3VXjy+EPzEVYTJiJTK9FqQ
bDb2zhfjF0zNGDjrm+RNuMzVkgr+9jj/2N6XBzsFBZFQYOqYmGT9EV+SyFOSld2F
DlMnAbbCMQSAKzIgP1FpdSmmAtlIynCQWPHEeLRVDvhgPjelhvn0aztvcdikCeR+
9fCz1xa1D2kWjl+6DW2/JXPi5nc7iMBMTi4N3W8HKSbT8HDDnh424kUd1Rxqo62n
VnzsLG3Ir2JXnvOTu1LGbTyeP5CBeEeDf2kCoWZzJG6nr+V2rD1rK5RSHRuGB4r9
Sp+BixVVTGUVE/bkUi90GhTNx5jSPLBxoVlv2VHj3+qcj3xvYJeEhqWKAARWA4gR
Iam67hZ6pxuGHMhI/ge65XWTd7YT6+WRRwXwLPaSSKe49XlcXMjV80FGxoWs4dF/
c2A17DzXmA5sz+tZbkJHTcflIcS8braSAtRLj03xHoBGNG/LKEGDrIy/5lEFR/3p
jbS92WOSkgoacgKyMRP0uZIVv3noiTP2sgQiWslpAXdGIUrBnzMgP1BhLl7WNLXr
yt+eg6GIvaHbbw+DP/YUQfB2fJjJfju11zo8/QyIcX6mOnuFc5rlA60zfINcx6ei
WnjxWgDri0wDeHzRpMXzqAhG8Ebu5qZua9XzXtCIQZJiEUaofeSspfH6LebA8gSk
LLh20zqIeNPGsxJfpMlCbTwy+ATthcJ4aTP8ymgyF6u/lSXsj3q3H+LO+ERjYk1p
KYGbxGR0J23w93PWu3ueTaIeZ23zuFVQ+FWYUE2GeEi3SQafnhw1Nqw6cNTz4Pw0
FNg/LuuXMVvl8yN9iKdXPVBUDHyJI4rHHMM88z2X3F0p1oojF8NyuPNLY+/NHRIU
qKyGelJi8w5dJK4z39bYnk4O7MaGN8XVsCmMvITvnUKZasyjYqbnJW+xWPrb6C5i
sVN2NUb+3X7m2BLQwd/iw5rY/wltn7epZAiL8K1QO3Vu4rJg5/PfXhQG9wSUjmpd
XRXmEUkeNZDGW/GWvpeX1/Q/bUAHiODvkvuAa5eu5EiRkrmS1tY0A1pzOWQtstQ+
2bwUZh1ZHyV4R4h14uiZ/MRwxZtqwmnR5JykOICTjS7JRGgCa3O/5p563DjiHQAz
yDuGP564G5TSoa7WSWdlndI/lIXqztbe+5A5NGU+EK8SKl8QN5Y/0hIweXC+UW1H
c3wuZaM9nFMw1mRsXvYlwplo6jTyPSTj96FSK4YtX5KOR4Sgm/VrhjNJ0oliO3lK
eYXj2CO9UnWxU2nFv8QWQJXw8REaKf2cvD7VydyErvaQTYdjjYpQxsko+C1s/MvH
9AuAc5b2Az3QbiLLyRVrtkEDV//za82TaYCS6n82JV1jkWtMVa2JTy6Dl0v3uweE
CJ1QBDPsdO41CxhPjEDANwy0ZAt/VmdQcolIisNWrtY2kwPSN6XDz5VgDePZiIWJ
fhc8FJDfcv3g/paezL82SAqexR06kvpLS6bCcJ+4qk4LvaU5EChk32rRfNrVgAYp
g5K904w42h3MbIlRt/1fqu2990yVib8Pd2GVKLX5zUiv0Lc9LZLCLXxbVU5AUBbf
X/P9jxCRIY65dV2shZV2s6LrSoSWf/K03vpIi1g6jcYfSli5yo8+2/iQ+BwhuC1u
TbusfdeDZ+XveOL4cgD5hRVNMVvT4DE+xB/5Z2Q5TaepoiSVHIu7dq82i4kV8FY/
4VyTeTLXH9xHjQ6zTh7elE0c8D1ooL1VL1V9mi7EFsewXvjfBABqrItI5KFB3dVd
YmoYdQuHl7xubXILuTow3Tywt+g8W8rRhSVB2EuMOAst3x2CjUFRrCOjVVjVnG+M
+5z/DdnwFBk4XwOsCyiBTxCYKKr7+MTB05k8tIZeNrC50rsMOo9mSc+K2ej/POTh
SpKCTuZZZnmYGqhUkNkPhLN7iJ0j/JahU5cb60gzpM/N5sG+ZKTVTEIq9OSwyYbm
nMj1Zr4r1nxpkxCRggl3j6Unjp2rV3UOBP7V4cB2eTC3GyJuA44vWgN6DRYhN3UU
UuZiAW6QLxJc6kl894dnlI2ff2a6yIIJhBA9degGJqjf8HxSjfjPd10awlpGr7rQ
lXilbGHKvcSDAx8GkU7/5yJSbFOjaPWOj1cV+cikjxzV6i5XBwYqpu17ipvnsaT+
USJ9Qm2vI+nu0WP2XMGVHYEDKYyJyLyg2EbsYwbVvHRMHHJV9xn7Vg48oVIsILWZ
TWiJaaOLwIvMQu2R5C5ese4SUADUGyeoTRzrsmZDOC6nfyhLvYIHN8C5mIWAbc5B
bAgGAGFWazTPWDPsWxQjBJpMdrpGdXp/UCHGqXadgbSXQXsya589lMN2xDRYYy8W
7Ea+jhQ35/gub60npW41M1Yi71dJxiZx/kfwf95CFqXLhfn5teZpCkUbLLi4MpV5
ztIogRw/OaPGg5ZJI9mgVg4gGjtkeysg8oieP/uubWyzU4jwoxaxXnhlVTTZFCSB
+ZAO4V1mJBZ4blk4L2z7w+g6JOAYGi+JSSyCCR1M1sfs+AMrMH5kAC5SE+5nLz2Y
NUBCjansGX5jp2m0Zj9i/B9oRJaDWPOJTzdHZfwu9PIlLrrFPA70TwOnkRmP949O
jZ2PNYwQgFFqCJzcf9dJBfBvtFWY4DlrsPfy62VvEfdV0gaQMSqXHUlroExGBETV
PMw8z5fzvTaRcCUic4kBczjHfTGCi0doBbaHzXAgaHCRGSldez5iAKRkTxoSw/WG
csOnI4K0r3yKOGWKimqltmI3FLbaWLXPzaA4Ienh/jGBp6xV5lcN+B/AOBnWLY1s
hOWBNRapZuAn/BbP82j80KDJ838wvAtrO2xLPfGFHh9XsHyEHeY88hOTNz6uxylE
JcNfNAP4hLKB4u3C29tjHmkRiNXBU8ITOdI0gvHljapWCI3MM2esZKcNgYtPrrjy
K7I+Ku10zIoDNY9bnLwfjK+JcBWomSn330xxIqUWQ8PDy2+6Oj3XWwpI0tOPs/0N
0X09/BorXMYbZah0IbdMAdl1MFiCUUVn41XgSVMjqh2GH3e9k7v0rjVXl0b2XKfA
k7O6ZJrefCOAio70r0NLLuWvHl0hJMLD9DInq/cbvz/4DBmLEE9bLxnuWGF1ziWx
ut/l/CS+RfkBZRRanGS+mp/+N4MtHb2qA0+/MMhvc6gh/ji0XJmOQZZXjJuHUL2n
NrTUtFLiIv0ap6D+yrTw7M2ptSPOSYWGqAsKuvYwq2zVEVOSX+3oUb1RPBawKUP1
b+9n+gBlJF1sv9tZCFo/lIwNzmo9KWsiI/VGOepKYV+SydETD67L2Yz30T71yvv+
`pragma protect end_protected
