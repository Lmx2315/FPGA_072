// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.0std
// ALTERA_TIMESTAMP:Wed Apr 26 13:33:37 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
giqFv23cwi1kI+CyS0MYqUo6i5gqSmmLvjbh2nJDpFD21uY2DB64pX6BmWMvXFQX
zWj8VG1YAiDbXZDzbZGZKe8gzaV41SVaVrHIV/Vrn5H4yhYoqUcaKclSy6rG7JTn
cCg9iYO2r5tzoMe4k6UEifqdBBlWt6xxal5cfZbC1Lo=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 71104)
tPImr9IP8OE/n2jtZCApmlHe6z4/221HtHELfwjX42l+Uc1txEJwLi/+Hvr6vIB2
lw177QBpAmBPm7TXCXc3KDYy1HBPKtwU8JKBV12tbRgSDcwxD79pR6U6NbMxA4gx
How5nu/45k9HogqL2PXv9x3yTj5QGMZSKX9UgD7CgpVn2804ka+j/xwJUlnxibwG
vpPCQcgmvDdO0urywIR7QnY2BJuhp050yIPuZ971LflOyIIEN+ssbCLQbCatRR1V
1XJ2cnGcOTHIGahjFHwqS1qkvgrX2J8RPE9dBfZndj/W82LDeLhI9AwzvkgS/Rkn
MXaT4ESObdYjl0Oo4oCvX/e0aYfN+P4UJglbsBLqPST04XZTzFKdsDqc6DrOuhSH
unK9nwR1zBhFtPw63Rpp7lru/y6CNnRduX9sGA9GZaPy9dmQvK3aFc2vxyMoUeOA
/OGa9RxP7PqcT5CrSDxO3awQsCkUgPkozck5Toj1rBwce+OMJwLNaXcpPKMm2UKe
dTxQ0/NQgzXlXFnafXD0SU0WEwc1jw1PdUz4iE8c/HduEbemklEn8TFyFW13tBhY
C15h45Mn4JjHQ32gLFE5nIuSvSELNyRVFXNwci+SgRLPs6/uHnB5d61bcJRPPHr7
ccnxIV2VCFt3Uz2TddCxWtkRqg87fUGCGJkQkBI9i8iwIbHXrxzFvxy1b2X4IvC5
re+D+nLKchkR3SU5hMB8fgS7832PJZvTzXwCto0AE2TertX9aTd5C3KNiNdwjz49
KY5ZesfKT7wmZ7q4Ft5JWWSt2kJEgol5zQ1KYPTEryGPZO5sWCdv78aPtAvWmJaK
B7Amm4V21kxwDcQx//3WdHCxCc3MiXuAO6RRNdlnNO22lK0FKO4bex5I17Qv/8ns
pEPL12cp9iCJtZ8bRLuV2oh3wL3uiRWnbpoy0eulj1dQ9/R+VOlvsUNSv4g+3RYs
Gjlv7hItJ+rQSkCGP4JMhvyRME/NLQwIK7ROr5kT+9iGB/K5MKfrn1ud1MVMcOtz
OYVCRRbgWkSFjWFBvQw2xbORIn0szOHtzDHDoSzttc3zjIfzfTuze4OKnw6M04MQ
kAcsucqtUFUIb5G6sYD+SRWJh+mMPKhY0B9kA0jSVvZ4JUj/F6Mwk31UQRyYcCfj
8Fis3g7PoMi1PEA8ZTobBvGry+waOBCMFSH9LN+MDzpvUdnQRLCPW7iE63/MG++t
oxLGnGnJ20wbgMVfTcLcDMCTingHks7AhTMwgeU1sD5rM9jZZyw5a3vqGe5zydAH
aByFPu4D+k5E7Yf+aE95hKaqRNgsusjXkb2lCbJRUFIua9CdnHS5ILJ99+xYWlax
tXrhuUMKo1KJXgXmTcntP+9kpRVW4gvEr3x1pb4otoqe+5ag6YVo502KQ+BZBo1i
TkC6fWMzVEi4EMnFbuOar6gdl6r074p+tsMPXklKpQRgYDnYN2Eo5aHutIhBcg4y
aQvIFN3dX41V1nARaVzRgb0MElgjuynydE09UaMLKC0hN0rYN8NVN06A9CpQ6ExY
Y3rwCk/2ogRFF+0jPzqP+8+N5R/xmaWiiIPKJsrf982rzq5+YaCC02/QQ59Fq1tQ
494FnIeZYcTUgnnkoTEYMuzKdAqY9DIe4uV2gtGyi87rVRlTuhwKSxLFe6t15iFk
ipT4EWc/TmgtdL6jnnm5cIJChgOGohJElYjQIScoHRCjqfceUnmhO6uwW+jpRTgf
YygLiAoKKSizvap/XmcYAFecjzYJm/WxpRzIqaALYb07jV+3SUvHsLKxm3Bf1mcd
zdbLQg3ojPOCWMo6wO2pJueRGZvxWNMAfjBk5rw3f2krCjU7au5fyPhEBiziSQ+3
vPyYAy0T6EAETttD07EbfPBdPwGSGF2UHfGN59hYTNG3F8DW65LF4MWj0/Ax5hwv
2BtHU6JgTPySHNvjGHWmwKX4cYSMnf4Bls9hy2pvLlmEFg53DCAZRmEAuc9Y5IJj
rBU13lmFk29ByrJ4SPi31/CTHhmkD+OEtAAVrbGTV0sR2fuLULClJ0FhYfP+XJtK
gExRkN42VlhLfb0492os9IPT42lqDALbAX7CLaf9C11C2QgZJbAVjSAEcsR56lnH
rxvJhAH1DCbKr37NDZXOXzcDw5JWG8yR466AQ+Fo2Uy+u1w1+Jo+GhQlqS5vEepO
Ll+pOAlRmY+rU05+6X6uFlq8CP5WdNZpaqdp7XQt00loy+spPC99wOsCCy2A2vwE
1nLtcwPXoaZWMQdoKViYrLSWJiqGNmSV95zb6BMijIloPjV4kPHjH9/UlvNolJqz
EhDhTlB8y4uSLx/LeG+OWRSH1YX9xzr6cX8y2CbHbPkCu6B50AiIn4LFkEAz9qoV
idT860V21EAFX/jXgF4b5bEuhErDcYoaCMF0ka/lqYEjt+KEKo9uB2XxFtrF5jAx
NZoVzU8un2Xbk+Cx70QtWAMgcZjsfoj+Adqqo9bFaRbdN0Lx3/dG4F1Tum+WJEeI
wlvBwNFWqJlI4yhVs0APu9S22FD4fQdFlwRPa/yaaP8bOWuGvFCEj6V2Ky+WBy0r
uz7LRHMUalK9t9V48bWfOZ6o7S08imBHaXWbeV3nkf/Ywsdn0rM4q6LsbHWGfjc3
DOcXYPv+9pFNQsQta3wbMPootvXAuxjm1YmeEhWyUbHR4PgjA8hvUV30C+aiGH1p
pyTWxgcgGXnIs8G6pFGIv2ArZ3KVMakAn6SM4TNqI49E4AwauXz40IHKeUlrWR8a
PUaP5NYmG5aRKW8QDfvIvHsAo97brGYRs1e3p5/F/8ReaewNywREtgwWbbQTsoRU
ZE8t9rsmE63Tg/APZjF5xt1WXLWVTQP7iuFEbEAzCdZKaDOtRGyhhPX6JrGFz14e
2QdXs+pBZ01sO2+564qRch5+1crt4g3jokmdlLfKo1gqv+VnP5zRJRF4QIm4GB6n
hew6cSRMfvvLdR24m4jwipiKZbkdaL4CIVVJ/slkgwlXDmxw0Y9CE9DXMMBg/38i
ddQUJ1H0v96PPyEBPVIDxoI2YoW22Ujav7svniNfHQg/naCEUw12+hepzYZM2GAF
x5XK6qodz/O6s7XxKtp27vkZddkwdISal9CIubCYyRZdVH5Toy7TusZaD5tm575Y
vJLXtGy5t43syxU2nDxNloDzTwU+/CN5K6ss6TwoToIBv7Wa68HBiOhZcTBqy/so
F0UD56cIh6SvgBUHOID2b9R5oYK7yAP3ItKb4mer8XzK6X3msDqBXBqwFbOoxW9b
9h9HCHHaFLEQB7fbuflpzaaUoOJR/ZgrmMdJHsqULOqGNpp74F8FmQzP5QKbvqzO
DrtycUKR3qDJEKrYDw92/0bjugfHeJOr2E3D0HfU21qVoWRtMabWFyTF/Aoa8FKO
PU1HPmFoY4dHrMQ2mFz5GpyZy4g6q0w8ijM8acQzqd+E+4+8V9k9OFCiGu3IW6ok
IHqgLrRv6iz+caikkDKH9ZEJkuwTGSlMl6UpkfNxHZB2E/igXMkzKZ83WsIO38/l
nBcal6gTAMy4vXHj7IhJzLi1yrmQ339ty7YMmAeyJs5rSPnAkqd8x9iuqH77i7tp
uU+dMGgAYHvrAfNIXO/imM5UTqHj2PgvkrxHIWCY6J+QJOG90VzFLqVhOr1ISwHi
bTjOpNfZQKzarcLhSrBz9VcTF/5tYishNF+FiQqE2X+Y5G4MaRJORyFvFGOqmDqB
zHmDalyg9l/pw+PPgdW19GA20DoxhVyIjUJ9Mele/DqcbgGd1dBJ4jBD2dD8Jep3
2JUK0Urv5CnPxme3KIynN3QX7JxP8in7ZmB+ZV2vCZ0tzF9NzFp5ar8vC1rRD0vx
p1RPe2u65sYKkaY8K8rzuQBT1vmFPxbPGlUXXupYtWn0Mh7nLS86S2jJ2Mw0X581
QUAdyFVet6JlmxQelhsPfD3ULG+64znRFJBoRyj+i9EUuJU1ONB6tRgzt1/VR8oR
4rCvuLwGnRMcrx+MAqMNDJlKhvihI3kbWRlDuh8mHP4X2mTy2HlVzPpDjUoOO3BD
2tLvCz2IdzTUjXxB1F7deASXkrpcMCkjuyZsex3z+l67LA9Y7SygX0lQYk4n2Y16
9XlOQi+usCE3mPGtEPnJzoq1dLb6zeBbaMv+kwXcthF5pKSLf/QF1OkD00fCOjI2
R5pH7nGx4oLtpaTBmjW14NUcvERpLh0QE7lzhTEKBi8vB1zM8MBhLqrR5NnuUjgD
uCs9siS/lVR4hGqUF+eCMrlhhfCPxe0RQFSNk4Hl8KpRHylmSnL14UmALSHVBX+u
b2tLRlW7kblgmykmPxyT1lWCSNCJNI43Ka3ZHy+ZlfTXOUrvrJFtQWeyM2SyRCYP
4uCX5Tee1e+5tQ7L5XeU51Sv5lq1Jh68y9yA253sAGpO5dMeByx8acuoUveeAfuO
aeT5s6xwkSvCdO0d51jpxFvz7rTHV8SI8+M7ipkJubj855p/t1QlCuMmFNneDki9
ZBfTePDXvVMkft/8oOEuA9GAzFm9kvN8cgfEHeOv8bZvN98T7o9M62bJOOzm8imd
5cuprQA28zPZclQym19wVctDQr8Rzc7j84spOkjRJuiF95kjwxI3dwedQxNb7Hun
mtJHdxZRiCLIBT2LZ9O3Nidqz/p6Yi2C6Ucapc8QAaYbZ0xnT3j98tkiLo92Zf7s
IM4abfqeORySPA2z0j2RBzKw/qWj05kVmDs+WhYMDT/NWR/D4m/UHz14tF6+EU8o
ND7AC8hOZz5A+l7rn6hzave5RanSnSNEpD1yTrW3a0fOWso+xG8d17k1caGz6mQ3
HJ6GBu30UiLjRNcsSZ2qEGOZuBKdkgbB/9VBYnBHm/sqCViM9vNmrbgFrK/Nyywc
6opcrbYDv0PQjfM63xDweQE6Y+nPEtbMWqLQgak/A/ajIbXRORxffaTur236t4Uv
dTFlgJBN69bqU9jjdz07xQ0fZ135i3+kP2x4JE2nY/uzPP7oT7aW4TTvFtPxikZ2
pazZkY4dH8YH/3G40o/zBLgas62X4+rMqU+sSoQ2oo0VsS8e/iCnoLeujg55I79X
XqOJhwhhFboxI9B2FkgRWORV98x2trqJsUwaJF/v3WOVyVRQe0sFm/vuFXjXEIaO
AUbQf9w6mkf9n8+PZFUU7vgei7L1iKQrIC+lS5sz80L4CDkUTHWLsAx3TI6Q7WdR
fkIb+4CRAj7bi2WkleZBLNoETmOZxVve+ca3wiIYFwaL64mpy7jVqzbLXt4+tBNU
DiV25J6KbqWFE/pZXbii0tT3k3CVUl1ZGnZJthRQw3Ma+YrdRuslwwA8KNT6qh0O
H+noQaOxQIhlYiZ/3sERxU2dCF7cYYCPriXsuRxDnGPgkDi3wzAh9RCRpHY1CYVA
7ONyKU9UYnY2PLOzxq7bHnihMJzxs5oiQwg1WeFAlHBXfaiFLCzocl7cusH2/VrT
ZfwrHoOYj3IphgPxiIXbZT0+7KuTsb6ioTge7ZrG99BadwvFcfYnpHNEh+Aku6ME
+yGrgk1gV92WKCc+qNaTlp1jsvXFcREvoKwtSh7MOkgIH6xdM0t7zNcsgD3uxklZ
7pPfReq+l39GtrvRemz7bWLngJUIcyL4INvDne77lZ0cqoCPYKgGVDdDPw9afezZ
9rOnD8wvsR5ySDrXw3aB78yTSN0ZpWBOtwuFhUb3g5v62ZUpDyn5ePXGnPgprmEC
gQeVwZI9aUsvrLKJVCqc+/VvjJRyeQysejsUnTnBCcTTFAMNFSzNnxICilmu+OHU
bM9HqPKzH2skt/MCl7wKczTpzJ/I5wsICOs+lFohzDFNFb8cdCy+O1Ts/7UwNwFN
v5hTX+FUPCaKQ3mdi47Cfvj1ftzLjjtfFgJDH6ttQzDUfpAlvCXQU/1sYii2GMVP
BJmjqNeTAON2WATTOqulqZXe2r+Od8Lb3rk5HPDure0J7B3vEJFeiHlK34t/0rX9
KJafI82fnS6wJSfyogVt42wJI/Njx/jJZOxZdHG6UxKsvhxWAWF9bo6SGGkTrolT
1QChss8G//QKdyjTSXXr6hT125xiAlN7QTzVAmDwpcxKYifgqbkFgRiFe+uH9wSQ
8O4BW6Y9djjwdsIrGBAzrQlXpUSnKoo7VVpa9u2XmoBkqoL+8U+u2phIBpadZu5e
vIrR1D2ZK8Hv+WFKMTUhJYDn456HtiIAPor9rPof0r0ZXYDV4o/QolVfnhzbQJu6
gotCbbVl/8RKdVCSX6d3NFToSGiqlx9Qyn2rzDaiW3FcBjv9F7KkvN5BOb7tntKy
Mhh5EnToeDRwLsot5MVw8AjPspcMoqseyc3lzxVXuE7ra+yRJM1L67XCj2gZyWQR
E/qa/PbaJ+ou36rRMet8NZtFA8+3MA1fJqoht0CefCfrCmVdi/ykZ7Kv5opkteXJ
0bp1gLbQh3K3mtra/5t0oYKwInuK2uNpbyS0IFc56f53DfF+I0vjSCpymP469m2u
bqU7iUHKQgQeDU/1cJiGbzanwrkfMfLudbqjbjBDRE9LgiHu7GHjqWNxdpkyl6Mj
p0fsZU7VF6d69BRQ+KQBM3cLVi8QUdLlmOMVpBJ/q1BjtjI6i5+gshn14eu1CdvK
Xy5g53+AhNUN5oo3WThmU8Kegij+HhSroV/HxGDDr78oXyBuIXQP0KpFepBUmsqx
kfmLa65iuDCtJjl30RibnulzNTOMNtCjtqVjeRKM+gLAXRkFuGLmDebw+P4Bqqzx
pVsWcQJaYbUb315FDeu++D3g5AVekFVEsVY2kCF2Vfz4LDPMwNqvPD7VzmBItT5s
9rNM1u9kJ2i/IFrwBj/6IS4TQvVYPISPCMbDUVFLXGF5Ge2uZ5mGqtetbG30RKTc
5Ljn+dXRGP0UIBgHGBLP4etJKe65apITZTTq3shdiRIZhUtOS8qfH1rJ3h4/pZGW
VGoipXg6BLcZyt0JhJMFb6XaKNRnMFxMdbH83JhjHnETkGL2RcrLAi3gD6xQqCG8
alv5004qgCvepljEs8X8H70jTCdU6xF1djVzk6UbRthZgvR+AseeTGUgIM7KXk2i
tgWDlB3enBgRjoV1n0E60tITTeSd4t8ICqxled1fmOrzR3B6moMXYpiffUC3sXRD
zDAfMflIgIfcg52ctnuuvn4uP1cEmIpOJA2Y+weS9GoMYiG9PHxY0DoW0hx5JrtZ
8zzFXbn4/jq2P/+/2zaIvAjCGtJJQMR8rwuuFnZWd5c2YdcamEQaaKp6FL4K6ZHx
cdpgN1lyN19oAbCVjoZk0tOQnlTbJWF0E1b0J3b+JzNtM6Bx/0BE7ZoXDGlwqQzs
Y8DjyRyfjBhygdF+Nq5wMYvUFnfToYC8tkPW/ifFp52PIYizDY0IdWZK4Ahqu+gA
NKy7nzP2utvaD1C1dfvNI4ZvJtTKnDD2kPywC+e8XUuSQlnoLaahhArZjmAIKAjD
1olAXR9d6PNXkG/rsTNCJeKVtCoCOdepm8hRV/8Wihb8tfzdn5LJ/G+dhXAUKjLd
XL6nE2vXpjZLA47sgu6e7v/Trx7ckNMA5WvlwJ53xf7TjiZ3BE3TH+jGleVcpz1F
xN6hUKadYdQ1xIQKp2Y7TdkdrpT3c64flQOlH/PTNuggoR8Wor9EmOlndnLw5qzd
2kcmiW7jmbbgyj192HnH6bQ/NT9SNRXqS/fFVRW7NSFYaJ027aJMlW4fwRKLJx2H
K344258erkIdMSBflz9A98Rhr4IRX+ypVOsj7Vzbf4XWo9ds0dIXmBHvR+TM+l5S
PewEE+RpAkbMP7RnVguJyh962bDfct2ThMDbyMeIvH0iTk6hRdgsg7hiib40PSq4
ZkIEDtwEaeBInoZoeW6Cvlh7x+UEw/a09KbFIyQxzhOzSdE9Gt1Kp+1PonN1pUiw
pWEw4ykeeI1mUYmEoNCv729Y4EdePNuPkPviPtUNR8/ibcbrHTVp0mGjnuKUlJKI
JI1qYd36SO5qa6WV6Xr8C99r5eQrnXe8kM85iNgVqcnLULiDqIprFPiml7/yY4EG
2Q28tnfSuPvxOMTxfME8gg4V0vUC1X2VBknun/nVWAfj9YKeJ8ZIVKFQBnkxpIdW
nNt6bFiJ5qzyAbi2jQjMiUkXndSIxIkbe+jCEDiNIAZlh7Yjod7BW9WGltDFRXwZ
oATaz9h9yKSbCey+qgIsqyZc7lb4/zgAWnotOcqQhvPsE/vO/xkDXCQEWhSzTqav
sPs+qHdVGS0JlWCTOmeTnn7euK04Yet/3+OIayuLXTzndVTZ6SE9k74Q6b/j4pZD
Q6hgqjk9vw5BwoX3h2ipBJDk4eUnr+GvGy2yoJDBtXSZVIlAujINVW4JcRjSHYgk
4MlOvLiX9UfXttq41wNoGNNUvGsXwL4E1lGNZZ/e7VmzPr/fjbzPSWwMAwAQj5H9
SCku5m3wJd52BSWK/yJtgImooSnbVpS+IDSVCKg261t/gG1u4Cz0FJoQJISJYNiN
Lbh3zUjnVf0sUQ4hVADY5x6wyPAdwkxwk6DEz9LmwxZn5ql8nBITBhLKq1lGC+D0
X5X7E+2EIQznyshj+O8SeLrbfR1494SVJvstK5BCg+GbArZELjhHgt9hwOdvIkYK
8fVMEfUHq8uieZUDiwKU+AvUH1/CnWN+88xx9vJlGyb5D24Do4tcdbiAMfYKfqk8
atp6mZxJ8DheBQCi9A6BY0YnOo08SZzEHxlKHRs/yApUQH/Xnf1o8/pkXShfT5V8
B1C+Tu0bFJXNLPBg7QVG2SKq4NibgRdujuMIb8jMPyYp4UUrnrdiJL67eTTzG1cm
jihMxzO//lj0gp7FL7Wba1p0XfYBresgb3nLiF4LSpKx8osbxI34L3pYy4gfg1qN
4MAZ560ApcOS9X5YHGjlspQyZeNgOT1kcyryon1+0Oc0KFJjyN7DGj74yTC2dFd+
hefb2QcQlQmqgODcOGUg7kh1zn1a08/LFqx0rQrwh3RbA8NTLUntzC6w96zZfl6p
2r9koDUDb+KYtRmKigQr1VHe/EZan91MWqfvXf7SuRV9z01bYw0uDSH1OXqCjQ+D
TunWu1Oe3iXz1RhDXcuxvuDwOjQZgHlFbUFKx704IwO8SCsnu6NccWSS3c0C6iEz
hsNojstfTe3zWZE8CQ70/Y4rqDrzJQT0YZ0pabQSC+N1MgGkozvNnR63+wEjCZex
MEOp5N7OOjncH4c4qqQ4NcaV5smKZADLFECynj/+0eVdh3nvz2C98Ld3+RtSv7/j
uODWHUwwYl5hxmvBoO2CRdq+glwahhI8mHvH1OedftypElnUQG5yoJaVIf+XCdxc
Kz1dehegqqslhoLFlx+ng8ANFYFrZz4qC7JdDIGw9q0K/FUQg1AMBhYI+Qa/5Y6M
zEUcTaF3gfh85gnZQWIutXR965yhqSkCmfPPE2ez8TBXEfpnKikwHMj0Z7NVoD0Z
0m3BvTAX5x2mpg0cNq6sA3FKR3cdQo5RFleRefaRaQsIOAeGqnzuZTkpzVeFIT05
4M3lPJX6v1ffPP5/ixITFR4fLIEMTs+7J/KsUb6sD4e5wlxJY7gE3DjFSQeBp6Hj
NjNi3RRQoCt6Piw02cI8xC01aD27ANvPPs/7S8A8vl43Ahv1WE2uN5DzsC4tfHO2
d41z5mYnkirXSYxpiPZu9ID3L0uy7l9r/nJIdD5fP1A1mdDTz7AhYu2BSl9Ld3VG
S+ZJCeQNFaxuOxtWilC+tqmn+EDxb83yj/lRS842VCj5gAvVm7YYfwvu3khTNDij
YFHJMRBkrP0TUOw7cO1dJ0g6N4Om+Jgp7qh2ZU5GoyIt0YUBgfwKFRPEDrjnKasc
gVuSU/5svh3C5NnXkyzuDburBCzz48mQ0qvECl2Y0bbnn9G34xKnQMKoE7sWeQWb
zODO/SKtn/jIU59I6XYWbqhXkB+Hys+2P74S7jcSWUlbF2N3w7hAk7Fi6xOuhJJ0
W1JTJA8JX8H4xLNFcd2iuQHzd7qAtyBdR7bZ4B86Nd/dwIRenIvSY5lXIeMcuQqu
AEpGHnbb+tvs347MxzgZHlzSxKcZvylIIwD1Dbzp6bhE574If9hlDK/lQ2VFPROA
gZIxfXYju0zwpibdoDcn0rpYCxrBL/XriwXe5TKZKfy56x5dpCAlQpN+uN0xlPtM
LVfU5pICk2Hf9SFeHAfPu8e+lLPhMbwDw20txflBUnX3rgFX456QZYHZSO3WroK6
+QxCtCt5kQ9O5//2osGrnl7a7/y+0sYtcnAeTioPxfETn+y2xJG9Z30rsjHV65pc
oxnToxJqPA/V3tosUUtkE6bbE05mATJAHqq3RWgOK/uSzL9CWjtXFNR2mOGXzXvi
gzADto2nufpiqMdNq6EyTgReF9zUz7Oz2jZuumgl/LhLISxDzOw0JZPcCoALOWLi
F8NDYsTTeibwD3BMbWusj8MitLDSygoTNf1NGVAWO+pjh/dwytxkXmjD8S06j/yX
qcCLv6mACx5zvymedzTuC1/iX2mG2jYLfpsQsB3OpaxrglpW54AAbjiTlY+1P2MA
Wl0/D336Z/iF5nm17+Pp5tuK1+9IMnK62eA2Nw7T55RTDWD403IpPEhukF2Br1ri
OQjQ3LufPw8Y4DlTBPZqE8gh7yYwge0PgxMC4Z6MFkHF/pUPGGAY+at/zX5zWTaq
LiOMfULAGGDGnKF8rPnuGkeDjip4SOBLF5tA+TuRaBeNAGRzQVvIJNwO/b7/7+rA
B2duNKdv/I8+xhin26DBzBONT4MZYVX8TBYSTTAA3JcrN6LqS+YTzwG0VxDZ/ZGv
KtKSyInoXfDenIYHs+YEmu+sSfj8NqE3aDze6CyyKx7n0CgF15hOl1phbCaw4KHr
ZTWfVLwaZ9t3ltZ3ZonCmOKqIn8RZMppScNeberr4s85FJ9WtIeG0NCsxBpKd8gx
MilbuUsxtC6rwNPnIf2vuiCAWr0zX26xVdyq/8PnW3lrbL+6qjcXD+0UFNHsA5pQ
dXuWtFvy3zAqHjCGqCU3dBqx2iTxMWzHIjuGK6gz+bLLaBlqxkytd5TQt998WkpH
8DVdmLgVxMltMcXdm0+I5UU4ffKmT9xzcLuNMfy27JfdfJ9rN2Q3EEeUN/icly4p
nNBFYL7fSFlvNZ45CbCM7HSCsSCyhpfkP16GHM1/s2ONDhkqM8xAWljjT9d3ICnB
CWUWlZzprqmIDOX0RQKCJ2FuHWgFkfLsB28btpjRsiF8aFOYPDAfzk/C3eG0gQc6
/vNRPB9HWJBly1gQ/faCgU5GcMyRTcPY7KQ3uSGabuE/kbexwWd5AHa/s83LBvLX
bCu1tYO41DVi+sOjk4/GnB02L9gH//L0zS2zjF2AiNdqEBuAx3huOrd6kADhkBfl
DdPL722F0R3TvwezJne38pMYdiWtsi5EFXRv0whJ7KSkiNGV1craJEqDCUbEGD1d
7p1BxkP7xHbozLHfcvxzsi9LUO7nsjsJOTfS5KvD2syNjD0cpipdjV1u1c8iemLi
TuUwRaOElzMlm84oRvLdgwOfCGl8AlGQFQa8b8WEDf5K+SKWX3H4+aXUpac88ipz
+IEXwqoYACWnyLAr5Q0MQse+SytPtBIhnFEsTWpTguJ4lKTXuyKkzdqpTOe9rF0K
I0cvDQUPz5EIwBzU9tJVXT7/5RRAQC762SOLGwvJkcBor4nw5USjXjMucQE6xsUH
vQCvC4XuH76mRAfI3kQ+lXQS6zKCwFNgw3ht9i79irrRibRLarAibpn5WQo5WRfF
MAqCm5E5NSSBQDWLD7r/jbpBJlgHwf9jh4MjApNTeWDkactVSkgsf6GqP4cYvGvF
0AsQy+mrXI9QuAafFlQMAxexBp1qyzlWtQD7srG+9bPmw32/ffhI+meHRckbYD1k
j7EJpGqPdAiaiO5hek7PoMQ2qjIZ1Vf1go4pbSUhtlgLw9dL51WQchIrO0cx0S1j
q5KGhu1zZE3wI3fe2OPzeDsNPsWTaDWdAQ8mc3tkp80FUSxKmjW4xBEmHqvvlP3R
N9hRTP2Szx8O71JrPKVRfbuuVfUGI1iyHeCmqUmO50H0y+EmIBf8NW3vq1I7FWXE
Z/ImFh9gIzKl0O4wPPSagW4MY/t9nZXapoYRvfDIem3h26idLXbbPkEO9gSy68sZ
ha0oWYYt/GyhDLe1k0uo6eWMNcaiPVeYpXVPzYVbDDo7dNAQSbIAp2FNWq5tYldJ
EJpUWPhplMppNRgvLoRd2te7JKZMeuJWPgmUcnXEqmg2QECkgny8eQFoj5CLqTBo
rOLc78etwl+0DrXcx+A8AZcv00mh14tFipGJ01NMCrJf+NupDyha7IYN5YcwJ3OR
KSNFVFGSwf17N3n/RiaqVuEPeMv6cnuosItlw+eDGwUTJNehLgqumscMCZK6YWKM
rt3/xyZuUYgkiM3kWysquEj7gQu1KGBFMTszp2Dd299wWKCbwCYi/zp6l3CrGuoI
iEl1vfNIjOYPc386uOg6IW+Db7Uz+LSHSgavLKHwInBzz2UiTxIo1KV87WWCSDTY
hMGtJcv4BqN2U7BVo9OvozXuvKUreJiB3dQt0e3Sl4usMJMDJ+6lm7JreCbUFTNV
jxQwxXJbc9h1uw2+liA2MXb7u4RXXNUDOgFwUXV2qEI5Gy/3cVBRvbi3avFbSEEE
ble4u/t0B8biJfpn47k3KBd0ymjHCwq4VruF9FHSkX6GreGN82ezjMNZCntKRVgb
8HSHZA4PWd3paluiWV0xBzM7+Wg13cWXdpX7LFeG/iHr8SIIJwkNXTW/1Fh5NLCv
9Actc/G/UbjJoHRHQsYCxj47DJ00EvItaBix8AzRc6ID9Y6ur3YM3Z+aP3IYGPtP
6XTjnEB1/EgYRojDR7evN+rlwsNoeE4YtNc7ECTArhs1hdahBAOLmDw+JBVrPBQX
ZZs+7ZW19xPpfuwbdzoTEjuQRMbW++0uojON1x5/jWSpnorkNzvUQwXHcZzMR8sO
b5UPwr6SqFx2NskQAmv5Mab/NEIh8Fn7EkQGeC6Bm1fjoNnw/zD5i1Tkkz60wsZR
jH5Ww/57qI54+hh3gCGaHELT7jkmuxT5fLfGVsGYCXbgS+eCbOafjLnL0uA1B36L
nKtMlTuSdyWysAou/X8+A6/x8zWgI8CyT4XrEy3G5gHXdj6k38+fi2wnBMRCnIzy
dVGuEFpp4kyw1xhYQeQrVXiMXAr7gNtckbP7bks7qMUEXjMNIqQGpgJEg/0njdie
IfgNJxTeS3RgJgoV9qvAd7rm2QV0arpSvBUUHW+m22LdUJZuzaDDWYvFPWEklmV5
qMnuLEzJFXiguNFXK15iyF1sN0xFjiB4/FhYsg9kEmHoKuindpeWS/siMctjNWtY
g9+SD8PYXhW1ay3F5+i2FvigPSWTvitCCHMoC1XUIy1w/ujlhV8+WzSc78eaoCbQ
chPVFN9MA6vLxDzBjlBZlIikiyhFGfEf9JQdlgdQ5Ix0YaJUBX2NvR3Wdx97Aw0l
U/vzd4QtX8bjYrlSIfo5BERe1pqgOTeSkTN+cCs4hXaCfjl8GouNMz4IQgfhReB2
+1QRHJTZwVLMJhqks2rwVCah2gHWKNI5KXN6Re/+hi0aXy4cZKltwrYX8ycXElOs
+4pCdEBa6RHgLotKserLjGEPDd5/la9o+20gg531fC3VPVDCmKrjo01qDgygYJEZ
lXHrs9X4iAm+hJFBd7xjVnDBVih10P7lPCb+F9nckuISTL/11nih9AVaBEsIYXsI
LrQ0pxMLuejVdiRG7C0vOkVIgA0HAVuEpStoi2HnJOSWrUB7m+m4xdtekEG3qPXc
DHS9NBHVEmrtNVjCdnyDOCUp7kyYKfvpv4qYHzRMeHkkNZuiT9AbIcmCyoWIIGrF
HTLhH28OXKum5M7CvshLlrw1LLXvThunx91sxvmktxM9SEjZwmfioX6xVQ9mmRz+
sBBcnQ36UTs1eMeTboDLyVJt5F28PMI99BKb15i23KRKp9JSRIRCMoLRGhQwGdtX
7O4QvwlQNSM318C7OG1Pl0Uw+w/8Mw+DLyEh+Ikl/8Kb5Wm0/pAmZ1EVz6SBXO09
dvMeo/SQAkIkvsm8J5rXi2v9rstaUx7NqEFEFG0Sqr2jAwSLg3+gyG+QuF/aGHgl
LGO1ML1WIdlgoQJ85+W6G1NVAWHmviYAW7nx552FCGVCVUPKRewwMFfcyYEaMNkb
ot+SIDaexrRQzes9jTpShtAmfOLT8eqvBHb9goQb1QJRUpOuLBD9ezCok6ZHBOtY
pMx80hQJzyjO4voK0RiDMkuMOofVMZi/GiD8+WaXLuTdzJzfUF57uzzSJ0nK8EfK
CN5sN+isIQN8p46oCKvKI3gRYWSEJNFxjc7QV3ps5knuc11sFI2TRQK+YudVk3fD
9Z1mvd8NlYBcvRV/54w423IrjK46MBuUA09Zs2Llcsn82HAbtL3amI5n1maepTnq
e18pRMBT0Mto9Do2EvnmNAs4vfWvVCroxvddq4pJqYU8P7HNFROvvJgS/XPiQjlL
VMfV6J62PLtI14OuxdfZzk4tfrB531fQeOywu1QjADjpMY+FY3PHk/bug9KvociE
WEl4jkTmP+jq03k8lNizXpS8jDyxG7f15vF7ApxeT11Rew7oGzcIOA6lrZ0Yd37w
P6iHy38nIn7OMjBVDBRNhzCf82Dj+wTHZamCA2M/fGfe9KsYYoToQ0QV8jdKcR4O
McjTjI/6iagr2OlRQOvjSQitMMv54JxeyKsabozgqjAB9vX+UDzpUs5p9ZgSJ7sx
wxGugo6tgY6kbsznKnU2Rr9hUPRVdY8hTWOM6n6pAFdkHJgI5SZPfCkuz7sZJT7v
mFTvaVFvpe9g2zPFqmxCQR6gckxL+xhgF6AGKHrkMBliDriA/E9SenXP1plMeSJ8
ySt3+P/TILmmiXV94shKkB4cC+qCmn61LF+uRzk2d+jBH/6RNPOcCfTqoMY8x1by
2vyhZKPXjoOoAEDOmGiCNvo1POdnlV+rhSnwzw6jkBQI0NiiQrpbuKN2MyS9q8VH
sc6S1o4sYKEbZhu3BGReK72ueHORzc6j8wK9D0Q9kdsp/zeop+LU2rX8/R7cNz7F
QVvYpdDbdvj9P7YzOPdDILg+nXJvBrFtfWwKGbcPag/pmX/zUSGr+nhUgftjNKIu
nx9CzprqBFQ9wK7A8aE1sLyg+4pEmI7CoQ3yauIuQlRBW8snD37CuWHKQbZdH9mr
O7xwczRnFtcbAEiJaRPMsG0HvNEb2EbQ6ZRruAPHAUSStWiNFwT5YTDeVYwqmQ95
/8Lefo85yR9lqdxmjA/hWkkRFTxnLrOI8mrVhLJ2r203sa1n+U0D4B4J+oyyC1/h
AtX+jV/R3N0ympITIPhgZS62oUoo1Nv/RRWZ7ZFXMOXm7bJD1IwrId06rCPy4k8X
xEfwRxlapmDI4117Tg0USRtf8fiEqR9xK+tGgJmUrYKI/b5nIp38m6DSaBtG61kd
ELPyI3NXcBMK6fCr3d03SMBGMbkcJLUXsU1B1BDs2rUeMmpC/66UZ9wwZ+0DzErD
qbQZHUy7C6QhBONHOSg902Csm2c9Zc9pKjaRn5lG0oRFJC1zoYJhcAGx4M3dMClD
ZS4FlMO5xs3AozQobR0sUQ5c82nQxXE8iCIbdTi6tIpuK+ctOoPf9F30aQuIUE91
FM7fVZ+RnbtHp3ERhjJh4D6AOpRcMsPUyxG9BYyN5kyvixVptXD5eJkRnbCBtNUX
0GwYVF1UWozlFjMGTwM6Rbw4pxHVgrtzFny2ZFGt5Z/9tlUuRalt0CuSSrL3mCR2
sZ/KVWEpIKvjxyqXhpm8/3oVp6K65po1ClSlufQb7Rr0mgBhRDiKRQw6O/iMYnD5
4jphZHr1laECu/qMR8jUBoUUwj7CUTh8n8OKxai71zUFJkywVygnEX32DJl1KK9n
HCfQxYv5BURT5bABG7G6ScQ/YSQRCeQ74D4+jPLKniS25kvwZBz1KMKyc9u66riU
pzkSIwUydupTeMJK/6FVKz1NPy2uAdNPTXguP5wKGJmu1gggThq3y4GoEXTwjWTe
lHzJ8fbtQmFWTOonFPJBoj8jgudfHwFnIp3IZLkOvqFKUkKDbFozdVa+oZuosx8V
1sy6EETEsnR0Wr8ySPbluedoQxrfKGValQGKVISTA6reU3gi9EdeDb3z6IkiCip5
lXBWk/dI6o+jYVYHqFJQQJXZiHZV9aXgZvMd9PslFqTDv+UVuCUtuMIx8dh9mNx9
zKOVInGK8IRzafjsuKBRMyAeytoXXEuGoGFOsYjF7Gu53e+EWmXwpwisUoe0P1ZP
lbrYKUroboBMHYbOYgee3uTJTpEUFjRgMWEisT3mYF+WMzuJbzUYaW/YOjEkVKsC
Xfda0VkSrXgQRNhYpEfqlk23Ec0hmozw3hbfgV2eXuCVf3oUylYO2TpmcwUR8NAW
S2jgvW2oojDS9PqYwD3Hh6KFJGcG1ehZtKHAXrtEjEL1U8zkw0uii3OcEXxITjF8
ctXZDnJqMVz1cfOD77oV24RlviWBURkLKIT5UDC+32VRCiMJl99iqWIzZ1K1Iqja
Vmo+Zx2oGoFyS3bCuVWs53RwPjhxWIs+497RAvZ/dT2/CiFlmMMOyHpmaxlmGdna
0DCXVCwF8k1RbDfoXcL74i2gB8eQjSaHFQZ70blFUP1fDWLcKYngMJi/6qUkK1XQ
Ub/tYopmdmsl158zxV50ReVtPXtBhRQKMbkE2165LNau0wV+uCtgsZttIayfIUx9
RBZ89pNmj8PrN/RE1EuV5BKh9CjjxTi7rMsBohP3bPlcXFVbfcuR2A2B6z8Th3Qw
5HS6JN9VgKBnIch22MIZaF1i+rgsnmT5AdraBlVZutgEQED1CPYpbccZvs033FGI
xnNuyzbi8NA8cMuSZEm8NeR8x0srmSNfs4IK1ldaScJTLhwzFiVLQmCnHCYQK/5+
pOME/8joknV3xHhGypdUGuA9U7jf19wlsDDWIpdgHVW0bG/hwH5joD4fQy9K6oU2
AlyzHu8V78l14J6pexZ3OmZEdnhDKsGUPxjpFn/YsJ0WtPtmEHxBit+ung7/X0X/
6Jd4mlqNyCfM0ZY4EBmqZ68h61ZSLdsbVI2NPjSjJMIq3LFnIyjNT+zKGlQq3F36
9uAoLwoqvdZFMWRA0btmf8wSz5fxqWpvz++XSQE7Yv8+fLtAJUVYmXMrxsadB2dP
vwdQyJxR6jihtAt6HmEwfwIdMYUQh9ao0Rba4zewittHKz1bzfiZFTcDfjHEwSgb
we5B4ypoGcbJ2ovaxGekiAZCHUwgKm9pUQ5Rdw8C+C0qbch3z70pkjG+ic+5FcLy
pIeRKs5XrAU+dL/Zax08xTWR15xbQ23CfVUwTV81LXPx+OtqNFZDiPCv1TAHPySc
cGyhNL7xaapVbye7hQdLieE0h+QMuQ3mqElYEhaUi3mtwnr7Aik/f1ovI8ODnB+J
6bCjqCRlw2E7WMro3yI8nyI3moDZGyfuVFsi67Uxsg0y9Jn+zTbCLJIrBnc0ok/m
XzWrsUHf5I8TKTrR2Xuihto2O6vMIZlc3RoL1ZjW31u2+5aG+6oSMAvjV0GJEcv0
PpQSlUfYCfIuRGJYdba/qHAiHbxoHXJHeC1NjSDAKzT8+5uSfhhyiks4YRxsG06g
p2fEzlzg9LkEeWKf2FDlgBWC7tVPLCtV5o+FQBQwMUZLPNB65BDyLjtvqcS5QBh9
aKJ1R6goBy3fX1N5go8uXWdw//TsdrXIoXDZ1T+iXK5/s/unHx9OGnNw5tYRGcRq
KyEgHtd7SvS2c4FpiILNecbMdKV1/moBBnJbeFS9LMHD0rSQz93meyFQ69vId/SK
19DZaSPl0a6HHwEJSuzezqs1a9jRKbobneU04hWFrlgkuboo3wcJyAKOgwEYhBtY
rOaqEyIjhLMeTZjOvnQZSs9NkJ+41bT23NMAtbULQsDiM+Xa20xF4mQMj9/QKeEO
5XoRCJa2J/MC8jSmT2yldyET7FiSctLytwvJHWvRnpHi1yyH+LV7vdYgGuR8YBEE
OSDlFizvSn4A4TQedKV0r9Jp+Owk4Q7TJvMtF75E7pGYVfogkBKdH0YSDKgDkvPy
FgTc/VQBi866iQUw5OOiyp45TodrcxG2+dFEvqeWpQq4PDP77sM9RosKGdaNGUXQ
hYrtJ//MoTsk0A96Ay2BLje3nA57JXJ9+W3aj7U5y+LvJRR0RAclUN4G1K65NqQX
Q/Io7hWnma/7PlBo8Ufxgi8BP5tHK/QYCC1asOQZIof9EHT75eBhdqMrPDPMxFO+
i0vkB/0AWalWhb9E8S7QZYmKcaDwJoHO8gukPlx94zTRqSQbiBq4u3aEMkXtEdO2
1qmHqrpJizsj8fyU4zcbbHnMqsACfOCiOMWo92J2zi/dC9ygONQp/uYX/ToWa4lh
unY7a3shX3gJs7gdOq906aLhXzPWENh+MQsr+72RkLyW9PAY+zr5TKtIuVeshQms
A+BEV0l+MFENRhRnvltJaQJLTTLh932ChSRioLqCLkNtp/smnZizL3CxCjQwTnHv
fdKatmPs452+ryjuxPgARqvEnk2KEc/DXBfaTeBcLm8zBV5LzktF3YC4t7ueryHJ
w59vzgPJLJIezN/ALWmSM9lZAU3vyA1Y0WyaNrDnlRH4Q/LWyq6fZm2n0MgxT9GT
2Mcyglf93UJEHR8GtSVx1CO96odErTVI8znj9Eeu3YKNlD/yCHTVZM93rNV9LNh0
O7+LaJz17+/QUw1CoGwnMDeekvgPmwOSlsbNcXt4Q7uyAFQkZS2uPmH0Yx6RWqp6
zduiu6FB2B4UaRw19DABmTX3nwUow/g767ZbjMxYARyUzS6sJDX0B8IO/qh2HkeX
99UiwbveX9uORBGRtAN0LpcxaYYR6IRYiQDvag3x2veSpzksz6p5wnV1nSsWlG6I
EY2mPCqshYVmHj3KAlz5exdgYXtB2eawMiWwzY3nnrr7GmT8QZaaJJBDuXrga6aY
+EIVqK+Jwy77X99YCPGWGg/3wGWkuAYzSF0d0CCHMjIGp7ywh7z77m9xmr1prAxk
jF56VUqrsnVVIxQk1ouVTTGaizFUB/b/gxdOSrFT/fOiBGFTb/zK5XaiRlan4GJS
vNcJ7CUl5kXK5pkN19cgcR3xR/l+fXHxER0hry4U4Rq9xBkCjwFSghAo6QQu12ht
J1hPzWfIrdoN0ClkqU04roi96R6pVkpVeXZx50DBEabpfij+8SjPADNmLYm9A8Rk
fz8DHOqC1POT7aSWLvtNOvhQVv88ohUUSavjB3OLM5G/NizrYcESohSJY2bsT5eY
3Y9I3rIizl3vGXFrW8G76sifBuGhNG5U95ZTYcbjLDgkrq5M5HmZeMT1qr0vQQmC
UfgSj3FC3ZvHnPvWtcxDAEnSP1H9HJzhH+u1I0SvO4IoS/zuK2GH+vPKECteXWsi
Wrh5nUDWyTAHwvGshvubKNl3ppqgJFLWwQ7R4EC4Sxd7UD88Auy6D+IBfx8JdpdN
+2DZrVRUWeEfWjmJ1k5I6SIlj8NcUmfbL2z9tBBCagX46PR3BWf5805kuszRm8HY
W3PCg7rCrstyzOWvZTmPfIceeL690+JpQ//YVE6Blow4bPudtSrMWV2fGIhNvd5+
Laf0Vsb2CMx4q52mzq4R8gafv/NMN/4frFSO5OVPu8o6vFv/UIzSD6o0zmwgVZoq
rVEA8Qker98SBCWJT5EhAL5EJB1YXfopJ82zHIhacpDXkDYu5XMEMzmzmgugcuK9
e7jl8CxZDnTOQCVKRRqo/LGIn7UFOLOpE1LYJ51MMeAaVHSpn8+ERMFuAUriePKA
VdtlZ9s0faAabshRlx7OTCtR1jc5fp0GA0Ls5F6fpN2WmG+2rEFlqrMni2TM6Ix3
HmYbIbmJy44BWDsL5d9RWulSYdh4AbUxbAHDAaemjFc4001JawBA/kla07fVy1l2
/QUetG8oY6l93fy5z4id9TfSvKrEFgxqal5oFSGnsrm/fDXMzcvuWYRHky69MdEn
/sp5uW5lA7lacegYIduG4cTSLfr+Gf8WX4By26KGeN48F1uxJ22xpZ4roKXolq7S
c/M96pr7UgQU5mFpQ0PUu6DfvuvJSaTwn82cGDjgycSvVBGSpjlZy662j6hvWlzy
za/DQMTORobggWv5dMnMNrwK/SauX+83VSCQcxZ8MStrM7eyUf2jLOrN2h0IE9hX
ekpgsBMJjfcdFqjLMqKMtc351WhIAKO+HxBvfDnzfTF+kajMIcbtCrPofMtszHqS
N9AaLrHk/vgLJVhX/ScRhrEpfZ+X6umR+3fbZiqISZI2+Mf0kk47vXcd7p3OLPrt
7g88Mojkl9UeVeSga/Jb1MWGkEzM8K1iqIxeHrSFbGOHzzGy1A9hFg9ZlMskuA4i
u+wp/zXP8PjKwWMoGlQT8YXyHHfJMvA1uTc/15cJLTPLrJxaqJ5dOPskNopABu0b
JYkYPcDM5IEP3bq0XdMVzC699fK007PA7WOWdS3GXl6UUn5k+mVjzt75AOKCFOME
ek1FX0AQyF7DF6GUG/2MbzP8yhFYVLHYgtf8DIQHrf8AUOKno2RIJFz7u9Cd8SpF
m0xD2uBeoxWgZ7kMv6V0aTwufZIXYtjIBv6KfJYT2n/I5DMulgvC0R2JofFJglmo
S/okFi9ZBRlHGzZlSP9amQxMVEDIbzsRSbq2MlCM7NPBOKL0CNq9T+d7AegUfRBD
eiB2QfLTHNh1aZB58WFTp/CTvvMbjJzUG+VRcWHGj5scSpNFXOxp77i28a0buFng
2q7GgdEYab8MKcjniTkrijTdo+aBsFFwXewtzc6M2SkOr0Vs89voRqbXeUcG1GuG
jVki7PqOTpw76SQsL9OdiJ6PDQh5vaImHcs+v+3JR8DADs4BMSNTScOL71tiFvHe
Ew8uOfHGy+GZqRwaKCVxYP/0BDkl7RhrQ96WYEwv4pUQsLYVhmgFmH87pkYEDzCn
Gog4nAv57YCF9nPde2ERRLFBFGAc72mo05QfJzayHkevzX/wfAXaeVeFHDAhKdid
5dDG92T0u7su95FBP0mCSpkBE0imV9G2nOGi0caJ7fbow0UvRWBcrDcI9VhErBrz
3hp7zUT6+fzNUv8V8eWGIdTGrkuf4MxubllsPbCdsNrdBq5ahaw77jpq4AgXPqA7
CN+Y5j2xJobbWPmebJD1kCfznnYebyBSlT8igr7dVREVy9KBUSuMJ6SgKFQU018b
pxAszo5G3w4UzU2iw9bJkKTtqa4pzSIyd6ocGFzMbbWl1WvESjrntWjqLkj3y09O
2mxffF6KpQ1YK7Lsv5ttbWL80jKTvjQ15gjT8EzAiMMMdBEwp08LPYr7gXKt+mLj
12d8Wo3pThRtvgFtMTkxMiafFdHMalERji3VlUrfsozxL60O4hTDw26LGIgzPWzi
16UNIO8Du92ijHFRK21wZAnRAecEKrjtOKP0/GefrU+vdzpTQphrOM4DZi4eIJ2M
YQ33SZlmA/HamMs7HemOSQteiONF9x5QUpDXTIlVnLRIE9vkdK7c9Uz1GMJvwtdq
9FCZI9SdhKbnVa0KkbRiSeBWSOAWiU7XUG+PQXfQbylipgEMTnyzveEAVZ/JWwfx
v/qZTVtqkx8j7RNiyCikA0hwpJSUp/TafOYrxLt3UyC2in1z08JYiXyfOthKpbR9
pjaZxf+M91i1bkJdM8JsGu4VBOBGIE5RfitHysAJt/sU9YoJPmvN4uGqddYBmOhn
CyaEx2Vxnis25HP8lj2bI/I9oyII60LVC1wIwQ+KZD2L/eCCHpFsrSzih+9wUPZH
Nkn3X4LpIfWYIbJf9sGQJe7asrcJgE+y9XsFtnokE6a0E7TwjKWV2XAFTXZswtwi
P5lg7Ar9qh8UwSf1/Z/uKMOVL1d8Z846syclq9OdvjBwiXz5fWPZ0A8CWWkySS1a
p5y8PVlX18JuFlp//SRgo8KUjizXZ8AUCf+CDOn4LyNnEJnievFgGX7jRbVYedJM
vm8FWDbAbVjyjhwzH9v9ZdkD7f0/XA3/7yDZz3KEtaL+bzSeWEKYzm3S3m9eExt9
gzGJcNEAo07BxZt/4LxZKPY8TkA2hZW0Kj3LHvtIUp6ACFwrbnCqYGfF1KiwS6NB
NBQJlSJpSWdExOkxE0YWHq2yOVKeqHZLtPrBRu9kWDcLTRJg3HZInWzkHwl3UeTQ
iz6JFJCSOLSP+tMlBrN0VK95xcdQff5uG3NFz+Ljp1yRuDYD6RI9OnXRiQm+s84o
LRha53gsWrtmdLjH4y2vH8U94GQ56tDh4+2dzCHWwJESOB6W6CamBWuttnq7nsG6
BXGlLIfL0hH5ktpEq9XFgWeUCj9EyV7bPJICLxmB9PQhTfk70pb6odH7T/iFxIIm
ZWiWzqG2TkAoKGJdNZzFgtYNc1Nh+nYoTg2KoATHR/rlgv67BjghWcSgxPwFPv4+
nuiLCS4+rTUdNoOjOeCZcW+Oe6x1VM76gH6Z4k4IbMKtGK8pRA7nrRhknY3LXe+z
Q6iAhjbfKzVVWeI0ghLGeRAYXtLvNcIZY4tBhr1pAlO7OJBod8tSLE0X+nFE5fIz
RNfhimz7eQt4JZhp5uLjeKatS/Ho8NjUXwZQX1SlhVpJ2VVJit/SrvBA5zxRs3Ks
RQziEMn39wI1WFkdexxNmixdVhPr2dJDrcErLZvqFklPSKZn6LuqIBGb1PhUBkg4
a15Y2QUevgws14WVDSboZkSE3A3YZ0hBAR7scF6yqr613uU+1HmXjBoaO45KsURU
3la75qrLSrtMlsnUj5FscfwnnxTjcsoQkaM4Em4fqSC5bHwo5PVqTWbwJt41ME8O
F+mOv2Be4RQD86YfruWOP697b/xMuKi1Ffvm+XOGYF0gMY6xd3yPSN8GgrBcqfwZ
xbE425TbMNTMieaJoP7SZsmJlyyICE49Cks2idZIQMTNjCBOOMGT81O/CrTZDJlB
LrULaZRaNzorgWJjL39tHK5r51HU/0IGchiJGX+8MsHey4x4ZZfVGIMcrIHVNHJV
Zln10/Q8JSzdmxcEEnp2sv6XiFxHuySvxFxl6SIQAlGtdahQ75SvgSV4/B08szwB
yuhztndJAPyvtK+8Xf6K1o9s/Gj1vbSod5aBOb3BQ83KDbMkvChrur+elhx4Lr0W
Jl5UwTK9yfuXf/uDr/BgC3joQdSGPvf2UBLzQNvg86LmpKH2Ys8Rt/gXDXubwthg
pdPiYIXy4jkXkTxWz/bceALRjkbRttbJ9lmO5LnZ6067hI1kA9h3xUOw+t7k9jNe
byDzJdosri/HA+lk2wO+UzE26Y4dBtyTqgE5WHVeeDR0T0I4kCeqUagEf2NJBmdH
6Pmn1VB5DVwx/tBrEli5yWS+8TqR3ACfjp1hedNIBnHHzwi13723CCaZ4TS097dt
W+mfKGoCMWoQyZpa9lfLAABuOavuYbGA2eyQKlrehgdZjlwJ8KLSL2cURPYVWpqD
sP5qWB73FqUMSlPmBVr0geZsnawPGAYehWZxBhmNEl4uMRt/Fl0OXw8Emkcxz9Vs
esmHtD6wkEnqi29B0qoVj0gaUxgOh2i8fkyPttWoRZXDt9eV2W+CiZ4nh1sDeepe
ubWr6ERZSE++Q1HHGeSeZhJlyPDrA8iWiz1tHg6GBuQ4EZ7UtVJB4kgGIiCfersq
CJmxjZQPK+ElXHWeoR7uag5LSuXr6KXaxxSGDr/ZFTSKk27eaNmaVuvSfQklCnKy
uRMRktV3TQ99I48QHxs2N/BOOpPFL0KSdIsiKEF3BmsunmANKfddXbgijjvVCXUu
o3C1i+XCGIvTRh/jfZsAlgXNnr3Kb1/Sis680U87kQi3uxUi/KVtOs64uAMTWtBH
pJ/cRIq9ZrecbnsAmUFGl/JJO/5SaXQqV4RQQ1ohqawFcwXfGw+3t4+YW53dLh1x
Aar4WQ8nGw47Nx2wFqBh4cX8BvF9wKmOBUN6JRBNumGNP6m85NlYxpRou0NdAcz0
IR3S5PgUARZhdSWH88fytOAWYBPh+9opeLR46F/DANxz0kQ14E/gQS11DEGET++n
95n2Mpj6gOOsvPYjfE23PnrnTK+VVTSt/YOFlQYV2g+1jYDqpUUIxWWWJT9UoJ6b
S2djlXA/K8EYGVn3/Qm0XlszXq1kzmT2WjiRFnpV1OcONg3kHaGoczGuIFJ5DFCb
FQyeN4v1QipMdlsq0b06kAf33vNCAJhXJ43obVtWNRFnVkFlGJq3Hs3Li3LnlOTt
xPkAYcSgvzjDHF4+CeHXsZIG46h/NCTWnuoDSHW0s8G5oe7J7RsY8I5LfXBqpqHV
DiofiPlMvxQBKREP6CR1fqwZVcOGZQSeeFEtTIyUv61JTVFoMwiJEmCJ27+99pqH
T0r9UJJiof4HvnWdezgBgYEZdUZNj7L0gRx64CdsG1eLdlh6g+fVkLAVuFU4RZli
Pl99s+0CDTBZ52NG9SsxpkclLgDfaWlpIUwvlJTp+FeNgSwRYDEKFch6oYLCEw+U
910sgTlA+fGRla/Bb6vKC2I8XPNl68LCxq4oCmrqlInfYLdXViAKvuZ3Tdet16Yj
XbwYNvfxCBmoAZzmqgPffZGDKpd/Hv5hWt8iVVvhuNTTGY0cY3gEMkI61kgz35bK
Y+GyGQnR7NSWk5f4lqPCg7g2+W5Ty1ePNNdcuhHHV2vKN3K+92N3Nu8T/RoWBBlz
AJtQPw/Dn6lnJF95Rn0BberDrSk+qwxuON4gzEveLe6vK8NUjCEpQJ8UtQltrkxV
cT8wT39B3Y696BP2JQ5zbuvovggqXep0Rm7Fd2jVCPv8xMl8xWN43ReAh/Ggm26p
zay24q2zAOATXpCAUj3/cIcdQA36/MXopZq/c8G7128kxcxbNVeocBOILfHqGqVJ
ZnSZqkfHeHKPzenfX9N7GQMR9v0//Dmii6Tmusk0npmDd9U0SZm9Dus/8GQkbTWM
1FGrUc63EkEJqMoaS9iVK+ZA1Vkip66T1Ts1acmTgTjG1BdYUXRHKREcS4Qk1n+T
z6+szzgFJv0dhktO5yRd4/KE07jX6LCQigmXQB5cKXO4OYjGLtZmPLJUQ7JKGpL4
ZsAQ2GrTz5qdVGhowyeJcANKBSyhuS5LAkemqmeiF1m3eZJmfMyGLTvHjQ7VbdvF
xGAevopgv8ilGkaEvaZQKUsSpQPDbMgt+cszfHfj7vNpXG0uq2/d+OB/coteG3Mz
tZS/+QhzGgEg/JGPPx+veV/ENEKwFx4NkBT0o/ZBe6osayKhtQlWRUylCe3r2y+N
nk+cGq1Lm2xazegzFFdlbIdwM2MzfzMllqZiCufHG77CyNQjp0Z/JCi8L7Uhg1oV
coqo6WBzinJgW3H2VMzjMoxfYtFmLO3VvffA34MM0FFq8dlGEzILTeS3Unz0Ss+G
qD6ElTjrdQhxZmH823gyRvdAhmt8PwpoyjWqfyb9P6yXHOABJclB6+FlC0/OErdB
X3OuigQduXr/vi6om/ekAfU+EC7hVkwbZSASLVGMEierBxmJ7LB5ZHCb7xaOdMqs
RQKb8ZF3kj5Qw1+fHkcGpaNKpChOq0Q/nevz1nLA0J4DF6Ex49V1ASuKrEz2zQY5
m5Txo49gXNHf6eT1Idrs7R9WZ1QMZyVAeOK276UaXYWnKFpbxJRFIsxrUG8UVUBc
QB6tn6EWdPFbWcF7WgovDob/+WF+/4PmoQWHSwjSRzadcHjCk5udiPNwNApJVR8E
oMF9kpfYVTl+wDrttAh0QzrCE95mDHME+2/iQGjJr80Q5NSf9LkC5zL0AZrTkxcH
MhbCAx9EqBqau9RNXDSDDKkaIDnfleQMFLy+se4p7U/YOGQsNDBv4qYIsHFy8JL1
0QsuOhW9kWx9X8LQRCKq5noRX7unG75n7Sgmez4BkwRoX5HkdQGyT87/e12veoYc
WGi6uFxncPRuvW3Gu6FK+bYhdobpISR6Hgc8OvILL85DePhtY9PUigb4csz/qfkb
qVB/VC241/OSeasI6+D1pvPnceuyPdBqZ70K8j4GtrIX6xm/bXHmc6W4c9TNiBh8
A1A4jDDSdNcuLALpY1tf8/IQ4P93LG9QmEyo9drEGYkuqojPwUztKjSACnigy0YV
MuhzeKFWaO3opw3JTXeyEkTAXqPI1tH3c/cxbHiiyYpHM4Ymt4xcO5eNEUpo145E
MkJK2eVKfx15jOej1iO+4XylAlIHURnK0s5b8l7aaSDwQBSYR4C6duaPS38tiq5d
lcAJwNaEdyfVwfbdGWHfgX7ba1Eirfgg7mWYFbc+bcIynX0eCREPK4Oh16UJgCa4
qV0Jsae+gO+ZZ7zOT80OKmc7u9GwaU9ol6lkNMoxv5bN4hGrWjdyMSdVH7y4pIe6
bHLs/iRZbVQQGg9ypDDeGVvt/BFr66+Vhe+VCJw34ogXszFAjpyJlYC3G5G4SDJP
cKp4KIrLZWx2PipwDx+Q8tpHDbuV2/EeS5vKqdrw4NplYqe7EJDpCzK7fp0X2rcF
n47TT+UTc6ezufzHPrxK1HiH/2k44UZB3RD40syy8U0toF32/HVunZWaO0BHV+YD
L9XNODqn8TOA/cRc8TgAWFGijiKQCVh6m/2B4+Beb3nLf+59wI6QpDeCgfUXA/46
EOENkJr4PPJY8gD5jlqn2ZqOgLArULMKgw3ss5IWuc7WLDEFCni62XDoILsO1CsP
GXFhi/fAGZ9xn4t+T+gBrQkoB1zAJY4z7WC7ZqOwYLNqPDzSDnWnSMuao9rCdLFT
VIjqJJO9xlAyJOVbpcNr7+rxwzLUAY+QHHrH/sTe1r3buugJiqEq+GlNn06NRV0F
2m0dA16Xj3UUjldrkSc2XvStM8xlpBNOYZ/Jt7Ouvrw752yEOV5JWgZHuJ/VXcRu
DxuaziPNwH1R/M38m8WfS+rNKN7aZ1aRb3VVgEdIudzBbCmun3oVCOxydyZubHkK
QHqaEDRMA99tw+kfRs7MH1aqJX0TTkQGZWsO7gSzoO1/+3ZBMDUXeiT2NyTa0lP8
b5yaq5bHBBxO6ZAoew1TjdCPPTaDGS3thmzy2SewuSMxKQAyNrT4FS1iY2Jpgpnr
PIqGsCQ8gII13Kecsum4UA+0oUt8EYc86CwdHJuZDvF2mDbBtIC5PLSmEzsBsD9g
seJSjnA0wxLCMxaseUVm1R2Q5nOACs4XdUyKbFhREUe68eh/elyeTgMxOChMNG+K
yY6TI5ic6qkSUnT1Cj+ewN42i7raaJtHC7QKQrluR5q08fdMmk53reVgl9Sxb/Wh
BuJKAzySoXY4l/PhFcHtFAd7BZS9LxvaaD3O0kyfNerb8CFuD4kkEHG2U/SNresC
J828JQt9pTwKghux0/7894ze4UmFRnWa256A+eh2R4mazt74/E66LVrcoE8ijvb/
c/8tZqTAUsbNcRFyfcSsIkHV6zcdqjR/hVRR5CaDHtodmzGYmKmMl0lg27xGrv2s
Z5XTtbeCQEmYwEQnv7QdzHNKNvFlLzrZ3ALCDW11VHHA6tJtCWe2Pez4QNW1bt12
hPPzrtUjD5e7PBG8PzZx1TI4Q5j9Ka6skV6F0iQBX2rwYx9abUe4pq4jvlxJIyrW
OXKXagX29SM9f5cjkyetrBycQ6hUq/BcLKzlBnLSPnFjbQ6WrINVUEWlGBvl0ECZ
MGjwc9EjqAbB0EGgVFDt50OajNOB1UlqRR8gO6Uu6Bj1zjwWjn8d/W7f35hN2f/W
7RqqNgpU3ChzQELSXe20pKCsmyETvdr1L4PDGhDXcQ/7Rbig5zDviqfNuFfyUbaC
prJWF3eLtQpqoYVTvjARso5nwFZy8aug3IBLoMz+KxBm17M4Z+aLfdSrcmDSqc2K
fGKGpleUFBMMaSCj04y0f5YUL43kiDcIikzzv86+ARJhPalSbLbB+GJFY+AnkSww
mpkSO1iTtx6ObRZ8gGoKIWaODIYt3WXu1Wo0lpmx1Hj2pgxbu5yDj7xFH5fWCnTW
zB02nlOzIXPO994LZQzS5UenZB2dV5HaS5La0eSTCNxcDrtbvq4t4iNINt9P7r7V
1fP0BKqbCdGpnjjvKTXK4TzGHpuKBozxxi8ktKtktroQDi8pf5YxikCNuGj3tt1g
6N0fKtbgVNhEsRcA0Bm32cHlajwwstkx7Mt82w1MSPKLm4THERY4+M8em3bruN2F
vxpa4O9px4xq/yrWv/MLWhBvi3nhg1dtRxbKI1oThJlIxh+sVexUpMTBd7rlFoXl
p/mxwgFu12qPF0V7eaTkBPsUvnqVW9UvB8krnYwEMd2JdbuYI2s2VmDFCZcrUeQK
qUFOR9lubBLug4y/clWWMczees5xCO2ZlGyhowR9POSihvGM1TYmXTVWIuyCoEfa
kRkmyfv6MlHZYcOLcKsvXXzj3P2eyRy5LIT1+YQY8WtqFIBMrGmljpGHUarI12m3
lj8lnKBPMZBin4GsrA7qAwpEo0Vk9A8VrqRFhxgzrYqmCVozIudvEr9+9vFdwgd9
S3P6XGlqdaMwOvzxsg3pBbK2LlhJpxYjnzY/Ue5+WSlWXXa42yF7t5YYJzRjJpRJ
NOOov8GdK+hbWGT3il1jv+/+aNL/1o+OEnOeix2e0yA9Ap5M4bHOxOeW845Pz58P
b4CZdyLy4qxOv/d0ETWoaZNnVAdENlfd9RsJrFwCucoe9VID8A+xYS+DJPbljbFz
lcMGFOdhfVoPjH240UOxwBTkqSILNZwkhJlsimCVdElIqqggqKhx1toOxLF3yOIS
KSWkCHM9HotteCMWAeX3TBUSw3WrgrjTszRbilFGvR5WycQKZH1zyWTx537LDSSF
9/fr9DTlwq/QXOAFs71D3yDLeISqCsJm8jx8dBbWqs6R3pQ6RXAo0ooasyzp3RhB
70ULt6f+dpZrsChUvJUBYMlW+fYnI+HrPOsLdC3vHHuQ9DaKa3FXgEhOCxLabJ+x
07DgCgnWbo6Uta7VkjCb0YGqKOu359YQpQ/cNf5iOV1O0GUgMjQgCvS8FpB1/pqx
pQwfDFcwCxEQE8Nr4R/TbSnFKH/7QrufMgi2FMrRRsgnd3uLhWPH+4erNrjUN9oV
WlR+tN/CAQ6O3czJde34BnFEw1TNaC+Ig1dSY9cObX8sGkTFkfVUcdrIAhnYG6Bw
pd3yOCEmyoCN78PIccHpZiWhuf72sIiwt2XFAQRbcMJSIF2pOc2QrXBlmhbJq9l/
3jdSaKzuO+2A55r9aLCKesDae85GqsEfh0TLEhebAfPhpvf+fXXYxkAbMxBc/JdI
Pz2MfJpvjGqWX97gbfZDeNiZrwxiOoEwRiNAvmhsCJrXLva/ev+ZRA0K/mO+q00E
+3iokSVvbQtyvglVvivviF6H9N03Fq6/ARsNCSP6fuN/dDZIVmpG/Gfqf79gtS6U
SmgH0HGUaaO2jTwrYyWl6STjuVQSj3xxHcWjN+oIhM+wWbu1qlmNhE0T0sYzOuLG
+m2ppQSNYI8+rqwRHNU1SGrT8yZttGCI6TwpVzesn57EiV25w/MMgVCVOIzhkhlp
cNUVSHu6HafNSfR+cTNG4RiwUVebkcpXDL2TDv26AYKVkCvndbZJE8fod7BA0Ni1
cKFD9l6eZ/H+M84hAs5pNYCRGsdRPgIqcZMGCl+3aZjfkDTtjBK3HPpP9ThW0Ne1
LefcyY2jNnALUUGy392/ire3i6MJOZz9rJ7+9cOO72mfg+sirhdHKNuozJm75VZP
xUce7EeizRQceT+WxspUY1Mu2aM6DcJRpgd6MV5qCwPbUe+rpJ0CpKkd6rT13SCo
3PB3TqQ+BDhv1uvSRpwfTB58TZfS57oyQupWRDWpj2mhWzz3o1/WW/iizH6SsgrW
TdBhrhpr8TLrjC89V8P62uA2jINtbzsqaj00njPRfROAEkh+/+rSgGcCazRdOgFi
Uojdh0S45Vr+02BPf9QlCYGYB5q2XHzh04bUWxKFtVA2eLHElNlzSbiOFZ2yHB9b
MnEUderJCfCkN4oh3sYL/pd8CZUcAJONI0JFknvPeK4+wijUo+3SL+imWlL+unNV
H+KDdJZgwj8pd67cMEjjWVsUdeqce0Ph8A/g/jJjdytF0FoEWZKs67PMa/Dg50Wv
Ujm8dUORD6kLYhnrCYyj96UTgWc/3HhA78UrWgiIXRozQTYEl1USZjhl0Ti7ov+Z
KxL73z5heSXceiCTNIgCtFPi4GpjNopiDLzRxJ5LRjlawANNOkyf/nQz/xPzYdp8
rjjNJDoQc4oaK0fhDotz2Jlz5NMdSpKvPEbkx8xGeMWRk5N8KSlK5vGvgJx81hKe
IoqqVwBUOYRXF1Py0prXKAxnW9biKOBJoy8VehwWViP8i9dnOHVOSxlLJjysQBwO
6DO8Vs3d1GvA/hq+l/+xsWxrrGycOgO0cRB9Yk1evcjT7+xsHczMy24UdmRRX48u
qGAs69rWct5vyB7S5GEXJTpmKN2xOqm8pjR0G/w7CBxxq4Xu8P/XnIBHChofpzlH
szS+idSKTW/CghtmQn2bamRTIov1VGuEIVYCYJw/DT/6EJkSAzNny2EzBnlf5srb
ufSc4ZS/sl66nP5Ea8PhZoJACIR9nQI8eygppe3dytbUzm7XZOfDW4L1HL+VRNVg
dwe3cKEDS5f4K76wsaSEOeFrpZshXB1wmGfZHtaaWe8ACnbLbaDdWcGEg3+l4M5W
LAGabNYNbUgLZE1bsi+bKzBuJ1KpAot/ttSB3xAYwYNSSMoBQx7RgOWrdmDABDIy
RlgDka4AlSo+0XSrGixyvskrulymLnA9mmPzImOLlBQSmllK2ka///PFCVgdbWsc
hV02CtTx34SaK8nbGviVghE26qRPpqAdjsZ1zKWbxK32WxT5J32v7hYcR8ay0u41
dyWe9I2/yPBOm3yICRLiBApcJymQm9qn/1cSbWDgcGxu03MX/cnrIGK+BmnUup4B
G96/h8+b3s1t2csaw9EAwKGIXwxi7SvyxTLViynD8g972/bwgjrrayl8xifIdY81
1UrfKt3Y9f+OGV2ENDSEifRj/zBhwYeEkr8BE9kJgxVJLVJ+1NGPVNmpyRqr602Z
f2jRAmF93z/rTlyQ40K5wE44rA/HhZhK/MlJwgzBiKoD9QtZyhkPPJfW66uUG/5+
81Vh19ciaWOu26LB7Jp0liuTblJN0Bm1AqJm+MkIfDqMrSrimNRH0KDPBap1EmgO
GooFWley4ve5O/Ekd+GlNkk46LgzelJiIyxH1yPQibzfSc3jZw4oNlTW/lMcaN7o
gAeUZrwmUYXfPz+V862e1UUPsBqZw67n3lZxasT+lFJzD0YWNO8TBEzEGJrz5xoV
+aAmFfq9Eo0XuuHakCJ92jIHYqZwxpukT0DMp9QH65mghpO6xuGb8dXP6SPzE2Ew
S3q8RQClvHroUN6PyRsCxf19bN1R/r1CiECN5I71XHIhZ5K3wEgHRGS7NeXw7v5c
hcsSNG3gij8FXdmAZgGwy4JxkC2IYXBhGmjW2jC72+9+fw13bXY7uybEHB7X8MZe
Mjct4ZTMhnKRmpoC1K94y+wsriAEOrinInvzWsP9kTjsR+wO0Nq0ijRgCQWP3d9G
/tU/XyB23/WprsldA+bQcMPB6JggQnqqF3ZyAgCVnVgzdIpzRXj4lH4ntl23+eVT
GIfJwDVEfKK1q8ugrETMI2gPFNNGwwTuld1ye1sQnFF6dssKWOczdsD7Exrn8AZ2
hpwmk+ewNzP3Insq6v6+qBIDY9SJeXKt+VpgHf6qvRMw0D5pcnsv08lJeLxv2QsB
k1YkqhmwTpvgyBSQf5MqBaVKorLlRPlSrZaoAFTTUPFexFpAFQWXxypvGvn/+lcY
mKZgKjQZ/oSu9DirVW5dorqH6T4v4NGj/Sn1HOBrHZA7e9bP70TBsGBrDV6FIWxt
kxcJ/de65xFGIVPiFUanPfZ5VOh3EDCUxjacGcQUaBcFiUUVWZjyJSvsLZEREYeR
JPD1a7bW2H/GJL1ti0rT7CuwbojmnM0alKfeyWH4tZP9gg3VVfs89/SHntHrPtzK
8gaEeV3CJ235+3WGt9oFjNejbGFqUVoUWBAxtS++F3LajaQ7zOqQuv73WELtQaZn
G9G2ftl3FJ7GYUolf8AzX6L/vp32IAaTAxYq5dy8au5qxnPkm6/KumW2tCEiT1Is
IBgyLMTa6YAUxgjgBkx0Mi91V3sh1kQnjEhb6N/7NNRd8uVcY6YQf1YcGhIoQT99
di+K5D5l6akTGSALZIJjllmpCueDTLPcl4M+bkYGQv/C8sZP/V342MGpJiOKrn0N
j36xcQRB+Vii4Zb7e9KqLO//imAsXG0XaTpFazy46NAB7NE4+JtTbf7JsGYhbGrv
agRuKoBfaSG+Pj8+/ts+1XbEtjRtf0fxlzetvj7b3Zn+LpMMJZhKuX3JtOx4S9uc
GT3dvmA6APL//0aSRYUWEg38lYQ98jhyQdRuGrs55yF3NjdR0HqVv6huexFsVL8s
L3SP5475+Gb6GdcyXug5RsZ+2r1+0g8Vr+FQEt0EenKPAjtQDDc21WJxS6p7Kv3H
CcZ0MP58GKAW7qR7nBGTLr4hi2QLHc7jdO8cMehGZXDwxzartdAZcjlE5J0tuifk
EOTLTFyJwmj+fMzKOw06ZaUN/7ocK9WOtVX45DXajS9zAGeWJSX08XwhHahlPofw
S8LvBceQKgNw83ip/aioq5gyauqrNdILTs4KcTWrEKDoeolOY70g9/aOuuy/IdmW
PXLmy7TEwWOI/Fa+U4oUPeHyGyQA89U0Y2d0Z1pkQRyK8BUUVPw+Jdk9srDPnKHt
efHcF6OUlmDo3Rl4FgP+YSEr6Mb1s8/svswnUBBKRdWHVTsae2XS7o8QSD5Wv4EG
gnLFt98RpAebC6S6yaq2MhGo24/EhiPNcZuwxUj3kepR/6D+R6MR24/bgqtagRc8
5clFwYUKw7pOOQAt+24Q46OoJAQNE7Uye9Haq2aJono6zps1ez013STmASIJ8qI6
IKjAPf14V10WmpFVYbspTopGUnHnLxoDBSLh2ydBb0pqFA2EnA0FQreJgGrxMRJj
02vvXSeWnOBM8xAez0ONQkasDg9HeoCWBuQbo/CbziIavUUEHNOS6HuyZnhqwC/3
dOL+dqEdRan9hfymIZKntIFszUWX/UsD5HHAOes4kM4SukXbYQ6YjtAQY72JWmCi
vm7SW+E5Hy2+adKflmOsSSL0p6537pZmuI0qOidI+NNwDrFcFfNmA3hQRFjZbEDb
T0Z+5n1I7Y8zf9Sm1tD/V3j93qE4DXGZJxpgsA70mZ+XDDYeRniA9WAhVIsh26+W
SBtZPx2J1CLJVCkh4+19I701WLfEaTxMFU+qKd9CLiJbp5c/7WCGSoGeWlSPDCCu
ruAeo8AJcoHfabT3bD1ZYTF5IhqW/J5g2meyGf40LwzfpITQCyrVDUcy4crOR90b
Nx9NSOBJQC1N47SRIAHat1+fRHDeQn/mrkGs5i0tfcgZLA4HubT0asiHnHJtiAuv
fP5NS+S0HOE/73jBwsOw8qBkrfjs6sDKvaEvTTlzkZHN43+MzWhJkPe0E5mYmenN
DTQETwklYuSrZKabnSOSicoSFP7Xp0R1sqQznzFAWSPblG3TAbPiWtJmd4DS6quP
aBX/HND0UBxLPqlyW46P6gmmXCn1pGMGGiWK9GXLbQmA0cF7wa9MuvcAgNa+gKLg
XSM5UCZVpa1gvT/GhawpST2gEd7iMwQiNraBchm9IINaVmHmxdF27ZIM2FC/Bu4a
sGV4iovOeb0X0bc7cP9auS/NuZ6dmLNPJKpCHT41q8BiDcVoozk0hFkBUcQYV4oL
2+AzW7JXCzCPNRGMjiHR6prlbuWtQDet1vPpsiVmOkAG3CA4CZvKmo/6CrDf+nLt
LuyDWfXYnziwqyOwTrQSJrHCZVHXq86PnhBfG1AIWIDMsjsLHVAs9hKH+cG8Vq+E
LB93kVvAO8GYpD34Xvlqld1TWA2lj4K7NrodjpXv9ijnNLM2+misummcKaGHTAq0
MAJYfNiT3dN6iLUaN7j92dguC0j4wEOb77rjGNiaFclhyU0tw0GehO6eDdy6Fx/W
3gHtK+mE5DkPBEPITaoFDEAmZ0Esh4PUfaueRyxXGSSUAqtym7RES13Lfxwhb1HO
92bCFnTjcpGNiy9rjBnmi5xvHJzcM7qzG6lEimZLJ04sa4Jo/cNkEg6hwde2Mtle
3/D0OKzD0xUxIhzpIg19lDMQOBWn+ACBpzoeNvxQhbuLUJ8a99CPpmeCP8z4Jtlq
V14i5os/aEE1Kol/PSN/GrwtYd8Xjl8DigK0o0bjbMFyhUOjrrmGib3asclZsFNK
rPQ9smruEpUUXa10EJF3g5Po6upc4oLOWcDu198nZTGoYfk6Qfrhh4XWg7saxdOc
Jt9ErZ1miwc7zFFoafqv2VdaycDFLVNbbJAS0VrDNN8iJja+BP05LTZMI13bGO52
10hsJbKRtTmax4GLMIKGDKArPSYnGivcE0o/dBm4NCughp3AE2rv8ipxoCWDScRX
FSWGPUKf4vIY6YwtbzAavSSBFU5fMekvb2S2KG6tYWIg639DL9lL6QVIPJMACUgL
epftZ63D+6N5LvXuIPEYdosNPsScN1UTXSd+1aK3HHc8CNglh5SIthl0uGYghrMz
nIxTe8kT4gCYbSzgLUJYY18GCxAjPjQWOFsJAKgXJn/HCscbF7b8WM4ifY/m4uuH
2E9S8+K4AFiY/bacwwEf01B3WpD+LRNbN5cQV6WFRk2T0+FlEpOMhdus385G00Xu
UkJ0yTnCdCUSEv9NVdise4KxeD0NGyQwGYcdpF11weyDNFltMnxNHq5O6y47mHjw
iagNWUG4dMQsUunHaeg99g4KWzZHqmeoUwyTvBQaxqxTgbC7rPkFF4mWFlkOzgH4
SxyWzxY/Rt6IxXEJF6CeRDf2ktLHb+pEMh+j6fwMEfoYguHuar+H1kV6B3VV/H4p
KYX+oTOdF3J9Bg6Latvw1qTBRG1V37ZoJYRvSqs+4pqmMBsJCG6j4GHc7nJfZd/H
U7+3AMqZQbgUEQbE7zvMDKknuWQRLLpSsJXQ9brvOAT4mVKyBLzy/lnG669zhHNJ
kI/n9S+NHuNein3s9TRnaRusgvYHOdy4Zmd1IGNL6wKn3jNo/ZQdPhiYL/Ky349O
Gf7tNyjM9r0NdHYNemQJjSbcmNyR1SSgI1qv7VQlJpvNDTNoKVCqNlqPm9EbhQkF
sKoF+3cqHuCzHiPWx4Ea/02HE98+qfNA+AqpCbPb2jf6umuyRy3HpElRxp+ZVG0b
kKqlvSzSz4auw/2Rfya4P0RxIkeBt6W6KBstV+CX8ms0NJZBXEBEElwRk1aCWdab
VIdDitksNqiKP31rPiyOdM8bQ8H7Ze/l/8pS2QLHkPeFzE1kTmotGOT8lqgTojEf
TJmJaFSsDjqCWujbHw5ecEk+qrNHWEjcePYvMHNM4sqLAuKcMqHY/cF5GqF3xGza
El8fYO7UhS/vSNGum1SfpufFtMbTL70rKJd7wNqdzldZDMpiTuY/G6ZB3k0c0Tjd
tXdwCQpMQMFFXDbWadz3TYWxUCj07AdC6Rz/2u/xxDA9e0WX+QYmt6IPbLLoEE+n
7SP2UloKlGEbYdyUheiQFeBHGNNi/sPv74rokC5mDnrGaW9FeSGrjGJCqPoeWfHS
IoUul8HrJNwKl+CsXhxdgnME1pHNIKguUjDn3C/mD/4d0bNLB7sG7Yb6HdlJtZqH
jmRliFVwEw8+5mxzmt5WrS1dH41jrQooVuoawuDod2hcewXgePxd2TcaB+PR6Q3c
9ktT2rf0D61AmFP7wOFlCM8G7QVWs0GaykY22P3odNFseQK1YnfFdnbeoSkN2QHS
Bm7prubTu2yHHJbJ3GXWB4CLAI3YW2eMbbfjgYvQ6Q2hNF45ghs2uak+7PZpvMtf
d6ws1zHeX0cIlFvEPf/B9M+qtWvnYCww0ZXM3Jk85tqVHD+03zav55rN3hJ8q1/g
BtMf+8FZkcEgKOGiEPcPFSrGr7VIe3o1DU/mY4YqT6OsLTcpIqMzbZSSqtPWkh4E
pPWIJImO3a9RdRDyyesR/h1T05kZti/DehufGM15kNeeUw0BtjkEAT+BO8Jgegao
4gKXE2oWzNi09EaXwHEa4Pr4kYpIcFhDYfq8HpvcEXLy3P/78A0uZ2fz7SsW1hyt
hALJ7uoxTywJCSJgoO1hS2xTSRIZ7zTcgLynTtWQi3QDENR55zKQLXHy0BO7t4fj
ybZbZ3pc+HwpNOvNxiF4lXhiAMYtD1D1PbJfyiVFhIIR07oXCv/IhjKFagDQpuRx
zjNcbC5O3+Lo8WhBG3SRwC2AeABMeS9DD5PMRslx5Evw2XOE+7PC506JLcFzvrEz
B1/gu2UytTFxwCIoCd6QKdHW8R/CYnVfVcjotMmDP9v00yBEwDKpwshST4j6UgHD
I4okgdfb+GPHXI9vOJ341P5Mc2DUFJrxgYICzpCmQTbAr/qqA4mJkXulU9vNprDK
a5dosScoKnA5YEx87pDPBEg8oNYldLYq+IUfVxw1kQVLKkqg+utI4oTb7aETWZAC
4nrftegmP21+81rsO6P0wDh764+oeLqxA5MrI9jSq5edo3BdwF4/I9/an8ovTnVN
B70BIMR+NnvZsKBSHfmq2wH368LDBsb9DEqT82QI3erWXf/EyN3Lm+6t4NZmLbFd
9gdK5ojqbmNDUC2W4QgWr6LwCgSxQT7GeRD6Ldy8nNCNObd7V3IOK0Zu0yMGSeFt
0uRjANgarBYyv8KM7tlWf6KEvN4CkZZCzc0KTSQCkkroS2ZFYAcG2WPRenKFI9/4
rZdNkwM4fEEvvqnogih1S41Z3Iam3dsaZOXKJyJKSG3/YIZ2JCVydkxbKoRlJY8V
SbtTiq9rA5EohQ5FEkB5abW8z8NOjrIHTkTPpfUE8ktTwNpYhC+0k4K3uTcjQ5Ny
KTRhjYK+q0Sw5D825gGfZWYxShhj4By/o3LVdlLXrIawKo/Oxl5j/eR+CngBHZnJ
am3p+NMg4+HqeA9wl0w/Pr4dS1RdLa/JPnbvEZvl5jvz796qtiDLaaTSaKz2Tlfd
y6t8N3Kzc/KXezibmz7P/P21B3BU7ZXLOluJco8aMREzKUf0v/765nf3fQuk3ePg
0/nC6jcxRr9bx2bad06T3D8rsWwkWNmLVr/dpDJu5GemyaLKni2LpoH/jyR+uOdJ
yfOIwAgGl2Rk5f7ORfDKdiA/mmfhOSGRxR0ViFSxqpawpqGBjbqgDv/YM3dsnSrq
IWtaeLhDbdZO4v7jJg1q+4GtFmivLhwFIc2AE760VACeACj+LpoVHdj16kp+iq8U
5tq9wKet31TsG3KxT4D7tc/D3zMIHqldvCSFJaHS+LpNXrH3BC3O06zPYGWnV39U
RzjGKe3sOPm+VC+Wrb/Kx4q7S8DJfvGmNxjsecg/n5mIzF359b4E2B9vlaeqgnn5
E0GyKzrP50uZTjzmuF1mYCnr3fbwdKlXE7indhy49ulcCOBRUHo3AnPu6qPStNKw
tHCWlT8x2MvSFqVOvKpzx+vnCcVZOidZbWNbwjJgewl1/7bSuy9D1oNgBkAJJdcL
3fuCaNrM8CZB7Isn8WmVdswkTnCiuwnIgai2upsYH9q6Mp+CIXxdD4Iq/ECAkMZX
ke2X5nj+TRbah5OD9WhmQ896JTCMyhy5p21/fcRafnfcq5xvOot0f9woXx/iCsWN
sK16nSu0J9fdVCNGtOZBUnT8usgF5c5VcbB2zk0AYlZ9lir4MVcFXOj9tKtiK2Ux
K9Bdib+t34UbReIFB10jGNlMrOYUQFCL1epgDfuSeOkFR51iPucriWVZUZJSECnW
xGyB/SbKLkgAPn0lfOYrmCdggMHf3FH48EmNIwC98tGKP6FvmZazFBgvdioDHYKb
l5zNn0jSXfz323Vu/YtEmaU+v6/iZNZCUTA/JJNfCUnQSztAr2LS1xqbsRkyM3SU
esG4rGIQIlheqA8UPrsNRzXi2HTKfCOn6LqbI7vdPL67rexBWMZFkEUT5vHzmq0T
k559vpeO0QlMXkyqrZhxqSQ3nzo7Z+w5kI1TepVKUcY8b/ge0qK2MhB2mkk6IenL
WNerFYI7QjenYP6hklKc1mVfl5JcJj9GrgCcwu0cQQjadN7Ep9dqkbzCc5TnfxZe
0SDLANPyohZid0FR+0drjOIEi/0cO0S646VbEa61/VFOxkmIZRHY6ZQ4qOBRHU+B
OcYsZ5281Sj3d+Zq2RQZ8qg7ihOvN9Mic5uLzLxfIeM3wxZuATQ/nwv/OmT/l3kN
t7DvI+MaEsPT8eqemoq2KlZjJXlg6WjyQ3xywj1qeloU32yg0BzMnjPw/njA0L4V
DVlfuTQ7Nq6VZWeTowXUClyGixks86jdgHmOyMMsPaBeL7776v+Ke7FZK8mm4ks7
BWYVJWEQWrRg59XpdYNITK6W8prJjM89jW8sWuTwHPJOCZQI6NtkpwGt0Q/k0X9D
r8XQlYAdZXrEZ9x1+48zp+kPvmaIUXf6unjI/3okA/aX4paGwqMGUCMq0xXR+6Yn
dBa6Cye31TSyQQkwt3v88C4JOfnyDEoIlRztXfGuWyAYMchqUbkkpKLr3GVHyGu8
1+z6Mn8EpNbLjkUIKPFJGIvZ3bvqUZfhnTZOIifpHdGml3p4fGmU/UKl7mPa5uUB
ZliHMZP/7SUPONIhJX9g+jVwgbA1aHNMimK/YieFEfyT8yH2E+0M+pad0s2SsChB
zU5NaB9FYaMp8xX9sr3VMrcMj/MhHC50V/YsIrf7i2YJxoLRITIkUxB+umm97iLv
og47ECJDUS4umHrVCKS58CiNCSDEf+9aHp6FJ/efWMw33y28XghVSt+RQiRVF+03
Up4XHkaKLBx72nPGuz9n600UEqYMvCXc6Bncvoj0937UdbTdRhOJjhUUXdEfAzM5
FfTzUZ19JQYoVHjkixODoZUPWgxMhqseGJsiZRYlgjzqyOsYvoTnMFofclwOL0/6
/X9Kv+j46DZqzQ0Zu3cTP00PZIs3sQiAT1k342wKNOrpPii4BPficQdslg71RsAu
/b/JMs4lOzjEMb3IJbp6VjyWATGSd4rZWObURBhdVMjh+djDbATj6C8Uodhvy2Yx
J/+/23eidkN1a+TTdvU3Uj8RKXyrh69BQrohlZHyxJP8r8ab16lJKUQmsciS1k44
9ACero4B7yK73Z9gZqP+OZWeixbg0aui2Wcx3uZ5lPwqnV5c3M8K8EawPZStIDos
Oq47O2rN9Qoa4pVsj4FkTe5cdVuKvQqfACU7ijSoBrLtTSiczuGVvgZBYq38HYmY
wyLyqYyyfulIXX72ka1aXdf0MQm8K/pSBMg0UGpiGTX6EMF0D1GtfXstoRTEVpYP
Al4QQYbOebHIj13Q/43UIyD+PTLPFqqaANJ5yXXxrqezQJtKyIjk2nMVsQj12VVX
wSutb89QXaQ9mJ3f97VBkWIbb4kmZfp68R5+Lx4Zw6SlgeWYfM9pp9kPonC2cLdM
HVQjwRjWKSdEwXB0cexvi6Lf2z5WTWKyjIWQBFUR+CUT8K3Cq5rAyhJiz2i4nFO1
sUO2dEKlJfbehsdpAuxK78TkR48U7TUy4xKhk8D6qZ6xcCEp6S0nyGx2ZjJ7VKT5
tzmpPB5QXC8qHB+IVv6MgZUxfAnSFpg3S451xTNa8Ux8UrygI/r5Zcg24eOMGUda
2vHz6y4i7+qzIJVa7p9MhlAo47ChnYQe6M4i9s5vcrr0vBki7rIqytoBKX8eNhzF
Xnrc9JS4BMnIhLNiQDODwRLPepDNNj2nfmbhAHUBrD9L1OpmKfWTIL9kx1QIWvxS
FWb65H8Ky+NQqxRtrRYrBE8h2QuYJMaDQRBvek6v6w5oRLjPGc5ya5irGeG+m3Wx
sxeLKBePDKjQlgGEcMEEiBtk5jDGnVb88PmoS3cf6SbM5jvTVGm/WzwMq37sK2gy
7o3S1HWQa9zN87vHUYOyrmhD3/DJ2WVJuWMAA7QpGVEA9HLGJSxlpftsiqXWdRfm
Idx5H0FXe/W6sN6rzMWrlkCH9G7LCxWX1ohsjRsbLGq1S20gFR8CvEZJQaARbPOV
Fddlp66xtigkSOrTL15vdQoUpMtKmwMvQAjBtW35QWKsBr0jw4K6zEdoA0dmuiYP
wlgjH6v61VYyqK/CpgbP5Xq/r5faM6YBHQTwJSGuyXPQqWr3/Ymmiv07vmIUfazR
1bW42KYgHn+Hj9f7neZ42Goqh5Y68UFUhsU+kTsZx8IyAa9z6rXMHSHcRPhR6xbL
gZzadobGqt1w2xLZcG4r3vNRHaoR6nQc/dw65iqxVQnxOPLbV/irSzV72+i7lVky
zLgNuggp8Pm8fEHzmfKqgi/sCwlTE9RXyzjU5sFEcCXW9BgeKjJmBwijVz9DmCwv
tB25No4ri6wgkPR/i9vCp4EciLXlbi0uyBEBwa0ACOblkYK0FZ/Umo+R51Ia8OmK
y7LAbGPI/QuaWpbuY+Faje1ZR51OkuJGp0+2bpDTfTkE9eiFBX565Ln7tQRHFnAy
PCFVZ1ojs9aCkrsB7tQKQnHA2q+ilVDVvqtuc6pezqsuFufHnV5OFqRTxK12wwYH
oizSxHvbHKLIBzK8jPOaTzx9BUWQ+AqGzol+fJc/NtOZu2DhqjSR5zusn7Ud5ES7
H8J84gxf/QfiIdSdD0IZ/0vCHLrXVwX5JYGD5C3zywLeXauWLVcGoVxXyt9ds3ta
vSDkV2cB/7RYCxsx9xqqwuSfKpMnqtbVaBbsxsb5iUFezLVfRkyNVYqUdFU5CrzH
m5psGXgQHb8tB9PHyGOLqe2uOl2sNl2iQEbJLuWPLnK9QBM+2JttIYXLxaIVWaok
QaMi53ueHsiHAsoFdiWVD/uGJdw3Y8LuK8eke426RbwUP/rlKqRDmTsjU9HgVgxw
Milo9+HnOUr3jA8drI8EZeMYUQpAuEjDXXVdVB6oJO2yb5ZrrwKaRKc2/Z8o/FgQ
RV2FqAwvTMvqkdQciOQP1dK81SGH/Z9CoR0xUh56adrWeXGuM+cF9yPAmGjkSJLG
a0JAP76xkEmiWqR7ClZWUEhiM2ZbbEDSKRdk9zSNDQVg4wGH1FWjFFYMA0q3h5c8
uTS+aDi/RIeArBaVnJRIAK9aFQsNT52aHG4Q2hqedFOXEuqS1Gl703Ni3yYm2OGs
KXnupUxt03FrLf7g9d5mVjtE2c7X41qgIIkgYZyyxX0krnyqNv3/7QRT4YmJYyWE
C3cD+GbBIpF3MXL1fOqP03HsaPl/jjAELDI4ocAQpBswXpWCMyBGYKqs+qs9z52T
ubbLXFQiCfuuxRooc9ueLb587vDOSyniW/zxG1+/Jzsh6hl+8BhQuaJqj7BxP+Rz
wsPtTx1zm4Dtgtbv71JjiZaGDViSFkAGjMud45RFA/uV+B2wGkjQxtywbfwEfrBw
jR4cKy4kcW2TO/I++pzwya59iRluHu2P8UJ6Khrc/Hx9Jm4gV47agtvByUAy3d/Z
fyepn7+cluD37xyuD3riSX8Y9DFb9CWbCK2qMOxYaG0j5n+2C7dX3YtrnvlMrqKv
NBhnhBxoRZKzb8f7Hg24axJCLsojEg9zGVRBDiJwa/YpqV1cWV+odenFJVe1hWJC
TVhpLD4W+YK6yL7lqxm0dk/+TbmYSmA5snqZcY9XdUFuvmgH3Vwn9S4iS5ms0+on
IotI0fBydtIr3KmRn1rfmQnLTq02zQ4pf7L9ETncA+CVn57KCULAWBJc8i0xZ2jH
G5C+rLxap8xn4+0SGEWzBFul0uwoIkz5mxSQUfuq15JwZKRi4xNtoSL+28O7Z2Md
g8vgQX0TsyT+Hi9mxk0BQeQ7jar0fbYAJjrneY5zW91x9j/LLSeIa45x3BbvFTrV
rAyHrXvhZmhgZo+V7hIK9EPBv+c/HNXOtmaovue62lkWslx8aQJ0ASmRnYwIajBK
u4kzW/LBy6soT25U/NmDV2MlVEB8DfK/18v01VmNhIvNgE1Sf2LWCUey90OkxwBK
2VaKcGB7M/3TRv/KCww9Enk2flnpnEFUfHRmFNJJzJwF/Zy2G7mtIbgdA5OqUrKQ
PqOCCvhK0Ge0BjfQvvb1Z7JTyR71MJkJ+SF9/g41AdqnKsOINULcp08W7s2HvcdH
MXNY88aWmKd/rsADjzLMII0EbUy6t4cQ0MWVfwIcdIIOcC1RA45kb1+O+4G4c28D
MI7r6Isj9Zrti0X9/D+UZEhpKV4v57j/tNi6RV4Ik4n8sbr+DqNCZiCjmf60/yBJ
1u5FE1ZWEWt3l5ynRazRt2OfU4mMQcdyYh1s37mjuPV7MHPElX9sTxTwCeDmFp8s
TtrxDCxMGUHVuw3sOLLUy9mfFaH7y2Jt2Ad+PRf8IzRD8HtEmp3H9KRlQHxfe2O+
GRJ/CdcG6Ev6N5LIyO7+rnuDmbWP6eEdoOU1loHo4QqL9ORZQItOxsHjOVkv9Wxr
bMOPrv+kKKh39uKR4H6kayCc7PdkIzQY+GiwEkqCSsyVi424IgQtiznYS8Z3A0xc
AyWQrrfILjru77lsbhPdcUk2YBNmT8a+wprYzGkmuuSmZ81+eoqEEbxo7VE/U7pT
f54BYOmNuFSUhiOPjh29rV2TFzHrOxGoqzvM/hDvH81gjSlStUiypKIfWXvjuXlE
mACq58fmmfYqO2Ml8r7Acznei9g3fbBW9ZOg10pKJ1t7gSqLY8ZAHym+9+2FVKFa
YeQM5tj0/tuYcAP3MuF7VbuIQWa2RZIJtBsrzDVXuUvMyea3wgWrwVZpbJrHJvsJ
flBmneiF+kqcKtRfU7y09jEx3YEF7tfWzYTMqNNXcS0+keq/zoKSpaD1qI+auN72
U+4H6lxZ+gB7//D20+HL6U2cNWPsbMSlVRWHol7P/WD4zv0yl9lj4fPRmpORJuZC
9Fcjw/LPtAzFMT0yS7fVHbQDMqudGOk0EI+QooFO/cgL517NopBVrAIj7xmUaDI9
vdWTr4UjOuYOMS+reB8MLs6Z45PKVQjJ7NCIVRhPoGMhWJC+VglM9n9ooh4jbF4M
iIrvtY2OD4hfIr4keDFuMFOns3ULoG0K3yuYZ41tf/73eQsX1BN2gcDE6ybxQlmf
7FY2xdH//n9pSjidd9ltR5r7wgpHrVbNZlMT/n0rMBm3EZunr1jqjhu5BQkAovTC
weZNd7SH2Zfbo6N6NPdcQ49n84ERqexX46PQgXLDuyP7z/9gB5/EEzNcjq4kPO3d
sL4tzhAQA0tMNehRTiC1YrzdvYAJQBdJo7bssWqG+yUoJaNSyP50hWrftx7vFO2z
CtehC5Nbb1CNv5VGrlUUv8pga/Je0O8cH5FWKhq0URW2YH2CvzU6WfV+ClkBXWRd
z/hqNkqzMqq6qWKiY7gTcq6xM9hJFT0WAloNI764CdwOkPgfBpDfhhZ+cnFAoI5J
stiYoXyS3Ks4cgSxGe/Gp8Z30tkV8hyFAtHMsujfSRqiljqHLetyKoterNtO34B/
20+6DeqJrpA3f2koZUfqzlwYjWrKkr0Wm7EAqEuSlrD/Kt5F0fzLFSJOsZJZZTnZ
hQkuB9Q80RdrcZ7Gldvm4nStMfS7Y8I8FMaMSdDE0IF+3L2sALFRkNblx58sH5d0
xQm8r4MPBbP2RdTLiL/H4C3wAgqCS+QgEYj3bfda9QvM819On7GQ/sbhp6PEV9po
kCpA8ErtnLXWlm8CiMT/NCnYZP9n+HSYchN1L9FQtDtwM4FflGqWSJPrO62QmFbb
9rFDGkyBMxpGAgkMJwRpAR4bpLQeOIDO0lQjQsqx/f0CnNf11RyEoW2VePpnmMuK
YhjEdOW77GzJW+ded4ow9uKM4mzcrAHdt+MecB1cSB83LX1b0BX99/+jcZMs92E8
anSQLhW8SYQuyWqukyl0T+z/qU8K7v54+Be5Sy31G03gcvF+1xgvBeSGO8NUPULI
v1LW81nDaKzIoi6ZdleVjA/xdfJXNHiFPpX2ehV+DN+w6O0JYiABPO7/xyM5sq4v
Cfv2xsZBgmOmf6Z7pNcbmQd4h0EFFLAk7q34+1ZRq0jcgaCFXz3ISQpRyvVcUrAy
jJCsiNc+XnNDrwZSsE5g/dYuNuccTycCsXl2PSFAsxuIgKdadZrzD+U2b+tACDXM
S/ei87A+Mofe5n4SujGAHYEZaljiHkOrM7tCL8BIXNap6e/eZRPyvqlJPwSowTQT
Cup8qOhx5cWq7jYtW/pRNsYjERkfw3ugfmzMPBTOceraeXUxV1yqOuIo9xzOdeJk
15krXnp46LS/ET6KR3o8ZSMfCtl5C0UA9gywze/Cya7NUavRjbo/e+n/hjRfUj+g
QdIAXxdCEZ2vxu97cB8pVM5nCnIvOuumQkGALQbJ867nKCNREOW4/zxJfClAEp+S
Tb8nTYGQlYqnGARCetsLVTLDu2M0i43nu8ch8naA17WElUalNbQoRDCMZBJlOSe8
RUQp78oyJOimGlZ8U7C13ds6vSap71nLznpbeNC+eLZkevvUnyoMk6SYQhkK9lnv
00ZVjbRAMeV414jQ/sq+SPZyYtzbi5sxzcgt+eKi6rsW3VWcmj3hW9ZOB2xozEgA
gPgLVGDisCV3Hu1+7kcELtJbmXSkq3Dnr5wIdEOYBYIii+qEsYk3VPoZb/szdQhu
c2+elD5ld/vlW496K3LW1nW2rtxpVM5TOPR6l97pn793evMwRXDOOaqOwh/i2FX0
rjqrEGSyaGSRJl4p4kA9ugnmfLeAlZ/W4t2gRhhKe5K5e8fsOq381W02VVPyYh7Z
2zqFdgQCZ1ORmgvpuRlTEiqHrk9TtdzbX7H8sPPSvrV2bpCp/A0U2zt6WNjOPq7I
w7EQ0EYqXY/MRCVkQnZ7fczqbrMTb4cut0ZeCRnKSNgkHWSt7tc0A7yKbCOFzU/q
L0EeU6jqoq1kaMqJx3Y/ic/F4QqJSMGwG2jN2xrkahwWZEB1umSFORY7bGeGj8lu
EccT5Otyd8u4tFB5bd3VeMGIa2iPR0AmLRdo0r9TwnF2yE8m1rsLgvCKY0OILJRA
LG9sZODct/KqVS9GHPhCe7+CVCKinLld7fRUj/a+fK0HAzCjofQ8WDLsJsK8oymT
OdjOZGityzDFA/pGX3gL5snQu34U19GPLEiruFgh3nzvg4y5O6xA5oeCD/EC+qEn
VMZjokgVaGcO+rPTeIofkgQyDPft4rX751baEukd9b+UcuGDbycDfb54MRXDEzKd
jROcwqN89mCdTNeWgzrqj4C31OKsKE4sowOJp+IhjLzc9tF44RZbFjyJBxG4/XuK
7h74QO/C47bPjzwsgtenKUP1eeaakmVKdHmHhPJS3w2axGM7BUkNnaMz/LlL03yt
RIVUn/xHVwr7sU727tJy6Qz7M40tePhaaW7bRXmQGyeRQ/gyxb1M53ckBa6JWmQc
9UESI8eFEc7jHnH/QEoPSeqdyEi79v3nq7N2YET0DHDKflqX5ctV0SpAGfyEkwZz
SpZpCc87nDeMALFJu3tUQP42w6zX1cnuh3y5G6E7e5JDdPUeTn+oygtr2Bjgw1R9
QcgQuKDMMfxDya0uepewYYDo7mf4U2hcakGC5lDAyYcjnUaJad1xl2o/E6ZE5Qjf
Q9s+ys+HCnRLbNGQ63R94bueQmWNx+VagaUYzbkHzwuV21Xr2zRxBkq1ruFtphCg
gE+OZywBs8Q3fRy+NhoB7vCe5plSunivz0df103KtT8wQ6l7/E0mRzGoeVpx5Bc6
8cSyydo6ek8DXnUCECieS+8mnoO1cr+Y6Fu9poK+lBhPvhAUywSvQCH2ugiUTI+X
C3cIIl8+Ads0BAFMVhu5w2MojsmwZUrEsOYmoGKSF15avsjvaAN+jUygF/EamP2R
dZCVntZLcGb4uzNOm9baSPEsa2Wm+eJDomJlOtGVzx2JfT9AkOClAiIvnTjoqKNB
1Nx3c5fmVaow+7jO4WkGtEDtMA/SD+rleOc/bNKvCz9MnHj3WSdPeRGEklyHIySW
awAxgNHBiaJWCOVwT1Mf12q3dcP1YmrQEpqqWy6yVQZoMDz8Uk82pw8RQbp33bA3
rhZFRg9KSqEVfgSH/izxGuBOA5aMqruyyqbjTomeqQ2qgYywI+918s5uxky2IAPl
WI+Mkp0wUWYernV3m5n63xvNPnR57l57kvT82BQOo8kLqI6M5P5OiroGMhrBE2Dg
cVLueLec8wpj/E8KTTB0Jg+MwNKDzTE2wIky/ToumDWuEHPNxlToCiwFVs2YN4fG
VFtCp3DufGpjr5wnJ6r3c4j0jIFbdDwLObxUr8SiDMiNFRaX5x3ugyMcWliFalSU
uokKDFePdDHbg199hpo2mtMJ/Gm4DGDPwpHg4YCDFtzckof8ntxFFbBU0I89OfTE
P9/3qpplr1jK2eDQfxeyoT3vp+AzQhO5cCVYwh+AEt7PoLiSxmRd4E/WCy1IVRtf
lC3JJ8hDsI+Z3UjpEEBWN2fmLFSBhFx9ar6b6Y56AatP/woKlg/+lPuRPSKK3HeF
Pn3EuShXUyKCUV2+0fOJxC+ZLG3HqCtM0SnpwmfaFnq8Be5wOmrAMxmHjjabMqPw
yEKcB6KAVKojYOHNwwSbNUcPul3JFZNbATcRj+dtg+HhymrX43cFSQf/ca27OCjO
SiKaOf7my8KIVMWB8dCSv50Vt0S5t72NsX7BtBpMiijrhYfwENdmNMueGZYxTmdT
yug9x9mQAOT5yDEKCkfC3wqIZCUEDuTRrrHa5i+QgU+chqV58NpXDtG1mpIin7dH
pJPHazhvVKSTrntT0g6pFlPBmSH94NLzkxlC5rR06ytlLvFYCDx45Jxg8PY4E4v2
RJyReiMl+Np+Mx3RwSHjpmvZZ+jvKFzEbxreOs0x4CIGtV/tMPidmpyQH/xmRzjk
CW21eQ+A+6JsPOFinMoio0q4VW1gZCqjwB3s4QRvmUsma8jWB35QdLfn58boC21p
nzvrfFamhgZzVov/Qs5cz55rogzXuPm3ndA2tn6p2srlq51b7qzwdEWOYXgzYLXJ
PRVEVH8iG/lEXvmJw4b1TWgZ6cE1SNlpJfrWHqTwY3CFrYUqC8m6tv+ws09/TOZl
BhSBW1aHQRKmI+5LkEM2i5cY14vNmRRIf2bJHayjKZhc02REa7aNxcDq/Auxm1XW
k3WnoWB4b5ApmWRnCqUmoemUWSIhW9RuXQ1adjZUmvZuId75ctJPTt6o+CVj7ROy
w1a1IKW+GnBRDDRtSBnGJniWEL9D2Fg7ovJXfnZ0Cg96mH1WqBXuNgHdNCZX+OIl
VNSaZWvaxVCP38rv6fd6+/1KjHDrmdr9anGd8qnHu8QhJhpLGynegZaRUA+dB612
/6PRWhaxO4SJH+ZLlniQisgcppVcdPHdDEHD4YapnqntTbtE45e4vmVNY5yiuzSY
exTVvEV1lyxLFv1y0FS0hONf9qBEQ8mcaj/ZTBs5KyORG3HZYUtyQzbKgaIRAuwQ
3CSC9z+0RoYXcakke4Cmo0XsCMIUkvrRDgvE94wGyE/2aBWBlnPT9xmv/M16uHqr
RwyK9JmdKFyZzY9tBnwJnR7Q1p4si1oh42cYYiZFVSkCLc9LT04x0hxDeTRuYWFi
mZdo06Htn8Ho0+GYF0SbobBLo47SnHpDpSaoiHoA7nCNOeFgDl4w2qosHAyssfI+
ckcgpii4r8gk0bjtUHDwWcrRus8hCCC3h2VeoLf59fc/1C1ZDB90/o3hPLTmlu7H
JdnLSG0VyPfs5Cq7jgTZw2Qp/FZw/Nlj/TIbUCUJgeesau/J3nznCVZ/RouYW3O+
9UGkuoHmRHGhZ0RFJ27x9/ql775OkfL9AEx0zn/jlyv223uh3VD48cc2SrlTBily
VNTDDxiCFqb11COlcSOQ3Yjl1UyNmybai4ow89IYQLaBETkNGYlkh72d8BXl/3qN
Qzty7Fj1SP848BsjblXsfxGbOTfH5WdyZGoL8K3Dfpe8cBSsYscdDluHgezxaYrC
IUdDa9g/LXbAq5GpFt8KhHwiN3LxVvTwI3HWb+CPlzY7ucmu1C5QxXUoKtT89roj
Caw2na/DKnz7iXSpZ8poYdRWyePMk3z3KH+LkkJDx+VC0X/19xZAeHZQ+jazWpGS
xIA5PBFQdXvYHFqIRq//51WnRiF8a6HWr0WUcY0N1A4oUzRjD7UAbsCNEKfRkXVs
D92iA2+9pCDx1eaxNUur4S2szjSX9Xxytt7dN5QR5IA+llN/exMitVsPXh5DcAUu
Y/agsyFG4zfg9ueNh+gaOFIspHW14cdfRoyAuBaKoJL//Tvivh7VhgfEh9ndrAIN
Uel8Al/CFWFeGoY5IdkvoInfoIgu77uNx4ptKvZLTORfwCx/jnl8KHlopkLJlZDC
DnhLli//UPc18DxEK+Z6bOzCM/gw739DhFuL5yliyMaiLz4ayiQBBWOvZV9jtHJX
7GwUlldU0a8sGng7sPeplepMCrI7OGjnbGuTY9aDNX5nyy8fJmf/UirmsAdcEZiz
ZX/qJifPS879pDGn+peNc+rYQknCth4sGLISOHPX0YTYWCbol7PAS2uhx4cH9P33
bQz0Ihnncz8Qj0yzWIKL5TEUPTtNAQikdU3gl6q6LlA1d8Q1HJDpKl2VEOa499Fy
a9/qqOIIQVopunFRLYS8WlfPpHrmpe6BAE9+GXLIAzS90oqLE3X8SwpLxovHdLfw
dCxWP47LXdY1PaK+3u0oR4BnzVZGSHcHAD/EYbOcG3IhQSAsojH6q5mx+XCWs3ay
TAUZBWI9NG4upcFBaib5FH08ZmPUx3eT9P5XodTXbFKNbuHJGnsDOSV5j5Ua2p2e
QyIxf3S6++e/sfN4+plKtkvvmqfrk3M2V93O550YK0ddocoSc8xDnQXkBwU8KX0C
+2WqWpSjtN1fSpWtDHB1y/vqc7a+ESC2mX8QTe9VZgmnvr70ZVe7crqc9zco1rxj
5bRW9Q5j/o+uNi0V0EFKlvvxe+6WTm5pl5QlNVVrdnjKnGZIFnyjRpqWd0k5vEo+
kT8Fu78NwS+rdaO3MWt/9UFYSnHZNgc8Ne22GCiMp0iWSUjtypLbfHM6j5Awecta
+gCzA/SkShQYN7eZQHcZ6RUrOdCF7oQXdmJ/HxrmCci5jZGOwttIQGx7VtHiI4ao
VAJ7LrY67D8aPTx7Lj3ZN0UE3XVgfyX3JfyRO9CctivqM+aqH7RhyMFrlhQbo3Qb
R98utOTax01cwAcpZPUrV+EXKaEE9npIfIrac3n72jIiG1QGCeiw9ddhT/WBFFh7
/lA13bxVhw6OAnlbaQNq0anGZuRJZogxbEHauZv8wptFWqJYABBGTvhEaMjZx621
Eho98TIM5zMctvKiey3DJdvnvhe+nwkcmmrs97defKVgZDMQNR1EL7duCs29MHkh
FZW4KxOtV2w36t89fXS/4Sg6r2wFvS29K/mzErwaOpum4ka2XK1UtWYOTZACoDU3
Z44rlJQlMcGYJMqp3h364eaP76EF4+B4Rdji/NCIzaa/DWU9YwYIqzNfeQL2SBEr
DZmrymN1fOQhpSaU19wDBsUReR6lxLoNUqWBcl9pMVpgCptNGDfCAV1kW+tISivM
+dUoqL2BaDxuvgW2x4eqZp7E3INp4YMGJfxCOm5D/TkWvaxS82oS/WYE50ZDXlZH
X9Jmjr09bQDhAn8uZUAa207qFbb6R456KRd4BAj1u8/p8gS9Gz0swVRZM4JylSyD
ifd7JYYXu7SxaHWvSvGkBrd+xcjQkRTp9vLgSiubtkCuiaWBe9Ntf7Bv48HAVb0p
Wd+L7pP0s/vVxzvtWZiLPoYI/xtaImOy71D87DGS2XayaZM9byo4sYEuYVLsn8wv
0Jad+UgaqzeVkpwcwMjwjn7a8R//LZqKJ/Dpce6CXwLMvitpt0YA1PG3NmPPg+1Z
XHxOMKfNT3w+O54h0hn2dJw55Dq2TIN7UpLS1GgBdcOnuWIbJC/oETn8OAd8A/tA
wuVtfs4j0yl8xGUaTyMXLqolNaB8L+52oVbbDv5Fr5rigOT5eGclqfkZEKm6t6Z+
h05ZMtSa3psI97ZMvz7IYmEP1J4SP8xTFGOxTKjIzp147O2invsiE7wuIWnDLEL5
pJWCZjYhUXoCKSBRpPo2MngUcuBE58HKnAAN6EANjEylxUSaScgzp3WdixQu62HY
lY93ZZxK4brY5i2NjymYz4WPbLUD+dx8p6iAZCfZspo1rnq7r7+R4jwe/ORrUS20
vdGWvPg4Q7AbRWq6ecEHa1dsX82XXzStGpgMboksHl4yye6Q8eDOvxED+oV5Aa9z
0XsdAbd+ormtaRYGSFmn3z59VZeDmm7I9cprA0W8IcYnB0IoEZEc3EufOQIBaeXn
d9ACy/u8tnyELt9+/DQ6hpB1YDgzkD+5Yw1EExGdotuOSPXvJLsfRRVxKy0pa5/5
0TsStUosCd+cdpJiXoaUdi9EsWi4tZNMWvF3nFWJk4/2FKGnLYZlQpgNso3qMqce
CxVU25qNL9xdkZt15PqYbgThZnRaj/1A7rfsf3hGu0iJikTYi7nHZm6EfQogKxzs
0+SXnOhAvQeNo1eKKnWRG0YBi3PKhmEH5sa1Whia0VgQuTQVnPxJid73GN+mHXcw
NJ2x+TUOiF6f/3EBcpOR+/mKOpMwge9srClahH8Zhl8bAF2QpMyEtfdEvF7MeVsZ
un+S+vj9IaXBIcmhxJBY1x66d9e3PD8q09pJuvXggsR8zdxlNn7osDdRNE9BAZv+
ciGTzVlovy+0z1+uHQ8m3X9bFMw+d/mDhkRnTVighcQzi3DKonHKs4P2Y1mvMhrx
TodsLK3w/R/FiF9L2nepCQMlJqPMtLskj7n4TB41QA4ti/z5zJ3W9fNvdorRqtOp
iZOodwfpfK7LAzPRk6UPfEV43eV0CDhyHqmMnTESIUiNwb6z8tj4QKVeJhvtmWov
ZOj+5cYZ/Mp546YD+ntvnIhJUg7hefMbBp0gmcckWLhqWjI9ndMAFdmwVRMS9ggo
B89au+ZhRySx8Bov0NrGJEMcTua+HxMJ4r20o9FfUr67xM6hf0dU2kjV01p07ALb
q3OQCEnE8hm4Thcxsx1FHnVyFS0dKPtwvXk2RiGSZpB5rMJi6RZXSiASkVJ0n3rj
qnyelk3Qqb7uThzhp29J9qvOYw2SN3QC+pZBQVeMVSWy5eOY650Sz6FeozB1WUj9
F7VZkZP5IQ7J4PbFxOqqtyT2g/vB1OQj4rJe3W1DUF6Fo7h5QGg4+zV+RU1vN775
VHlPzu5zClt5axDTMAAC5RcutoGA6f6HUv2saVhScbjrVanlg0oZgzVs0fEHV4hc
sZbwHmbZoG8/wsNsN7YSVdqFZu62b87XuBYHSd5zvot3RotbQzqwp3cZZhN9LlpH
U7b2Lr9fYDMapiiMZfbKU9kugM39VU/3AnDxiCecPVMsCXDftxm6ZCeHcu5u5gUT
AYOv3spEHYUzhXe2Hf9XkvroNORcYFRTIBL6G/2cAtu+wc072n80D4DFnwJa05qM
XBb3DkxhlYvn61pEhRZS+vR0NWLTy6/Fl7MDGwBArh6ebt/NrZhsjm8NmmU0JBCW
YnMmpePeyiH8k8TVAqi6t7gXLqtgh9GsRqNXPMcbzelfbRodbGiUEFj1Pney5aRz
O608FOIAnJXW/FOO++ZXtbrVXCBIOed8og8RUBaLbjDRqcDYdVAl9WwC+zYpcaGV
sqIes3xfRHlpF4vlOpGWYDD1jwaG/aJ/2hHS2sujukubVLj4ATwc2aPS1CRKtNdj
f1PO1jA2JLWJILFKD/BCJ3j1B+A+2mAjHavwhwb/gd9d9SEvhFP0G8MzgNpmLb8B
hNXYWAyY24W5fdWK25721CNDgkLXzMKRl1Vwrhb9G8pXX3foGdO9tdYOlFMQezdB
wGOF4pDO92odBf2kJ37cvkLSkXyGXkoKmZ7r79L+keHvMRToEMEO89zb8uJ0blU1
c8Aztt2+M5Z7UrRn51Y4IMmRirjjJ0elaHWov2Kr2nREfIfoYGA5AquJh3dtZQcV
NgPFC66enyS4HS9DeKEcbORan+4egIVtYCbrbGn3te3KyGH+1BGypquqLWDIlKx8
XpK+FzzEtpmzCvyd3kNsdaj0v2y+EipEecnnjogpNwGDFf3OXn5KqCct5R/SsHqf
XfgwQH9PnNe2PUvsh2roQMSrDqBd1oXyRWBep+Zym+1rrjyLvNH0eWL0yDt3Wxsb
HNkyCEwpE1fXE07jTT0bUUOqidMi5dGtiXsjIucp9e1fjhmu1HTKp8FXMqGpbgYz
vyDdZBaH38+exWC0M7vtTd8zEAE7wMY6PteTluqtFJuLBZzgv2DGZYsjZWoHHnET
i0wp9ZERwJoUyiX655TzBpq5A3QNLw1C1Fl/mCwEo/XozLPv/Ly4aEJBJ6+IXUZx
YQuPX620N/ZugLpfrla2fZtPP6enwbkr20YE61vWlTOmaj4FgceLlrrQ3yX8C2zK
fP0/ndOD55mayus4d3Rw6oT6sbUxUbP6nE/nFSnvZEDHklhHjj/MBtTGBE1XBpcK
taqm11VaoalnwmJ89L5+vjUAX7lfypOiVJtQUsEKt3AJQKEe8gxNA9MF47suuAtT
emqUCXLM1h0cmuXS8fcJVzYpYmzLtJ1GkxqFs3djIcLBYG82liWywT5PGM44Mvmc
3C37XytRXQCGpvjXUQ6x51KA4IqpldbNTAh//nbyT+FT/aakj3N6ExnCEdeKAuIt
VW7XMcPxwBxaoD85yUgXHPCIpb9kqlG8UJM6jmI9dps4PbEz3lKtRsIW7pA2fIXp
kZnauC2MrxTAOypxi0S4+tMXrDKWF23eOIk82xqi6kAqJw/LSETM70c82GcxAc2f
JxUP5+E6mjCxzfbvQ2fcs+UpTugCc0/2DVE2VUHSaX6XQfd9Uegnz6FPI3RFVC76
7TKPF5DnfqLms5WcFE92VkhTBgGKH+/l+81DQwIoBmP4yKp7llK+InseddQE7yVl
CMaX6n7x2TaKdThSM6FAo/IToLKbrRccg4+OfoDG3pdPmvH9OjwJg5yWARGjJfv7
xhGFaYHANmexDuhVEPfZA9rU3/mt+rn5hfRE7nWB/30nTfe8JOdT7I31lf+lTksx
F5qSxtLNbhmmNWaatWCONECY/7jLSboZaQAvSV3ywRRd2mb5uz3/3oL6kZOqf6ff
6MRdDsC4BuHEr+RJ+DgGB37vt/6exENZDxHortNLZ3/yIMhUEeakEdnSW8nKiiPE
KsbqZaXn80NnOMrV1e8m73cHxFlqfLB2NFOodJiC+l4yjxip/RAMeoNAMD9Aa8sG
FdMgvaiJqIy9Vf7OhtotdQUSMextzsbA7tRjDm7WsBGOChGm/6v1RNZ8CWlsMJRf
wPOrRBDw2i2AaBIT2sS2cqJhu5PMRTnWYuBQgHg2hk717u6C3U/PfkENv96Dzsq7
LB2W/ug5qVD/fBckt5EOGOnkdgP1m0LALwZuD5pPI2Cvp0oc6EtdG8vNsBB5uv47
q3w1yZ4L8qhNGItLIZLUy65UeDwD1SiKHXw4dE5niobyEIGxroL1dXGSexg2gIHO
2ah8rcFZYjc3nmA1uzbNYvm+FYFY+EGyxgiJc13Dw5GehVElGy97DRzoXkqeEKcP
hj6ugiYtwkWA9OsKcqro6JBhyhCch9yBBhMuXvfB/ankdarLhFU5uTus7qFhWj6F
+AhSg8q8lO1mev57+Aceh6qamGq441iahYQETqCwhCMJXuE9HrLnb34VEtJW+zha
ZQRE5ENbYbyp2xrwIRCUvI4Nzujwz9LYNBkTUkS634HHC104crA1FHQbl1mnt7FG
YBgvUXpyNquC36/E/tdWDqwYVH2qt1qfcROOGmY819Pj5WJvyK6GyxdbgLVMgK/P
zJVhId18k0hd42Ls9ya3XoW4V0Rkg5UKmTJhi5gNPo5up0RYsfGDD+ld8jJn5Zw0
I4zVbI5jSFRg+CpL8RuazicPX+UKtHaUxtfHbm14uPK0FoIIjbUbL+Z0aow0cw43
BlV03iNceCY9sTaj028UWUvIUrliKWEDVs2e25eFBXi/TkKUZWallp2nEzOZwW1Z
qjgalpxzXy9eUaRFh/yEP8HAWjhmXlrdnC4o6a/69wdxBxpRNwILhAiyUVF8qdPM
JGxsMQUMr6vaGVlzGNhhmlZYhqgnj30c/o3dIvw4wWFlfx0kpsiP+/fAJbduIV4V
73DyUtuFIkyc026ZLFBJVXTuapkvbmmPDKaTYvPSHnya6sr3RErvzaqpB+Bn4PCg
3xNLec76YFWN4vLtsfzn35O75SkJoWjdLKlfYJwxHITBzs4ZUHMiXbYNZTPFLvh2
ggqnAez00BJb6ZIBh39MXRuLfCpEVyTlvmnfS1vQlHP0ab2Pp9gRNf2dTsmFBlPb
7AaSAb6D6IusUPRBMhqf+l5I8e1EzausQrNhhZ1hWYvrprNU2eL0BiMu/aceS2Pu
gwh9DTO6cOva3MywL23Lpnd7HF3e01UOz/6zcp64ixb5J8Z13GzHf5qYTVBnE2k1
iS7mG55uOPV3aJMIMEZlVTh8/5R7hhGqOiJXzl6ZS7HTxrQ7eqEp6/4fbG8SsCsP
AxEgB4+Sl3aWYMHNxne9jHJ55NRwKzPjbdJI9HY5zv2Kj8Oqi3k9AtfJ8HOPQImS
b+mu4GcUY8tnywAAa50lEY9OfjclHrO2Sa+mEN5anbXUpKZvk13/V0A2HMvi5dds
nOFWNemVtetuu+R+G+PrUwtOHht1TO12sQV6gmsIJelXQfeGKGVeEt+bZZA4kS52
097hueUDMDRZiBL7DY4jt0AHn0ZLL20W3W1mQM3sUNaBlA2SexwVNhQyPgexhIzO
Qj7BWCieDYFrTOj5o02GaIghtnrrhFnozHfMEBCvKXRFRxbA9CefPaJ+jeUh6AdJ
La1BRmfVFl8CmZtra3vfqHfwWoo02aOOXLthwxDQJMJOqVh+OTNJBcH4VceNK+pA
BKy3/Lcpz+qUH9QeNOlraoORsoGGmjtAJFOJcAHyVUak1/4KzkN6jRRLvZU11m89
QlkGhEmP8gUBTk+nVj0Wi8eAeSFFNmBetJITdGiZAVJka9ko51ql4mRrkp9wPNSW
0TarApYnlNoT+qZ/3nGUzW0z+5fyEOJMrWzsjETChQqXIRH+2/JR1d8QHLvI/SjF
txBxfiTMzgLCVsjtZYXfgaNu5NkPW+dfol99fFheVjeZ0TsWfKgrc3CACipjComD
JovwJNgiAjYid7xiylyRkyDQpg741C+17bQgZUdhZKjtP4J6y5phoxwdToJtGIqV
KMcz7ERvALkO/+aqAZizknOYF/80fp7JwR88iTeIiUPK/lr5ZdvW9tlWUn76ajYr
BK4zStQO+V2D0fZ9O8xSFDHSZJzy4Bz9F6tOrl29PotC8ejDAuK4wC55drjkKZz5
KwyQdabbVLajpNOkT/HwDsQ5J51tLQZXj9kHzY6yula8Pa4xt2iebShNf0SJeyxR
SEhWL5ndWipGguPCkFQiT9nSzJYl6xUGepP76ll/mLiKjpYphV/tG3rIiL123d7/
vVWEwI49csKi/S03E9NCNpp0j5INHlSlCZA9WxoArYdm/cSGeLzLJ6KURngac2O1
lhUxpqMNSty9hZiiSEItZmKF5ws5Vpa/h6P3s1mzQrU64moIXY/YOBmIYXp2kGd1
kHKgdJkrbhbwVg5G9It+oO/HMZCA3vHRa6pYuEInVFwS+3ocoLLaL/ibTzKeATna
90nsC2p3Izg5oK51QvUxB2EANy+FebSQwxn/TyY2cU/iglQjELOfnkvwfyb0oC3c
t1ykxAUsElxhk9un0AERARiq+qfa1wljlLZtn/delUZDle4InrU9qBh9Qve9aU1g
ySlNw/o+KR2hAqZ+uHKeacwxzK2+oAlox46lfDumZbY4HI/q2Yif0vyFBmF8r/jN
XNEPU730H+ShKuUeiXxFuY2ZpU8YOTLV32tqwy/oxfpPPftqmfMZRH8uzsxMhmOv
iLEuE48Sx5OEZjSgoz42tB4Wh9TtaDtX5nJBr5Cvop2ebI0g8HJ7ytPiRRsVKJMq
cUxcmZtjDtoELpqawW66a80k+OvvlsQCIlr5wPrcsGcEW1SNXqnLgxuLncehYlLV
KTsU+Phkul1cko0YoJ6413uzrLOh3lLwvZwdH/v0J20m3s3WQzzZylwiVDW5l3yZ
Zd92I6tgStg6TpsCl7hLp07TcvImugz4JO2n1XQF2OPyV3v44//yZz3t+whaQunn
RgEUlNGveLAaL1fVclHLDvhvLCvT4BuxuLSNL8c0eQK4jqGlqpAo+kksLFYr06kI
IPGs7ecbyYVtktUQuaHhASQOIOyrd9f2Q0c942D68HuDL4hn9ULRTSop5UI5wqDC
wyQ9tQ1TFXvf1Wv4LDzw75YD8RkqdleeiKm2tsiChSC6Au2iI29XNOZJuf5Q1VZn
xjscoDwFaRJn1I2h7xHThFxz27DfnocSqqI5Ba+CaEs1kKfJIZHznKyB+PCwMG1n
o9kdZS8r0ptRQyo6xtyajrCLJF8HPIfvdjv6/+/lllrAHWzrL7gwjrS4dKCCqNMS
BYM38D+LR+znqTBevLiPAHRT3ZgFh9Z7N28L2UXeZq9UV0VlPcq7OmwWSJGJyK+J
0Gjmc8v6SMSCtXogBDbi/u3fRGeO7lmgLZDdEzqkvdp/LS4CIZSW9x8DqYy9oQl5
eCl67VcPn7xy813wKZoi6LqzJzaP98lleYvqQDWP2v0e6vog8tw9Fgpab2N1/9vl
Q4CiHXUaa4Y9WUqpdw+z9A1jTXv2VsQpPm1Qkal805VUgO32Zw5kgQsxbwUyke1S
M22LXXsl1z57O+zVOPkAHtDpIkXrW8vBkw5JoyWDIyz27Z2IAkweh6saEtPteX/s
hXygbha1MmV7GdCfz/k6xKpbJ/0X0K5MMJV1kwPYpu7JkEjIWO3FRaw2I1+hxpro
ZNgs6PssKEmPvpQyzQZDjsaKRue2J0BfOYpJgNAuhvksfZaZ9HlTn1dw4aML5Qsb
gNoP7YBw0yi2iGfVv579taAxzILEdH1hbGScglFhVUdH/ROihCOc2sMsgf8uOU4h
NtvgJRyu+3qYHeaRBjo/VgdAZOQb4TjYkvwvLP0itajy2m83c9nOQKPYXUCJ27tc
DosvM+TKwZCECipFoilCaPVaH25DTw85RY1sopRcu/WnoyaNChF/8Uib+2SyTVmC
Jx+mdVXWupfq0j/k7AtVOGSECrgf0h5yarNNEfGcWeoTCyFdk5lOQLfqQ0kAlmz0
yh7uwkWWVqp/b1sqSseQ7zQlTi4av2j+mvqaobe/U+XdY/okHanzXFtiPbcAGvkP
k6YI73KRN9+v7iDJSoYZsawsE8BpzwhrRzO/xQA2fSqRfsy7MeWMG5ejQxVSYhI6
qicf64H4MLgN95YH3EA6xYAjZt49/LTBE7o9JGIyWFJhWR5kWqbMb7E8pJPsSMTa
wXjporZ9EH0jXfwE+Z4afX5LIaCkDL2nfnV4FsYSQUCxV9gcayyl/BKkNhjGyeOH
2aKSlm5OCtxjgWe5A4c+VZ0HF1qFwIl1SmvdqsSId/m2FRMo5oXlFEDs+Y6j6Dw7
vdQvdhMq2SWQLL846QUgSKOvLCNi7RKoq3qPsaz6nECGmIGa+TbqF5AxQLOrcgZQ
GdlqoSjcW3UCfDzLq4PpwKIp63KjfD7yUrDhgwwyRd1tAuavf5Z0FyfK6vph+Yf5
tXkEkdWg7U+1C+BcU2cBh8afgo3JYOOVU1SM+qKjiRyKv/HF/JMSFfgndl036mkp
wBSnJAdvtfai0/E81yRapuaudvkBWASrIvHndrK/9tyVLp6wcST+aLAdg2ILnPVe
9GP5QVXxMcNevbnI2884hMLK3DMpxvdjkfvJD2lzX2Ytx/6/ixA8SSnS7N8XVr03
OxxKxzdVC14Yqr+uCTDUyf/XqVQe7uQ79Ahq2B4H9agdiCPu8mzYEPfC6UXzLgs+
EKynH9UOdahPc5bA5//X3ZPvJRPAPbx3oq3HyDzDr/6pl32fxn8zc4gGpJvIXRPS
1UCOQph5Uo/4YMVx9V8St8uYjlFB78l+7MAe5agCy99eS0MWEoSXjbNjlW3sjMjy
pOVJAB4cZlurLVr3ojCz0GLQd7gU/FKHJ2ZUce8km+GavuSukWIoJZScQg4pkn8I
hTiqyxP9Ip70VGhBXIL31xjTIlziYyqyWTSx2DudP/wnxbOsRF79PfKI9Cd3Nv0B
UKVXqERyL5nbo4KDhlOG9QP2wSy05jR+aORUJFVejeAFFiczF9X/H/FUk+MzjYGO
eM0KZRV8/PtInNB8MetL6yDaek0s7e+sY7AC4XGWx0YmRMrYX1Stk2sJpq+YGlX6
8mTDHoi4p+QtHeYJRWPMub1ZAzaVe+bFQlt8Y+dXvFbumTqwt9mMtD+o1CFENlPy
wXEumLT5FdilDhSgzV1nkVkTPNYG2CvNwyOC0e4Aa8I+cnKh0s3TcfU3YGpaFhUm
b+YtcfmMvxZbKiRr1pK5Kr/TeCrkt5I/6RBZtlbADKD1EkNO9v3rdtrAoPhSqxdx
9TxI2AlnPRW3f2ltcPbwE0opWZ3LtKPVy0JjO7KwHieRMJdKpy+IJY6d5R6J4vaT
AMgsvKTtp8mkF6BNr/jwx0UjoXyz/ke1BpI+DUaehR7x4SdpayZZ5KG0oxbdDD8+
M0GNdH3LxDqSrDBxUbQPnI0CeNxh2uyAqn/FK7OLJ2BuW93ssUHjjCOTL74dfpNl
I0DXDMsllcv8Ei8ukoTCdabyowklIL+5hsB+8poVCdayIKMwukmFwWbof3QFfsUu
yd7XgrWnM9dASnVPTUMPBvLNgCMKwnzjM+aIf0Fh1yo3yPW8gaPCmerTRo4yF4iH
5mhl/LdLgE1kX4wNVgY9R5TL4+Y/kh71FrSoM6a5sNyPgsI1igalUkVsniz4U2Uj
MHS2PRyLZ+lS0rKypptl64bER27q+5PLHMBsHefr2NmAyBRUDv6ZZ8KU682l4QWv
s6KdpufluhvVxIYplGYi9lBTq2K93NbrMscrAZBYBPqsRmLh0lPlxI2T2QYcJCWd
266TSK309cmjJbbsSb9wwcZ45qh+JsHHfHPPAvi22OIx66vhyKW/pDnd36tiL5PQ
d1wVK6K5/VrWwCM5Rw+FWbNQayi/6XB1xeajtMKfdjReG8MF5z1+NzxrTcrZHXfC
LAOtKgzXJoDF9b5V3hx+jiHLIow9Sap0lY1eT4j33U32YVcGMLmhtSCMFeIIwLti
6q7dwUGYuRNCCFLKcsbDdR+Pw5ckS3M5QmlNS/Y4bYG6BnmsSlBPAuL0kW2Q/zp7
rHwG8zPUTUypn3+7Q3mum8MOSxYs0y/gVvnaIvJ2vo/Xtddxv9zBzPhfYCPxKTXP
6I43O5FsvbXh5GZ1vnd1eaZkzfyzdacZIBk8teluVgKTbxxRrFrDq5YahX9SZ7Gf
ctt9ebrdF1S4xxuyYgQYkew7UpPIGCr3oA1q2trQwZ46iQBEItKZPGIhveYgy+22
53NBewdU+Gw0UxMZ/deYN5k+dg4rH2/eYQO6daLcuk7q1lH1nDCgKxIlu1pxh16H
H7OXmJ2VnPx8VcJyJsaCZbAAyYsd95S4TAR0o5X1V8sgfxg26zZzCEZVs0RfAgX0
JlX0EfK3HnG/jCatp4BOF+d0LCheaniDsyG+KEajvagW8SQLI1BFv/72iTkJddBc
QXTC7FstLG1Dj9xRi6IA3Y5SowKiQ6Wj9IiX20QpxwKV2nnHsJ790VenSjRZAKgz
OkMbjwnagP7XBcC5zHKSsXyOeEgzRtFXb8gzMTdDlsukIrNBNIAJbYB+NXvjE7iL
TU5CxQBwogQCppCOBG2y8ryh5BaS3E7vmCjavytIN3HmCrYSZYfXcYJ6vNqnD/Be
zvo6C3DkjhM4XFPxMbe5H4nRTOg0S1DOf49x/HOEwzhjCj1GJ2vkpjoMMxgexKSn
lVAsntgm3hyVDLTwC65GpOp2WeF63e15stitUa7W51wrlwLkHisULQ02X6l8B6GQ
614rxCLrjx/x857HJOhKzE8I4W3UHDqm9+TGqnk3QGZ/pgA52WB/gJXtXiPDv2Wa
Cf+1cD5t84Did8jB++XYenPGsY0pXxwb1oHgXv3YSzrASqMwyzEfy/rrMikuYJ9g
OWsx70xFn14CvdIQroaIrOYOXTH4NZG0k9tVR0uW1rpX4PkzV2uznUQSgppkBW4k
JJ5VNvkRwcKIntjteSZQJZu6Ev8IzBqm6cmnnwQF92IkAskA2vYZar7Un90NYtwg
ybhPcuBAJjYdRrXP4xlJKW8zsZlCHyFzlG3TDTUYjKeke0c4CPFBVashaZfzHKgS
uJCLmrlgzyLURge16y0vVZ2CCXV9dVaVLC9XnUZUv4EzUkpJg7jPqC2l5PDjJenq
rq86hWRYlulUAD/OEFQsTqHgdLQ5hchzfLw/QxD3A0/zwRA3n1l9zmsF6q27b71L
P1Szl9WftQSeHdprlFFGMV/Y+4Rgub0c5p+3MnXUh184uOhmbaTQ746dZLdqxyJq
1ptMp85+1r3WghT2J/xfp+C0KZUxAe8quWTtUUpfbSnJfxpuQmZ7xW5a6cp1sfaZ
2Lhon1aaTVXqmTGEiZQmqvhCWYqT1jR97tQrPB8p9TNDLwfDHuLzBF0XHrWM0oit
WjBXUjy99sj6NFlhAcOG+i6ZJ5VqFb5K69ska30Mgy4T/qfw10hIu3LmA5mgKGKf
aVp5/sjZyQrHZ08RoHLaxPyuPdzDWAA590oQOKa+1wFgDyZR2kKqsRuL/YvRp+uF
oK1zSaJuxXWL+8BF8SLNeRZRLrSW4iPcgzFDUVkeNlJKm1cCrL0fm3UqRctEShY8
8ChILvaFPozTr8L8SApT/PTe1tG2NiDrlLP+eqLseK3vbIoE4sqdlWLUr72lmvxQ
i1Y+FNJ3uMqeVfkW5ThRR6bNhBhAJ+RABrScG+K6d/9sIgsXNDgQ7Q942H0BYPNb
EnWHDNuzhGXDQxJTTOWRkmqtf/8slrWgFCBuwqBWNLIOx+/j+nsjrhaXLC8CxJh2
P5IQhUwPkhg3gWSxKZiQQDkzS8O2zEH5/nve9wTEAe5sj79RlqV8JvFfGpx3rcMh
wAyrUtepGDnJ5tWydvpn1+hO6t/ap39W8Suznt3nNefVsc+ETkqA4v9iaHCBNwtL
Obea1E3yPreTprMJQ83+Tgs+f8plllFO6yYUa3oGXa3XJ/hPDTaWk0ZMe7wmerkE
M/BcOyCY1MpoLZFSRNgeG/Q+3Euz/Hrrp2YooEV8oG1wvmv5AF27RjWM2QK6COPa
4LsFSxhLoeULIGAxqS2fgw/vrpsZ4s+apf/KJpgYsUz1DHBirA11qIwAdmEV+7sX
+Th8opVmHXZv5ecE6pWiZ0SFD6bkGSHHAaJOVcXPVcptsYLUijG4uogqO2dARfK6
YP4OQhdU2hwuE82atQ9mGrIg9D2O2wrTsyObpzb6PVUyiEDwtbZFALD8465MWIYg
5fxfoDWOazuhGW2C3B9/xMbH9VwjOe+0cjtbgHPASSp4uW+8wf++SpEoCAu3Dd15
fdbij/wkmg4LBP5H99H83IiXUGuYx8GNJi52giiIuaFthACsKKDNFTFq2on9tYrC
TCP1FvEKsnUHLpESIillyHTRYl24hNk8Vb31L4YIWhGNtQ07YiQUf/HAYYK43toQ
egxyUJNNZMQ5hfubEdL4XjO2dCLTrvGLqVaJ+pO58yrpyTjg8pR1k6OSMv1rRNQb
cvwMdRWLwZ0pg3978JoyVYSWfWytECkJpf7RzIK9EgH8dZ2KSvw3UrCn7v1I/aaO
LFKHBazDWTJIurB8Zb1o7fHUMxHPiVw2uuEhzYfAnCr1QRPr2drjdnU438uWHQzk
wrKOHUFbSqChr32RAtWn9omzOa8rMNPEp2brD/OXSWilmXnHD+h+yBpWzCKkxWjl
Hf2kXGYaSWbqV8osH8HabFpdF4k5e43Kcwyykaj2SKlUPFlLraLjo9FxSdS3S324
MlV2pvHxCyHi/kDqPF6Yc0j4Q3EsqaOnmh4bmYuQFDhLr+W5g6nSPHmLN+mKByXc
b7WZVphOHbhtu8z8xykpWsUGhocRM8O5pZNJhLJg49LaHdM2mEMtosfWlqiWdY+D
bl1+AbluqhNAsRww9t2UgCtwXvM6Q7ka8VornfWviTUFOq9HQ2JciPPRWrANtpn4
eSgdZJeC3eSCapiCQXVg/c3BFPS/sO59BoMX+7Ap6WRxKePri7OKWhdX9n6VZJTe
KDYaQKz15D9R0YhTxIBmu+GsebaLQQ9akYa+T7+7VeUFFzZNTOX1cYswMCAm6sbO
Fgbus7Cad0EInjjEzySybWa6uyGzqz4iBzpchFaarNar0no72pbQSIhM/dlLSyB1
neta6RSXmNEJca7oDEF153/b1eEpiwFj2abvd3gBzCG8SCIPeT78sQgIqPKHIMke
0KXeivrNxAVyc28cARYq5Sm/iSRs6Qa1BvSkjIrk1Y9pzt9WZF25SMdID/E+rT5j
gc3D9zcOxFjlhrtbr0FKqCMXmWwzaY0RQ1xihOLzc68Iwg/Dd0S+C2iGoz8IZZPL
Lsusd8JmS6cXF4D55d7z5FvT/v8pWU53JHAvoKSy2BnEp2BYB8fjuNPmaDjk7Pf7
BeE8czUmWRR7x6Sc8xy9ReHgNj1lvAek6qNwxqUZxWnyUw0o22g9krWUpmIV+kPM
h/fdFDFuuMUe+kw9Q5Rv5z029CcGvmK9zl+NB4U5LhvR5L+PdUFBALnDl8mEenka
g33Pn+cH7V8uxQ9n1zkuGlxIaJ64LUM0tqF1oqd8n941QLmuQ6rMB/XMJ9txapdj
/7MGqDKJ3USpF9W2/bwQh4gO3mMSj6c8orz9OHfwTYzaNoNrWdo1Algkf6uxYUjA
UDZ4zOPcjaxSw+jVAfmzMOXBiw9H4TjolKDekrrFQwkuBd9QiG6Hx/V7VvDsWWNn
x1POzVzy2TnjK+UJw9Xfgn5yjayGhmWSy+61kp0DK+EoiBcnO4Js+BEZJB4gQkbh
kKxLeci2aF8uwkA2N6YYjFF7qEQbWs9nKPwrJ58ay4rg1j/3ZpIoxPyEO4GhznTw
ZYfNQffwY49hyWEIlLXjbxLXh8teXmlVjQp/bZuHnJ8DdkHcqvy+W9iZEknOEfNT
6genC0lNw0tdboeWaGLpnTpVsEwoL6few075sjaFXNeVrDI96ToteNjwKXwLZN/4
wFR1kU1CePpayIj0Q+HC8OnlYlGnvrWJl0qhDPbI3YP0XsaVfX+ndN8/NgX7w9wm
5x6Fs++3GsBxulh0DrqM8XXfK2L2+7AQDA4VAhXkD5Yfo366RmNzNnfkAGk5oT44
U818ie4WdFWVhhHntL6LgY2gyEkD5hDt2zrdsEkPE4R60fnYrj3HtnQTO24NdETC
dlIAmLGSu5OIqI62TJMK3okiHrsdbD+S5wggno1f5htGZ/fiSJTbFEOZFJJHCR7u
AdSnloYDNHK8oCPJS5l7bg0IRFIng6j8LlG3WkU8UWueKbKrljVXGFk2RJdg3bRI
Mto0LQF4+l803u/ADvPrYETYciPmAkPE4ujtHJ3Mx1CSC5QjJJDf5tWTprJnlaW8
nljEPbfHmwi26e15zsAB7rsunRD0aVprCtnn1LsRplttod9f49Ef9UFTYlVoUCqn
YlcHI8YjnDZu+SdYOV68brg1529aSWAz/Oejxo3lIXzs9yw8xbqbL1CAsKiAgt9f
r3gjhjE2hhDBJC2U+mTGeLwJ93slhW4OLmp4haa+Q7pV0F+aH07FEk98B8iZV9fH
ksI/DE2SIdYYRTo/Bv+0OMuwWw5TBoFTKXYEy22Gd6ZE/K6vq8N1n7ul/TJDb5hv
WDSlnczenPicL7RsrBacFAxCyfeyPMtuZ9epM4hrDM4co6OUF+mXXw3SxQZRqnrY
u/AR1z2MFr2Jkp/qKAAKbDrpqYycmv0Zl2ZNfikttF5lEwvvVWlogSuRzQ5W9s+e
458l5e9diMPvmX42+3Wv2CTcDgwgiImTN0ODzanZ0rW9ZESquRP+RYCTeo+tc1aC
SMlnG/47ukDmIFAyH20UgnBBQeiH2O+TsxOrLIe/P0JuJjUdbSGkkQmXbMzeA3cQ
Sv9btSVzSpLDRhIm5EKeBky5Vk0OgAfbPzub3DvaxytiA2T//NTRIadoBIqvq66F
Mg+KZQyQ1XUJvy33P5YZrYTcqbZnAs7OjAmABpJyg4WAIBbhy6XrPQbrOw2259WD
h8s2dA7SMsVa0ORY4MRWvkDVSFJIkprNAglgVYVQa3SDV5ZMGxrdGjlss8uQwQkd
nXDWjXe65N9j/6G3dGt+v37K/oRRjx7nyHRxJ0GbwCzpST/NfyqR/9mpueXwRV/R
DsoCNJy+fWOrPi4IjpikKuWRAONyEVuETrIyIHl+76MmVrZnCp3CaTo9o2nfetMP
Cc7uqO0c1gyFjMgdJUHP8tCCJIti3laLUhxO3sYxl8t55p9grKwQFw6CCVL41Uo3
/OB9KpYdJ+jO7tKPYGHQPr2yFXKCBfQW/xGTFhreLAS+Be3vfDbpgnBNmQjlxGDW
4OazqNl7A+9MOqpF3PuVceYabjpDvOlJpm1YqeVF8vVcnBFebaxHWFM6xDRWCFCm
bEi1QW/on7a2FtgC3Oi8q70A+u9dEYUeuhcz/rh0ZDzLZ7f5ouvhi36jTD9xDrFT
0rOIhaVJS+s/gfk8k53axf3m9sXwHW2VnbxGjh7A/cIUE/KQk+tQQa7w7qrCRnD0
fXxOFY+yaXvHmWz2TTnQEBulOBlHmiB0xnEhzF69KkNCNr69FiCj7MZC+7Ce3CaI
ueNiTWyHUPHGP9GWGz97qCend9TNAb4PtqsJPDD+EQ1lSY5cUAxU1KAfLxjvf2cQ
pKldTnDRPuStwUCZU7MfXv3oTRriWQP/t0aDd/rWO1r7G+vHJ+N28O7I3LJgpjDx
8j/4kS3otNzU6J7ME80GsEmfqtCiYTxFl4lUvx/jHkYkMz9bUpdoO7LUrit1YYMO
TzbSymTD4aeYhgCQte1BRv8inHozQ7kcWhkWKCbI9Gp4Zl46G9pKX5AgEmiW6MHz
srBOmjeKaeUqxStsbuOHpgPRu8M+OWfTftpr1wY42At6Ltlc2O0hkFD5iFaNUD6t
MgLw31XsxPw2GrbLlyrrinBidcRkCG8OouT7lU5w5NeYTQPk7vBbPbnIjQRMPO0f
UWb5yRMX9mQSvqNcwhka7CmPqJbgRaQgT8WlKb0ccQKn9NOPkjBn8bZhJyzwthOV
SyXR+fgDazkaClYy0Bkt+xr2LmzuZWlEdK7zWTmspwf3OGc2ZxGqNPMqgT8E8jbd
tGexQkgTWqYPeGvrQayX7AQDeXtq/88F963mfNPu7/hAPkuIGX/5OitWD+NNAp3/
urHCpoeA3QalXjEKM9kL1bRzQO9oDhRnjSKT4vZ4UiK9BRWfoQmnlDR859gAdAKF
0XUhnM9CjLrXaGHh+IbzBBNetRCN2L+cxC8zJu55V1b24xliEjLfqRiDiIzsOawp
ihR8AcpepP0OPLKKEoYgm2yuVfuuK5DTHIpznSbfmSu6wcMhs310kzeaANyuqo7T
KCNkE9Zlsc8jwIYi4oftVKqc0h3FZlXxf3iEW4C8M547l6YE6z2JmMfgSMtpinLL
adiR9UXvTYaobGweAlfO6gz32eaUvdEN9B9AXxwfbCv1kSZM8xy5zQ7m3MpGlc6D
8i2hXUmtZ2MM4F9FuNJo7N2kOgp2yRHcRc+ktrRntZwgmMDf3i0umWZChEc43T6J
BfL0sYgLHWF2Jed5AUNix5bjk5q1x+1pXb1tQmQ5UrxFbrpBJxMnc9Sk6r5grBG/
kz4m4xJBdWU09LfkB1C5ujKFdloe7n8RL/LKXNYfBlhYTiTFDCWEPUEK5np3p0ri
tl8CgvKyxRec6N//HG7Rq2Xe+IMg/7AIieJuPlQR1AXpmflcmK23LzJbIFiSQpSo
c7wRXZ5UfS0j7/eMTvcOU4qIjGNmkp/7wWtv6zUbuhewNGUJFMo51XOZQn6m8fDt
6Do9Yh0UhLNbXV+orqMqAmoS0cXzdDrmUU1jl/WOgwp2ljQVNoQw2mKZDVjO6ijL
CgVo5/zUCT82mlI+Qr1qfg7Yqhrf5sTxzLUTXL98/hPsbGyU8zWQyfNuAcCdgv8e
c9x6lYlS5jUcu43GU4Y81qrr3eT+5fiIlgJlqSqt8xUS4JAI3BkCmDqOqgWLY4B4
P95vI0ZVkdah7McJmuiUW/H6d3ki5LSk4IWRjFxC05AH8WM0GFg5o9vDTU8NmCLu
m1t9HmJprQ01J3HiD/8PPUrA5f62ZuloZOFdmNVR/LjLEoa07hpYwYIiZ4d1wtmC
p1OZ9BVofzwUEi2eRlx5Rw5oO806xWiTN6jsFKcyQr8Fz36zU3H6XIMX2dtdSObX
bEyT1170dPppTlr9j5zTDHkU6zhrbvvoBDrFtGi/isazeK0JH2Wyq7ovYg79UaIf
UoGU5an4BFdqFTWQc+/+jVrlrVnuQ1r634fvhW91jedaktRjBrbFwcq37uc+AIiL
zyCbJqmhQq1NG0wSksleQUp+WqPNIOZLO0iJZLWPifr8JBiHw9reffwbIK1Gvh0m
8Z3tb44l1cv8CbP32GcRbpiqwFybwSvL+dc7K2yzqxRylUw6KalWA+ipuU1iB2UP
6Lf4RrFqTeITTOEmscHhYgElInCytVmngqsLXBL3OPoT+Zf1MvrjkA6CQnt/UUlP
3a3JKVmaXo1OXeSx/8h3M+gOonwAwXHZEE3mht6QviOwgyuuchzqKszt+4Xp40k4
UKlwrxYqIcm3tVqi5LKG1SODHQd3wGPTNziMgGeo8ShCGFxcMyBUiTkKyciz6Dzv
zpXqxQMpfZWPpVmmG4F2KTAyZjuDyK0Q616DaKuzhl08FFnOzIhJH8jZyQs2UsG9
jEycaVnCuWEhUb+rykZ7UMGctpGMq2Jixq9x3yoQvc2zoZCm8uJUTf7cOn3d8caJ
JjHCxR2uOuIOPcqtfxJSH05mbv0iDcGYRrcpOlPq443g+MO0VLQGMjQE/2Zg7Pst
4MqmYhzz4zFCGqUZRYpcxgp4n9YJWZBd8KKjTid0FrOcWkuzqZqTtA2mP2/EZkmX
lvNppAr5ZVIK/Nc19qQAFmn96Im+4uz3Xpt5Q3rnySqSCe7750qh+vOb9xDkoxuM
TtEf0C2lDlJwYPY727+hcr3J1stkEnPHu84kMEUj4THDuZqKosfz5uAj479gV20S
DmTeIEBfDdpqkE4mZ3CSw4p/04PuNkXbnTLgJzD1JmB44jqmggK7vPzObiU3y9pf
21iFU5aEDxBM3/MwpiVQqGq6MaHBRywiAUq5kq/jVkGVZyrJZMdAC6JK6T/QGe5V
5msKWxZsUbFeDYMLQxMbXgwfvzfa55MLUsYPhX09vIXIdc25LF7OyGvN/ExY1jyk
Im63M1UXG488rwmXWSutU7CDkmqmJ+LutiIdoAJB0ITMhIPUMasVLe7IZASmXBsb
/XX9IyP8IuEd8VLKeTlUTiIKHd7MnCoWYICUBFWD47PmD6Atos3/bCWBuZcKJPsG
K9SBAt/edATglCBSWnsROSakFUajFlq0E8lXBNH524MvM58nj2g6vAtq6Z/nQ26R
eZG51q3HhZpdV5T6SQHUAvKoZQF8hWRD1S+/tgDM4BUiTXKS4caPtaSRs5Hn6aOC
SWxDyKMBYlrxLa0Hb24A6OP3MhYCLtrOSyKfwJIKqK+gWcKuMiTRbWpjqIpMwPiK
mZ40NCeaqKdPkTIwIXSwyh6syltF0RqoJBIheErKxxVYYRV6pcYJNcM9tlZoeqtI
gyTBOrgrlZZZGGw7jBkveOGidpY/VSO88QONX9Gz0OCbEEmRMkHPxh0UP7NBCRLu
XMYVSmOEVyxGvZyyQs/9yGEVnT6G7Q9Nf77J5xED92ZOls/kwAPlcuuDoA6QaAim
hrLEnkhzsKdNShuNnf+ORqjOLBaxJp00GjZZ81ObSejR7Mr/joO52eFGdYZkfzdg
sehRxWl0XWe22UOmF6Df+0DDWmGyBywQ+LrkJN/kr4OamwBHSCgWhEdDLQ92ODEU
R0+OhV5ZlQlJjCxw9uytOHf8qQFIKgFaeawHr00ZiVr5xPJbqcpEAVMbPNMNkMHz
Vy1fgOZvSRpWf5r/fsLLjkMRGgNWfcAlEeC/Om3P8jsc1krozzEiFkRwmGk3QEmJ
c+t7lkmNf6O1yM5n4ndqIbOeV0KWVsXdUzS/jrRbOmS0Q5bD4NfoOFJbYqX9rpRA
BXZFOVjanopHXWfROMiHF2xt+pF819LIBvb7DlJjqVhziUZL+k6oVKiOS58oxmJx
TtFXd8qKauB2Fy/oQaGf1BRlHSsPWk6q+2U6Qf5eEmIjI6xz3t+PTN525+zq2/ZA
xExDKhV0HmqXOfm/IFJerUmK8aUKHg7jM9shXCfiI7vDyISwKVSGyi8V3dxImCfu
f2fSusL5DxBTALEeArXH2XLXnjLNI5i49Uq+NVGJmRj2poD1UePfKvYtkM6Jm4T/
0uWydBMKwnhzpsoKX1Ioyp8dDhk+Et1fuPvLnKzTk9gvqpQKfeHyjAvOFrVrHcCk
3MyO2DU0I1AopSTNNJDmqiLegY/mNhMffa6FVqGM94FVOrV57N3XXphKZB4CtGW7
43awRFqvpV9lNS3A75kKoVP+rjmCqRAEt5yuCVI/trAWfvW0H+BuqIJvSUFoMcn+
2F+1oLLIzm3sCGDSKImRnrnf9Xx1OayugKCkhCKvK4No91zk0JazVZkNdN4Q+9NM
7lYI9DsXdBD4NlYSOyefE8JaFzXWhAf5HMKT8QdcziEdDK+K51McxYf9GPNnVk/K
nvNFaLLbXHZepag/CJFVBlJAfRMGVPxhZhD0bovjQi6B6W0kUbU9ibJNaznT4tvK
pG+IJ3MgQnmd5rcqs0F3xlHk4G5G0CiEXvDqN9w+grZv8kJCVQ2yHgILaAuxoHuZ
bRjFnJ+x7iGe629seyeg6iOrOlQWeZeoyHrBA2T9OR/zETu3aGg5CqKC/G7ReOJQ
qFq8kHb3YsyPfBZtdBadUlu0RQfjwuBkqifm5j2gARNjRfvZWdP+vrvwoxX7kIvz
ECQtD0RFrSabug4K6U1TO9zs/FWH8U7d20xo7EY+oUiOQcQoJPGXpBCnSF3BfHgH
vqY7tnQdfpfkkOSl+KRLHDTEiQtbFoaqn5WMUjFsFjP2iJWas9O8QTNGqh+K7oVx
VZdEZB5Ymu0ATduWPZFFvMm6FA/jtNv998842sacMZFK3VD510oinVFdG4iA2uSc
OxrPJ1fGEBstLC/ZiPvVTzcC2O+uHbDArQk6LPlofFPniw4c54QgbOQmTeQEZP+m
xUDFrM1zUrzKswbjBF1xRDL/LgP/HCAY/GCn4HlmtUXgYr9K4kxqF+IQSGZ9RUY0
C7+aoiYyZ5nl+fweysO/+wupRIjOaXexpN0gWvkDcQYypPKEC4hG0bvdu2HLkNhp
k5O/eSvkVz32cYl6nGZlEwN0SY7q6a5Rv39rJhMKvUYu9EBJx0f35k2OOnatqheq
0ogAMIWzBPq8xl9moARWrseHrxLiAMaq9KqJbPDF/rs68OmS6Dl+2b/NjT7TKMxV
6mHSBd4zUwAuyM9ZYu93esLUk0T96bymtCIu5HxmKWWU7zBL0OGJlZ+n26b+a8sk
fOy/GTuvwD4Ew11ixk7q+XE06gx//c7b4FAI19uFyRYL0YQBv8wnRJluq3oSarHK
ykrDYt23VKDD+bPgD2j/GfNGoDbMlFqTGTRB+ifowtAOffjZ//sf3QONyMJswBD4
YuLhpPZkpZObnUS/1B6DaxgbfHAY4War87MFEMvfiO10ZgZFFep08c3lY3rFS4v9
W6woR0Uf/FPeYPga7gc06J6bs8Lyt6xUZ5AsCSP581Gu/7cFcpWibMMUZf4RSg9v
6L7CBP/xCIFQ9eT1IPQ2WaO0J91h0Z0GZz5Sizqx7BVEN8/FMvQtSKcfozFdBjS+
xdR0o22cqrThUxsPIpQzlm2bt0B/E+NiOG+KpGweXTRTDqiBjOE7+9WLNt1B1HhT
Gv+MbBEEngYBF3lUDmhqTMRUMtfFsSsFFtod9W/giiIGngrdmJrbjxUytZJuZeX6
qxSXweCz/xcvnAb98ZNj/0btHrSY1UqdbEbAPETnJOEIIgG8G/PMLTD2sZ1z8hST
1+pytMkm+VO1IJxTKwn2yo/3DTbk64WF7FNh6zrVNJaL4OXwi3NdcmfyJlJGNYx6
rmu03P/4M8XyJ1lXI70QKynyKfZGKZtibaRbbgrHb3gsSXpm78OCp0vWQlg+FmfL
1bULzjqhPJXwHXcIW2FzZuqcnVNQegcqMXr5po5eP8/5NUmyQ2DuY5gNIFMBScXD
OPcTNLm4tuJKNcFM2Q3MzGvuq8iUJeb8TTawMBdhBKt6afwlwa2onsvyGWMV9MAq
hqLnhQIUyw2n29FrgrKWKUo5kg8QLESt5UVj5R82Pc0CU4z36qvgmOv7sLYe5epj
Olj7KcRT9ijS4CUa3uhjIPgHUHlaavnlULPwQ0XjOANr8s/DJmh4JZn1DPg2FXCd
H4ax3k55LgzY4czwuApK3awgsMe8DlXTV7kBaZWXipqkSIXMKsGpfOHtIsm9usB4
VR9CcgV2PcwYD5Lc0IdWJUIR2MdjgW5omvM7r9IOHa1XNOtw+xsBrzAkwdaUx89+
1aEG7mXRv8E1IduDL+Mxol9qvXQ0/BgIAGi46TtjtxVYYfMXBMwkH2mX3Y6pHTE3
/M+wQL8/6RfuFrYCZIgSJeeGHfMxWO5ro+A42+3c+YnRCE8XEOp7KQ6kPYSBXN+n
D9oq3TeikyTQ3WBrjucFNLCh+kfUi5rz2vDBrB+SQI2OsE656s9lfhITAdzqrL+M
A0Lrps41QzFV6aztgj1FWr4GwWIxxm+y1qxc0EORsVOuh0FnUmutkbgnRpKhq6o5
N8yjiHI87oqJ+Al9q8XHcGGebak4F2TxbYB5kX5JzPTE7v/m7oy/Rd4XpD92Cxrn
nbYtzMIjMJ76VBSRktWNXy/a9W4iPqM+xOc9TLh7E1MrEy1aQgbYExrCn2ect96r
R1u3fMGk7h+tXNd9KSenNCmnx1n5Fdjp4UOkX/evZDcGAOjT6vlecMhkWAMUXPhl
3VL8BMzdciqDTXUSqfAGb6L68uef0hvICNSSyxXcokm9/D6llDdwWhVbM6AH1ZMO
QVUSz/GrgqNdtvzvcFxEKmlx1KiiVm5ENYEvk3SeKtJh1UlUaMuuenC2LPyUOPDW
k7uXhqj2z1iC559qxtt7FdVkYso8FYnFGjAzNEW+FL/HzUGWpolxV7K7lrInLKC8
MYMPHDC7El4NE8GT2AfOr112heiFq4Z6q8Vl2vx27sfcWlR+lGk2NJMEnsZDv31M
Lfpy0VLatPW/0dRANwB5ePbuApBk9LA8wTX1MT35Dhz+hLCizCWZVt71rbkenytB
u7JThI+jDGVWJK9zTCcph49Q1FREBK60RSxViSuRrVUiAESucVLDLYGaVycxSNQF
3nMGaVcVWZGqjfBX1ctXxp4RAnp1J/pAGEHpet8/rdSy/nhOVL1UaOinPW5T8y//
IBlyxNG21Ndae5hQAsXK2EFNfAF46sMj0Hk0696wvuPHJ6h9zxHY3qietzxag4pJ
n26zZ7WzoarUt8M9wUyFuS/Z5pFnAUbTeXxtz0SdvuWjGIFH8B5ji3VnTmidsl7j
B41wdIy1+n5O9V9RAVCIRv/86XvyQrMO0wlXVfebJmjgIaZt4uN9bEH6/2hfnTrE
KMrlBir3D1Mb1EDMchkOdxEf43E+izL43Jl7RL/A1r0gGE3+bPJerksCTbnf+hvI
qoyWXKspKEtjkpZd9wygZ6SWh1CXMz9rbDoLkTlxgY2uD8yaWZZlukO9qBlvNT3y
1voooIWGFWpLXBEe4Nxq4P9h0vwV9YDiUf6tAg4vGSzl6nOgNlsbFMMsOkUH2O/W
1G/4n/j9IZg4X+8CmbZN0agoxs6RJv1HGG0LNGLAKQ9Np2y97/KUF5CaI5lCa+YK
5DXpGCQwp2bOQn3ytaxVKoEQbSl5p6aeerMlHP/8ZCD7ULbL1KF6HaZiy1KBW4Qr
oKTuUZlWzptjn89LGXzFYyftzC6Qa5lzRMu/K+ZT9IWgxyAIAK7k8/HEzCR6Ct4U
6n7W6JRSf95roX393vbUnC3JGiGE+0SOC0cIFndDlTL4f+gFq4Y+EsJ+CQkeiyhB
r1IgsDM02Mdvo549yVzyqf7f5FJ/GrW1fjx4FEVKC0PVJia/2GspwGd0RJln5ur1
04mT2Z9dlkTiJn0iuk3RKHEQw70ryYNBellTE++9IPQUEbw29LXUi1FQuMdOOaLP
M5hZY/UzIvN5NnRoeiZTlluCI6hfatrwT4Yk7XU/kQTnF6etnOzwQbPAmnkTtV7w
kK7gSL+Nk2/CJ9cpIuV6vqojR8Vn2BDsHZLD9w6s+5BhMK7r60ckurjBy+2Ioeel
FjOs/yX+d3+rCNojv1feZ6Nz3gtrF2y2GyZzzhsGXEgBwwA6C9VlqHbKv3p9gBjg
jjPVHD44aayYVE+8lvOJzP82RUkdr2Pwx7mV5SRoc3NTcSTP81KFDq/zCW+d+nfO
V3MnkOMCgtoUxXHNbxoN6xat8droZnjFyzSiG4at1ydg/TPkenydZWrdI3dml3Wz
yWtnPDtX5GwG/B4Yxt0uwmWGiR7p4S8bboRlCmyEAywSmCBeImTGmSqh5Dr+5nzq
4sAHEg1JCOjiUZgjKZoBlHH4OMklmMPdoUkzW7Fqw52jT6zLO6LbGIkp9Wu0cPEY
pOjftpOC+BaWxFkovJHsxwhzKhw9jmi8s8Duve4O5VE0mlMilk68IJ6JF8QLK9Ha
ZtVRYA36OJJXzfeXl90NcWK2pwtRI/N8YsFwxtToGRp2uxd+CrPihAOBPgLXGsqD
yhTgRlqkuHqVQOZxS68LfxcmXESTxtCh76inZX3Xgk8+Ptbkz1HHHNYvXoVV11St
LLFCt0JB+EzB8Rzqcq5knvMr9iEHzETKK+YAKiDJlxq58edIiEYa6/dpnqd6uq+0
CdFVlYwXIasJ2dH3X3hHAL9fn1tRslRaZ9AR/YPa2+/oqcZ3fLjL5yukRxN9P0fb
SWVo3OL5wP99BQvjTmz0eGU1xQru24N8mf1hHSVh/eEvkA1SSjqMrurp9YLY8dgU
mHE7EmIWQcVLlVtWsBprxFHg0diLD8iPDyYXlUUXjlIEPPzRKAV/1WVpQYU860e7
XrZ/Cfa8ltgsYsM7cJe4HmydOLIxuJTS9DtLByP21KKdVrT3iX01Z5eQ+WNsMAQr
Te7zyB5xD3pP3TWXaHHBg8MKu3WDKg3I4gIdA8/EULOIzQvanHvlsdVWo09+1p2q
OUszge/EKQ5F96toXj7WNQUZzQGHQolS2XSBXWip6HvQlzobNudtmI/x19jYwzub
fqGCmH08VnnzWjQA2YJEubTYjFevKqqk57BRPRFIuUJBWnOdmM7XY2CPZtbNAuGf
rB1HWbF6T45dhCVh7WxxKMBigH/Q+lJjYQKNHzdoRfdEvjoTlxj9hUAIr/eV6fg6
eY93ed3rvqvygSTb9WM9peK8Qt3idY7Dbbrj5hvVdOpbkv1zJlFtTDC3yF5BrESR
3l1rcIW9K537mhaSCTwO+aCqFN23aL45Emunk4n1mdb1LbI9mit67BhLOcHhEU9L
BAIgbWdHrBj5ESuxt1gm9M28Swvjmp1dy928mcCzdvku3kaxI6vLGE26SZUQXVns
GflqGj5CLks67KYtzi8hG1UNcfvBtAbj2OZADVnBXt9j6tZglp3SXMq4B5Cyd0w+
z8znN8uBVhAxYsCYRdLz0fpOxPXrAdYv2QDsFTMEn5qhqLM9A0t+OXzMccsqyEac
Qk+jj3bhd9CAsDuM0Xqv71gylOe+jHRJkwO82oLor+dHTdzEsXoMFJ4X7KAhosZ9
YjT9wEslL0HBD5YCsyrdT2pSYDBRxn00ykpZYAkCo5tK+YaL6+Hyyb0XrcDbtA/3
TWuUV2QrNmvqPjVEznWX0OboK0NE85M0M2hDJucx1BM0ehZ1k9kT8EVqmxSQQIuh
mBkbY0fvaet8swLP3X1ZgxU1R9QIuB4rXLtvIyqHeolOWrCYoZAs+z3yqzOfdEfj
CxwGWN5e5YpX8KyhldxvqSpWtwx5xSoToa1Cyw6ddAA1aUL2ZgTUJ1WS7VgYAtrO
qAiE2aoxlAl1IoNeUNxXxGO1wxtVzfXcViR/7rhGT5vTjg0gzqcDN8Htt+MCv56G
DGUQgAcPETRUiCXDw0KrdcCuJTFkdYZe/1Zm86IETFuobMbMK4Gxm3ZJvLDVd+xh
da0KJVnq/+ovhz9FG5Zf90d5b2+zIPVzbUkMmkmO0aOpK8MnvmUlN6tKh9lnq71s
TwIH9UF+lLWbn/2uHdEyW1sYEa40DQoTP6nyZ89QO1sbt1oFdR+uLLhNx7ptdvDc
87XtofjW/zfa1ElGmsBTXOr7ZB00NOgtwziOVr0PzYrqf43Oyt5yprkCXn2z+xxP
Yfi3Cbdp8jgv0cwSvRUDx+JfzdjnitF8yiOVsct8ST95MuF7yB4UvlYfTQZWCW8j
syX+Jse5AExpUTF4y0gVC0XBMOMIoPM48KHtzDoQ0l8KoQKwPXD0TKJLStZtl+l1
+MgzVTzWRJMjMqV9i7dHLSHuxi4dqY4V/7q0TBxq/8qV09HZJsBCnf/Jvt19FRw9
R06CkGhst1eAkz4TpW5esG0Yj6rfv028nUu01+WspMfGcE5pkpCK6S4mwnnnsc30
FBpkZZsuHM6UbjWYH5RnjS4DKihCoSe6pEnY/5THUXaUI7tyZYX4hS1VBYb9C4DV
qL0C9QpsCZ2Ll4K/nxg9XnFzWdKmwtqmQvg3JbRD3R45ummX2s07B35LhaholM6A
IpQD2IMXF9x2XB5RjzLYmYaoZhixuZDUBm3xhyiRxanvdoqNPuTNCzxPqYjbJhM2
lFOshUhW8YAtjmMyeZH5i0b66li7mvEjFvsYC04CVYSnuZqiyXqV3LeVPLpJSoRr
TCfNQdS+Dk8agmNTIF8MdPQ5XfwBUhISfhiImG0gAz/CJ3KHJXDqJv4jNVcMZomh
JaKVmivbQlCBb+OoPy2Vl10qAUceAVlpfmS7i1z/fnUoZPqfMi++aAYzP6hN5l6X
R0BEnu0B8xbOChxyv5LGIkYZbW5xWD6L2X+5ywLfHF4A8XUS7c/KU5IdAs33Xqh+
Zwq8FVpehCv5+0ZLc4RdpQfrH7R8K682fE90ur+MoEbMOgE0E3mgpKKaHwPWb0z/
OI5wvz0SgBz63LQBnkPJvuAh51pwjUHdeSkpfBR2CW9S0oS1WPVuB5EsL1lIPAak
yz8RGDhjpHAPEIpQznnxX294omA5PYA4lj2w/8e7G1+yJ9k+lDdd4E/73bxtqURQ
+gA6Xp88WmxZhMPocJxjtVkFVb/yRUAQFLUeEQtizVx7RBgptCoY2uiSScFscA8P
HVfDZurT4Kunv5H9m2Gvoe3refFlPCTW+zpk7i/p3lHYsFVyacKVMfancBURQG0E
bzRgWIOzanBV4lEyYR3NHSO+jnKmksuxpzi3MBVAn/zUJq4wKUII2fR6t7wRb9G4
s2ZSSWAjQHOsP9o8nYT36DG1EpS7GmtxBXyIgJb+LGvXCpuTFZR+c+qKOmvSuonJ
FRNiySyZ6gaeuH6bFiR/emlrMasoQnm1ZEAgG4q2qr8NLXBMjvE/rCD/AQ//L8Wd
3L6EX8dx7gdwBNtkafFAyq9WywfLWa1hoCrHTh8MPvEVgUhb8pw8v+qrqRid88zt
FXdgBE4NQPDtbOuc1BbxXWD6jq9uO64Zcwu0Z8Im3voKVIt0VkgzSNar13c6u6d5
YSKoSR6VqXM0LRIGpx3KYiJp2L0JnyNbWaG55SB66Cbvn8D94V8MfbBfMaTZIZoO
t1GfKNS9SHxfnOS74luKAQmPBxOT8+qZwuv9QG3SwVj5UOyFF1PbIpoC6wJSCT9q
ZnlG2sboE7rzpnYY+pUNWhdFc+ZTb1D4vI3YGejSIwfcdERCNdJjNoFgDlHQKJ2F
Ok/3D57VzSr38dR4LP5VGmsPUqIWnsdL/y32Qz93n352VwpMzyVaGEdWvdHe5k6z
Zjq3aKcJCXaLhuktdtcsn9B3VEmN53txnTH5s5ulPTNQHM5davOA53Xgs318RRgY
gyY+2dh6Jkvru21S6N1+CJOGEsxsUWq108qpad9+BkrDmo47hBsqwdxL5AHmPE9W
0HWuWT27HP0S/n8sUKklSCgl43x2fCqEzHXg9kJL7QEO/cOfkHWo+4/uJZmI5hpc
qjGnxq0llR6O3szj+LGDxXj62hvzU8NL/qq/zfrvoMqOdh7kI1xL8JMaWJnOEkaP
DCizls4in3HqtGt40mhoK1nsHg2WQKhfg+GEHOM028ttl7pP2ZOiAsPyLcIpKW0v
FKCQBeE+fvul2SpvlQGm9qiKDrJP8E4taRjAbnXKIQ90E+au5qxl9XmjFGWjDuib
PAIdtgWW/4ZXY7hLJDi2/qk4kez9jQf3rSfpPTJvekdNXzClZOR0Y1HQxGfq/QUe
G5qygxSAjWetDMQr1+bocInNJKY5QKJTol/8cEBSt6CLVQ7ZtLsedeLB9YI5YahH
UY0PKAk8UxivXvD/7beeE3JwjKCMBEiLLh9VZEqHheGfDGrJWTA7LpSG/diNp/31
vNMjas8219wjH8NTEg8p5s5FxTeehvHdNtN96Qj4NIlcRRFYqgQLmpOBJ+ZSdgJZ
LJQ1VThEMEqNC3NUwK8u/yV7hdNEaPQr3iTL+gNNGdOINsLSltiF4+AVEgu63DXb
Olpef1XheHB0xIIfd5LeUHd08Zz3YCG33FayrV/4U3aCfqHZNHvFD4RJVg6Sz/jM
T0vTfU4kMTWWV8TG+fBH5tz/jbCDkXQh4yxQdA+0p41Tr2c11eR7uv2UsKr5arfg
RZo3gfxjZfnFPsac4mHPBqSHU642rANPo7Z29TW710bi0MLCxpEVptKCvYzueTgq
K+igLgEB9no8EqSeTucF98xxVlPXVpZ/Jqb9bvPDjryFn/sWtr4YGQfxnQwl3ErR
vDHCicTxYku20waPxjMa+ZQNTAetipZXFW5lROcoxrP6c49mDAT9Tm0gbXrz+Y6i
qYZEH+wXRH8NcqO5CAcNkMhHzJTZdU6w2gRP3cO7V7ryU63qrenHOxNzzmI99bku
/7Hlgi28V0k3pI9JajYqcPxZgwNOCB46FXY7qCXi8VbWvsg/e6lCsRew24wz5qom
RMbQF0riLJBPvS0ia9sISjlcX25C6Ow00U83oNsxkrbdsWjY4HWpFVQTig2iPUIM
de8nnpu1wLm9JLsP005+sIKlLYHxR0trPl62+bpf93HE8DoHOg6dR7Rey01ZN3tc
YGlxeAJY9xQXuBUHuOVV2toNmbbNFLUQjPn6kjFRtXlUEZVFFaYCwIK8DAMmuvY2
d1UBWoIXR1wDnp6HGiOnHe4kkNxHu0o2MjzstZGWv+NNUQD+vDMqym8Crnam65tB
1x2rwX7mR6NrZCfrvszD9J2FDKqAxaG9DefJ7oHfR3dFl0LycyOTTbk7gZH6W6FO
6b5fCopqJajQ7MyvLUHfYqWn9Azn4sV+ZmWVP6TFQrSVeRXoVbTti1yJNl3m6zPy
WpKU4MAevvr66gEE2QBCursUt1cvJX2QMHINzVUkFA1NUr5mPGnVUx2XfHghojTv
ChKrG/5plRx6647umiMgivNfLmfWUpYPtlefMbuYa6X/+AT9kvfShWigctS7fE7D
6k0ahuoQ8y8uSgH/XdNUr2IeB4DEDkz/bGAGoy2NiLlXuR7G+yAvpzeWy+tHlZCN
NVFITYd4KJmjwUfrDxTZvJP/vJpgVZBtETqaUUqiFO3bjRfk5XGldz1xUaQlOEnA
7CxHp44CmLuPuy7xZj0BqNOSBy+ByWS3M55ELwENCUS6+m34NQGpKOjGIe3YL+jD
WneujACnQjkahlKjTxq+rQhQpSZAdoeyvjmdcxhfCSFYna2D+Xrn8XzjYdGeoHCc
1hzWPti3Y6ho1jmHT62WyosNDUWHbbtWvKJjiLEsisOFJE4q76HyIWRBwbZ27VLM
kru4FIZvzUOb3b57Xi5IeaB/jUzPmnul+ti7fEAihEcUcjfSU7XoJerDuv6hBW7i
DUWwOjToDdjlqssHmP6nKWPQaGYmpHPkwNXNZo6r3vWtaQlz4uMTJ+MyTK7iHOco
Cx0Ev3Fm56nT8qNXilTy6PCcwcQqhu9vBdh84/rBCOeyqiwRvKt6Yj/Td9TcNj4b
4BG39C04KOzQkNA/1fZos20cace9dEv6wzpvo/870uCJ94QhFkDMwAjvWB+5U/F6
oQnHGmcLaltGjNZ4CY/MXvHEHnM+ynsX6xtZqHCEGEUxOioUe7nkSQqh3e+9MxAA
53oJOdijTw8ugYKXtmGAqDT+ea9NioAO4zi8oJbBhLSGfS3OcaIHciLsE2lbA1SD
2b034nUzirDkDAClaYHvBgMhzGx0iTs/6vToAzaOMlCfzAC8dqIGxlv+FYitcoTh
bPu7MJHZjp+tZL8XZQFhOffWmQXXow7bkjj5Db8atKxUpW1zZNK9a9VOGzrJwy+F
6/+KUMiBTAy7HF58I/42PtSKJmCgCvu2EXPqR9Ul9xrL200e2lnZ0Oxfi6KSGY4Z
i7qfK7M2wcz+/H9uToCe16khlkRUAyZCyndS61/lGj6rYayGgoU2GhG4AkOVih5u
LXC8nCr8NImyrnUpDz3cd704RwFkD2Mi0SjCXJlPckP0thSslq4qvH1QrkRuPtDz
fZV45P4egmc5KzCgGgBq1rHQPwj2Vh33Q1swhRzhVGzKo/VWCsRshn9YCI7oHLQi
GAvjbf71NwIQjdXrKccFYeTTT40grWb3zitkfyXleP8Kgs5FEPeKhJp9/Am+aJn1
JtB2GnwoUyJIfBUWrE+mthQUK/n4f+Gc8UizRUI2iEAiqroyyIB+cExvx+zsHWeK
9uudDQ9+yNO+n4ZLMXtKAGQaazj7uU4bPuhNQRszFAvwKYf94fjAJKKvvMwVxZF5
hUhFsh7oqeX6zJqOfgCfODXiP9nNsilb+YBXaFZZbjuuE5/OunvIuGFJk8Ca7eqJ
PPQr0NtafNMy4CCSn0KOCJVKVwZmpxunGvaZWRjxAjqBpQjIRHXXNErBORSu51lC
Lk0f9YV+6HlcVU3JXxojUMMSO/2wkQ+VKkS1To/pH+t9vnk68NHYVHHEcCwgYJxR
iQE1T2DqKo/Q5zEm8rDVmF5UzTZpifhYDYUgAFai9PB4KYjuycinMHgsuW8Jay4n
dvYVbipnb3Ce4WULGjUQyROMYbrwofmg3MNQFmsRcwggnbH0jYVd7WDVNZjapH2k
UR2NFx6Dt3XRFc6V9cmxObUnLebTmRjS6B94JrfQ0KhcvwKDEe10ehH+0jjivgLn
ybcjdUg9Ux1GyEfMT075oN0Ji/R5hkCjxoN1hPQwl177XQuBZlNGbvRjj8Vgf4wd
mNA+eUCmI658r6lqz9UVXsA32gAj7Klq3R3W3bWKmAffDwVOvozHQZ4HTmwtdMRO
lEp23RgTrIyEQ+9isUYctOCcnRS6xsO2O+pPGlDHIlTiAxvLFvLSbHQiI0ZFNKi0
BNmjIhAM/ZOPA/9vWWJseekufn1se4uIse/rpCr0YcfKoL0L+uJusqHEHyXVNs34
gVRrZlLc2trv+Oo18OkiSAhs5wA8W4lhtO4o930xaSx5tQxVptv2LCWORlKICrNg
uMRKbhOxXTk5wfFYJXJR2CYQo+3L4RzB5bmq7+IXnLXTTBMvdr4ACDmJclwpA1h9
XyqL/9HDbDijLMMlYYviU2Th8OJVcZlXc6SR+6PpE+M6nsRUPrteWJI+K/0UyD6C
jyNxxmsyo9H4p46jRHmNF+hP6Wxut1sPtpmw4DZHGGF7UNASGLhtLHR5STWp7pyI
TALW1QFuDXY5v7rPgn25Gk4bt3ZrYRtWmIXaS2ytGw7RoZXpbaBNlq7Z41Avhpop
1y9BgmQ7gVipnU44PumrzKdUPqcgn5GGouxhKBwwnqlxXnZhm1pd//mHUjXcqnxg
vbo0RWX6FO0fsssOOp6rWBKZvOMvWTwn9Y1QvibWUO+tYNUdaIZnHgpQMKHaI3OF
vaQNZErFnFmM+uulcVtFQmuk5ECtCLCejAMn90MH1rmieNeTryoN4/hjPqIEgX2S
f8xOxl9LSsMO1bTkq+9qBpQ3tzYBjHjZOjQ3XMyPeg/6bykWyCVG6kmMfEONjKBH
nLyEuvp9Lg3+iiAW5lzGxVYU3KUKd0zv3PmjpeRLL3gfGBFPBZos4Hum6W1mWKaU
4v/HbQPOjtyZ0jC5D6jYqr+mnjZaDPzpk9e5aeLpspWb0s4B4qbwtGtQpgsGcKI5
ODbWYv549kRsdXGjefQRiSGbpiOA3OGn8Tj2AU3PII75OdGEerJnMK1+zfBdqIfg
9lEenVFGATodVKPyrbxR6qPfysmbHVpVieoXWhO5UqaZ0EaHeI5qlgbxw8nnh3Lq
65g0SlqA5wgs8Fwnh4KpWwzAls8GY3GBXRx5cN5dylvM92GGxVpgjvwK+3EZ1qHv
8s6TerZiksP9OVneXKlFY//ZydW/RUuKbOOuIthJDozEFn+1UNeJgKrrvarDctjd
ck+Jxwf8I5Tq1+HMvqFsas71OHdzbq0X6JoJnJhr3WX4pPLe8WTkGTORUT1e95OM
EsLYTa0rn0zBlnBOlP2BG8LvJbFwibpJSHCrT42/M9c+th/eMZKV4HwUGQgtGcyF
tmy0RbfgORxK9Fo1+jUcsflo804ut95Sn13sko+cNt9a+cIqBKyRgGMAzpTOg2be
Bdwy00fM42a3Tx5LSrrwExVp1tD76UmORLDXX2IWfmqfvFOnK6DRg6BZhqcRLwTt
s9Le/alu4HUj6PqXMvD6y0GcdSniyVW70GpDvqace+JWO8TlgU2+OMqSv0H8duwc
vNWlGxfLd2evfGMUP10yiToAj1uNQd8PRb1rKbQtb2z1IuPZfymuWLBmtx/TkavW
eYaDJHz28t8mGURjRV1SmhX2/ME9icT4woFKlQZFpo1IEWU7aYo3fyQ09cFpOR0t
NLfKAwt5cCZyjTv/WpRH87GgEz8GFXKapI8wQDCJSOOc0KKme/wKVkQxBHCWM0WR
jKO3LzrAhT0oeclZypg/SUx4pUPW/U1G4LzfCOOmQIIYtkbZ9dNXVLzKSmj5a7DW
sKwVg+fIpq2LHjXjOy/X0GA3uQYvsYz4ppY2sQ4UeaSiA41oouxAokEeDgEwX1WE
NELv1zzNprn4UmjQpYy5Vcj+lsKTD/IM3oFdu5uvXlZNSGjfzWpKtLXTFtQahUle
TfVrSGqhp4dQkM+WltUIQ8gGwCWr8fgvt3+Et1pJ2TeS8/b0f07JGYZanapFJ/ja
RUe6hVFLG4N+VaPDpAiKobCyWN7KZlDPQd4eh+unj9+tfV6yIXPVqfT4ZZWkzAGi
cXXtI2owW5FIuZGUIjSWOkY2qfEMCEOVyLJ6vGTG4Tg/gT8k8Z+yYanzY0REBp00
SkgZCMqsmj5+ClVQSAsBx5+o5oZBqnGc8lQStmz2ZFBbsVYdXw7LYKwj8GwVZtmF
qQiIdc7QnPEsEHThDIQ+rUhpl+yOAjWju51LHyT0vC6GTNAsKW9t2yDeboitA5/h
81UvKrxGeiEQ0LmtD/L1wklVVahR1rbOdFywe/KokYxyv5PR2o/5fo0hu+xLVDBn
qI3wbktbXaFs47Y6rEJMUCsr8UrxTDe3MmCc6ZQH1SztjUMzcu7Qn3EZci2IlvnQ
fk4KgDxq8+OPcnMm96vDKgIZH35ZEmW9Hk1tv7pHGuBiH4T/A+oIGur8ojl/LLKf
B6jJaSDnb542AfOJdWJdSjtYDcIkzX3Kuypfs18PBUUUnwhW9kyxiZTDxkJ89Jg5
sCCXwYWrGK9vc2q0Nk9Yb+d89tCdO1/WAVHB5Az1eQhNTzXUa3BbmPL/jnzlXXQz
kOcKD41toGhE+imX54ZvdMJ8Ri4Ju/sIkzJ0VEeH8TX+HBnYUkUVbjKlmH/Hf59k
cRnSGuEYWKcZQJk3J7jE7FpV/I46HEq/8bPRCibd1zQ94yLhY+SVPwmXg/dJqEBg
q/GwV93Wo3Q0ov1fUSprBPuBbtyQbbEdIKNW9P974N9Zi9zSB+HLtpVsL2TykmgE
8bU/1O6NXSVQM4/fgPIIoonOgLHx3BHYOg2dlU2JXUK5EU8/5usm5XSruYA/Z60f
qDJHiT7BBy0Ms7sKyfvQGke9OP57dUDLdOaiExLepP3Rca3mugpY2gCuwRDKKbeg
vuhyESKZ/+t8Px5EulrSarfUaEsHHTSWNM8OEr7jdSYIOop41nZWTuWwkvBzDx8F
SLumTLMBJYcIhmlX8vAgHdij305Cawz523vD1uLhF0oX2g6k05NwQEBop95rZoOx
VXsssmYOMzlpVmdoK+KGrG3CdPHQho8wJU7xS0XRGMBy63wKULrxY0LJtqki3ZwX
e6fQ6EoJl7nNwSwm239b+iP6wWNYS7VfFmb5xoMk+IlcRNuHOV11JaszIdtTNH0U
+aHdMbi0xg++jYDZokSqXj4xlpd5CT1nukr0hCla+/YxG64Sso9pqV9cJaj9UAMm
bZUuTvIJx5vXJuroO/Ee/6n+75jmwFAaV24ONITevdUx+DiFLY06HpLFQCax8ZcR
W+G18cdAohSDDFNc0cpEPEfDKH9iCJ9PGktPB8vcFIGPdrED4Y42XIIA6ZrWef9M
IuVKXfFtriTgWEM4PIyGl9liTZioUULKHMpylZuZikU1HwXpaC6JDIB6WNL1w8TM
CT9Rj8LH39PC28JrnI/z4vgFYUOlomVCnw1Jzkrb+y59F5Dhh79tD65XA2n+t7F5
0NQyGTb3Y3UAMPn8It3idYTJwcFqAgG7aMD0NBjxVOmz3bZkFXjyO2JOAVvYgdfc
grWHk+xBmY/zO5175wy0jQve9FoWQgyKeWMBvormmPGilEK3QC/kgOF1AI63kl+v
2nQ8zpB5djmKdh4Jt+YWWWcWgv6H3TdYt006yIuin0KSVLHMimTdREJnQpi1MlNG
HDmDxYL+FFDbNT//lB3Z05d25lcA+Tc51CFQ1V+jA0cDUAmWQ4x7Bls7vnkjhiGT
/8DQ9kpuw/pwj4MPzfkIFVkiHQ55ndLMuYV7B5IdO8XkUDee8abNKInNTwXy7zd6
h0HnONKLQqZadEGVCak+sZbdAKWQXxvZLkltyCLH1n6hvVtD/MqjRAf+KdHWyoEU
ymEJx4VLBJkW7ez2h3LHUAuPY2IkGV21YW7DajClTXBfYBQIuLKa0jsW0HWluFuf
BD5/R95j/QXJfPXJzFC5J71XD6/zW7v5Ru12DJG/h4K4b9ueCQiT7Zg/EUT36N4K
eE/PjraIVIKyzJd3ngBqAfy9O7A418M0rGsakCPqq6jbZjj7VnV18DLilpvXL/oG
tH/Sw9K7vW59BKvlamjmzWSLAlr2zTDRiGk5bRkiBd7HFojQpoZ7i/8csgL+Hpcy
j2PHgtIB5s4R2WaIJC1t+xXvvKzULOTGDo6jPpTVwqu4fiaW0m2ssgNC0Cy7djfv
jpx83fzeSvVS0KEmtNm/rsIbvSPuCCDrdZmTRsKjyGpo0drDkcAydrhgldPltaYv
ANiNxzR6SZnFXUBkJ7SmxJ03bdeiSXkZ4r/jjQPnb0WasBxHQ3UabC5ylgpZYDP/
ha/2msIRNPH3lO4t+3F8XqrIEpwCfWCjQ9cwUAWTZ2zVopwIQ2PRTbs3x+3bLopq
cYKs679sEiC9iScoTFd6Xg2pwd8Hx036JcLEg8MnH7/f5nkqe4RdnPB1XtqSr2w9
kYcOxMOatsW6kjdkj03/bV4oto96NEriKbjZen5dJmnbw/G++dkTN1xVnbQm6tnz
dUCPe7wjvBr+jR8Eh4gS+WWtQdacM4JTVXaahZzChaIozqLGGzdvO8xxEA1DK9GY
7Exszj4VZaPPt5Vvo/D1PpHA8aeVpzK1A6qcrsfsqAWSRJvGAOG0O90d3RkF0mlH
MfEI5JSUxVn5AFivETMLpFI4NnQD/AkHBWNiAWvxt2ElJWPyIFOgLtM+ixc3OnjR
z0ICATZITTh3/qcWjGK+T+fn4MjQaXBkxaJsfa15VxTpZUIHztlntdhttMg4JR/D
lqm6+UPSSBQofmnJ3HSKcXX8eLq5/lIWwAM5ZgNc9X0T/8MmqZRLJ+6tIPfH34Sp
wZwPLZCiekr+2r2iya0/Eh3B+Jbh26OAvHPFCGbGXLPo+IytHqqFluHKjSM/8n9m
UnBoemqd6IsZQrin68x5tBgl/uxpRjMw5aPavP5ik1v1etPgFBlOefJDkr6BSGij
Ss8h/DQqpPxw3+Vb4VRt+Gb4cj0KGZJaH2Sry4/WjLaa7j+nInSjEspEoiKzh2VW
urwsS2NPUJO094jmMgsihQvUadtvrcSw9kxkhAXaupNqIjanhqiE4aTh3AaUOj4h
fgFPp+BSSPxyt4pReMd77IPwr5QX5ul4pxgwghPgaiHCJfGIcZdMsYYcfRMlhj0E
B7S97N7pyJyfkjsNuGQ9TiTGWlzRxZ6ic+reOIMAoLTZ/ZvNNXLgZJgywgVQnRni
jTpq5nvwOcATZTRygCZG8Rlr8QpT6VLRab59s18GmV77Jfjp6poxpSDcfVpa3eI2
YoK2pi5+24FLsZr3wSlWrkuTBh+NGB0Tnc27SG6VF4CHwHG1/i4chMlDAzbV3kvw
sun13nq0IrvW7jhozCeg0badrgyIWDJzVl6BVYF8e2V5p2wZwKCcUBe+4XKTN01Y
yZMALzJmNGkVDifN7IfZETPvaZXACvGo6P0H31d3DoKM0zqMjKChvYQsOWMRsJtG
rgyu8P/bOSc6cuPUT0YAPhcebolQ4bfwRutzMmqN9kB2TPW8FNvSoaktMYGBpUci
i1QECBZtqWUbA3atPKUAOrnTaHAP/FMDNXJ04iEChq7u7LclfgaZVtdeK+tru8EV
LT+E2qguEIJ5WxOIEzrJK/pF9q+DqtLHwuMcirAOg/WIYO8GUVx61XrUb386cAuf
1qm9HYD+I+1Kif7vy3hmrQN/OgEOHBdWDTF7q4qpMWdVtI4VU4MVrZWLck021JGg
pZtCM9uYCPTOJbNo2wXvMwKMT8Z2CqT/wZDTyw601XuORAHi6x3SS3T6g0ufRAt2
GleXn4o3If5Wbe6pJU+ch14vJE8HaNai869B+Or0Pu06ybh2F5NS3o3Zaz/t+EWz
YpJRZl2cal7ebYLneLyju8qMZqA2sygZr6NBL3ecg1RVuw6mAqoMz9lQCTe/XcJM
1rjuTE/1fFcPv69wDPd1DLWIJljW/I7zkM5YLvlm0FbqKJu4t6gbUl5NacvO28VH
HkNqVDUOBppTqDaMO4/Nr2obCyeLzjHl7sgMxDRBcfMf2b8iGUFrVRnpLHKcN83L
TOI/82YKCB7twHydiwonNPXhizHg0ftpGjh6oghOczSReJVY0nGREtnqf6JgvYhQ
4pa5Loh97UjK7qfd7BXFH2YYi0LS/Tw9LyzPMHPJNVNy6E+F9nxt1uEvJyHCIm3J
dfoGf2XsDpmfOZ41OYul41H4csaHtyfkvWIBExAJTs6hSeRBmaxAbWYDvorF2ktk
LXxfax2jN4rBCO3RbHQNrB4A26Mcce74lCHJlsNIAD6MFG8+p0Q+DjwmwKdpucFN
LQGQel3Lo0D3YPSbRILN6LZy66HrhS5equuPQ4U7ZBADLuUgjpSr8l0wZAQ9oRLs
iu1BuY1z0PP7vFgCwzTH8Njvap9nL4A7LSt2Ye1OZB2P3ZJk+Ss0UeXoEwn9xgaZ
mYnXHz1+fpywX8GyLMlTMw/yPwcNFOpuR65dHg4VotOkNh2JEMXd9i6HC98EAfGt
8Ayx1aojkuvNpEugGBP+Z/Hvp/3f26ah2pwCeHraKB+tdM31XoZaDftaBh05rDoY
QQG81+g2FEk46yR4d0zpYZyVUzd7RPSEkrBIyuvkdGf+mn4DvUXzlf+miSDH9m/d
VrJznn8MyQcBSH1R5WtyGYU2lH6lC1Rl18h/TM5zDzWoGko7ce5k0i6MfRSpK9qA
B9R/nSQgxyeU4LUbnOCD0tvj2S8jz8SMzCOQ88a8I+SBexFpE9nqnojT9eCyWdiu
/UAHCLSICOES5ePzZYvIzzs6cajAjCwsOVoUMMVfQrH5hLI9Ob3XEBB97QDkf3si
IdYxn3lDdRg2H8+0m3GQSmjdLrrnNq/yJ8OAIsxe/TVuEVtfnWdPx3jxUXv7/pq6
3Syyy4F4ewJZLNPFxe4IwiCNVgl6mDcON6E8OAJQdCiZOoVelL1CCRqHnY7fJpnt
1Gm2sV2hQ+lmuHQdNZo22fKxgv0tnYwaJFukt0XiXyvmpPHCasHJClv2FEMTC8cP
+pgPyTua/p8waUAZmtWXydqwHAP8MHAwIJrrHONSPdkdnxMfW7IqBDJhnIhY8SDG
/l1Uwzoz0NtyKQ7SrVoCH3rlUvG8pJXeasRvbw96V/rGQwTWnZV/9ansnPzBhTOg
ix+bwC24XbBAAs2T9X5DMBNI8+HFi9RnNYhxdm3wW4rLwZ9WavGgEsTHPz63l2KZ
B/y6VfJ5yfR26jvXX1Q02meJp6u4vHdARQqs46oeWwHbVdC3IJVuHKV4pK3GvV0b
qkRQuJKibUbzwCou8H18higeWxCakU/lFR23pDLVz8268/rcWJJC0Q7TiHBrSHc8
Oa0Oe48JbCAl/TUF6h5AIdln9kxbt3rhDUaORoftwBdM3FSbmqH0Ri+c7JJ9R5w5
W+70kaDTfdYh7NF7rC5UvaIiLlGp73SsJLyG9tfZtPyiBACSQ/Ko61Nt8DeS1A98
E1BSdHw+HaT5h2cJ3k9kN5M7MxQOf+N7OGVlH3XeLOmyncZ3JUPbJnFpMe9WTGx6
Yl1XrolfJUjWp3aL+FmNpppXZdw/ll1u/a2XNTfF+j2Jbg6p5//PkmzLmqHXJzj2
7b3Oo3x4v69dtuwy8l4eAjZKFQvUetsXWJAfYjAuaQ3VgQw3q4O4TCjeqCoyoMjT
WdrPnSzZ5B6qxw0rmNd42+jbz7A2jTixaxLZ+L8CibRQNQOPV8K0IlhN9iXdgmQo
7n4pP5tMMAdg5a59LosqxUydNhKBaFWMqEQBBg6d3Mp87X38Ed1lqpae3ceQhruh
a5iBZnyMl8JgVBXG5a0+C4noDhZfK9gyGwgEw5tmuT3mHAQ8DMbeOxIg0uVAk4A6
GXVlWOBsF/1ExAn73076OAO2gewTi2CcpZtlHfX3mZgZS+KLRWBd0osfrMps4SzO
sI2uyi+Uye7PFKfuMlia3rZsb4d0PzK8Jml+IRbhxAP3IWibGPQxyMoFqjkQN4F3
L6mW9CUk1alZ6zfleeFqzuo9hTcU3Xao+efDeMXm+/2yg+UigmrBCVjQFfQwX89w
ekDnLYTdwTWj6FTyz9VzsM+GFuf+j/Cmi7/IgHviFC8Qlgiv1fk5WVXn3QIsR/5K
UqoFfLn3A7L78BBHkWMgPADTpTDQBPRG+WSOcyODQLWvmQ8TLOGoIM8tv8e15oDQ
Fqf4euBnyyzBPuiSKIwDPozttTUPn+k4fCu5trAYSyXhqrzYWzsKa6pngCi20GZ4
SDCkzkOCZ6WL30izPTZHOgm59umirGNsUFPQI0o4WZL7h6LNaj70tgv6Puh3hFTB
VNtH6BH7RzAwRI7oBv55QU8yAbR5+g+0dwli7H0lRBU93WvAf6HN2v7q3J0Dt00c
sHJtsu3c6gibe8qOSl0/6HvqOxThlk2kGA0ZMXXg9SxwwVaHv6AGv176gPGvo//e
JAf5MMVHvzuTaXFaKviDkUEoG7/yldxOcOMhF0fDDDxmG9+WW40wMH58GFsebQqx
PjMohr6OibKLa8474T/gasGbPj3MPu4WlbMwsiMkfjcJ62lFynD5nnroHvZe8O/l
l8HCRVk4+JVw4rB0ZMTAvfUmCLHC0h5M7gsxEaYM1nswcGDRjOQRqU5sf4Ne+C2P
4LCCco344erKSWAE7Q1HbR1W8ngKjjNUO0Y3Jvh3StSMAjujawE1nKb3f//3ydxO
r7DQbAZefsOx3ldD94ztMAUCaminnUY4ZmyknA9B5QGgJ3NhOTXCJQcSYkRXOIS+
mR5i5UEie2179RtSjuKFCAUtEBHTaOIkdWdHjDdsm7u0F5ImoMOvaZ6+fFZy8VoV
xJMkv7FEguQ1tNRzu8Ly7qAhPZrR8RTM0FavL/1FgaUUf2rFMbrG4cyg+Qg+CtcZ
ikPaTS3OaYQ+vO7Qk7gHCstDFfYwRDm7VIXplhtyFgCL4NeWa5n1WPhInvh9bBc+
XcvJC+lNEY378W2CD5RqHxbliKhH4NOBDI5P1cH1tEBOmbWijRQTHfpajGjeLRgG
CejFL9aulYwbQipgMjvwWTWgQqu/AhmrRjgQifnFWHfMkZdz1B678xgMy5SgRRAo
40a2qBezBSF8AYgYrW04IRf/JjGfBMPpc/XnGelTMXkChCkGJIvy46ICZflIoWYl
Z7gMeYnn6sCP42ujSstV/hOEtCKvGRY6w0TQsnN4D2PEhXygMQbUrbeizmW2WieV
UQYOw1+PG9cRNYtI4tsWZps1heYLvPCYEBxSJfJyK65Bj2R79B1DdyRN1e1Q0m2e
sPb0SgYymCv3kXOSPt3Djvy+YjMJHJFcJ0QODYP0qExs0JfuY1AsdQfftckEGuhv
aiy4h6WjWeWke4V29J+UjLfSz3c2gjlVt4okq+MogpiuFt8hFJdRRbo2k01E1xg3
hvjYFQV5PD+gnJL2cCPrYetZF54/1b3c/aoE5lGv1kTxpy156JXi/Qw3yDZw5o66
hpnPsrKSxszvFLKoot1ZFQjLoupfibbwpXaiUVrH7D/fgGFYPzRLH0mk6EezYGxc
GZb0iSmS30tufaXx7LE5JmWwlDXf7/6IysW7BhMdYWLVngTcN1WoY+Ol3ZKEX3KR
Q74pQL2ar3u20DhHys/tk+yMpgsGdGmOfkwMWDaD1M/zKnLXhLUz20ZolTMNFqXT
eAt5tNuW6W4OC16/YZlhFNzfGggfiOBP0I1AR1zwXyjnQ4SHmsIrDwOFJmRkkdge
o1bL7k9MB1ZGkrdmSjdRVG4OLn050tHy1sqO5bQHobkv+UiC++wHNCMBdiu2BxJ3
ScUt3vS7ZyfrphuGZWR6vmCqh748U1DEBqxHeaorPT9v7LJbyqADOpFpfJv+DI/G
9CmvZzfF6w8bg1yPy4ufC+f/uUk0tNiyM0mzJYOo/DL0lxrZjfnuIyeof4XbDtIk
rS2TpZ+2Hz22k4B4738K6DUykDikJjNlLhjDT3NriYEkfGrGh4NaK6bwU08ZlEQ+
qQqhfPYWyICabCWyJJEqXQeI3Of0qKr+OtuTpzWr7Qy4XwVfQ4XW/UOl3lpLggGn
OBI+Iq0I415wuPADLKZMWK1ZMEwkWULXFBD2tiQ8/6oBfZHjVe0U1/oEM2saXCNP
SUqe3mijvxlZ3cNihw7PTgrpyefijlKJi2mCAbuQR26B/7b3I1nLa55Aeri3r1Bu
luKbL3cz2eUOLgtnPlIbCIdqhXKbSvazb5WOjElYfTJJX2b9Kz82FeRzX5Fulue8
DA5+dzRFU7HIC82P5iVhAqTzPSedBjqbLGwTUG1uetsjbgPUPjtNKEoGU8A7RsR7
OCyPy21qbUkG+0meQHHjirfNrIdfLvFxXW0/KKwLigpjk7K9vgb2ZPbCypyBFATK
8GVf5JtFTHhZxNWXs24o7O3KcUu8iNdgPd6qEEiSKIi64Ysnn7dUi2z6OvWwxmO7
UrZYNmO/DPyMHNy+j/hhx3l1rZ8KaoI2F04dYXOd+o+dkwpNH+PZsfApleJNKDF8
HYV0CNwJIJtuxiMQ3GmYDLvHCMjdG0MQrZmOKIia0YNmwd/k0aI3vgWHbN7vgrfR
QJoBtIT2TUlqedgw8ZU4hmyWdr/hHCA73yCsDUFBc7giczNE1ltXnZkFrcbtKHeM
4nabMhP5cBn2SwY13m6IhkPpxF/RWcU1sPgB4QPZ+OvfLEMvviaF/JiqKV4XNs3I
Nwt7skzg8zbjcYUNEbeiLE6Sh5q3LZ3PbNtRxfVB+MT5NM71+CMWzqJH7L6sNR0X
Sm28vylIpUZk2qYq+2jYIKvZM6mvlzLy5TFOc7HH3KUHOz2X6az79AolY5wN5JYR
/GbRueot7CRH++9b6HxqSr07FtWKO0RhWePyWIwDjTuhayIrwcHjCFtUrryRHAlx
e/G5CEAW2NjmU0MLe71naVhebp0WmjCCQ3Kp+edGnXIQvF9rHAbptH9KI9/UWqhX
agyIi/lTiJfcN5PUS3rRgSweKaxJKKtUD8c8VIAofH+fOjMAQFkyppRZfmS1U1n1
uoF850bZBmxrtzOaQDH9GkfLkKZxWv6vKke8vGPtFjkuUfCFoBIIx1s0YR5AtODl
OQt/Cow/ONDhc33L0EmDlfJ0Wh2Xk29n+Y6lpszFz8UGzg6vq8L8jVEjyKxnzS28
1I88fldY8g/Qm1PcrzszhBqAu8TdAF2kEQKgdzV0t+DI906m115sK/EuPEmzzHMB
a+0Ep9H1KTCKhBHTaUCPKeMDx9YMZ41D9M68pMLPe5Oi7tpw77PnEea8ZYSnjBmn
UDS3bqXNJW7e3kJ2zpHU/JT2y9ftIlrjEtEbpkLpYselFY3zH/viKOsY474nil6u
hqk8oF4OxQynE3Vu9u/bkSOnX1KB9CK7Ik9Pi3TJBeB3pQJKhUq50/P51PzuGCmy
eBjsbrPPrretCzbLU2mZoRncY3DcnnqpmGIvJ787MGFRl7HYN2v3Kju0S5UFCRPk
H4B01vGoikMX7SWo+8VELc6k6BaXjJVNkzmDA0A/f7J0uaJHKIP6wqjqRorLn8d9
/ygQB/vBlV+5TLDRapo3lvAM/H9t/ejLyzy3Ojje8uO8T1Hg5GFO3RMyLJPYAaCo
ImlFCXIObi1r5J3KheZZDMgh0T2EiH4zD7oysbuKonomAQ7MVYGX14IoKbmtPOKp
NKMsI0mMwqvgtSYnHdXnH93M5qbvajGolB74+9FNgNTXS9hzY3PjSDbg7kM1MNNT
VA19oqJYciEuKejxOxHp5tZ1wkrobAHfQPA4PbJtjwJ044xirHzFlhbq86dZz9DG
9TK8/sl9k2g+6mkbWIzjVhHWWiZ/oMwMR+FfJh3hWB/Oy8ifInl6eZXaowSfq4Rp
61qlFa4LhO/Ecoiq0viMqEjeL4FkhBXrI5X38IwrA9ttoV5bODt0ro3R2sQ9hgD8
UI+7yK48TYlaWP/4vibrX+kP8rBqDeu2v7YelnKQGafG8zBNWEMmV/LgKNMXfXBO
APORJ54VLhcoed3wVptq84Ivzob9FfHMdLOGJvo60LeNQSzGkvqDPxxVmMVODRaW
YqFktD3Pd7nEFV2M5y3efTBhFuMjK1aLPJHqB6kCeHrF4MitSpM1pyYEr2F9kjxs
LaE2ABzF5U9QyVv/W/pC+JQxp+zOFUPJjoV2s1qNBiN83VV3uA5uLAAUMvU1Wn6z
nQ19KfSih0iXQuJs+frA7NF/FPtE5r5UoqvMpHIW6Q5kO+YWcdTl/TRABtVpched
IuZNccldqbu01+IcZ0qO8F/tpN43JBxnegGrWcExw8/SLGHpsggR4Owyo2CTxVds
ddioa0k7USQM4iyFOIP2tWIHPtm6FnrFS6ZOR5ab+ldL6PsgCLuk0QNBz9BF7hlM
pVzHlPtn9ULgMB36Bn47MhW/kFmKVR17qLDk1ZkdDzcnE5RsjbLTac1uzYUTsB/I
WMZViwJCd686CfeR+wspBVkKZeK3f0dBKtBYUnrixjkz6Iz9/+458CFlSY3McjCE
S1Vi6/CgTPqdRS9dw7CCDuRzXINTHe0zDeC/IsciElaebv1xzabXx7RtM0BlcIGV
bOvzk3RsJ8d24i2SPSCZtTZrslpXR7b4djmHtK6dG/UU75TQ3jFri9wj+9rCO/An
y8+T6Xp1qK7/ZhgmiOPmywzh9QpU0pXeS02tH+T3j3chuGNi06va2AFrz0yDzuvL
O3ZMfpeK34fGT6c6b0Pq/yFhJLvmPkuRv+j3DP4wmnraDNqAfY/BIE0zK66Jq6ct
LnO0KLy+2Gj4/Vgs2ng09aXurrczGpRb0KsxSJJsCcCKbpqrGLER9qLov7se+2Br
5gyNjVXxvHq9BQG4DpaeoXsXjq343xOIMlNIPnzraBkpL2/WXfwcsjz/cjbTFRMC
EXQEJTYXVTndQapvztXNx1pM5YwbXf6bo9MtqyKQZn5dl5Ncy3VVbh1wHWzVpYmL
lwCMgjH0hleQuWsaGMbYPFS96C3CdScwSRIZTAj32qofrqGBz75ivb6cStGWq/Wo
FgC1DeEjs3RO/nlP6ih4BUW59PTeIQSXQ1Mn9BcAc6tYl1hYZNY/4ZmSgXp2N+ND
+daI80LaKaZwb2TV5A5W4aIqaAzBHSXn7TDyYzST+B9j8Hnw2Kzao43dZwOwlPwV
2TrRhkEjp+B3L0MNykePJN7i8P+PKGUF3S4syz2o4vz5sr/oYlJZpNw4Ap+f1Akk
FIO87LK6GdSY1IrZw5Ti4o0A4AlPAx5NJZxKw21emi0F1HlvsbttFYKUVCpUWueT
eq1y51dlkxZhnCL85SO7uX7agkzCGmq7tZhiQ9B6SigC+ekHZZHPlAT+9Ab42dRX
D4I0R6+qK8L+j9WaQUyY8WzoNGHG0tjOAvz/TrSJofrtn3FTShMMrSoGvtco5AsA
Ewc/ahuKtLDhftRBo9B+fRQQCGWQ1+9goT7tpnx6X+bAfC2OnFvWEeQr4TGioyxl
wBL09s3R5+FBlgBRRIf9pWa+CCV/crMZ3LXeYCgT7wVQBuzOVjIl4VjS+DAxjGFE
1WQrFNerTaqZ0lC4lEib8zjcnX6t+6L8IpBTHylIXCnN03eq5lSoiE42I5yjD/9Q
Z/UFU1i1woFdP5CPSl2VCl7vAAoBFszIOls2mRwv5tqmdJYdc0UI31tu2BB70b5j
zz4f5NHpDgc1cHm0G5Y+1QEowNdpzW4OkkaW4OThxJmlrDHdmDzHxsmP/wQDIPYx
gGaZEIJAQxzwEZdOCfKmfZ5Sk9EPO+9bAKr73bxUC/flogABp0KyC3iHJCyD7F+m
AbOJStw83o7v6sHPkrcr5JFufGyp3ubbOJBsGUGtN67ar4AI7VqY1r8WRicuSR4F
vmXz9fxAykm01/Jrs/v6TDYutQcyqGQhJXw2CJXPGJLlaI0jP1xhwGRMAGtz8zgT
0uwAf86SiQBAsC+ai4ZRK2KNlgW0FFr1ay3d6P24CvrisjPsmg13RbcSmX02wo5p
SZotomnRUjzKfWD/QaaWEArIJJ6PDhSa1FipZ+5PZF86ydS7xxFpeMyqi9KreIIb
v31MSGoXJJNFDiGHVjTIXr4AVDeN3VFsOxrwwBoPIa5WicaSpdETzIUKZsO9Rh8o
CUF6VypADWwIpUo2mWNvWsDf1atSIS8ukzgKzNcAArp/yeMUn2vJPYkg6BIbVhI8
yQuzQ4gkw4fkQzVSIkbYwFAUrGwDf37fc6AA3CFpXLqkN5JLb90PHiw+QToUFgOl
lHONXSIqTL+rhR5/TiLsqgqA2Dy6hmxkclirjFl0ZgmV2DTDfQHstjg5hhCX7ajT
89ZoNI7ZiJl6JVomuGO8jHyNL6BOg/WXid0d3bif+1ji57w3VXoJFyZM6Qtb2VKS
tFV864UgxmTyCH0r+SFw7rTlDVGCpDSg71Ly/ymBfq1rYUzxVelWggFeGqBURMYP
nb0/sTcrpnNWhxFDhYeQzUeAbHVwY9H3Y2fk4Jr/8c0bJaxVixAxpoFSYZGRXhtZ
hvx7ZkZGvoW8nnbNFbwD995vKxzIy9eBBwkvPZZl+dnUw+zPqRtTch90azdV1rOj
svxfzi/gVhaPPfwN/G0TUWOhSgeZTBexpQEOz1oya93f4fJjLQeDUM/o2T1C8mN/
dU07SjzpsElRDBKZAJgpUXm4zzJK5c8T2eX0i8Mm0Yw/chS52xIghhchHdoTeEIX
Mj63QIKZ0V/QOROv6PaMKr1ewyCaJb1OySmN3aZbAk6JIn7CyRqbRjzBvnk/fz65
OyxNlOrzxqxphZzYVmLbPPlSnhQQB/aXIpr2zCvzYfHHN63V5h6hqtzSw0JENnjC
AZCkZDmuquUYG17A0dWuM8GhCKuFwoWqN4mxZbyLdtKD3lYXWP4XY2L3OmSmV0WC
E1LAbcNF031ImQzBe5y1x0Xbt55BJBxKyrsjQBCh6/rs5piSvhDPToeyO1Fiit8l
XSFU5F9ePOMJ4sp+bJL1PWVyg9+LpfhPJzhy1v9AVLWs/iwOKZLNGpGpiEoORThd
hQ1shqDLzDvkUnHHWtC2TqCHumt/jK/KlGfGOSD814lboPTRmVekabFdJafxShiS
v1eg/oxquKhxQimXMlcanuewdRqzzwucu1v7qTOTEV3x8vCB1U4is/sVNiMkwqzN
dF/u0Ce9ZP/nO20dplqztWOS9meOuzC1M7uaLpzlPyq8DxHhElxDbtiwl9sDc7xW
cKnxG4Z/vNiZRMw9dy7bBaTLa4cPOGdKYI5v6XDtUckRF8aowrmOcXlBWlKwcqpF
ZFj163vHBRqLTSg0pkJOiqNQtchsDQPAXr6jhi1X4r2ikm6klXH6aI2oEdbifEkO
wYdHkqZR9iDuEZNZUv8q9on+WjezI9tyKhg+FMGPsQtHyWPp8QSBdjBINdjg2pvj
NgePMQe5SslnEI+C6q6dlp3kTkrHnpsQ8Y2zv3qDQoszYBs1yr3CkDTghKp24xmQ
ysoa3gCpm98XgFO2DQDClfquKq4baADYcUnJsT/XXeBnMK+o7KSf6d/GzEE0i9Nh
DmKZmOzd/FnJyhIdEozIlQ==
`pragma protect end_protected
