// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:32:37 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
VaRc438jKY5su7b2g6uZXyv4k9b5aPPYIKlIyVTwLQ+g+krySyMTeapUlq5gCGoe
JFPx6stjUdq5iyzXNKFCuiwN+OYGgIUZyNUMSM7wVoJ3P+H6V5o8ATOfqPleHBhv
Q9N+II7Xxm1CqFqQ4CLwrT272GBM+VGDB7SgWbhRLpo=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 71088)
dW4NFgHbN7xShdHQ3Vv00Epyilo8aYoGjXhlIgHdjoD65ZpXC/i4DBT1tlPYgP0f
NMJS+o6v5XgIji0OsXabnUikQc9xNSL5NAAQnQ3bCM0zI4P+o1DHaL6DCzLWctRI
sJA3Y7zLjDKlYRCQtrXBrbFbK46yLelCHfP484jX8KZh0k5T5R3rUxocHfVd1sBx
2jQIxUkdkCBkhghisbnsw0hWaIgpjqSL5OvmW1N4kpVjXQyWb3q1wlgebei5VwOE
UjRuTGC+tje933PGvg0k/wFZjsi1M7qAMMP69W/hjLGEwMuGAmN6Wk4QMfIHGA+k
HU70Pf9MsUgNXeYpsAKSYrldlqjDEc/Q7l4PZVTS7YYxZDMAsT3ETFKIeOvXjnSI
44S1sEf6nvQyTQs+C06SFciUDslj4FuH571ifXzo8Cp1DFI2OAQgVQZeO9bIWhwA
HvJoi92I+EBVoWcwWt2ylgpxW4H4geaSCUW9aFoqLnbPqkfFMG5yWrLJmkI2vl/5
J0VQKTrBXXZa87ADT8xFjmpv9VulqxunAnguX24wsiwQ5N2ec+Ryv0SP2GQ+sXEx
WF2LpGXjGusj+yLKAXy+8jLicBk80g0aN9CoMdG6r6AR9wx7yiDkc6Axu+8IkVsl
aCC5lUBQsVkm0U3GHvn3b/GF5rYRITZ1bCJDPqHYcPJnhw50gyrvOa/XV7bCbQtO
EAfhT7HpBFiK17B3ugcVzuiCCcFZ3VVmzvbVi9gLtnIEG5ZPYpK6eFVAZ6v/2eni
xwnSZeFBfNPhq3uKvMbqNuxmsvOgOwLxbwgRKTHurB186bovzDiLSQjPCONNBHge
/jQ45RAPZe1yuYzIoKCnqiNuHMYw+MNR2+VVUk6Ljq38ZFfYkQqcqZkC19dYrl/1
GtUV8AMsxTOkNBrRCyVpc3m1RHTthwuKJAdBNVv52SsP2sRKQpXoSW4t2uzuFQDB
Oha4SJqD5ilzmvNw8KtM2knDau+guC+qXMpsXg3NtMvWeJS+pFHKZmUskJ94lwx1
efySA4RcvD9qoyFXj4Hey2jYjoOHRRFJdbJ/rxN3Kivcfgw8RmI/69ta9ALUIRSg
hIGYo9ZMgIxt6B4RIE574TzADhabpOQAPR0L4/rGku5TTJCxvk433ti0wbdYLWgX
rudYpRJEiitYwQ4muvolXTqo4N4Ng5DfTzIjjQfvMgZ9yf8LvoxWNPdgxsUvwxFT
dUXt/11QeL4cMr6W7OQr7txyBNyUXS+ChgbRNfChUj6Ht+6dATJTf9dHjQ3CCzds
8vgnaGMYKQFceOFAO65c2Z1WvzPOKIRdCzbSgYY+rFlFdrwS6yRJ1K/k3j9H7lqJ
ICb28UwydRJ4TFYlWwcKK47CMeoKR8zPkYogoptcTSqfGW7rSLVM48llMjgXgF/y
GCwlUrtIuqxBo9t7tcNIo5UisPY7kr3v5l2xdOmEViKkQHRfWokFormboYFG2rU7
5AoCtVT0CxTjzt+2pLgD1rq22J77pbpxV8vxVqmaGTlFjS9E+rYtDA3OWgQv5dMX
fi85P3WkPHaxDv5alSNNpH5r74LCOt2DYDWuEgWSJHsJSqi5B7kou7ydIq88SHCZ
Kso6AdKhuUTCQ0JqUBE0J9ZgTZe0lnyYZLpJYBTPOFeVFS6IxbAg0hjY/Tcqpmkt
dtocG9TPzNpegiALemrBr5Zl0mbrk6hHLy/rVjodCpd7W6ctv9h2CNptxIqeU1Mt
iRu0UmxsDM+7FtteSmGI64ghTVNLN2gRMuef3vs+MvSek36C/4mARJdVluEovFYF
QDah18i+Tr+zsTa7LFvxrhr+qZVeOcMrb0YjYCyxWL55XHWThUm8DYJZn3i7Xy1y
jC0yFwvTfUnHzL98FCIDM8wcTpwEMA8uRqKFtN5XvRkMQ5FAHAiNoCy59sMydT76
YAFhpOJafKtdVoeEoNBlJj3vtoMIe7huv2xm+M0bH5WWYuRsar4mfFQIoolJEeyd
7UnZXxm9BKxCxwiz4glkc1NIZ8Hc3msIo370KFAR2mThrKlbpKamEuWK2LojAalB
cYv3VXBA8GSKhyz2PVs70i9kFtlqQL1TThgpmWt1gmzKTDq3RPIpfDktasDp9O+G
RV0KUwpoacuzuwuzBOP9mwYbtnbI7IVm5PrYeFYa+D3S9DJ+/7qrwSDL5XP6Eqq4
8TbCOobsYGX01FFOLp/dRfCOtpCCm5sSSualvqGkTGoLsXCq0CuKQ/mWy5fAXL36
/TkAJER+UWjZHy+IVEGLCeHjCWUXYakyXDqKyJFQQ/3hDsaWGz9yz0+gIBr+bdzV
5xiKnVSlRpGABFmC33UYNQV+fzu7JkmAmpy3ELFU3pb7fqSn4hHdwVNmtjkv2/JL
B5MAoJuFQIkAosNzhj7vjKPtB8oIdhAz67A86bK++yP/+saIgfE8m/mY404Plew3
RnTYqt5YovKpdZs9kQU+Zx3YTznUiEpBcfeLci6L1ArcJlLCzKTtnmWDAKFKZ0cF
XqF0mxZjjmZ9xDQEl/Xyr060zx1KTq/CEBNS2mCwE8Dvg1kPoKVdOqr3dQ+3ya2V
PACE3XcuZJ1V/Z9K6UABpuT4++4A7b3SILDcNt6njunJKbG4M/8QWIubpTu5AXL+
gXoTDnt1OdXz3xfqqO0UlG0ACZNuC/7jkUHhzcXZFjCxhip7wWgCDoTycHPd7r+R
qUWHSRMSVWCmeur8vwlyJpo7Fv+w5UQZ+plVdFFOC0kydD2pXi1ImGi4m6RSOiCD
+UN2gALBRC7eJMlSpN2REFnCDK5Dgm9jhxVWsYOVD8p17BlrvJ/LWjMam/oKvxa0
knAbQDr2AZRCYIQCLWvGpN6gPLTTn0T4kDGPm2Vvo/xXV8e/G8/K9fEfEKnrCid8
rRxJkxpPCBUC+c6Sqgq7LKJ576SXEdirmiMj9Kt4F75WNzFZ0gpsXoaFF6vt3Mpx
w4cz+YKesdBqvAjm5QkaT0p1wsSpP9I610vBb3DK+vPsT1RyMUaAXfsmQ2icV03+
wIew8OPfGvfmu16tAh1mb/bMGU8xx/r94cOCcrOmmo3akxNRtpwlHAiYxuR2kEuN
qYw9CPxjZH7fnzJ9BRs39SLhhzY8DRRP/baF8LPGelIccfGgpmA1s7uXOLfXG4Cf
5IALDge9aytXuCxroVN+9n2JGDDX4z+EioONu0Vj2d4VgwBjhiY5ZAREqP9o+ixx
eisaAaB447qy91jUc5iQr9DYXi0TWU2PEapLHsti3njhi/8/ge+oWfFTHBv8P3HK
zDqlf6tWFtdF2aA6EW63eiloRQSvyHYjElqu9cKFVqF4vW5YQujxBuqqiu5eIYYa
aNZYqeJWJcawz7w/H8GntAhZQNfm0mpRX9r6brtZ+kZvSEndlkN2o4pXdSTVwKpo
QWBpdU+DbZ+e6nFQCVVOrmTvduW9E2GtNgrlCj0QHLRlcXdgOzlKDER38y1cCZhJ
aasAV6eAXOnDWi7FGhw6b4HK4TcWywNlfACaMNWEVgf305r9YH2M2XnFsbI1eXkU
f7SckJD87Mq51F6ElCKS1lqtpdpCoJHNm4Uc+U2kzWr/XIB9jW2ACLGNPecZgQDR
+E23BfbGOQtSA0p0AVQ4mCrs4KAWaJCEg80J0D8R1rlRCrh7uQ6zG7hghUGYoHWv
iIB0+BHFvFsvgZto2SuWCTcufzlbrSOecQYWIrpy6Q86mzEORrI5kCFwMzgacgm1
jY1jD7sZEJU/6jiYDZymYCF41VfgFa6XSzX+GuWHULNCCHZKbxlwTsvE1ph7Xbiy
btVtTwi0EubiMiSQc+esdtQk2pHTUBqmuMd659gqfigo2Yc83QifECVJ23UOAlhl
tC/0WdgHDO/eRVragrNuoHNbl75rAjhBxThpeWeKbhZzzw4/0uBbKXV6SHuoy1lc
adNR1ChchtRoAwg4YD2nUl15GMyx/HJwbAhrJ9jbp/G0xbsmiyfy0qS59LZCHfiz
PUs7xFII/r84jGNhOV8tZR8yUPsK3lOfSVKmKc+EY0T5M9c+Rf1dp220KBawpv86
LH+M9MVZl9YEp5795LXg9RQLi6K1hLc9nETV1U8+0M/iLEDQN+g2FKei3/zFjxMV
nf6VcPG5Npmmgv+nEDjIq6AD+5Z2di8vQzGMp9jOpm2TlorYuQ2oydo64pYq4Bm2
yayIJ3rGMWFjq1iGofxpAqbmfOLJo4hn6upvTzmLV8XxWJaebucFQfARLeS0bTPS
xI2DHqBm62ZJuvBJ+kQ3u8AdScXZUSFDqnUROQglpLnVPZaa9n6c3kyJN3VSyBUn
+4Hg8l4J5EKf4O125yBHiIwyM05s7n3QZ2oY75xZp6NpqQ8wSCLPnVQlnZKOTOq9
6Xyi0i61SYUnDHyAkGh5MM4HItpJEqAsbTFx8LOS5SEIU4S68kX5KmwBxJPkl+gq
oYbfRrP5B1ze2Y2uxUPi46jHApgSo7pA6vKBkO/fdaGKxt6HoIVQwLteTGo9fkt/
jm2p8PvysnHg6r38FI7q4koRFXilq4pfZvdwVptDCTE2xzTetG/a94ea4GuO1ZR6
aih+beoK/ZRd4fTODzoOkmjYOhU/aXw+Q1bOcpmvMgs1eFlmAB0IkOmNJkS5gXuU
bMWfwbOFxNR5jtT4/fREv7Z2xU2rOpAHNQbwFQRGop5S9zjsn7tRfeJv74rtNP56
VX6l8+VDLokoSAl+kJBYpfGZS1tmflPM3hgI/gX0jmPPtQ9EQPz8nFg16L1jK92H
b7EyNpYr9EgO4sPx3OkrNmNfH41H/8bIYo1NXk22xKYubQb7J1Tio9Gt606Qgfod
kcVYaerM65BCYblNvfDG7JU7y8xatZ4NVLLaXrBeUlKkhMvslD5qXaeNBMA/EX4N
X4kv1Veb8XB4l+6UOzBH942sTFjd8AyOiUjkh+u1DF7D8JUUqUGtREdMTSG+XhHp
CrUKEsVjL9uMwB3N6o54GFi+ABnxFr5Ntx5yA1NbgPbxzb+RmkD7Mv8qsrCr+Fe4
sR1op3tILmRZuBCvIYBmPvhIsAQ+LE8cM0OkKhawfF2lK6lwRw1zulO2hNpgBI/a
t5RBGWoHE6kdSF1X/noyClQDavCK4RADxbodF9vRSwgbmkaPBlUuLwfJ6VKSI4oZ
f2A0hEeMi+dHz00ieiykKu6mEWFu0st+NC1BXFMZOyv9p0V0I2qitJ7zygYhJB+c
IQG9VEmmraTuvbaBGhBGcithz7xvMfqvdBMMVrtdrE0Ebk7iSZsJy6wuBOPE5rz9
EAzoyR1QENE0o7DahQqR7hPot/B8P6d3G/3wzof/1aNQvalpz4bOtMZMNTokBanb
T2au2WTE0Fcguqi9vdWqgmQC3YaiA7lP7ha7useYwAt40L4fxNGLOigVCRib6FsH
yFswIi12f5I3bKS08wF/Fw2ziKN2UpF/2VnyOQf2YdXmgwh3Z6Q3ftqJSdw1omKY
XQACkjrCxlCAnDPGkmfQtrMjaz6L+TY4QmPiw1EzwBd/EvHXjfEJmFJfaCP1UIxK
vaVv51VM0EixHvIxKwDwpmQqTgC8vIy/QD7d+lovujABbS3RIC9S5cNRv2IIvRzr
nx5DpZwK2F5w9eEnsuZ8Lf69h+KKbqGl2mka2OKcO/02v/v4Sd+irwSkLH3MlGXW
YjHXZetfLTBehc3RO+GrerpEg0arwa0Rqzc6KQzwZegiDPf+bmuNmS7iZEEVe+wL
05qLU7recBQyNCACkb1/x6yA5cfH23hYXtVWlsX2kmbjhamKxdzYyaIWqwXggtSX
8ehxnvxACGf5CxLgLviVOx3zhoIc9fvu0/d7KXQyw9OxCmX+ZMlcPfSfi1i/Pph9
GV82K0LU7fwjjb5qDJ7Dxb62IHAuw3l/uyPnLYKrwd/RPEPReMnoFmf+VG8HBwb8
2Wv7iD/W+b51o/aRW6RkxXmMADTy+A56IvYWSLnR2OgocFwudUmbTcu7j5Y/7+Kj
KE8FkL0QnGNu9Lm5q+tEoj0EXsicAtrhKLCq/3j55IdEXNtcW/ySZCRzN2LVk9mT
w/iE4dPHn8HQ9TrN3tlQOBaWn1j8ewkbjjeY1aIyQS+wNoBsWyL6hPHc6wysdhP/
S/CbnSuxb23cqcalaGzb9cJEYin5OmQ60o3LWbgdHk2yCbYu0GIzW8g86epYlkgT
AuLIqwkn/RX7f+lmCjGMpW1T/QS/+u7dnD565xRxpbWK+fbumvJDBftO6aZP/0N1
P4fmsXl5nXmuOoA352Ku7eMry9dQL5q26eACuR+ylCIcpGLl0bjusQpqGZ+faYPc
KNg1y2MtuC0lVZs600o51zVPgrpDKaLb2YFSbvKUiq8Up8Bcic73/Hyv6UTMG2Rw
BDT/BiI/VBmq2u4MpipS4WmGPDysBlzuXVQ3mby2sqI7rOAGJwwAfh5Ww0PsUJY9
pkY6aRyiS1oAoJMJvTQ154OghY1fQIZheqaWqF3IYA/c5UFma2RmlJYnWMCsE2TJ
wWZJPCxsrHLtbGApmVHJB3625BreoR9VQO2iK22Tj6FL2b3Xjx4TWDi88BAU8mHG
ImOLqDCtXOHUueddqmAgGXG6tNcuM4xSRJzeTvMOTewzc916o6F9DQe2NNbOLIgf
FgwhFXUZOYaqSFVCpxb2h3Dc+bGz+jz7gq1HWrQ4aRQSLobIlGLuul/rpHo4Xsit
qxl2LOx6wZ2iilqW6XIrbdMvWwXCloF6Ufh26yxzWfgM4kx3QyymlVGPdLDgP66e
FpKQFh6lvpic/nb/bkcuCkT2Yb/feQxlCv2bJAm7nacDlf3tChZdnTmVcY0q+3Ha
ZIZuXH+OUT3lYmhSkDsTGWFEDGlUhlXb+t4HmnTkMwItRu/H9cGWSEoGEGzCHKMw
SH6LAzuiZA1iFaeIO4E8VuEPgFveR2XoEmu4h3IsZWQru/kFjvgzER/qiSLOQ/cA
mmdgr+nATYxgcV1I4c4kL59I/pvqvTunhh5T2lasZ+Th0o1ImmY+LAQ/v9bjFIVS
FVu4Z3ZnyjqsEKI3cOG4aF2ET5fGmEEFsBSVmQTJ9JwxTTqHpCSJT/zqcf6FisU8
zOxz+mGVRJvq68njAEPDx/YrB0FKvqSDYDVe538dUzC76z6BrPcbmOTXB+rpemNw
lTduOyLNhnIxst/sQkNUV+wOc/b2I3olAObtJkdy2cyQP+NdY55laUvV+ktVUpys
xvrspui5M3goVx3B4oTM6+yiFn4e0h2VNp6pXqp1KOuK1OQepEC1zTbDEQJHfJjI
iIsD6VzP99bu8F0mH3/zwdOjd25CP3i8w4Qr348uhSzNQH3rmK7lv2NbhzJb2Oh5
W8QtJFzynEfoKTcilZ+y8tbmHpcQQstQ5Blhyv4OJr7ipOz4Jv6TmO6v6d2hyErm
64JS204MUHCMv9l+VdhndFaBrZweQQNsikMUCl5dNnW9jdeT4qDN62kwKSZwi9uh
GH84AYXcoshJdXW9WAs8BA9/fWBGhDLuSmC6Pw4VwGdG2QP7KI+nVwMz57nidXTL
hklzn8mDmug/V4rCSzk/XwajaSPigz5Ryn8V3f1M0LhBOIi/YfGrzl36fP1FKhV4
XsxbqvdhwvXankHCf6Uz+xoGX+Xxd/WQr7OMabAxC7TltkMa5U+7yQTHj2XwjmqK
tYcqSgTusNdu6LfOyP/UFHA2sAt9aU7384241dmO0+Dz8BO3Wmbo5HKb2UvWskkm
8EFLkbP/hmI5AF/NK2LVak3w235WAMYLA+jNBPbZXhMljT8LVD8VwDPS51okSWCA
9OPg+UkNXjds157dfa8l2cP0sFabwX9L+MCq78UmzPsxHo44vMKTkRISkVa40Y2F
g2IkJ5rES4es4qRYXB3Xt3imzPZlzF3XQd+WkDK3u6hZ07gDn+yGNfXtWW2egAHp
jEFi+sAoTq4C3gsVR8DrywOibWb8PYR6o4sxG9GyVsf8cmAPp3DYE2pfH4RiIh6k
eX8q2fjkEOCs9HOCJ18TCliXh4t6J+otA9O1C9SrBYuZFt2fcHJNquK7jLZy55mT
uOmst2Lm1+uUe5Tkp6IvvM4jhpCQPPW69OFspnJcJqz6NZ5fa72SaPjzIcHewCKd
14UNgNBhM3aI2XgIS0z4RKmSHdDVNB2ijuoK3Bq6sNvIbg/1ze0+9BwXFS/EXuUa
zNT2QewwyrBoKvOiv+ensKR5ry58ERf2DxFVkeNd3BOqycZXk1IFdVScdWkLg0CS
SrI/Xpum6bKYgji7rMHR2ifc1jtZ+WmGMi8iOjMKq+hS+UmKu26yO8KsqEAH7nRS
9vCykmcwnxhWajDajIA0G6o2CMBSL50wpG8rDw2dEmuDdC2JlU0fhDhlyzU3WLhQ
d0TXzQi9PHusVbU2iVqFRBYFWjW7DvwYeEnBla+XS07Z3iEWg6qDZiCFSY5xyK4M
sRhmm1ZYGA6laYfR9/ITSIi8zY2hJjNV1NI0dO23SCMJbVxtANbUekUcUQ+dd87+
qcMH7IHjxRAus5cxityobpJVEJiuyKwXOJb/uxyf9iYHFKFjfo9esnZnn24ODPWc
MM6mNRGGFQfOYJYXVJXBhfOAwB5RWkObCAIx0tzb4w/05hNytdJE9NK/Y8wN9wGu
bnoXWPM/kMek6EXtq4fG1AyhjA973C9ZRqtHqCi+SAOLWPUclZuWka6ePWeqds3j
b1AAtyT/zX/HDyJNn2kF2VOm1qocOE88r2Bme/439c6u9Hfb3hi2MwhYhfItahZc
HA/6vfXAYobK2SJ2zfq8oV3DHlwUUlZeyFSlfJHeExaxH0in/Wvm6ay3Q6329Uv8
a0easoySPcHDFKQ5NVhPO5gF2RlLnn/FiN2MYDR1WLVmW+HPZxhQzQYilDIyrnWh
jSVczzhJoJrRxl+VnvYAjdrbHO4uaxwhQQWV5lBFf0FuXNNgf8oxZZIN8I1bVGPg
s+3is1axG0BRq6MilkMVlMeDiszpWAd5Vtx8TS4eWnNBCCe1ilbTarj16d2H1o52
X5jBHBFcIzqyoQI8jfe4FbynElDZNZvL6KMbDy4rH0Lkp1rs3Y7FTydt63bYdTy6
DDGc90OSKZXODTbNxeWqLiHMmW8jfDtLVZtks0m/Vt5EIHPJo3LgbcXl69sqL5TG
RbOE9U6YW8eR2mWaLtw3MHnOjKmRSoFBCI8CTjkn2CmK0sJRSZX/6lj5KjshDjZB
iScfTN5aOljx+3mPtKU6YI3oozC/tC++11Q5PUSZvi+2QMpQ9AbYV3wPFg3/zrq9
CKiXxSPVbQG9sGY99z7TYrjhwW4+PU/9k4sVuxWJeF1mgUMuUXchd8j1LR1uleR0
dYhebzBpYh9Dzwv1R+CmImwnr26BbTmAP4EbXwt2OJzUFIskX1RnucW02vti9AyX
twXGxFFOclmreavdXXFIdspjUmtBNYAD1cMKIMRNvw0sBnORLaEB/tON1RiC29h5
5BcMYv5KeQ0MGRInXvrIPrMuT7STCldHJz9qF6fd2otbUQNdqickojRDNhaMXJCJ
2l0ZFTq6w9KN+V5s7VNG3RO6mfVhz5sYkQ4qdWOVIBnAVaXabBe1uPZl8pig0Mug
csEdPWfdQMpoLLOOHiotzZmkLHfoo6ICDE4cYirZd1dTGJHCe5U4PhgnI+WB1PMA
1QAS5UbYeM11Ky2gZWs62x0dIWk5pbXmWCIlkd1762at5KTK+jdxpygApWJ8kmwg
Wu8knvsUx6oxWIhcHYtrRzVcKfcBlCDwPblojlEtK27T/W43cHFmQ8o6dtMHomPA
Vgiapk1Quu8YRFE1dppMTGXsr+ZwzNDqbhnZ7QTeuwcsEN0ei1RPjjJjBmijxCC+
kd0EiEY5aCSaEOoZi44TCO1DrNeTl/Ud474pBZ04ljbK6l6RGfUVDfTC8Af38C94
dMLp0k18nijwOI3RRJJFfpMljhoa4ZdgzGRNw03Bs5l7SRJjQYj6fvKavpUdfjhW
9Tu4SDAk9fVo9zbCUndQbQxm+jeeESkJbyPxhJ8bw0FVxBsAn5ozSGf4H+5QwtV8
9vwGknkEEF9ZjvFL6TuE31tTsUrHtmpJXJ0A/T2zgdfYbeoym0oWdJ5EfIMJxktg
xVk+otxresFdMlOe4QMjdbNdHVSziQZjRug1GDfVS+EmnNlSberbaKDKFtr2/WxI
ToHg99loamJqyL9sQ6GpofgKa62vGv0wK1TKQsdOekfc4uQhw8zHoDGXdLVDe+eE
HSkihoJxDUkRcv53ZxeyP2Df3thq6lrt13wkx6KEbta+NXFjhgRlEniAl32Ymoe7
yCkaCbU0TcJgkk3m5PmpgvQqnCik6HGliXwJyQR7qW3ViGV8qiYfqCW3SZEXxfrz
uMIas1MP06Q7+KE/S/kTRYJ2qkuzx4ZR2INqibuYdd869B3qHYUoxg0r9iTk6qcg
WUjdr5ib8WkCfL7UYuDkwBAHY5l20XZBSkd5TTnQRdUYJ9AT7vGAzbOsiI/zlcQt
oFHUJmMV6go0QUxCvv6rMN0oZ1vTTrawYptOVmDO8H3vnMeM66BP1XnBIQKBPIVZ
pIYMYBef4tbmcUZOUcdLFTpTazdAX10meg2GpV8oy423Ai3Pp9uSc/MvbaV3/r5I
DMbXw3EXsK9U9Tq5jLiNAlLyhTLgLzQ3Mqo48JKRSFug+DAmLUnFwPmYTZnMD2Wq
gNcrdbbkAduBxAIIEF3jzJwxKJxgqba+5/M+HZx2OAYODcV/sgZjq20BzaehR1wS
BO7nANMjADZPYl1DrRwsbUgqFTo6CydF5SE8buVjwxro4yuIuNqy7O0jTvdUxIYp
znUVgtelQiPd5l5OHcfeGLHzkJQyxYpqNBl/iPIDatIvoWunRnLghqqekZLlFDFv
IRurOE8+YTWPdzUTh7oPF03CBr+AfbQQBABNmwdKP8og+8HoLz/t4fvVEssrQmmR
L2DA30LD7k+7duYd0aXH0wO78m7uOz+LKzSflQmZYQPif7Bxvsgd8yGl/vUDXPL5
kET1P5z8MX0bbZA8J0sHDFCK+zdQjPMGYpWGY69PSbNepjOgOJQRQEuaHs9STXgb
NtaSPog0g1yn3B8zAfSHmVF5iZ1AWaaXj6tEHmZnq61Jn9OwCwqV4M5AFqjEkM4t
KEgmeaMg1ijwTzxsBqlysfmMsUgMGO7ATT4UXN4obZvYhkU3M8DGX3WEEDO0ml/u
JrnnxzeCHOZ1ICiLaR0ij7WsdNtchfiD95WmQpKCfZCF8FCElbdzPlbcnGxZmDdg
f5Xs3HYLw/hh4bgI4Gd/DmgRHWljzYmhy3cQ+L9d1emiOcGZM6cL+xiUuYnnknbs
7eltOfo2B4C57fVy5eUTLUsPWPMcU88kKD/b1/AoCxyAPW2A9za2DK+l0m4VMQaa
qJ9jo+kl73Gombil49clbOm3XmjNRoQ6ljVRyKG5E8U7eWYdCBNEja0LHMmcYKFt
Ch/13wipHpzI4X6MNv3l/hHgRUmLaKrEEnI6X8scQUbjEAEGUCLNkWlbeGYLcs3G
BVu2tKaL01uPXdBVVNrGkRiZPrcjp0aWf24q9xUSgfZ+iheEb7KntszNjIndGFCp
AVssHRAa+RT+2Cm+5w5M5ZLeIeoZ/yWONjCpmbTn4zX+jU08iNIiv/Nz/8/YS0Mp
/DtBwz+MZ0d29WAyxEMn7c6EVSe92jhz5bhSsb1KdbHjeWStAEYY5rc9tK02Sxjp
t33lP8Kzr/6JTSTls77p3DAfSQEEq/MAGtikRZ4gIi+Swrkw4NTL9boze8CwfhzE
vP0JtumUhsH35Fp8EsBHDwCwMYwuZo48yNMJplXijJUzMfxlo15nV3eWKW+XGMIX
AvIYLvfkZEdG6zW7cwctVatZRzFDoYrts/gw0AOKFOG1M3fis4I4r2Quedw0S38Z
4d6snNqCwHQkzU17SqMaaJumFpWQ4PLqZfF9L5zbFXQ3ED5rIv97D9Mf0NSplFqd
jIMThIIzVLZ0Kf0LcVW16aX5KzNwldu0MOrnVEftuEn2MrVUny1Xr0ekhwP4mAl7
TBZQAB4IpScfuDDCuU1axaI/OK1ePnwKaos/hpwZAPV6cNnKdNPYbeC1aULRKqcb
VYh/hlwBkgJOb9x4M4GA1mDOWu2FZLlJ6VK27dGfWHSNVHH+yF9rsXWSmKZoHPsD
MLl2M4WmzBy1YAshhxWKCw+wEgT/bHly9Eu+xQkOnXEieCBgoByhR62g1zKKGFFi
LkSO/qHZCSCb2yn5XzFPf1psE6Wtt0IFRScjE0IyW8cMjeQxcrWo0R9H1YMV48m9
KgIe0afjQRXV2j3Lq4SPWQ+NfLVY93EIL+LCGFZuyswfOD9i8lQKCuQKH4AXg4uR
WQZLzxIkm5g9dSHAf5GzqqqwRLtA3Vmuk7eLfNynQhMCL3Qdh5VWjn8jy2M1fWsS
lF1enl0+QZlVoxGI5a+DFIu1AcB+ZH1c3xyrjk51YKU0RhjZKTx2iwXwUjBUalft
CfwUMGgWPJYnP8Omw8DLJfgwI/EfJZyDLoHBr+wOT6uLXNnl/HkRdjJh/rRdfjXR
0RfZRORzlWwUtPZhZUrXMrIFrHpMo9MMe0C6ANTchp96/rSd7A2KSq1UBoHFNnyR
D0ft2wlbyvVG+GcXQ7asrz7pgvDE3WHAiaAYeRlfZDiZGQ34ucCGNJ7XaP5WtU3Y
+cW3mtZpywT5sxIvCmCISH4QFi4JNuFACICaYzkIw2W+LLd6sT1VgqmQbhySlRUy
XwYxYk/EjivliDZVntEyCArd1VlSBNJRDVKLhCavixJ0fQHgg/nO/6vso6Q88bjc
FLzCL9aW73xgXHW4bBK9/hEBf6cnQhxzK5dLm/8og5VqAZPBKhXbXh8TTBnNCkx+
8LY2Tg5/Yt8S38YPYQlGHckQJijGo4UNDhZEfrdk/xy+fdaTtbPvKE4yV42xJkyh
Ui1zOPE1tN/DBIWC1Fu5MWnVvmhsr9YwRN+V0aStKGdHQGYMp4BVHXMsd6Rlz0g0
0pdS+8+ec8cylJQWUM4O/qmG4DDBIjadVxHF4SNYuH7BWqtNLbpS61HHwv+H8wJ2
miZZqX3yBsSZj4gs6U6bh4simeNJ4YRvMpEUr/k8DpY8edQKf1Lt3mbe+S/u+Tr+
Y0a3MYtXwZZcSkk3nRaEq/3zJ6LmGKGfkwp2oI3ZRRg9yjZ762p2rev5HDE6QYAx
FUy7t9mfLf+xFjDmrsDZrWOWrg5VLk3VS1JlAXx+UnEa9aDR67wVDhBK8tw9L6UG
Zwi8Kv/rvQo7EzEd4c51YJHJQLb3DNvcz/tdWHwql6He8XeRi/2rV1YEf5DuxdOP
UusKBYNo3J7sQ2hwokTwopyg4R3+7wDOLNBCNzgABiVQrnUr05Rr372lJ0jZd51N
69P8wIK1pOE1xg+GPOHEXba0PHhM5wroeSbkt/y6UMfk175vQhryWu0HoilQMC3y
YOqPNCO2HHpa8Im2t282eapJsP6oHftpMxQZLVMq36yp4tM6NFJwlq/8uQu83PIV
LYXa4svaawq4JpwjxPp7BCtOPtHelXzh28ZGjmks/WEK18hCFC2vVXxzVpAt9I7q
2tOwd+7y86w8OPt0UEQGAqXENFDJGGO/DWstqNzCHIj0TQFE5dO8fmqWyvK4M7y1
M1qy3+ua8QiVFhsWAUBkd4YRXEVOdAtt//W4i4/iQ8IPFUAkKtThfVqD1uhKfDgY
KKgtzne9aYy9sm8E7Zg/hTWbKjTj6uKLGEsjiup4OilKxGng0Y1RZc0nIg/w2t4s
sOrpoSv9BpumQ8nIpDt+aca5tJYgpQ4MlxylPgZ4mbprUt8bMn8RHeaiIZ7u7jgS
d40HEDfiZhaOUvj/rMOT4s8mbZ9WviD4bbQL2Mj3xWVvrQkdRr9FexdC3jXlGF3/
vz1miwY3pR7GIkkS9Q31ZA7nmo49VRmCdhLfqnEBGSFA7R4/S41EOW3OQBtMPKpz
4hzYBwMKZVvt6txnnKWDnwgxT1Mvz/Zza5PbIdekXlNzOAy3SLrIR4f8ozix/YRz
BRfcNvLqRJTlEDSEJR9iPAQmwSbZN+JUUFLwMuslCyIi9txwEgjOAE1HLzquD9oZ
mPafLkztYwPsaSX8WK8jtJ2LZDztSLnTiLbt/bHdG6Fv8zR5SPLF0Llt5tl4rb2C
Zu+vuHKVBkg47Ayv5ljy1HAVzYh8Bfa3dFcvSJv+F8eOH2eYAK42RleDHgze3xzX
OvWUaHCNjEBxvnfH9jHXXS1RnTMmbVSe0qX5oKf9HEkfpXIqy7yB2KPqsM/ZGksj
X/vhyZo+nPUIcZ5WwNr0xUMpnT4muKpV81IA0pspeYHogTGGFVOlhhRPHr2NEp3c
CKx06mcH1VpxiABl0y0ILulz5FMLMa+D0EnGcDEOfNDrLBvoh+EWriao1alV20Kf
ZolaFAYJCtB6Aq9lQ3cPrkPE8SfqodJ5JvS3uzcXkbXyHwWolV5fZ0tAensBbZgL
2h+4u0pXNZ+LbK96mO1klF9sShQcDcu6bs4SqDdlvTTo4QqDDu4DuUfPyk3Txq9N
7X2VsWCyCsPo1Vp87IYcaw/Cv+KjbYv2WfWP80H+h/rG5AzntrOnKrO2JDEtWz0/
zDuWp3WNKmYhvPmY1+JW9AyMdxr+reFMg9wbPnxQGkEUs2wT4SpRXx0Sijpvt2dj
+4nzqBEiZwURIiuV1nY3dZJUPlxbePturbYZqAjBs5gYECYqCxWYJg6Qi8a7PfNi
4GRYYDq1Or50JeELLJPPWdYUuG/rhAgiUq1JoM6h6WRxtHR11UF6pwuIWj/D42C9
zoPBL9iJmIdGE4OpV7gBBsaPv9PxRXxK5nZ1dacQUj+HQ97qe8lORz2i/HqYk6YS
sK7SffGQnpuZQ/ZxpfosjZ9qpES6nfOdlvJHoVSUKMzdokMbHsf8vsefuXxKIIe3
iQdQCm2bMAzPYniScIjat+Ex31qAdp4+mCeJmWN79ppd4qwY6YSW0dJKjS2VsWNs
4+R2VkfLrxmHPumCEDtFWkKjQiYsRUW+38LXyo4W2sx3n0ZkuE6ORjKgJlfQLalZ
Nlt3e29JUr+t1CcEID6WvD1Qp5N+OOgZWkNlPmpQE5mJjGN5YXQ//kjoOkIlknYd
A3PRSZ5rK40H/zETwByZoXYFj6hj9Abz9kZgdWMIQsHUHTbOJcglwt31hzYDmA42
2gKRh8u2Zo6e57EpKx/BbMvKyV+rfS280nSJ4ADaWm5Vs6Wbl7Hm2bY7rvpWOjMw
Xp2V5c4JTrdv8G2NUldXTN7YIPgYqFjJDWeTwg3lHY7oL/xGIXHGkGp0IqTRwKUo
QfvW8kLQe7rARfJW7DVH8LdEiPhx8bRdflq33rsWMKi996oG3UPbNM4L10L0wQC8
tchZZSOhP7Oz7bmObwi2/VF4skt47aOVD+iDLL6loh0YlN51vQMPmkGSQHKYLjBf
GYg7pOCEHamCBbI296l09vEsfhE7Kk69ZmHdHO2vGnAV4W+ZqhlavFKDM9vMpmRf
Ge7vteOIHxfUdSELxEsiTv5eboPdj+i50y5uh5pMFVD17YC5uv+pbJ7Jl0TUEQid
FCjxMPBAO5aqZfRAzS1qNfBUde4ITR9Rr5flRDaYriOSucGeR0NYYTBMzlo2PZd3
T1DGPuCO2vdc8Sk+VrUP3e0woTJYdOdXC/DFRSFis2KJ0Pj0HKzFcwtxU6N2Q53Z
irtBhubxpeYE259sHxff+mJEh5+5F/fdF2DShBV1IFe8KYW8JZelHyO9k6Ad4tDD
QRXvU+8p1/2sZdQbQBPu+pd69Xka14gmIZsEZhMQuA0UeMPdQFFiDvKIGwRD2Gmz
WhS4igDq+1xInkjtp7Jgm8U4FsfEMAdUzApBm/7WYqE4LlvdnY3MsYydGGhT/tTC
UMkykSh1fkf/FwnSyV5k0RSCLi+6I2q8/HnQ/i+JYEyMNNcxO4xTkLVyOuc9O1/j
gQJvR0m3cqKKFWxkHXU6z+FW+KLw0auKN44xsht3EwBB3rwqp6hcW1wDOdsSQhch
zDXXKOpabTG5df5qQ5iP9wG88fB1jyDMhCqXmG8jbauFD6FallCtTxeExqvxMl++
NKxzvox0C7nWDwqI9bLHrqh5rO9WOdcdVNNhv5yUq8/5wvotP0Hxmg0WPKRK4n2R
zjvG+hlhkLfaHNnW6wyX0uUNynw2FtqoRG86zALm4inLgYorI9YsolEJUo5cqFD+
2R3elGUI97Fv/knUsuc9gsqNBoQ5iJX9d1X3ZzxT3YwVd8d/utEGUOxMROWFwvi1
t42RQ6fC9l50GT2ZvTWYWO0sDMt0kV+YM4R5z2UM7aNJVWdCt38IdEe1Xm/qwfrs
6q+M3IpvkMJj2Z3GbRHEE5pNghkKs1GREco1c7+8808TvNsI1jQGuym4z+cSjsDb
gGdAQsIwQPBI54CuJ4KG0rwkGKQJ0HrHcoG0qxyvhgHfQ9Md+zLUQM6WEDGJH1p0
4YPaauiwUA7pVxR6LkMo0am30D1Yo/HAOYo4lftPd0q3aWMta2yJ0M4P+t61k5T5
ThYKHJcWNVm+i9GJDfc0SGFGQUhhj2dLeZh8095sVs8Vu2dIPYhHc+bYZ8MaetMC
q2JEGP4RfWVYUdM0tpMBMG8ZTrXghmA9yq8OFaLbkeQGDOFZXbEFPulRMAcC8V3c
RfHRA4K9MgN32ChSec5DxrcIlS9TwHyo0Rzir/5XlO5iUyhNyVUi8F+jw5GyIHMC
dH0fAgr9cm7aFCHT6AvUw4aCEJD8BVa59xt5XaNNTuzq7Jpz7ONiRAykejnzR62D
sLK2gntORz7oGI+3Yqacz7MzLxbSAfZBnERzKN0JSyrzVoLbQJDwXTJdpd1z12e2
EDL4foN/RwcZrP+NrNYiAmssq5lpkc/ouNodTSTwoIFMZPQw5w1VUf8B52k05OEE
6q6Ra92pBwjoqtRGtLMojQPlNZsvtYNjyOILV1axZbwlYICNoSQONHXrYZ5FhhAd
Y0XZy46cw79S2W21CL5yKhCmail8YGOCJMiu/NaHmTqa6bVzdP8bckaQ2ocTjeCi
XwNpBzTkdzLjTy3TQzCfNJf16WAQEuyZ5BVHFdrVPRFzz1Tk1eHCclrJpTJ0ITMR
jIaP5M5zJ5rFvSZkx5w9cq5r+uqTYRf5FPYl5xn5TFQOJ6qyvsglPs7chj0W4Jtc
TZ4bYJgveWcMvxN8pu+KCuhg+NVgSzu+8vzHnNmHD2iV9YIOq7Mj6mN0KL8+qLEb
njZezfFFKeuYBeYx9ZsanK/WS7Za22/jA41RQ3MK0eDRa58zZ1hiFa6xoAzl+Nfk
3QkNY9FtJW/NhKZFu0xT7avnT797lxAHRCwFzEiGODVZIkSFgK3rLICeqH8ADUf+
FXmO0cnVoTvZl3xH48w4uv/1cd5h3xt+NUKuCv9AD3pqWJJKL0xO/kEOu40tly2P
K6sfpW9FB/H5Kk+elkkxik8WjDu8kzHQKeG7v//u1mOKAG234ndr+lEQcfLAJ1GI
s6zqCM0G4TkAmFNeKQjqVvxCFQ+OGItWXGB3ck2dad7hsUSbtk+2eOz0KxNnyY3J
g6/r6A4i30qVQpqHhdjXRZc58jXsW0sHct+tNo3tdEPUaYle4gnRAqs5QzZ9vQq3
4aRNYswMv3VV535P6s7cUIKOT6BC0sGl63Ow7+l12AQAbprraApuvk9ELVy85Pr4
0D8V9GjPNgHw65IyQM5XbSwmZ2qWAjE6yZbPA/6ycWFw+3N8o3wDXImDrverxz83
dkIz+ijsuJ8lVbBXsrHSS4zzMG+9PU4qqz9eSxu428RO7hfGakU0W1674yfsh9hW
4/J5xKnzRkJnqTfrABjTSDzGXm4qV538VOK0+6qDmSxE6S9D22zwAtuKDNX1hijS
G7OpJpk7pBsaYO5mFYEe7HYlDGXYYQ1fVkVYlBq0hUK81+YH89R34mDguYDI+yhw
rv0L4mC0GYVqFg0kDt4lysCqOgI99ce2MK3s6DX9GOuo47vZD1Rcm2j3Z8m9E+cN
2VKqvIq7uPDv+YJ2pG3r/rlQLvnDzxb4GDX26U7MiLyrccwuUI5UeNYJNZb/xwcM
dWuSf6B7IT1w4EcoEz7fBzjxzcJ9ZzxNdt5QyobKDNHCtGJ9ObdrEEuWp5nSoFOS
TIWkhnnLWdMu+/1cEvyReVxRA3XRQs3NnPy1qYGcV2QhyQ6J5FeyCLsi1inexcrL
XWAWaIG6NmT6g9CBlZYxgqtcvkQ64aOV2xYtrQ53VH7Y10Mu+4ZpCicI3QBzvWqR
M+rHhvQwy4R1IMc84ZltZCdpjnbQdYPk5Y8AbIZLOUUjnl8kxmmdC88RZ8GhEczO
Tp16F/KlP3+PQeftPsmxaLoxqezou2A3S5D4NlpkOZ4yVaomxpt1QttJpVmy+GUq
che7MkivjmTASymmFBZfoobaI3bKT6dLTG/Ujhh9Td0y5FQuptwHRYqyYGVX1kNW
beE8iJAmskqu98i4rCzj+s6NasLkCC0VJLCEnJJlBsZRRCYyMP5xrFfTuTnyQSlp
HIKUBiPsNP8orZdPsRZhAePWIy4bQ/1yFFHl10M+hLWuISDRa+CLapjsRGedp5dY
GcWh64eiSP4DkyneaE1LrzDg1Sr/FrqdBg7BhpgKuCfwS/P8NflBCr9p0WcVUGgh
TPltwIM1cTKFvaRTWTGzSzR7ulRleACrWlnxqw1KevAACJXbo+V4C1fOk71V3t8m
H5kNIUQdfAmCi4Vy7gwKpqzqGxrIdYydiLrolzM/1f+52XjxT/yd7d7boUvl6NN+
zvpdTI/agmXi+TFgOxmCCw7RPmmmnPXDt6ez5RzYIr5zVa49nrRk1PTH0UrVtLKh
OTtNSTPwftxuBKsESacyShsEABYzcApVCK5QJMGW9rpEd1BXS0AX916/E1Bvk5zm
hM1+E3IVXYr1vu594kM1HKw04uhJfPUArIt1duwikZ1QopEtriXHZ5PZ4FEUEiFB
UOSt9QI62Fs+JxikUAlFU2o/HNkb+9YvZoF0FQlbEOrXfXm1X3yBcC8PR29mTAx2
CfoeSMKz8pR425x++rtT0At1adzkNT092fAFl3nfzEj027LZxMaGUhgUGlE3g2PH
xdzqo26zMXW6xg65jLkuA7C48Qs0wfghJIETSu/rQLRXFxVSB6rGNJxxWYVlIr/0
4uhh0ho5M5xa9mQu9vWR4wlLe/qABLyfnrBoBgvzZvBSn+32Q+V1uddveQagZcXz
b6EiU4EMtkM8khpoepfJVkSNUlHfiyhYFlF2yZ+tpTQUHhHFd966CY3KetYyzjFc
Zze5dbLNRUn+RweVg/+wwYzIkzoCLN98487VNhhcBXKW1UT4LF9rqASjQqqJdN5a
xZv4rrZxGVzUf/leocXE63XA70vZYmujx0iEza/rQM8R/ivmZZlyNbF5QZB9HI6K
K/7h2jU4QGUiOzxgKvDHEn9cK2T5bTLONfAA4FiEP8PXaleNmmDTbORfmY1xDh7E
grMwxcBee3CEaELbPKfEg23YbL4wYl9hLsHCECVyyKZfN3gsDjKHnLkRmm/OMkRj
OUJLtpV6+j9sxJAbDsoe9RkuOxQjeVNeB+Xqpb6ePoyVX5iAW77Q/9zFqosKM0HK
lwyRg9yH38yJHIu/Pg5KuAtybAIW/Ix2ER6M/t/E8c53URB68CoVK85V3UJ5kOx/
CwnAPwExDbvf+me7WHRyAehJqIMMbYocudm6I0QMgPIU8e0P1cOsnGI9rRw87Z5q
0bWsJy5tcPjMp6oztpzU3wXkpXOlpjb1zgjmnMxF/VZlDI78B2abo+G+6WqmL8LU
8ABOG9H4QxSmJD8Vm4M/GXy9076dLp/GzRB49Y2OvC29GgaaCPBZEoFGK+G6PY3v
ZfmrBUREeXPMw2SJ6wm1bujGLifI7MzuJ/LnsP0x+p8yVIBhnNB/NoqgpBQLdtNn
z8+WND+IFKgWAzKbr5hwEhAtEaBlEMxeoToR/uyvODu+ROUeUmCP73A1+YmO3hwa
gYLx5r/kk6pbPJVd86eBFsYqzGDcz2NsBQ3c3FfdSCOiwOBBE+Pcg3aNskZEVsXa
V5HdAyHbOq4b1e7nWGfLFXfZeIHpFk2KQkiYjaV3VjzaoQLSmJ7RUNwGcULYn4RT
EWIGcA0sALwEGCEZFNxPCZTBUrbKO9CF5FtAYdJwVmJqAWALueCBWhNeu8GBd2RX
KdU9Oz3K46eOsHB0kmOOwFZq+Ve4jqCaXX2M5cE8jYZTt2jhgfNXhvca8W1fvJ/k
InoVktp1qN19u8CtfsCcFiDYaRAy66N86HYx5kjnl0GY8xP6WgijpSMWRMLJcgBY
Vxlpx/jYjCTxcnnQEKFfxIt8Y3mT12xRff+BXHb1VKIYa1cxTSKOw5CvfKa0+K0h
99PYXo/B12lWSWnmYiAkEZyLzGynS4oYUx1byrj9EC7TF4+uJrxxmfxt9WU1yQMB
wkZ/TBrDqQyMcc8pN1DvYd+LpqC1CbtyE77OUJkiRA5moDJ6Rg0dBh7iwnFHGlFE
6uZ0B5zUXabtgo9ozjxKqJu58SCNqilycNleX1r64AwLP8pWFmRXo6sns/9wsK/j
uB209zURlDEjTxVxs8yr1bMc1tY67SoqPo9/1ZS61BKhOXs/u5PwcV4d7UT5zGPH
IWMavujftkihfSwaejasEN65Me/6HxmhwWveJ8yK8Pt6nkEjHyq+pV0MgbegzFut
uMpHJ1jsecbFs9QKeRwQ31upAV2ItpGq1SNdAtRNLgiYyR8QPRGZF9xe8uoa6W7J
is/9Mh7SuYoOv/6xW1szYe25YoX4zZrqmCH6UI85TRja3NBr/T5w/uWEQeuTp2dQ
pv0ptXY74NQdjF0l3jshLIlt3DExRp0vqLRual3P5kb4+jdfSfSLZFXxeR8kVcBL
+VYSGOrReleusVQ/yBmHGs16RKRIn2AOb4C07F3Pre1rzDVdZFgZGJUoMLUQLxyO
YZ8cX/3KXUJk2DLGc8Fr7BYT1QQuuJamwbg/29RdAVNuEmESaqQDydoWsuaV1kW7
zVPKoVh/3xO2UFXrH1G14UQuIeC9x8d6gRTaN3JzvJn9rHqlIAY81GVmX1ICuV9k
QRa/Qj/GElcCqBaRuAmaRCiWxqt4NBI2wDWc685wPD31DzZ90aNqOtQijBDFQMqM
sWcveIOVZtlCOjlRmF5S5ISNZkZxXIq7KIAcRo7rBoMVmP0Lpzzwl7q7eFoR8xLv
qn3B7vxigpVsHI23WAW7GPyGOOcuLqOvDjMpfCaATftO8F5t/QNdh/3vflEF8RQM
t8naVQEb3cYLXU5FWMZ+E5D2g0JOn/HEjS66hASkLWVLMGIj22XiI82DFZzPXvQ8
fcH8UZBfPD5Gn0VG1lflRkvnSOQvmTg97lEftAt54Qf8V35RhZiqT1sdTqK+5Hz9
6eLL+hpX7P2DPIK2khnPJYYphFp+atgiO/FY9l3AynhUBHsTKfEz95n/+yUMmHJ+
ltXKobc5+EAe6XltJRyyWjvDTLFKAo9VVSiVn6PPL8gyWYN2P1wJ2xfSTc3RihHc
dz3O2xHsFSfa0voAhO1Z6C6f/ymBisWHCD+7c4ITVS4ikVwCIbap4UDKEOZMW0Um
zc4a8Gy7DOQLKiXcD5qFqtfb6byonotOAFzNMk9iAZLUocF79ob1HOQjolK/JfKT
wW1tQsJKlMeJul0oJshNDM1NNCdUPzLq0hN84psTKDQ6QqoeqIHa60o1FiApa9l0
cTxH3ML9LFX7yYsGgzN1eC9zlLbwy3rN3cd8uA32OTbhi2wh1j2Oh3QOk6dsdQJD
Wq6bTnZ//kl1mgqn0m1MWmOa+iEI3lWIuXZT15vcWJI6AIg/dPycEKI+uUL+IiNb
Tdkab1iNGygoOvMRZh0LAK/2hrnj8/gxbtuTeEb3KWmUZv+PZB7BXJPCoESdkXfD
09U8iCCBhheUfeOTYomprKIC7cpTo5KgK2RrtJ88s0/acAP9CGZunDIuEcVrIshI
qOwe+EdY09q4UQ7s1k4jQ2u3+wXaF+pf1LUjJn71XhUzd0VrO/X5qMfhFnIj/Ein
cKXCoJez2BY0LM3As1n00ZGQRiQezSLhFza8+2YPLybCejRC6pcX4CTCzmoBi0sq
Q1hF1r1cyB3IC/YleZkKmcS0AQqzeAr9AAi6VqXDTv2NqI/AADm2vhvmaDjC+kcg
5YjxeDnMZl3V15MW5nC9Jv5RK8YmO3/V9hvw+vl5zuNPI5jkadqOYCIL+yC5WnWz
OlwG9Og0FS8pd1lO/GTuPfrjbcOg21uiN6My/mOpG/ifnlr9ut3HNrvXX04kaLDs
wQ4MB+Zu9wvh9ji7mzlus0vWsFiXm78d33A3nzyjwm/EmLqURKUIwU54TlcWjZ7E
FjvZAQ1+Fh4KpoRpHJk3aXKWOW0Ke3+VwPYn9SXh1FHcW3GDkTx+tWQdfk/C6XPq
B4cJNRG29XtzDzuPn98vHffqyBZCDQdf90ilqCR194gRWu4hau12rLR3g4rCIAIe
0ZXblQInBt6LVovGxeDdQiaNndJNhKJfBbiFg9qVMQjq/Ubw3JH8iBREFOo8aYNW
tesEhjjYU2diEeraE3wC3vcF3k789Id+smfhpU59HY/kPaePLugfRaL9AwiVdemQ
Dmmm/kywLXlLMXgn0iWh5AHxs4sGXlTpkdMBu7TPrBnmqO67lo/+P2XipRgxV4g0
adYT4h0QoHdFZ3eEdsJmWnzeZW0XmW2KrfnWv/xZaX1R1ij7EQhFMhAJeYg9OTaE
3Fkd8y5hwROH5MTUXXwW3TZjteVEVoVMOdF1yHe/kYrFm8t6H3Sgjb5KaOomuT6N
IQqyRz9yqKeOiZk3TF7RgPNgcjCUxjcqWyh8uy4Mx/thVXTelcPXF3b/Wna7P5g9
tLAMNTsE1QhCOjcc1fdc2CLG37A4IOLB4WBspS1kA9Jvtg+A5DBD0yzfziX1L/Yn
wqm2OiyWsANujeyEhbYkaccAtSWRdXN+5ZKADao0p/cP6l45fdOT2pfdnxEdKflY
0FGINe2A6rfI9Df5paLDODErC2T6dkopGdbmfVnmIw28bBMWetPEi0V5NJjDQns8
MgKaHx7SFTNVCdIl5xnXNHHgOCdBWEd77aAjCi8Ix0yWHFsAEs+TUp8NAU9b5AbQ
8kiiPjNCW/C4hf2qbWeFcTcsaNmTK55MRbtdbopVMcCAY2Ca2JvHdR4lRPSzxIKL
SDq495jJpg9E/GL3r67yIJ1fh/KdDyzO+e1evFr7oDBEwGv3qW1z5ixICgB1SKV9
2j8u+ofJzlfRsvqPfb7Utbw9qCptvxVxdSHTifn2mt51mWGJ0FAQ7QpSEmFrGPRX
iFGmEyxBs7RvIvASyDmTcdDmBhWrnoXxI1RS8fbaE52SYUE9IqbF+e8eByGfqowl
icUfVdLP4FPojFGhmuWKMTHCC0s/DG9og3GWo26R+smkpkrDMrS7f6us9+rKHOFb
D30mxeuf5beCANeQmfL3hm8UvuZ40GxzhrsRFSNSLWKmqmAp0pWJKnMZNCjSGMj7
Nb1leKSaxbsp8xrM7WkNxtGie89sIv+q770fSNxjIrEqr/5Za7+HayXEhK/gkqwt
xzjsnZP+AXFhQRKNlmFd1LVuTVpiqXsGfuMgIzb0+HZfzfHFATTdMgFMHCsWUspV
h9UI5aI6yzzbUqsmLuhsUgiCA+6VrwVHWu0HwnBdFCqC/5+EbjU7yZgssVGuV7Y0
mYtaYjTMBEW2CSSC4XxzIK4ZIrHpE4BD7tRyXQ1GtrTGtLfWtEq2KYKOMvdjSTib
DJ8kaMZmlPigQncbxba7PuJZdoUXjKEDqIm/89qri8fbWM8blCj1iVFfGeliyHP7
zvUytCOj4vCnSMiBNRluzaIbscdnoTgp0uBxx0Q+gHxR/BrRJh0A/NXwMJe9A7/H
zb/pY/2eRlvz73WAPlilpHWb12crYBcd/MUJqR0Lr40haajtx3PkMNe7LmgFAVo1
1b6wrxa116VFduKtWPPAZzHd0iuk7IWfpnoVrYkFQJlxr7+47Mvtxjox6Qe9bWKd
kqhxoTwOO2w0zq4sr3MqOM31l8RJH3IOcyC4gDzNkuSFri5hvIyc91DuvvrzyPhb
g6Br44HbV2qF2iRa+SdQ5ZGvJdgMAo+GnUGIGN+Raf71OmWloVXOcIt+mVFlIJ08
xv+WZ4/PeKzqVuOhaQOW/yNG4ySLbe+7WNPnsFzJG15ymoaYMvY7tINsp+m4/zvL
bmE3X7jWGwGuI5gjRytu5SzjDaubQcUjXO1+uEnHBeEaiNX3xnlPiSkBMlAnFwlx
7lhVeWNhrAPkSAQtH3IDM8/cCUg7206EYi+vlBsr4kdQTXqnw5meei/TXptndgY0
vfaJ9M6N6bZ0THe5jWf0lrCrZfjWOYLOEDcUV2U/nioyUHUnxKGyfbJHv9S769CJ
MfZOrwd50mcavbhz6ovkVRpY1yIh1IgzKx49elDwL8dh71Mobk8eYuncE/tTfTpL
bf5LapyiyWqCq44Bs2ZgiZOxyUIYmHJnOZ09dr/fmDHeXuQvclObjqJFQVgbuRV6
t/YEdyPeA5nbR2ZyQqhtQia1UkklbQgpVVakm2QS6Kg6c4K+w4qii7jwtEheYgyz
wqNfbpbyk0omAioL0t8383rfxnmPtjRm3pGluLPSFbckMTu1jBOD7SJEosHsqnx6
msEvvvao2ni1ife44290u/g/Vc/1kf8YDqfhMEfXqYDM1RStGxgHTMMuSjQ/UIrK
0iTD+tdHJBlO3tmXhHFZz4cc3P7Wd57cRuWe2Ph/ojMP78igvCH5dzVUaqpUTXcV
KmAVMyp7zhS/iR3aEzdZIlyjHcXoTyCwcz/laUf/DnD6iWNd6RE+vFw3B4OidCEy
AD75U5kg4cuChyBgVSDk5Bk5U/J2S4csG+z8rCqte8T8dtxG2axKOZGA6mg1bn6b
dlK3ZC2JGuB3BacbevQS2f20hM5Pmcv7zlFLNf0a1ln7d1oiKXVND+4sdpULNYXX
nXfmryakEnAUu7429C1w8SKtNaMNo9vdLObhI/pTk1oQoKGQgGZx4EEg4vAmkM8l
oPhIUVMtjATBeLi2FYTvCTwc5qivEqfjsTTgIkMQNdiGFT1n+IJr7aKw9Z+XvJQe
F9c2cgxaaqZNj4zkG0O6WREqXHHl7UbwW/H9XYk4BHDamicRqqWG+w/YX832gWe4
0Z1MJm8H4ukgj7gUP4iISEJ6lPYXh8Z7ilzZbAY1QnBn0XV4ipHv0P7GyOuHJwWY
/Rv9XXtmbG79p+F4Y38MMxsRsHDABHp2tuRbRbfkx3I8wzkSTp3WHp6kkIBvYcOE
FaNPhYFJWu5rEh0LDblT035kZThecg5oPrQb4eSg3gL7Sq8xVlf2pnbVv/YsmZgz
uEBynmoChe7OXR+hvbUjyCBUhp8zIGP9/UWt3/sQXyC78Lm6mntP32qhMWA7fELP
/pxhKR1CCOjLC5C1NqDSwvSqE8sHLYGQqI4RFnQMkQY0RwjbpwRD6qsC/vAkmJ5S
KCm55QQkQekB66qavzyn9Rd2UL7au7ZNqjOCV2Izgc1bCF6rHs8JhczCyAukW1yg
4wosT5ZX/zxNKjy8UNfUKqquzkAEXfJS11Hbm3lOFx3kYG+S3x2Ty9OoVEXdm7QQ
CyGQVBKJMd9xHbShorztCCRHz1NpMFoBrc7XQyT3oxnaz1QfXUZZdSaPfvto74O/
MUpqliaUIHQ0MpQZshZRel+AhL6rLrSAb2l9QXVOpLzMT/pmJOstQl6sS+XQXi9L
mMIyI2mo3lHzYSxdC5kiIBAkgVqx1a24/C8qMSE2RhjH9LPL4SFBSU+ECmvg+1L5
hZBJKJT4dsL+48qJeJSOol4B6zZjeOp9ugQbcG4EXD8XvP1B+hXhQeECaSQ573Z7
Y2wW0Mllw0Tu6Xxr6+Wz8GBWuDqbfpr5rQd8VJSG4FNOdAVCZSHbtjmsorsPVT9O
/Peg2rgfnIlyLMpbXVtWRZfUgMKFajLIFsbWxrzNkqvl/V7UlKAX1Uo3S6hzdCPV
SeXEYxn3l7yot9ZUS/gPE/kGPp7v1KRwXPn2iup3WnjzpyO4MxHpEtG2uFofxo9K
5bFe5aj/Zlunsff/aW3/3R3zwz+wx65oLldI7xJwrEKGFlVXiBeGtTOx2BkTKc9d
+Y0pnMwb+O9kxEGgTXnsDc5lzZPrGAUyz6QwNvgrZxBxYwlz2oYZsHIWfDOp2LjM
toyyt1xCg4VNzxSf7SEz96UyI+ioi/cSGr7137qllpiSpyNIWz4r3tbZeqty2gx5
+hUPoU3AMsnBOa8AoK5TheKnFBGTaxzrU4IMpXOuW4p0pq04nHYO0R2GlTPER/aK
reug8yvx0dE4IyzdxVnKB63YXjmP3MOK7480Y0qBvy9QwS5nKoQr8X1ZuKPkLF5q
iRbY4Pfs8N3rSafkz1BmM57lX2k0lVR1vZbIJwUEpcofxrSU5sgqJ6QZhEyLzmBE
KA7aJi0jsgnRacEfNsLBALVZhA53gWqKMHKJVJwmzFPfxUrcTHs21GEngVL5zCkq
tHrhYHuWzHvvcyWtUAMukOQl2nrBmLONDGbe+7TpClPxNuMHFg5gKkmsHOKnPWlM
wGmc/zvLtFhsgMSfKRtCnVnSWK17vlNYPXqLGGXY0R444fy7OScw+vvF+nSdjsOI
Aa1vjt+IMHdo6flEp0/M/bjmAcndpLfx0b+e1nZTL7xb7IcWvoic8yIl68kyTpCZ
T3eI1SKLL9IOeKnKDzFETlg2x+hfkeieH0KNcvIqcSkHa+9OLw3YLPurwsKqa77W
ytxP/n0ArX6V6YdNWQ3aM+wIy4u/qjAajCH62jv26I3xNIksHW/MSlLOA3lydwpQ
yxByyvPMSLE96RiZB+zGZ+BAanx4XUsqbRltPnBh3haCp4ZllFAPeeLqPpoDI+OH
6/OYtD8fmjH1P/INBgK83ivdErzCy4pIbp58+Tz3yHsLYjbIJ+ghmmghEGtbwQoS
6hdVVYhLS8Ax5xFB2VHIyDwslN5SrIT4ydGrMNxPmnL8tts+HJDTiImNWtuv6PnM
nLtnybZ10a65Jos/UVikc3uNiDc8mHsNmxdsJgzG5Wfj+l8Zax4zZdDhLZdKCI7z
mO2KU8yqsmYYbMj9HwboIr/N88Ra97ow/bJ4Tw+Vz5aS7vQ3WOvgWApASlgk3Lbm
r2TB0Gt1yqSgtsFk5XK3MKhvuSxqWsUfcgmjit8ig2dhgGOh0VD9zSOmqYrCkf93
c38oUl1pFYgjVUKPSpJokQ7jQ9NJcdDByjwz3pJMahATTSoeGhwBtgcWNU2Ew9Xf
tkXFc6s5A/9MtxF/KES47kc77aSeq+/Mt9iDR6yeArrWYqXvz7qQkc0N3Yuw33a+
kyUY86fJ3X0xBMVm2uEHAmQ7FRzMoHf/6uZe7sPP4iG3Ox+Z0SYhSgVVma30p/2n
7Vt5EZY13eA5NYF+QTgjjVsVZBwuRiFXr+TK1UQUkXCVeRCUu3KkTIWNS+12/p6G
w04VpsRq6Vq65g/nqND2nChAKH2JnYLKedDaj624RuzbKDmprJ1S3xxvDdqhQWVs
a8jpqcGn7/z0KKOFE6nz0TUu0CdL25NU01ZcOyhIG3lxYvJ4Pz2RK15LaEAviYST
aKonoFtWR3b6FXbA9cPyfyTltcq1DC4WmIhBUDLSyHOJYghPgzPNXPdye2ym0ITl
C3JXbUs3q5BuzG5I3JshfkTiD3vC2M1HtPAGZk8qubPrkoWBbOW8TIICFAr+5Bum
GIuz2tMaiYNT56tgHazZnSrFgSHfkflZBeOHWMRfou5Pf9UBA3S+PV8IblPpi94B
r/Sk6KYp3O1tMDoXLN8Mm/DjpfRxX4A9NUqX4fUrVyxjeyGJn7+5bRAlik13KbgI
uAObwBGDY9CN09gn+H41C1OtrQrSFp+Z5H50oz+1csChLerQVmmuJwVylBw/GQK4
ArtSbesjgJ/92ZPjrmbZ5QfB4Q03Rb4AfoD5I7FvTPy7UYSMwnolUOeetWI8Q+af
bb0mTVvXndBnYBlW6F6HSk11kSvxOrH7uWt4fftN2rrCoCgvP15R1AHvj+BsuStG
CsYWiC65zDSy4/vW9sTrIkYZeJoKwrqvSHi9RmbFS3jw8Ce2cSuDdAARy/kOusgV
r/ULceODgFvsBiX/5GnxDPepKE0ZQKs7p+eTtCHQYii5sCO3SdWmZx4SGGywOJ0C
OQo+EjS4f0mJtOHoYoGFFxdVgbtVXcarth0f8/eRHDvruM785j2amLfCrsm53ba7
6XcfbZUc7jeVwykvzbfFMqejgEsMKoEA+THZRHc9n4ZUAgf35M15IiT3xIcFq444
8e/6a5cr/v6p3KJR5SdTeV1Wd4EsL99+87+yci3X5mFK6dI6yJY/1mKnYyy4VyjU
3jW8vR1JuBTD94rQLL11cGYtEYaVVIJFd7p5/MrRMGg8fC0d7O8gSiVK0dxZj++u
2I7nKqDL5TrP0OiVhYM7as/MMh9fBg9dxWFzjpk3/eToZEOAowQNf4rAGxjNYBV1
ZE+5dtRThMmdjgUydrJYxKMQv/ZgVLisyBTZFPcpzwIFV4n+ZdBEBVZiPEo6aHdU
fllDdkCy+cBilM5Vm7Y0Pm8THLeGXTmi1koE+qgOe9Szk1DgAjSZ+iNwocB+UtqR
cOOQdGJDOBkFo85qM1ZYMvKmq0OiKh0JEhuFfl2+9lDR1AIztZRRENo8seBosTT8
nCa4hoaMdzfZmU5pgyMmKRBJTrVLfVLbxoJsjow+PeTikxPIcQZBc5LuPiq2Gl9Y
jRZ2GUWkx6fImd0a8CzoYk5QvvstIAVf8T2AmvIivjnEcRXjZneMdkoFUBKxaSNo
w999MGtnW0AVnyM1yvjxtkMz+Vq6SkHYrapXn1IMYlkUFeFBq0VOdmKK8ztKS9e1
uqNgqPsyUOLdKItDiYeIf9yC2DJ75UIoPTUBT42EVGOVtEt/S50k0dqvcRKnTi5u
lK0ed08/x98XIksbiwTkzMS+qUzuwS5hHFQPlg6H+dfxFd17SaviS99rpY1jHEXj
VHqcdkI5y04iItVoPxHL6/Bs+T4VShPhTYlCX3zxBHLC0UMw9cPalX7FaGgSP+zt
qXFPXmaAq0nrzY0oYC2IQCc65P1fBwfY3vwi0Vaf6BX6MnGskISTdw95y3RJCH2c
BMiX1VKI8D9cBN8BkC56FQ9L4JmNRvrvOK+9SAkKh+IOyrH5JnaCYrLd6ujBBDU2
y76Pfv1MY2VQ0g9hKMUd0oo0Ow0tX5+ffSR3PsR0SqGSKVfMTJTx7ndanqLPRvcI
R1hmGINh/o0OtIVB51LHIfRQJnlgDR6HjQ0cA6Y5bqUuyjjq5lQFQkcnquEmruam
EA2YCeQLN2gd8KkuDH1TIe7XlT9pALsyI6lFxx7h4pvV+g/CJhZDsGIvwSoozZsV
aZHJXD5IvohmVeIZgPnHUCrHHT7nA4q/5KHVD85YtsQEmy93nDw7Wl83uOttgelM
aXCI+WgNSyxkPBa8Gcowz0Ft8jdX2OUvfcibTsLMfKLtEZQfp+FyVJ3pzTTWnlRE
1wav/fpz1t77hwHcWQ/bhgRdr5SGAZn3K9eucOoWHgN9GitECLgSW8OqX9rxX8iv
KGH0vDulursxsNYHfjoxF9beNdhDOwoansAx2FH18CQdOdl8BH7Jk65crIitTlWZ
qqkx3D6KYAIPJCtYr7UhJY4/wEgerptiWMWCHNmY7pg69nIG6UJyl7a3ciOQBHSu
VzzOkRDaz0f3ll8yzjVQJuu0XTzCEsrh4oGLewAQ9Q0Lt4GIGe98ReDjuox34eP9
GJkLjcLsr6mIsjHxaXMR60nC5gKiDwLkKGYm5NJ4MNMv2nVkfT6ktcjXLgYy//iY
IAYD3jUwFtE26tWVluB4aT/zpsK4gfKaPmekBN1GAJ0U5P1+EeSQy4gFZwFk/fdb
O1jH8oowvrCaa//mR31I2BK6Wtvca5dFXzXh6MGNv9VLgE9ScLiD6ktKRUBQWa4k
Imd0aZySNIT6OOqnGW6U5onjzd72yfdMuDmzVlKvklXKNboRCp6mrMSXc0WsNfCo
F8tLBS9Z5P6VeMcNbs82iMkFxcuIZTxkEJaOC6YoEwv3MJtIFIizld/2phtn0jRm
e7voEUP0bVAxJUrsIqIV6Tn9AyIc0fQR8P8mqW+1VihwX6sbxzFFzkZkOlcQNm8/
7IwIzVlwpAc4JedumHBdpmaj9XTxC/CLyw18yQCjpU8gA25ILsEjF0sK+8zOOTOj
Lj/AtZri+mzNoSD41Y+ONyOJVOoSdrWzrC5W1rDnXXmK7pXVZ5llfPUTtuWeUgmx
6W32BpSAxA7696evqrtqtO3ZzhSufugRq4+ngPdD/YXGDdAgeBe1azvyYN3JBIMt
3Aa6nIri28q6jXO+85wtgtG7QIUGu4yvpQ2BhMJQ3Q7z9tI3Ji7NmDYHhwosdELH
95tBSVQa4lecdSVi61ofEaStQzXKcFYPtEB1lL1YAcPFXrBFRPsf/5a0Sc4Kou3p
wI/B6MwYMQ0/pA5ItUzChUXIlDwKYmRmar0lWFQtjbi0q0fHOS1cIZmA0REZpAl1
uv5VPVOuTs1xJ8A5m+K8/djKnCtQv2g0af3sALwwhPxaK5/n9Jn5aDS41nuRH6fj
6u+QYGHx0OxeyiV9hPzP7mX4etrn9Bh2T+hn6CTxFTq3fx3uuj8iC2hVXuMqI49R
O/CiT8o2Kt/42o2oC7rsVxqQJ26zjEabkSoJOpgst1CkaV+TkAo2hQ2auiWwS/hh
law6Dtumo+9JnTgTpmGfqzN/AAwNuDtTw7cGOfoiqoaRXo19N3v0VwbfSRlkZcrU
CVSE4gkj2aPWFq6MPM9Y9RyWhJwV+TkUZoSdi00gGxHptfl0A2XkuZ8HK0cNmiQa
t5Ra6aWGG/G8GW7XP1grgPxPw5nQVcQ2SKOVtI4wOXRNcYoS8Mz7FdH7CjCs5g7D
lQDDbMF5I2ssqHGixdwEKEfAaI5a+w7JgzORACExsTv2h/Lqs4yPJGrZ2eIEglLi
+iEnhPIth5IzRmzMrkIZX+u7LRbfoyw+TKTsnRAblB1PU882rHNzLK8lgWx3kxG/
r64xuedL69DVvbMRAECElJ1r6tDA6UVVsx8cmRFrfzOPuOYaLOfkDhfXrA+rZilZ
vWqGfhJyvTDoD5EZDaCVVpNaT3DnAvol8gU2sF/P3JbRhtOxnDU3RdZedWsUJvdq
66tfNhj0hRVKA0qp7Q+Gifr8KWMCTw0pEFdiRXmO42B9f67Ohq+si0k1jCggK4KZ
qcKt06ZO5fh4SV4WlJMQoEbTQpmSb0BV64a+Fhji8TCzdk6JjiY1CR6oFDyQVUow
CuPKxc0sKgDMmWqY20+zQdNAxFNg9qORKR2+K3i7YoS43ZI0Kp6203To7Sq40N9u
DFjzr/iLGTd4zpAeVJRM7F/hv6r8bzud50BD/+IJhjVs1/YZ+pmNDTojEaw3N9JI
6z2Iol+fiDHUSZeOfSj/DO5P8ONd8/HHb516f+6lnUkU/AsQBRh6gP9aNjy34hIp
NF7BlUnwyjbOX+qJXJB/SmpD1EK0/FWPki1LBav2UDpnc63/ZwDmV11jxmUN6hUS
MN9sfslC614EUzpeP3tz1AwUKRRyKhMmfMc+3+gm7iQ12MIiO8NIC61EYsVJoGkq
2iGAQbgD/Omx9WbbzDA/56ozGibhCar+HIVYxlaK6JPSZrYVACbjAZ0bFPNX35ak
FF/5FzFIDuXKk+wkDI+dhC2PDhbT1dqK7J+XebR+dJJeJnzuKckqz8eUNhIpgupL
xy37YVlhcBhT9GuXPEaBFqSdiZuYVBEGUBE+VLO8QzR3TNBdHfYY4wxRjHvA0olN
dwdvzgetRw8qkZ6OLSCmnCqfG4RyXKmKi8U2RfRsS2cQR2AJMYQQD0uBckLVuqST
vzS4aZJA9hx7hDVzhd1UfgMrM07n4CtbtdK2AEX2mz0g7fJXHiUjiPJqKs60Bey5
oGJcH/1mCxrxG6P63sxIqpsLtw48v2j8/Jw9VwiLTjkAfP5AbfnlrW6rzS3m24Tk
fxlbh8qOK9OATNRJ930fi/5H+iDBx9Vp8ijQXQYgQcyHj4H2nJE6hBAUplaO0at/
PSrGfbOkUHU/H1oRJBxPPQNS+UMMiTRaMwDpfTTdllbGIzU8yur8Skli1c3LPEH7
ghJJolz6FoHlRmtLPber/atfeP0x2CCSDLbRaFZcDWg029kZEMrJXeTihDbqDeNA
gLsghd0cajHHnhKb/9QWAM3UZcGjCHf6M+48PMBAiC3DWlFKvYR+Rct20NKyhg7n
1NWnIseFtDbi6IZOxQNwvJrB0QtCJ2S5PSl6LQOTh29HP0F9zeGMUAJnnYts4EGE
vT/4/KKq6skQL5SHKc14KSl5cnjAHAVZ7IyaQjkCHgYbi3LvheBxri9QXs1HXpk2
Y6qGbgYjQKJs0mw5UOr/3AeEAWHJ8IZnirc2PZ3Jeyqw5GX1v0nTR3CtZetkE7Pw
EmEiZ+L17BJNd/pmDtyZ6pJGzOQ95XxdNQBhzKtDrlFGykfv24ywbzKiftStLvcm
mqZBBpOoeGzXDKUbfyWfzqW0vSJfH5ZJy/AlykTsV6/Wbv7BFQQjLRw/Kn5zu12+
ibt8gIIDIOrinIGxAM39EdZwRJct2mtnIulsWoQxeTUaxxOjBcR3id6YQSpIB/pa
jmLg3+OaYwbjLN73Qe+SvmcnqeVGdw2MlX7usihaYbq9F1GOlnWJuFAmHB2MOpRk
i9238WOHPYrKWBZGZM3MAvZsHmwGQEsNuBsVcLqUyZB6HHLrjG2NOezErnwtkrL3
59NXO25EWlN/1rMAiLbwaCF1k1R5P70lFrPcbZlwd/tI5rSGh6JJz9ceIr0W4LNO
6kOp4mV7HARvI3p+R/k/XsyyfSse+BBFKgfVZIL5dJ4EEY+egWPEhjUvhx/pg3j9
2Ti2OAvwBmvd7RkJV20h3oVktF4L0W944nYmgsnTu1xZZnG5lGoxwUm5b8Xa6La6
5yRCQTGH1cruP0IzM6dtX5Ilg8KZzpbK4ZOXIBbwvnrvI/k+h+wnaaK3mC/bvrSm
DZdF3whyEphGCq+JmyRgV4pDVcsbzvlTgTIGmv3zfygp3fYnZ7KcZBShUt7Uumb6
f/NT0NjGnDZU8UDgcyaJeKnInRcoB57XC1n57bH/j33S1nnBBBf+6mYSjUs8Sjus
526KTGEUc+NOzFZC0vWe0QcLczd37Tf/nfDAE+RPWp4CY0T4F+ScRfI0GnXB+kyH
X+uIBOLmg9MRXyeO7Yo5oQ3LR2DFD+O3eTzc5PlNzGBnFqI86EHyuShqAE9xDMqf
l0/WnerGPit5gdyDy4bw/lJkD+M+qkYxw+nriGe0DhcUe18h9S9JvP9kkLGIOTWt
JupcXkKlfdWpO7hQJ8SJ6NpELhFwrYkIlUsNCDZ8Z7J7Q5Y0w6fhVFqrnIsb2G9G
sMtRViFHtL9d+YqM0Znb5t+VZQhok7HsBGLdvx+D3/dqqYDDgvIGMyQhp3L1NHiw
pJw5OhDhAai62q9gPuMfUzXXpzT5/QHp3NsPokQATfVVx9j7kuZOO5rQ4UXek6mS
XwStp23SYpModfzmkCKcVV0uIei7YhSxWL0Z1uPtrZK5p31pKAJKjE5vP9bn/kOM
4iLea96Zrr+l/jok8kbQzADNnU+BzC2FYufvM+mWQ+8mEc/+/ll9DU9EjYszaOV8
Kn86Pzh4cq1WH3GRW6BHqLeNFFdvkHgYKxWReeoXTjFMUlIJBce0S9f/35qnd55I
mptVxDcrBcEd8hfVx228J0uBvqyaOjfnRsqdAJUXC9B1tb8I3Ok1t7h7on+1+u2c
oXFSQOlGy3Z42oBju+fULonV7uSuERrxDdhs2KeFphPf0JsLllE+J1pVniE/O6vn
5S+uykxXuyjVTTWrKz+8weD1owNWIxH162myfcRRkRKVvnxy71GuKh5qi2T6o4vA
nbZM9RYsDJk/cEGIt8p+PsAZiqu7YDiYulvtI523ko/h5xBdIPdTb3y+uLx6Q7BN
0x5CkncgKf9JJKZpAnfwcGiUZ6Ze4iBFMrx1eij8B3QI8of0qjL1nIJn715O44Gn
LbSpRwso1ZT8G2h9q7i8wqIZug3ozipMITDXYlFo/JRzntgRXYUVO4GRcmv1tpTt
vkCQT+PEEj657ZLxXedCN9DxitIQprUGwO+WpvFXxsFW7BPsCyGED3ysf5i8AmDV
Ty1XWtC3ccAiDfbUE0VORYwChHfvlhDJt7uYkSiSBnefu45B8p9SycRDncL5ST+m
D9Lhrek0SwxP7tb5QMWp4w86MFo7dcGt5AkygzJN1WTCfi1kNH1hOaPWGBz29X4v
JIr4Fz18aT7W7tgkKODOKLy+V1xvno4swKSq1K2gnt9404rhAqwcgHi3zYbAwjJL
tDmUl2WIgA40Mo3qxsqct8Z3xoPjnK4GXiBcy3Thq0xfrINj1BND6MlaxjzqwelZ
6UZO8Fu+08i6sih7smfs6Mul84CDuub8Jwb8+CM7bljYnecjNuAr5+sQZWbW8RCP
HhKl+GNRdTtYSQ/D78REtdW6CqG1gSNRL4ZdcWtrntov1iQOWQSqFzB0dlIN8Unc
7OyhInuhr80CB5uPv1FP67vu1bOBx2VWgXP8P9L9TuFUueRIcONIO7+3ya/JCZ/D
PdbW0RgrDIuhaE5OqWk7tuDnHKyLprzUAa9I+i79S2iRm9jiD3yjkBsRh50GzvU1
v/IzO29sD1X3+DcbULRshj1kMGiqb6VmsVyMwcuIyM8B6PW2QtpLn1t7OqFYA1qT
xxRGrtE2feC5O2xDPIquRjEyxCzTh7u3CccxMYEgHZjlhURtrTTQoSv7O4oAJzWb
0SZEPiCRpSr66VTlz35N/200BnBRWrDVZnhBkbXTUzQc4tUD/xo18IsvJdnyY5up
uJQdsmWr/WZ8t94dUKeSGClWABWmiDKsx5Lltrqy2HU25rw/Tb4gREwRF2WJtJ5x
ZuTKWLdMcoUUFLdHBHMDT5VqMGz4PB6QEdArDv8UsPEHUmawYPWllrWtlVSOMBUO
aA+xsGQCbC8YnNBrpbzz3A8TaOOzsvKoGg37EzLxM/w8MFoPhEb+srxlqaulxWlw
pnI5zBsN6tpLVXVSDsm5oXeUOi+gi4p8Rj5Xcpb1loZOGR0+aXgJfXVB5aMo3NLG
baX+4aDJiwgcRZAM1nzhwgf/xx4QKEFsTls6Sg2e6CaPCF/6sXjFW8AtqJ5ucNtV
/2dkDFeFS02bSy3Bg2rrTJJ7Rn9us1trS/2WzpmxjBUtrTNqhJ7GJf6vnNH2wuYd
h403tgfcijWdr/7N2blvxICDyH6jVovz7kVV7vkINombGSDRbpxBWel8r5x6XdQT
kozwSau8jSuKC0PY0SutNo4sL3HttwakiTNgp8hrmoXxNzHfUl1U06FoNtr3Kvxv
NTuPNJSdfr5tff5xX1Tx9CZ056Ysb+Og70OmxdlP/16E0Bcj21RVF5X86b3hEJ4t
fQLWIdS1y2pSro5O8s7pDWGsk7WzmYyVfx36Tn+g80DP7Ayk0symA/IWA5ZeAl6T
4d89T8lbKtseExG/Gef8pOCw0U/vqk/Xz5FlUqyOilTuupCai6TV187ho4kKfgev
XGpCLD0/xqo4c0f2tHb1TrAsFqVhkYOTYQ8f24cpsbpdlx48tEKgSkiuGIpo8SkP
yL6Qat0Mow1vRQqPta7Eqlg854H/L4B39ilcO0FfxBLu8iJ1fkVwOVzqN7Uy5QeJ
bY36MWBdJuzcpi+CH6ilHSZoWCSQWWldq9gpyGxQQJVyRsaF1v4mURPEv2nQG2So
dfUI3uBDjPwzZJYdmZDy1Qf6rjktOn1euce43sXoYeIIlR+bRrZJCt8GKwIgWzPh
OeggYawmMaebyihm3HGC6epwOpazXaen2VdabntFRWv9NwE3cc6NCluBTZ1ivkZE
q2vg5KqEEewzamCaJ3WT1TaxLjoxpKkqyjPond1TkcK3G3tGIqr9TFQF1L6gpvMy
0TAq+Div2QisKafqq8wJy/53leDQxaaK3pl6z/aYQ0pypb7kS9hIefLuh6UXJnXo
wxNYRs7jImCNyl4Y1XHKdIkM5qathuCqyBkhoqa4cCwJuSvxiSqSPBy9kS4/KnX+
2sh042EzguStCuJwu+EMCA/xHApGGMR9kZPXYP/L2srIg6p21DgWe16YY1S9Gskm
Atm3KZDdbIAyR+cpSPF457uI7ekrPom2PcJRTdjJ8FJW+NfgPplawmn1MKy7DbJR
OKSm3wHeTynocH8MYEQ/zaJYReCKDkqHmIGPER98tOiMIRI1VVBcupKL21dd0BgL
dof3JZstnL+kVGhe+T2mGPG+eliz3/DcU4JSnuPTWJkeXPAOWURxw3/XeRLsfuMy
dSMumDhEAVKfjeWhCy+Oh20/fiEMzLRzz+6BBW2iZZmzltrdR8XcTFFLSwdXs3NO
D3JbnZKqo/EODFzaWo1qpu4nVftQgnOT+SpIKGooXwArDOzyxXsTUP4R5iafnDzK
p7/53xUM2jtQaDsOdiYXn8oufMVUQiZsR9K3geAaT0ZKe6jOrcAaDAruhmgNo/bb
Wgt53OJpB9IYtUvVChUnYDld3y4GPK3JavfKVdP/JFqXIwLtMLkTxJSVriAp0uGD
TDz0XfzpSobvZn/TtlTX2MpEHuFgtMfd7WTlCkImquRg+OXl1dkSYBq2OiZVQXee
NaQt/99JU4JtEpzSBip7/RZg6DneIeGXaePBL8WqajZmpz9ymDdrSOhCwvZ7/ADK
7eO9yJBauZCNexA1zgo9vSSZuSPCwK7e1YbuLoSPC0apP6HqOs51pzABgHuIMlWu
9ryFqSrL3t5wyBYJ/deMnz0RcW43L31VyysR+AeX3ZvSwOJ/oSleahV+Lk3mXIuF
YKPwNd3UhB4wrBTROST4GicD8ieATG4dDcviTYgUgovfedRCypJrGUOC8ZBeGN0F
tkqLd1nV9LUGFo+Lcib/c0E1bYRrA9MHpJI+OfOsCWRIaX1ZxZonDCJhhI9tlCG5
K2x1rX+vWTS4gCTIvzXQaEM1Q6K4bnOPPkcS3obpQ6drq+UxvIBlqO/IC2iewxOc
pcDKMxfqZVuXi9nD3kGzywrRxfiP947gyp6QQhtObV7MoOG+iHtSqEU4jRZQIYfr
iIvHYUZpAXzxHhMGiSqVtoWkpADd9VWt1Och9sj46RAtMZv4KZhtwSsoa2aevTlo
0zBHbcX14tzJPecNI9Bzo8Mh/9rJfJjhV2zEuIbaHIhzuXnJ84Ovfaae4rSv7IwR
8vOKgPHbogwnP0Y1vW87Nobh3Zlexc8WZ13uEzTX3BFwXxEOcRuK2hG6OBpCIuHZ
I5fZD6YMeDYsdVnZrbRnecWMHQx0WRaMmfZsu3k6gblCaLAMkrdy4LThPzkD8jg+
PqGM3oyjmQeOn9s+Gf1V89rXNkrKwn9wyAiiQLDTfhN8cpxtCpjY0qlx5voZZaQ/
dtfKzLgG1R+kDvAKw9WR54BPCr6zzfx6aaL/BHgDWt3FK2ICjnzRSPpe5Rm7+Ti+
o5h3YffMi2l2aToWh5/uMi2Z8z6GiYd3VjAgV3gB1HqMK3REs6nNP8Cbxqj18k/D
lnl66wbVpyLoTQBFeXjmSHcG8UGNJR+bBcL3+bcPo+k05ST4hhGyOm+mJcjE3pQS
yhtNcPK9HWuBB4+9iNq1FDVFUlt3GMrEkubAcM0AKDwWjE+vBsnMqKdd+REMbJnz
zPYnitm46tXV0p4vS0TDd1BpUkvqyeDQrO4qDB0tTtxnD/flIXHV0BcchOUdtPlz
V9iiuOFarQRXQojCwktYtRPrSILrbU8jn7M4g2bygqCZ85PVgMw+0hbSsz+fehJx
/UuIhkZDB9MQTA7tFmo3ZegNqrZfgSokpmRrj/VydgQBXrUAqyltMSoqFucogZI1
NhBEAQ3yK3GzWoQAthloyEhJycy57IRkjraUx6wq1yyRaRdsxEjVr8sMKV6JBo5U
8ZG8mNxLUpcZl9GVxJ/3rvGT+Cc6N79iehtJ+rJ/Ym9A9cbvhHiHwLWkkkD4OPEl
i9YFEuL2xFnKY34klXBxwYM4Yw15JEYaDJ2RsHUsNSfmTb61DLX3qCvpVlmD34aq
VomY4HHJOPgYd/TFt/2ddoCXQH8o4BaFAO4y5wI8+m4OCN/IBES0lcQrPan6NZUs
mzN5o788S2eO+oUpTriWeOGdEvyQj7ProVdCRkVy8bAvE4VVUaCvOhP/ieI3gJsH
x5gMMitHFa79n0k26+UQxIfUEtZSIAqnlRwZu/KyiVmxmd+YGjGVfkx+NS1Ozgb2
up13RyxVHKnD28Mzw6OI1DI3cOCS9TY5SGXkinbgILiKDh8q3dLs647qMn8Kz0xz
iprTGVMx/LNkxm4mQ+wWtWFshm/oSjUau2iaibdlp0/4r0Pq4l7mF9+M4wByE/Ap
WWYnxNrdG4nIRy2i9nZBL19EOE8w7oZZK+YmfrwPJ0cTb5v1wyS+1jNgs07cWpRl
u7Mrhf4CIYMlytISVpLSvzY4JNF7NrkpCm4hgIE64Qncq0en+7XiQztT7/yH6McT
gqiP6tKkyADOdr1cfYoaigZUY9mMTLSl66C7Cx+JtRDcVk0Skpo02RS2o1YADObx
MZfVH2/cQTel0lRcd4+dX3Q+97YaqTsQG35yHjeaMQBnJVqL2Y9a+05wznvV3/pN
WBhLyUUbMEcadm4r1OvUXZ31Xy1FoD/Kny0AYdga44U40T+vb2P6ohkb9/S+jo/A
0PN2xTeUfTyRkWMGOeam8e3gX+q+61zVEZCARa3HAsfIIO4n+Vp0M9E+T9K/b5Li
/SUr2OAA9RVbj22x4pEJKsK3wfRWycnIVj6OaNbrLjqIO9EHxMnfyU5DGSA66bjZ
zUI789wo4tb3bIoyTzWVaUml90DsNLy0Gm9lCRuQWmLaKeGEjDRP0Mic3FdFt65h
Zxk0H3NfEiGo7YnIrU2cCZD8NBVdslJ+S1Rgjq/hXZ6rLWOzFF4zSZYUWYXBarLQ
JwtEnNaExGpy/v0Fl4rf3NBhziB9xDNRjSqVAUzGQhuMU/CP6vtVN3dq6L6uXpt5
h9ZU6D3fxfeNF8HIpwKB+f3pDJY9SUiXgUvkRcNRfGM2JkielvPRhkbxP/wBuhhz
fiwNXN8jEKFYPfC5nM/vyLrcj7Jf5I1lg8pATfsJK320cmIXWgW4Nqt+mAdJkn9q
9o1nGHERf0mhx17C7grQvsg2ipYqa7fMm9KbH5KLkVssrJN86IPnXOT44QcNQp2h
Qae7Hmtz9sCojxTrWs2Zpxvac7wowB6uYnOC/uGn+wGTqr1fh6WwueHOEjw21Pl/
iFKmG+LSvM2yPC6lKQYpcdYD157wtLmz3p6bA68X6FvPSlOze2/tDdF8m8KyWkKp
+aBN7BPP98YiexNWPm/IKSLNONpi92d+NXvNkNlsbaVjhSr80qan9MpjTeDDq7kY
SeHrCfI+wqh+/qcBNLcuuNf5BY97yOcGe3gaENC/Szyl92IVsgYdE5g4KKy48pRf
ltee9sPyM/TqNdBsSjLE2WgeFRbeosBptn/v0WYf2UjcyNVIWLT1qL7Ze6xkyaAy
saIDBK1+zKIlXZFkSFC6BttWmiJeivRGu3faCKas0AHvqf+2KkoDgfWauWbeEp2B
Qg4tPRo9uRg/ECoe0qP9WZ7MCdc+9+v6j8ZQ1M9HAVaqnSLUijNZ+EV1UMtOJiWU
0qhHnnIYf/Pys6UDxm2kxL/qG7DMBbm0kVNiPduIQIfHLl8rLJfJTU9e1wkONTXv
Cya9TNR66pCFVlmdWyRygUBOi0Onqm91g+gBBJAj6AQ3LCSzL6iHslmyZm4tTnPl
hqlxdT+voDeS9SdyxTNps4xAJEAtb2eAg02+YXwPPVdPSe3Co5rz+aVACiVm+TzJ
0KUeyV6Hq/Wpd7H4LiYclTlVy1S7Gc77S4qYkVCG+9G7iNY0kEQHR5JTUF1cwRq5
MNwVlBJv2bRJaiH/k+s7LxT0+4uKJ3KgJn54RYfhC9erSwDabgs5hyUlIOUh3x1F
dngb25j4l6aUG3wOelthFPf1ZKQwzE+IAe60/NVRKq7R0Ka87/5E5uRZBiovDteg
/8do/ZS5UX6jH2H3FIj+1ol+B8n7mKMg4jCGiHs3wE0+N6U1wGmTJBfAj5i2YlLH
3jhIKiOzOM8ZXokhgNdxbeK2VaGmWaavnYQTNih2WwesyjCLnYaUN/So5HLpGrjv
sx9nEEfQyWGC9paGKdA1zIw6wDOOiJszM6fuIMTLDDgqHDOnHfbjrThMVJHXU/NB
J6uxOvdnllDcayPS25o93K+kWtXaazZgaXVabuf36blIQEV+C5aahGLdwi1spwSu
29Amo5NdKmnKJ5Uek3q1Tb39lM7XGJMSeWPzUTm+12Tbhi89D9XBEh41x4Po19Uo
OUZFAiIrsDssAH7ZbrRsDB2B7rbSgKV2D8NHK1d0wxZrN8eziRxGtLzzjXbnkvbC
tmWvn3/Nbx0P10SES4eOA7zJyk1ISOSxQjiJJRfn+13TWdBDFFBqkRO0+R9CgC9f
aArejwytrC4LpYO6X9gshiVm1FKv+aMIHm1axWwPKm25sHnZuCKFbiVCOSCqL+l1
UqelOMQJXCpaiWEpEBoit/mr8ySSkICfS2QGGBOql9GEUIKMEYoxAKy5bt908XSK
64bAlHd4Z0bRgPG0uW1YG3mcWGXDDLT9KafEJW4k1GQYDwZCwBLe+1H5dGWmobDn
pu8f86RsQ/6OItiLezl4hhkIS6OfEnCSSKa+aY0Uz55haOPwHSgVbMG9juf0AB6q
f5u2EgGBKfcPPiozoZ0d2i7/avSDbfIfvFBDIDu6Zeg0ggK0EsZ38gERBa7P/d6b
wB7fMsbdVeyTM3qj4ITK9XwWPssze7Su9Opwibw/qkoPKqejZc0tcGndFD+KcQ+W
6DLWRR5RZ0HgzSLt2UQeiLuRzLz6P02EEiiEudUH0tpfMswDe32/sABsmITr2ppV
3ey0gW65/YCAXDmJ5tI+y85Unv99wUssW3iDuaRkG0Vq6J/d7VqcisY5gBNCIx0u
CrNRyRVBvype8Ofl50ZKbvBhUv3eHSiXLnYDa9ZVZWmnrRSUZ/J0qvhIY8vbavD6
R/Y8YbC5mVT/eBd9MAgZ/p0NwaMZAqGl3e1ydBEYJoucRvgVMuUjv2H02qAeSuoz
Bx0Y7Wa0x3lGAnNUHxTKr13kNC0LramOFIQfk0g4DSKwAaVgXCOZiDdyLCMUrTrl
C3hzjTe+RW9gzfOVCfvE1CFF2WiI1TyGWEl+ZDWlcaF/bctFEJ3zYHODFcfn1DpL
7g2OMCH9PbOQbOA4wZcy8QkPAIdUhwYTgf+0G0b1yl/bTIhvk2XxogCie7+crLrW
khHsqAoTiNTANxszIktPOKCFsAvhqel8IQ9yZmZw1CMe45vQZQjPT8GTyQdWpLWW
Z0sUxIfcA7/QcoughRy8K0mfyWF7PAU4Z66lED2tftZEN14CEayf3O7R+W95SG27
cnv4BtWmdOQOqjmwKOtRQcseeRRiDlaV0n5Q4vnahlDR2FrG0n1Iytg76AwdfoTG
vuumIOuFoTo4hG0W57ux6BwyqsWtG61WTgwqcMBu4WGIgeGEJFTAKeCXMtUuREEQ
VYJ0bD0z1uYNDK7GVwv+wnLMB/lcwCALMQV2h8U4CtrrNbUz/Ubg3JAcAtgQOLzY
8lYXKxIGex3cmrTc/DOEeSJVFUD7h0IC4Mz91moYwduAoAog5NVaxNq3+E8hozeQ
jaH1ZPxSOeysvnsEhgW5ve4XzNTx8srhgxF1f7ZPss84uhVI5MPBVdCOPinujxXE
faZH9vDbTkCLGc+l0/Z8M56F5oG0tm+Hqo9sE2TbuN9jz5CCGqgOJE9tmFdFk8+4
qSme99kE+bZmEioKCG2PQy06otvAeoZLsumHW87t4aE2T9LowiNIdGVIvHJY0XgB
TFb/2uOGORta+An0xLkRl63jvA81ukfwKUw0Vdo4Kt4n9CJoORzPuQZoSoY47sBX
XoYD58+zJGpNm0/eQITJYXZNc/wsEzKeJcXk8CMLLg55kGs/fRFctw8wnjBMQGfd
NfZMfI2Lr+5OCcB0S5i+E3/qxjqRVut5BMMJCg0vJIgF5UmMCylpcLPSB17+Gxxy
40DDYNDCJQgh0BOIAQB3MUkvZbZ9Dzpo08fVkFpn32DifThXEPf+l80IZr4y5kab
Z1NdDiPnXaT5ZlKh1F/c367vcZISubLN35Ee4Qxrcx6G7Q7Bnmzz0SyVtvJh4WwS
H5dhY/WUdqZUAXNwdw2bYjl/NPZmMYMLP2bUIzZb0SEb7W6j3jKVZzzaZ//1EPbx
aDhZAg/K4cVn6l1UnKuTQKC0fqX8Szfpuh4zzY7MBCEsDjdVLzViAmctJ4Vm2LOh
kUtgVuyflFg9zGqoeogCepLJwNeFRpNICU/dRzLEGvS1Qu6A/J+7GfUdr6KjKLYr
z2yQwDBmTBkWKnIDP/QQbGs85JcBt2ntjlxfrragzVWNwO5h+w/D6LqBo4+dqYQZ
3Hq1DOO1zbJ1gN2dG4rA2HhD0klokPCxC0xmko570s2j59XnMzOAA2uHaGpA2Y4S
c+Lbxfi1ddl9+4OiZB/FBjd38/iKrbOJVW1CJcORTli/G3cGYrGRGur5QndVsaJI
806bDd7Zz48CKZPvyA3lUc+x6NxuKBYFK0Ua8lcgzDKi2xtcLrVHeNE296IWTHCm
a4V2H2oK7UaZyja+V4qA6APOEUss5Rafnp23yxS8X0o2qJUbGeNkDz1YUuek+o88
F/4wbkCF+cs/e7tMKPZd1Uo/kDdLD/lehI/Q2veSkLNAxnSyVyDpe4D32uZJbRxV
0jFZC2vjDXzgID/DjA27nWeSifeuMIiRcaaYNf3qRKPHDOKR/ttel8ll3pK3NZmL
kwNICTXLbyShIwNsbZ0HjeSRupP1Mqbcvaw9xZttD1IH9rlKqjbL7LviFshG7lgf
Uf8XiS/r41+5uyGr059LElHB+vmsfKj+ChZEzbVvIXdOkQOLSXD1U8/1ByJ/VkQM
5QWyz54vJ5nufgwoWdwJgLp2irE9KgtZ1L29IOjHD9a/kvhoVbT/L6v/gB6P/hgF
BsWgpKxKHIs+SFzhFXxNky7q82pBrQL3+f6P09pBicS8gcNZPAmW42ggbxUeu15R
1Ahg/yme/hbQa+XzQobHf8ddSkzsxcrIu42Z+PB4LgOIpXHSzRlJE5TtWsdV8WxL
/O2r1zxopaNS7Dvv5gmgsyt97Trj7CWp5hexUdsKy2m9EcQZ6+UBQ6MY9OIuraYE
qfvqMq8exG6UzaDfM8sGzZINVBlt6pQdpiutbJOtXnYptErStzrkOHfM3qjlnswc
Pj9RH8J11PrP3fvyjVOCK2LGOzx2MjF/uvhb28SbUdEW7/hercbRQ5+CRqLPLTvH
YG+sC3uU5GnO+CNXQsgyvVVjqEzGy0lN1OtYfFFhTfGoCZIg5A7ggVeKeSc5F988
xFxdg7JTG4NYzAB8APOPuYr1qI0oQT2b90wZVzzH3oxY+gtXcZJwlNtAOsNl76wi
/7xUfMjp0BwN65GML3+SUwB8Z/1E4U3DHU9EaZu5SpukDzTPAWa/Av/JwCrpNvsX
9R02+4WY23r7A/lXiITRxkqViGnUrgo8C1lUROhdwO9lAqAxuyHtirR5WExWsbIf
oJyryx4v5EAVje2EM6cLcCVxghgujZ2t9d04tag/w5AhRXlv54eObtBaSuMmAqV0
X694f0wC0l13ByXAKWJODkid8kJcOu3oRLl30c2cF6ksHhGRUl6fguDaHYqDKvZM
9DfOf9n9aVNsTPJApEP1eaKItUOF5iVJP0HsIg6lQdl4gXo0ubwnOpDY7l5yBqlg
DW7ka8FJDeNSo+24nLZyXP90VEqmAgXsaYQcKDovU/YMYjT2UyDAz/ABOoXqTw8r
GslxSiMjSCp66c1pYzwja9LkHJKU2u29BxXYTQaMFyDaDpUjCBMb1tjmjxpaUXcN
suCvni/OcQ26v5rSkkF0OeZjnGRD47C/ESwXDMtCP2cPKfePjHlI1OTrxsLPTiDS
bxuNvkviWLJY36LcAEOu1WsxaTF/zDCFL3kAo+6QiG94CqT3UHdndtlbh7Lcs2E/
Oq4vACGIF7HwSSp5G3/UrHhigGKPWC8VsLwXszd7uB9M55dwAN7eh+piEj2Fzu2a
a7iJIV/UMWly18WHOKk/3HugHNVHeszhGPqPWTZRP4EDiGknX1uyUTsyZYVMcxp+
oEK1UJMEQ0FYcx12PVLH5P/0DGuKxUMWUTMjaLTdZBLTQsgom0l3bwlsWbk+AIPa
q5l0K66AUiq5CabII+PkJqzlVEYT43cYNDMfDQ0GkVIFHctQ4RhQaR5eiUtQc+k3
R+UNNw7HACKrRdb68dLT9FVLHZetnxiHTbTjH/1cH1PGdMKRSDhOXdXL7AD/iIyw
3/859Cly495yy/CSuPzOCTHU52napdrlzki8agHdTBDokmhtu888wsm1nDLN5Bgl
6bcKMgzgHJV1w3xdiDmjbjKq6VTvfk2OzDS6qLdoTJmmePtnEv5Iq0waNRd2TAZE
bT+my7l2hWoKAL0QTArJO6caibFubl2q4LOgR93V21bfQQbZx2dU74ZOzqZIPNCY
LbSDUyccxhvjgkUqLIKbTcWxKxRUmKjNkg9RsIGFoE0M0gNibGrr+xBXZw9NpB6L
g7xAHuSjX4GLpUwAZLyzw4YcUJcmSzjSMxYn3wUaBhk033IyKCu18qyd2wAPS/bz
2f15wg0NlK5kmk5jQmhJk+6Nx5QBtEZxBQjgoYkiMBPiUfX4dVzd0L0SB0lqiv5F
sbde1j978QY8YuhCLm+Hse4MDJS/PKQ8Kh5LFsfzKCTBPoc1csVJWvtyE/TiKF3u
ZAUCfEHHF/C/UvF5Sgsh5TVnPAW0yqxA6jGBpBif2WeK6Z12+JvWAo1I2vFDZu2i
XPTh5FtOoJ7c1Ow9tSupJ8mUiK+2VUoS0w066I1akZJmX6H9LZwjrS4UlyNUZNfj
hHkJw9e5hluyuQHcHSS5gv9i67R5lfuGpP76t7dKFTVYKOaOrL25Y3M8NkdvmB4e
vqUO0WLJ17wMvhwUtBLJwerjo7YQ4AnhSDoXl/r/BFJ3ZMq67fa47hta2Mhin8B4
+F9MQHzoshZ7s1oVrw6FQ1/oweWxHDIa6WVW4zqPSiwHj//6pcBV4Yp0s1vsXIaV
mfszeVQHday+jDToKmyt5+tyimVNLmsG8oa2RaW8OIOmf+7vG4iNaTbOI/83r64P
hBCaj3Zaw68UsNm52Uuqw8UM3SMvwaBeXQJdn+inuDruNtwzGWbDe/z3cUEYtIku
R1Htn1dd0dRab6qe8g25hTXGv0S2n34eKvGV3D/ik+53h9e+Lp1ot1CIlbp34vs9
BQZhCCkTHPZcvklKxgc2jRpa1su80Vnx9/YomTLnj1DOmwCmXRpiBNawaxG6j7K7
I1bEWD/Rqr8Ri/sPXe7Zd3wf7r/WyO8q02u8+QznLmrAMAJqjQhMOV0LV6kXXnDY
lJ8GMLtHqFytnNV1cGKXvNPAh/IVD61zYWgSpKaN/ULkEvEJPWOfuGW8Z7LJTqOA
ZqrBcAIzEJvQM/qyq/g21TW+b0rRhNmteEtrbOhpCsaP3qiJm1fVjpKvehcjCx8d
kG52kSN0ujAOgKAWy2K79BjjHasNBqXb9zTqaJ30DVVD5jqqUEajck6KOHS1fma2
cL7OBswkbR6Lv5w8cgvxRYsOvonYxsoBSFOY7GCasYf9nKnjca49F0Na31bUyXtJ
03RyyrO5q1MjJTflxOusNmidhx8O7gv5sTpWlYC6ta7BSt6leN1Sfb9OdRfTzDZa
b7uAERwPkrNrwKyuM91+9iS3crJcfUXMbMdHk4iF3Wz1S5GiMOKGqe0QQU71Ps/7
S1ZaSiIm9uQu3N9h9n2zlB4nCozd+pIrDSlAuWHfbBAwe+Ee81YjWU4HaMCs1VCu
F/fBjDh3H/ShddD2o5Fs5k1CobJRtNBYIX3U8WQ1DF3qvh2ZXdtvcfwsIE6g3KRv
UJHyPK8gWO90QiIfJNZBbigfRYcPA2b6w/7oK4fLSqzsjl/FmiCpdt2oYOQ1zpMR
ceP5g9opXbhdka2RPX14SLfz4uJ82ABDssV9oMARL3eLPkHTScsdT29VnBQfRCQF
AYefX5Akh8v3Voy79t9Vdmo8NRdxdyieIsnkRtXsuiiv8KCKJEB9/OmfJgsRaySM
EF0icRS6SitUaIwRXIngSfmaDtWyi5Ag4aNrild5Lq0VlUXC/zisNUcSfofVbR+N
iiT2/u29vODvzgPZo+kVqTUQEfHr73UUyc5lBW+dnonl2+KfUYGkI+oLDqxheRS3
96ZsnLN8nTX4LPoGmGWwaVyz5DA98lqMXjzg9QI0qEZFybnY3VPl0xiD1TUmSpi/
nEEpa92CxK3kx7H91dQugeub3o3yoPpgiZElRZYgOpgLMGhmV9YMpdXHGy5p+Zwx
DJcdgBZvGmNYLwMyfeSbMVEhkIWMZS8Ssbianhgk467XVxZ7xcO7UoHRCA8c9xhc
EAYXD38z5833Gf1TJ8T1kOi4yOEj7GezMKyMjgQVLUWSS/KP/dF9Q+qYk9Jzd7s2
titMFv/Ty75YBf4x2nw4aqgtGLiIbOx0rWJsYWeWeztJZpEzzSx8HJeFuqCxP2Nv
GEEee5bCJmy4tvQ+T+YZaHlQ5dcgQ/HRYFwWCsncB8dyEDOwkqrCtIOZadaFqVFu
QkYMbRVQfPF8TGX36hdWFGDno5ncYqoVkScnbhKfZaLcCskIgcFJXgD6znxVTRm8
y7jJPlHm7xyPtrGekYooVzRbjiw+THYrcMFlEY9fiOalFIdgzsTSw+fD2zctC4ig
/qbfbsjr7SAn+l1GpJxKVgFG1WTKS+i9HdG8sDsICUVv4ACPzf6i0eizFXPZlQlM
RU2c6EanFzjZNi34XgLgyV4Gy4UMxCXcQMqMsSOmzNlCaYxo+2iRuiYCjl+jF1t7
hMYseEP6mC3zsMR0rzTxsZpGSO3ZKs10oqTCfsdmN8iGTg04beTUIXEjJbSQmahX
uG1hVzIlHDbyVy1a9qQp7+fUC26/Kryl77LneQwfQDy7JMSO63LM3GXBmtldIIC1
nCdadtOeIBXwMZRZYa5Poys8ul+uWfsxrPz85sVJzCGKmgTu87WDtpK+HGeVeCkB
Skt60+c5bg9UL0a+emXtRGiaURhXm3MofQ7ERurPpZZg+XnkRiccSGXDHjqXINSj
aSE4vFUwANUgyIxe3xUWASjHm9Y8rzBXcMTq4pJLjBzSQDf/W9mcusFi3dyOIgjT
0aiEfhmWcywDDAtblHzDzJ10GCiEi5OVQBOEHbmtu4qvUOu9XBtjacoxGLG7oE0N
6/iJZrebQXNmO8axB9/RZS0gOJo2opwmjFfHSIyve2w352H6sCpeHKNjeBvVwMHh
Q0YgJXLGL3MT07hTGeJP1dhgcBDGUTFv2VIZYapRbO0Xoi96iaGYskHSYfAwZxse
rP0bfV0Ewne3XNgvM4TEokJMe2saDTwr8H/rcJW86zmouwdKx2TXXzYyr4D8X6cu
25E6rQAf+kWq88XDYiIyunIYADdjyr6TQoxm90mO5a1ojJaavhSTxQdwQUU7eQ27
jl5+1V9/iEq64FMO/7X0EjeIyL+6unQWNKZ0fvAAFhOnqh6Al2x5yB8xxYQtkamt
QRnik0KX8ULI8P82bft+Pb1mbev86Ra7JAHOfEU3+Z10LdiepOhilJ7k8c6Zf/9F
S0KzwhlYRPnpenQ42ckLxpkErwrBhW64cQW7vP7qO4zTS+u2XqfpzDx/Jz5JrwJb
Z4e7NnJnwXhqt3IuvBZLLxU4J96Ns/z49dq78owZAd6aH+wnv0Hcz1nn8HFUWsWi
rIFRmBfIom3ST4/aab/LjUFvoEP2bCUwndr2KPvPaTH+zFhWM8TqN2HrhAyLE8t9
8KtYHXDNVqSvsbML8jI3/4yj+3Sn1FuY2dJHH9o6IFRVuFF6S5LcXGkcluOhNh1K
aP4Hzl4D0XmnI/5XfGQXBh6juVCcSp2O/JBjtoO5tg4Yt3pXKk5lQCFLHqcSVAL7
enZtT8ndOOe6BeAQ/qE7LeN/TQMAnmBdBTWACEy1gHapgHuH1SGxM5/W+NAfzoNr
YO4qJ72ceH5uck6AA/2AiCj5BCFPuPYSHpxdDudVPq7KSBvl3+TP0oCZLQt/IdC/
BlVwN432Givr8mGILleGaqDndLC0I++kLwIqti351KeWfCIyBMchjmv5RVyHTcB4
bTOV4FQBWWOSxuwhlsdDfsegGFZR7P0pfh0RLVtG5LUXxSvvnX17kSDufsFLWIoX
VkgG2VFqswOA8mzSJ/JlOhPknDlILaJ1UoVnHSHfEG34QqR8dk3aAtluZgZsEGoQ
22+vHIG7g4lOdmgY3mMD1Roiw91UOWfSEZ3hanS5/tzpR+D1XnjueTB1g2r8rSuE
zi5CvDSLJnaaLTttWQgcMyfRA48PzviI20VYJyCPN0BC77tWRiLU3APVugZt7Yp0
VBrncxAe0esRJu5DORrrRqZ59QAqhE0Qdr8HSGzs3vDCGoKftaG+JjU3SVhvI5jd
Mr7SMv4+gMhG7PYioDA2dDLKykifECiXIs+7CdyAYwHoOhT0IjalZfafZ9D8px1n
30bAs/EuO8gzxOIN4buvRkecmjC/EuYz5TP9IxG74GicKZghRpkPVGK1k+3lRffL
qDUvpn7zeRt6gmqE0yEzUT0V7mde5j7Vs+7zQQbKynzB1N2GIPwAnHTRCeqy2P3M
5svCiojojYlvAetdikmFgNCFMWUJ0M1HwuiUrtjTCl5gzv7TLT/vEPuGPZOuccms
RW1E/f7May2qKID24cqCz9oOWtCcAJIL51FTtds6nsaf3XSgUG452/3yph0McMRN
06Xi7SyHp0VPmbOsfqyrOUjykdWQDNn+U4cadvPylYny/Y6QGHkYQ12w41hAWaV/
jdtL0dNcJrRC9fq3KPYCjPFIcN8mlS/nMp+KswPWRwkTle6QrAaAfl2VzZbakasS
rZqHa4M4IIUTWWSsyr318qnxLUh2KETUgxyl6mBdbZmSeLQhAq83rCP7pfDNiSwn
uVqZoQYcFs7TUjOCAIRLxFXHNUtnA3h4zxqH4EkwNtFxzmdjz9eDB+k9iLhkzCEV
cWrtlo6UDHzDo8HBtGVg9cyIVdddtW1OMP1touqUQuQlnZL1vLfiQ5Ag/67XA3VW
2BXJpVxrBH4TSA3vRrgPmG9ZlK3Z4bI+1E0molttCKZDxf47B8rvlajhteCc4zsU
7TJ3G/8t7aK349kmYx8g3AJCyCnK1EDhkKInYNuam8ZfIGLngq24og2NeEEbetxR
qM3hx4xSLePd8yjoxPUyNTJ5ZZf4yPLHJdCuEIKyqKzMJqLtrNc8kf039G0N++CT
/XM+26+IeeGNw+IEp5R8yYIGvDhSn2OIMOwKLrlKqzoOfc/WWtSVl8nbd6jtf1mh
dgJm7Frc6DCbK8PER+FEg8wlLBOIWY+Gsrowuv//WkPEL4l94q4zpQDGkIgYX6DH
JdIWLUynhMk0801t/J6JdZnhNx2L2kpnUzR68R493+zpEoC5HbyiP2KBxZUEw/W7
NziolwHLJrK5QqfJXh7yAl+1HwkQvIOYRq1i2vz18zSe6zTmIl27GBaE0xwh3rMM
b/3w6Xlm9HJCukI1xQ4SYdCEuxeNC8QfZUr9DLW3n8tV/z5O/f9EjL0UKYg0BLkj
Jxt0nhRL00uUGeTsJbP6HxrFwzGsTvBWnuU8rVvB9ODHPcAo6L/IJXM6STpEsmm5
kIPvqtfIDchjIgZIP+VvFggnBp7AgYHNctpbODGRdZBQe/0ULJqyW/ndCCyiaN19
itsc9fO48GzOC3ut5C7psZGKFU0tGZq8C0Eth82geU1EXLHrtgwNF636fGB1htz6
JowM0hYS4cEhHEskAwKrCxq99rziDiHvbxB1D5xj/sDZDkT0tK+yviwoZlH9b/yQ
r+6PFTXiU9ATykPMd29euxHrN7C5wTLUdTmkPczUVxrgr37JUtUFZIPRi++rM8Xf
qLJVnyWrE1hUi19TmqDaSIQNL8D5dW2owfY+6m1OUN56vLzQjA9v2/HCvvnD3cZz
dgwfNb9A9it8lhfkVmhrVL93SYynYQYoJPh6KT7yeeIojxGGA5Yua5d62q/JV2zB
v+5gv7iTdkjRI9rR0JeilT6DjFpNj4IZBMrS0f2op45haDdPdU7yW+d2s4VntfB7
fhIpFbvXIx3b/pHnMgzUMnNAOdf/0Ck45+/yX6LF22hBjTWtzFFEGckXLt40Ome7
uh7FdBbL+ehSqGZLouQtS0Jg8I6o68e9nfUZkznkowScR2brKRU79enDoIRC4Y35
Bp+iAkUCbXDvY53xJzz6DQEfBGuMazVURnkmZx87UEi6mWHMb7g1FtV0Lp2XZSid
PDJ/3ZMsSRfQdrdzdeLqUBck8hfNl5DebO5tLG39U/XObXbL+tmK3L/2pb6a1LZL
oPZNw/Q8o9X9uj75sAKHSSoPJz+ftWWb/657rSbnRcPTjrvEbOQ1fpIyvkBGN9jS
xuciHybmyL+7teEEpBzkxFybc4p0C3YIsKicyjtWG00BM2N8U3rN+QjsF1dYNbyH
4JmD3EUXiTCAR40x43hWM1mWoK3Xzr5G0Fg+1hx1xJgzlldKlCjzeZdLbduoxuXo
/MyKFi9Fu92gQ5+HdztREE3skKgNQSPLrR9SxbckoTJDDN9B4ufHs9nuCsOydQXT
sadl/tRDDJaOTiVZQRLJkruQMTMFuG71k/nRJPos7YNnfTKQkBA1rV8VUDv7L0ge
qyfL9yHSgKxoMswur+4FZGC2XDbo/sySgUHugOIjcEEbMWY7H3keBvZZRiOvsQtf
Ln7J7APamnDicRWPh7/WDX0CYjBu0c9x+ShXyIMYKQ2CaTbiajVq1fsw08uaWUxc
GWo2APu+AjeiD5yCkgvtCW0547MIlclfF5dLwlEUUOYbMaxPtyxwmCGSpdy1qrYD
d9Y15MPOeL3Avyy1pU2J8SLIQ2WBN0uJYuSZR+wgaSAP3J9uvrvmvCIpp0ajg+og
yS3zTQsc5LpgS6r7ymEF5x00zEROqOF983jEilD7tB+jyLHHKySlV12e2eb+HilP
/DHI2vvVcCyf2c9fr94JQNmSkwDgxB9cOUoLQoI80Dk02PGywLqSx/kcxwBcXcrW
09Iz6bjL2zw979o5imtjjIVnjXcOVoaPh1XX89spbEuSl63Rod3YiB0dSWaw/kRO
LOai5zT8GlNaM/pI5NEojmgowrdXIGGAI0YpC/aznooYrHK/y4vlX4omEFx4JBa6
oH1Kgnt/BfBvunt0LywiQjee9kfxCvdIbl2afTX46zA3UVaW0nBxv+Ey91rOZHGa
j0sNwl2gjR2TzQt8a9c+6YCAiy+L1RYiZXuG0XqlQFwwPmVfRRtMrOjXN7FrM/VY
r0ogTxxhF5jw00U1gWNY7gPNSg4bg3lufK0WDeRMImABIGh7SzzGUywTZKxCVI5t
ZPWAf+ROjby9LiMwcKCfN8/tLrGdaGAeWHGlWtXIt8BVDVwgp+ngRp7VdlGbTjSp
A9Z5Ooi/sHyc0IOv9XKVIdaXyS2igGFc+Ev6Sq2ycW0KfTjkD+QFN3bSR4U3Ua3O
uPrrGelLvIOAHsEMFvq742L1fQ96q56fKTN6UfA8r460lAOKV3tV4b4nX3sQuoQC
TWSPoTauTINsK2ph4FsGMZBm6uvw+SGagieJY0UHcNKrIwSRT6gnBGqQLeMdhafR
6st0G5jGKkcMky23k2Jp7ZYWGd8cVtL6VPCLVYspXmUEm0wEntcGnlNVzc7SjS2J
kz9ooF2iaCHxpC0xJUfYCG5DHRTn/mwe6oFL/+bxBJ19bu+W9oDZqweTb+02yJ4f
SLPrVf1AxW7jmjC6+8vGipnd7mKgx5iw9OWDugYvy0uaPxcOv71MzEUkpFaioI3X
AMmexqS+13lKZeRJM4UNmlcj9PB+C4hPG8HPsOUqwdG6CSA7mgb/Bt77su3Stoq1
E91r0mISoFubFYECq4ABcsH4avbzXPfTR3nNskGi0NhEBaT3L6TrBejJlhSdJ7cs
ZP1oS5ja6Fwan4JvqZSYSIzTL7gus8XGSXF8OzZgdu2Q3LMiJC6VgqdMkeF1LqRZ
1j3LyzacELnFWNW89P4k5RhfrlGYnRZ4hT91yiUo7bqpf+cOobdeYalIF5JtiiQl
gfxOcTPZ9Z4WZHKZaoqCDqSQDY/QDGH72kqZWXjRhfs+AMLHFScLxHi9QI0Opva3
l9Kzs4VcmK5C0ZBDt+qmkSArGJVc+F2sH2fpS8aS4fpcg8jAqYYx//Ur1Ud1Dzgv
+KqkTnecVWQF4dW+CCPrXVmc/xEW8PkuXomRBKQSoWhbnDwkv36Uj3fNmOgKjqSi
4nEJZExzRvWxSa+huAHUCPQqyw59YA3GL5eAIql9RCvViwRjqp5JIalz3sOTTp1e
PRttndU6+5Pohg6HS6XKHDZKYe/QAOQrMICk0j9U8xAnjBrntFqpSAOiBiucvY+a
Fea3CYJWuj+aN6FEb4RTt9evL/t7+VBLKN8pqFV6DewZmvJFHpgmRBzGu7uUci70
wh1NXQlHkZRoZqaN+x4Adcf7+FyMkFJNSKGSyB385sBzn/mVvoEdiJ8F3dfc7fny
TunJOfs7Tc7LQiHuF8EhYOUQqvJFfQGUaJn/6bu9KNqKYoMNrCIyk6hauazZd5mF
lVeSVWp5MlEq4F5hVwZaNm3wRFOeKLrEqH/bFdRhQbod31k0abc3XTTjY7Le+2WR
gVFvGufYukPDpiXpDART359TLoPD9CGWNtXqWJ5C34aHN3YfX9YqA4KmK9iuFFVz
9MgBu7VQ6ZpTQZC3x8oGyeFX57xW1DtOqc7L4vjSY8/UI+lDfZKlLRzYEBl3z6oK
8kn4u+iQHW4jpQN03+aCb7pQ8RYQQ9aNT8zM1Ag7oBZk7a0PjCVJ+1QEPVbakf76
6XHqw5E+KK6gpiFHRuRaEhzYqTV9OdpN33/kRab7CnG1HH2vmhZ3zjqFg/07czr/
Z/CDwyIyv60YqczCegdxLpCoeJSh/x4VTfUqOnzT4g4r/kDJqIpVAy608KxP8Ut9
GP34HEPvxxOUNAVRUeGL3mge2yURhRH/0nzBcOWR2was3CPu8afBQgnAn8llYiaD
OMgyuIKvQHyaVf5ot7ebAMCHnzqQ7l07mwckVHnXYiVBeL9YUydjtPE7EPlDSp9A
KEgla+M7WBv0f8z4X/wuuOs9iUXj59flLif0Sv9Ft4iOHOuPK0t0I5i4UKS0BqVt
enmImM6X3yr9ntpVFLe8DAjRz+gd676MkwN/e1Unt4eUd7ZdofAqkEpJr53cYcoT
3AnB6FjOMGAJjPIjRb+RWa0Lz3KMC24sl3vCFPC1sgeXt2xZ7fwVGNEiPp4MqPHK
jAc4eXW13cfcN/0yPh2JJ8DULsx3S/6Fyc1ZNw/ONWzgmZlCwwZNv8P51eDA3Run
qKyuHHOhkphV1hM+MpQ5sTHpGRcuNvJ4CENXl1+Aeeaq30Dw6ud3EvyLyAbRvUR/
ebxTx6nLRf+3zr1s0DY89yF3cSEKilVgfRxkY6c38z4K/7tjBI7jfSdozzKhw087
VN1WAk40yCIMw4FWFFkZWDp2HA8NceSyRni+hUWO+XXMlaoIC8G1OwkQ5+8azAyp
LUQ9pMjXPOA7ENMS+zDryc9YD0pYZ2muy4eIpAi74/ZCs0RuMJp1xu6UrDF33NLO
uyms3vx7eAVks1szIQ1ppF5Heh2Fjv2iPf+BySbiZMriTNPiKywvN4Am/aMIpfMa
A1V+aRggAzFTjTKmnHosszA+Z2gi+ak2ZwAqEMC9zzTliyv14w3KNKiLqTe5+Kzo
YJ++d8Rsn6Xr2ia+4abY9O3ZzmLz2K+YEOmdQsQbVp7YPQxG82KY1UE8qdzYiqNb
BubNxFYGe9FgIKBM/6NdDAUy0iDJooKXbbg8jD6gItXzcxNzb4WsXBFafJM+cW7l
yosELahOhRSgLmqskjZVZweWpWmATkz63Nwk810hkb0VdLfdia9oY8nmYZPQ0JjT
n0sN8VlVkwfwyc7wDMU11Yhc29hvqjVNt/Rv8F7f3sX5TJt4JfX0kemYLwr/GD1E
usFUkJmiIHlL3nnGTe2XioZEdkH+6bNgnn5Z/7q2OoNJnH9TI2B96zgzywneGeo5
Q0FOd93U1cfdV3wQDdy+AbvxsRCXZoc0bRtEwlP50OaGSVoGhSmMcEDtPnI/CEoL
bghTTJLcN79hjtbaF19TVrY/CtY7cQF/zIx1tGGlmCFEQTE9QwYu4LTfYe23nZky
bIaTvDrFq2qGNIP501rJDkQ4eh9/E4bikQRC2KjfMsXAbSu8z4+iWT9sZvn2lW37
fKNgXcj7jFMkYJb7SkzSNVdbe3NRASIA3/STBSeE4fNi1MmD4VFAzXjbKjvA399D
83lm73rNR2bxN4a6Xvx7ZchSE4krxEsrPhVVH+HIKw4MCe1BmNc7ViA+jnxU3EDp
Oa/cuCcNiJnAtGAeAXCHQEIRJWykY9Q1YPb1WyGqUlC9npAQOmyx9c62uNoOOjhS
zGfWvaQqE/iBTgs0aDoGU9v7JMjfKOW75iN1kphoiH0ZfHfOWDHH6pmYS/h9vl56
yH/e2kiYcHgvnHSlKqeKv7rrQMTsI6sycwLjGW5jupvVsVpafmu4C/QAcCHqG8MH
JRzpQYTWIFLdVN3Mvo0QqNyiMzj5BZqSIgzFgxmvk1LXC0uokqs4URAafBX390fO
oDaiSS/o+It/CBpdjlVOT2ytG3CSV8qV9gutHQDT4NlLKF0UfqmDyl1tuuu9pKKD
Et3r4DECheHikF/gCNV3E+5jNrySvhC4+2321M7uVKMjFgCLjPA5Sy6tBF6LeoCK
HK6YPwGMMDftxnGNY6AByFRYsKHwRukpSrcJmhmxlmmy6RSyIFjVum89WFfHCWTr
4/Ei5fp1zCy1ZmwL20QTdRjTdK8qCNz72jCpm8S1xJ32YcnD+4pJhFdq4rX6eSPy
hvjugfekabSgJosRlySXN7LvZjmYKF+VhTIsLFNwnwEf9EEvKaIxo+UuCu4vqGyE
hVT79DwLZpQD8e67EAfphiyG7+ihfOS+0p8UOeDwlppVZwC7+FqNasyIZ7ik3kTQ
YqUPE0h07795XGDfvp2R19dwZIeZdVahQUvzmo1EteqdYwBZD2Cil/4E3pyIGNaA
JsomoaGciQaqQKhWJMqzuH+JYtqTFNeM2hW8iOtrevBRMyc3r7nqPoID35ynquUY
imettl2Bkr+U+pnYxTctNSt7ZukmPPn6XFKJCxASKSXyNQD0m2kZYkQdAx9AqJoT
LH2paUVexWTc7c2DuJxWJ5UQ0rXBKyxL7RLeaRnku7X7OUunNZG/bX5wEQapXPs+
iGwauULc2g6Ains0Gl6Wz+hwoYaR77vmNl9Sn+NoouZbz17yupOeg4wIg/OWenea
z2KmMa9vk+3OYeEEBL2h8aMULR8PzFTn9YLU6jBKEXm42oCwbZFVZAeaCB73qSDc
ba+xpdks4skxSIR1AaBYiEl5tPSh5zf4Ji+BhaMVOwA3xudtbQv0Ar2BT4t5CtZV
glBeecS+2oXZ7H/cQnN5Icv/fsD3fO7RJfT+I5VSExu8QKm7Pql2JXDdy3JMaVZo
gsWOtRfRHYnSd0c5NWzYKb4vpLlKdTj1/cJbdEtW0jlO5cXPkIPHQyZnro6okMMD
8av2OQsJly/O6IKpx5iPbT2Eu4QRmBiwE1S6CSOChGdne45zLpEng82wgk4OaX5u
SE+M01H/XeZI4+QFvl5GDEfHCb6Cj/CBJxNciH35Vmys5EVE+KFUF1wxKlzOHOiK
HLvyociykG1yZq6O3h2BaApEWuh0SeigGyTtE34xMKoILUjoMwHdQXJOPH2RO1VK
L81iv9P3mulXfy+u9VvsyYTxQS+YgOdwHh8PimXT8AUCY4Z9pCxAesz7BWRgmuAA
nNnyYK0icGcrso53OeTiTav2/hx4vLUVDWRXE89UkPOk6GsTOwis7RsOWCxo7UsH
RMPJIHpaEoCyTLCb7R9NgRjtePd2v/u8Y3mH9cK54LVEvU6NudMZno+Bv1oXs6VT
Cq37h4vZLWcZ0qZYWAJP/9+j4Uoe75lVT8Z0cc+dzKl5qtdaGlfwUSaNDEn61LhE
St3zSFrthFEbKEWyu10YjnsgtF5Dbg/OPxwVa5+eWxIQ8cXJir7cFJQVVesj+E/n
9+NSo+2/9JHd2GP7ONsk4RiDiV4kCAsnXQjl+VbBfb5xHfXbmXgM06jSaqMSNLCK
1rcMMO01tQlStIN+q1tXKeUNt0TySlp9cKVX2t88BMEtXufDk8o551JLen1pmEFT
IVOdao7cVd2yk5As9iASZ7i/pjm1pqemEniIwsW6Uy4nT9HH/dglmkK5wicn5QB8
TSZ2judiDxGubkAyT6bVzKIItlOk76T42MQWa/Zrj7rbr7dVhcC/2GrEIPr4Gh2K
REDrvELOYQuh3hk5XPLe9QV2fzwm/W++9LEtHRbGtVorIvRjpbdb2i1bQHGAMtvk
ZKKABRLuTebG0sBv+zEdWfKHSqsb1Z4pjVH7lrzYeKJ/oCozn/8QVpDoLir8BbKS
ZEYREUiS4ehxjzN3dQTOBIwNFkJyMDRk6t35Kf2C0yeif8+S95ZNycqFp3Xyo/S4
NoutEFdKxJHOBm4PLQBnxWQKHSV+HFnzKphU70Hz19mo2wmtveLu7tvRjAyOjKwO
uymgxuz09tmytw/GMojTqQ3yWhk1W/9dhbXQvZA22MHWuJUvoZ4CZE0QFFUqH9DI
NaBMzwPUsw9oQVSRBQLWaWkMRXJ0ngWPI31TRMdNqXNa48AsvKZgPy8bKo31OiVc
94adLgDa40c7fqhW8+XhRMHX59WMglEFqMQPRAc9c4jIltlc/+kp//HjuQLYB9Ch
mY76Ui01oNSPaUXASNQkaPvvRE68FTA5uf5g7wVB/bxs1DrnJlNX73XPiqJPPGBR
zi4+xvwEgIUuudeuTl6tHlthUkTcfTJVkalYAXxG/Zf9h1FyLB2LSzAdmBL+8dzv
RStFT1EhdwtQvorV8dzorwQTqOd0R5KYb4O+lRxYIOALGDiFhJRBjlyRfo1B4ieV
EwAza7EIHtTph5ueZP51InulcOtzvL72wb6BlVfHTBnbAxVfqQFiVAOKryN5hyxH
B+4Uks7XA6fcPyxuqs8eJ1f7+6TCeovlLDKKO2tpzdv69NXi6BXi2bQiqZ8IC6vL
mnjMk8pAMV56T5qnJIs03D5sKZ0hzkjyoNdPHCveXsHVcue6aCbTcUrbWEd6xgJW
6iAcrHAaQH2lLK1jAhbL2bcjvEj4DqVVognHmUjiurnFjm7bQI5lsleXnnvPFad0
mqf4tH9yT2YyACEYTnRVQZ7lApLHBSTTO9NzElukz7kEXBy57UKOh45NPOnnYzfa
CoJsB0uT+jsWsTU6kgrmXMVi6alK+xZb8bDLSNpctoP8/TKVZpN2OdLLv4KoIq5l
uFAjqDDtBtQ9ia0ezHcw7jIjp5GpK0p4jCwuGE3MJ9VCHUO9lYP+pMtRJOWn3PSB
iQAULE+BEnTUBhm4qTfupNPmlk0yLb9cAWqxZLi8xA1d4vy8GVyF1SfcacofMkdI
/Qi8GEUwdBraFnJ+QrGrqfM5Tuns8FUVIHzNqsUeFAn9w0U+tUH1OSz0MuK/b9gs
suRPBY+2MO/Zf39SilX1LP176/yRfKwNmXnmGisReJkAXmApgwlPJ3EtdlF1p+Kl
PD4e1KgqQcaxNeKOXKBy536ZU/de76Uw7E0tdsGzT0ErUzanG3sSlVL4o384i/qw
TzwjpewBkHl6XS3P/+T57Y/q7fqQeRQ6WjGksqy6s6nLW4oSHM+jI9atkLWFlP33
oxXY59yrYFi0xEHQfg5J+lFfK4gJkwRKYctAMqmsonw4WryZ6L6LrL1zHBgCkm84
Jld9zv6DExKXCR4cKtbGy+j05RUnkaXBMhQiD6zETHoj9BhDK9ezb577KnH2Whmp
4MNGrMBmbV9ui+xZvxSfNtpi1OL+mqVOOaPjc8e11abPjDPEUUh9kY6qSaEBq/QL
MG553lzGZlmF+3e176H9FDBjE0Ch3iopCdmkkwtQZTkbo++vXCDRVCv1KLbXD8yR
wvXk+LANH+tsC/82J6BMAcAuZ7KZoxiN+ZSGEFJ6IuXVJiFNr6/6P1YfPDp7/iq3
kSXyz2Bhvp0YTOaPHx5dvEQ1kDv+ZOpluWLNyC4/sATOxfjPumFn9QK+tYBbETj1
jD+BPhJlLZFz8uhjr4TuG7GUeR3SDZevsnzLaERpdfKy8KIgjZZ9m8w5nTZnsXmK
2GHm337AUONpyNCDLP3Y4EsFXFJERrbqjbd2vHMuBKuPhhAZC+3u0LkYIDTLPAj6
TFmeRMJ3g2kyJXEi5MMlMUqzg84BH3fJ99BMzzmqybSORVk9Nto3Ni8ah4OvBDVo
F0/C4e7O49LPiF5ZztP5Cx7ZyIDS9wAExLBfABU8n1HlDAfTP7wNcO7Ik4ero+nt
FUPFLNYqQLNDdXJqejvBwnTFJSjzDKbUvCkl9bFEuUJyAC74H7zA8LxQygasB3ED
hLOvzUR2acKb+SSLCg6lmVGoJyOeI27ZAIJz9lbJ2Ld9iBPKrOshHUySoRe0n8Hf
lbVDk7uoXCEf3kJd27bFbL4KCabzSA6t1Cynqlmj3va0UJ0iIZjIIXiu5YHR9cir
LQU85Nlh0hmOHkEjMFuAFVg6YS4ssgxbd0aFLriF2GNDJn/ZDRZSUQLu6zgyjizS
Uz9ADv9Xw7qAeAq1XlFYVG7N4qTPtzb/mkwgf0ZvX2HXY62d7vARqP7bWAHWOBeU
A3U41QUDOqM97nWzAzek/YFMrD481Qm1QUbcdyxfwdAsm9BCXXO8rAxNFj3evklc
Ry5g0Znz5uhCB3j85wNdYI+2tDdAc7aM86f7ZA4Zr7Cvtbm9LGiqLYZHGt0qvwSW
Ga+yaTJzbc4YkTZnqDcI3a6ZjydzXFxeJMHPq0iTFjZFf+m3t5fuiRGgGsluNbCs
OP0rJ3c3nQ9Bs2BBCcWnTvrHAqR6DfDqCWkobekIalFIYRHlnEEDghpnTwcOhQsx
SzTJQmBHh+lL0YgV3Y3gIwhH7cFcB9CoOUxvzQTVeGN7HhkdtmlKz5i9y7N3w60N
eH+7i6PPqE1OVE3bvf0YV3B/z5wR0p6ovy8GkUnNDTeWXnCxfaVjVmNqAGOchViV
7jk2cCPo06d4aOYF9O3E75QaTJ7fRt91yxYyY/BG7dl5hunhCer0dgNB0hkA0PYr
fu788aHnbhPgQ06sSrd0wW20biOsJERKinCDaeqkTuF0FzF2PygrkWrI78VQjjx/
MdftvufRgrWvvtfjas/mYDqeiusgWDPwV6uIBw6FV5TzF7gq+t8Z3kiyDo4VGwcg
Pif/1mZV3twFn/f8QNBRgrIyw+PRL8LnwNS7yXaOC0IhEC97ttNXs1pGB33z85G+
240qmZX0QKwBwH4Dn+aQc2hQaGiMrx8ORbLl/K6TrbD951Elb1ej5ImAFK0u3gPN
WOICAvwSecLkbuKRUvijX+AhHk4CQyzIskOv+DbmLP/0RtD0MuSROzzBeCZy0WEp
cWfS4l5ARKLi3W8x8NDenTRs4GOkYhLFa03MagfLWRRTmIGs4SoQk/tVh1zNeCbq
oldAfeCbuLJ4gSlM9lIjbxT+2Qp41lXTtokA7o0T8h0YumdQEh2T1bx9Kc6jDDFy
3buARMGXcVnr443tgEoW+ka/as24EwbcYZJVXcamDZT5nAe0yu5QlmD5sokvahbu
dzDcgIPLs/kmt3GhH/Eg031K0GtiBJpl1yFEVNnNil+qFH/MrR7df1NER/SWHCSz
uOFc113r5bqU59bd3LFTyIbBKCJnuAEapIq6fyhyOqtRtO+tsHq5G8Dr9yEGGgho
aukE4cwzuRDi+jCurr1lMUoJTjcSaI6mhj3hwUJq3gu0euDcBwSkfhn2fwijBQbD
DrTgLTkXSNckYAQGYWtMkeq4fXPdu3ozR6hvhp3NPLSLBlDPupP8gh0sFPn5sQGt
8ueOmh2RKNqxCWn6Fp+qYHlqDwVJ5mzz4Ip/Kbb+UJI4fLtNCgO+uYjFEjg/npwG
ASK1gs7wVGBtqW+T902OAuYdlNc0cLe6EdhBFcv3n5lIwgBHSSS/zc+X39TNVvBH
QvqZl7bIEv4sfU2fIbvwaYOli0G9mIi2yWWpOeBJEGzohaWj2dw6KBhM7HjYuEQt
JEQeaHdFAJRWglURFPDgDkDu/k/ypGa2OB9plewL9Edre7X6U7MiDJ90OP/85BcB
xHWlR935mVvFWzvhMmh/Rl3xAySUdlIhrmK3+UVGTpYvqb9BzI6RHbLHfWtYXZKF
NUQvbvVUJrQpq7UWXq+5tMla8zaz0pUEr8K3a85cAoimJp5mAZ+DEqblD1bjEeo1
2SXhu/CcwHFZvFm7bQ4ImUh/biVTG242FgKfG2p5X6uM271CMHTrRnJ9EambC0kx
ioL0rLOrv/x/k30yFAL6s634udE1tSkYsMuNPHf24e3HSzzWjFvOenDUBEuTyjLG
bOAQ6OIZxlt9JgfLLpg2cokKemwjeRvsoLIhGyZgf6J+bdRVTFy3P668AfcpvpE+
UWx2Hm+SVpssLePyqcARXkHQ+oXTI9aw+/kMakJmGgbJNIclht8kcwi4LWyVf6Zg
yB2Oncp76Wvs480xjClGUnx7WBJMaHmRo4MtIhKVjwJX7uUZ05R1Fa7sj40Do1U8
povUqKBTrTI3cN3fIZ6glNgngfqekFUiFJBK+NI1wivlIemr5WFRVQI3FyfRLrl0
drl6Dpq0XdXJeXAZKlytq23ST4hxziiUhh4eUBj7DKSqUvtjlR0olnmNpijR+ySi
dG5G6ARUtLnyRjSGSdAd0XgDf0S3Tye3JQiHMuRKfaQ6X9P5+26jiq5nAvf2Y7yy
kaISStyG0qwppMSQUEbSj3Vbw5Zmjw2C/1kAMxEVM/pXvkPEfJL6ZU+1E6/uxTG+
uE6LJEEZqw5w9OU8DooZSQGJ8hCkT1B+0MjOMX/GGr9B6KXXHL692tuw6LRJu++h
BbDlLj8abZqBpsfnuH8WyVnTtslj8rJXvUo0+UMMY2gJ9sQfKEMb19Ddx4vETk05
1mh5HiydpizQ/roZ9m0Y5bMpSbq4NnCYaK0vY+umtSY/HbHzCn/Dvhq0I0IHafOD
8Fz9jLrQifr4y5116on53kQk/v/4cRkMZQoy+039/pN9jLu9FVJYT/U+VWxz1thk
y4NHOYGD4tFrea/IIEnucCB1WGT8V7zZUmUeKEAcg1RRC/Hb2FXtEIFbHdfhZvR5
dHcOVQJEn043KxqCjHc9D1eziRNxawHsx1UeWNJ6qAil5r8WWpm41rWhMwBuHyqc
RSzVBjASy09kuVQncZHHQRIMPSFFMLqnWD8RV/+98oT7c4JAg0KBU7VRuJ7z0+h6
ActKS86jv8FnYabtylWU4LCXl7OWa6hpycafXTkcS67EIPNU/KyKYozcaXlvUGUY
IP2s2Ql0ZmNlggT566JepOb1yGEfUi7AihAdYGj5c5DZHIK99Yx6cy9wXddq4pOf
ECKz6HvWZsvQjkFc4uSVfE/RoGm1wu8DEJp1C/NwHPfLKRzkAM+mAPheyDoz2Epz
MBLU9V4WiMcASAw987WoNX5FIkU3XUcVyMyl6xJu+9ufAXz2NMoOlhiECIcd72nW
zdfeGq+qH95r/nPrG1JxulIYVd1v6S/m8q1rtfI7QrCGZd/NIz7YpPkB0FvHPa25
/rT1pSmGXfGeToWG9FKLFbouV6ZZuM5uqvPqOqlT+u4MsddKf0SkoaQqjiwNNiil
NoO9udml4wU1+9pJd7ML6f81fGf39AwCi7/3x7++0m66Buu70ACC6bA0WMOsAi1c
cqfeqT6m0ipBNPscQxqkkPPP/KoAHlslhePnj6NVpDK4nzwSKgJFh4jXfnZ1BSHm
ht74OrAI5AKUdf5b8VdlgE1bp1YE+UoQE53wS4OFPnfDEiSAWVRGQBYkQdPxxQx5
pqI1O9yfO+cdeVUI3AcgwwvmdfpRHHOsiu2iuUiTFfPUusiUNzC5ZD362MQidNK1
E2F7dRcyJElkJaW5D6lJE1sibfyBdXLxTbSLUR86BV4lhA7x4LHBf7YDT4LcIW/V
2OrSRyOllXvxVyWB3lLRkGietnLMshxm1boBELROw2Q2sI8dQxmFMrppGVzMH69M
2TcTigr8H6EGuQNOoYqQS5aRmwdqafAkkOlLzGtneXGsVVnADzX0aP16Q0I0C7Ri
BKSGJzxjqeL/L5Kakg0SstXthDbM8k1xXcsrTns0nB4BQuydbJIGW9DcnP55jEbn
8QS57HV1uq3aDXGoRYWFuZ2YnLRJVlxlg+nYXfyg2NmgWGsWnRiUIchX2Px6b/Dr
f2rICu9lMRd+kbCtUwn6V9jYUFFYoVYABskM+Z9nQre0y0+c+J2IVFq3qC/QCA6b
cZebKbzLueTupnV57zC3TZ0zrMSG/tejSAUiCZEtC3Y6vt5zGpZkGj69ZqAqkoto
ygi0vdI2Qm/roPt6AEveTEYMceC3Ber8dlT+AOBecmMlGsXLwMI39z6sbJhF9/kw
9sb5a+I7V/ke1Ni+j7wfgopm++jhut+doZus4dqdj9p7lsNULScGs3nVG46xwAW5
98rCWR3QJKPkP4/qtCA2qQ/7HVLGzZrmniF9KHJ1BRdA4v3lp4wFVnvvbaERWgij
mYSAne9FnIoRZ9MHg8K/N6LZ3SFI2tkytAJODswzDunkkHM9zS1s+syXAkaivTua
vPZwx2MUplrtmIvX1KFz+46xWW1gCnaqmRsnFY6+xkR8isPNi6a/TMoqH+gME9E6
eNI1NzWNqOJdcUPW6czOKlbXrcOU+kTaqKEYn2a8e67T5SE1nt/7t7dLLmLh1zO4
EtjceAf42oMao/BFKa+LfXKc9GmnplrSdM0L5WtmY5VjjuigFGLrrX4tPPKA7+ED
pyYQL7KOGgeflsMlDwBEf15WMbjlDZhxX0ZFvUvfA542OVPxb9r9CpkxTmJlj+ta
IT9oxKRHs1DoioJ4H+w2JJt5eOrq24hux8TD8FujXAoFyYs7Surf2J4Pl8+SSq4e
8Y25spH782ZEff5FNpZzI6oWWmbyUXsW99tAa61Yu53GuacGHmqKYoiM31Mvhysa
h8vJ4bdkN7GxIAqYJviEhl4gZYNgjfcVHXvkD5ffSU2lqQWl0AmOQ8AgE8V2R8hS
q/0EMsXD/7MkOC8A4wg+N2X+lfqkcK4MWZfhqf7sDmiDpiY/Jxgf7bUBQnH+BtqJ
9/44IrLC+NOPiiO2faA0CjlT7CZDvUHhUy/e5jcnZJUvSIZlDtuVAKe/pIAq7Chk
eQGDWm5CFS8X2TLq/99MP1ib2cAmDDIv6YcF2k9ypxy1tWMSLMV7ezMQLBjW13BS
bT5fOvIJoHA5/rpdGKXQJxlRxnR1ejyygZzdFCrLAFnlCb45As4nVltPo1ooSok7
nHkSqs4oGs+CGMPuUmMMJ5Dg6k9QlMjAuQWBmZnzpQErEZLhtns1RuXA1LfVQsfv
bXhX8RHxiakohBX4mhPQn6utqybTbMKvr3R43RlrFhGR9yv/xhdk4cXPiRhDPwU3
Bg3ltH81V7onf6UuA5fP/eI81fd6a2h38r9AIVFDDu+24yJuXA/LU3IHz7UUIAUz
vGlJqMmYMWHv/FHaONdeEZzvmaKQcoUCHBTpfJWilycdnmHZPGYPDUm5zMdaG6Oo
ONYnYnlg2K2dJHprfxekWk7oPy/3vde9Td5UvZ85i2cJwgNRwKIch/sAbNyuM67F
oSggIktQzM5nisggJlHRhCDFhvcDGKXm0KXyxpwsCvA+Qieig5PTv9C2jYqPaK3/
eugJcqg7VGX8IV0syW28k6EyjDniC8p3LpQqE8i4kndbVfWiZsa9o49zTcKc957m
XX7be4ZfFDJx9KCiXvkn3b2xGJ9Z6Fp7080Euyi6pMwYDSxCEHya/SsyQpmdlEXe
oZjRQXpovCVnEqL29xPIwkkn0q+x1LJITwudLgEOmQvS9QFGXazbijwFhnGYxmuU
1B4hWaWAhbDB7HeaXR6rnIcAkfmNkBKLQHL29fw7kNU8seSWRnd7i6Aq1HpYtdCV
6NGy3nolDmeilC2WsC6RHvQlxDWYUdgLJbC3xXH9Mhx2nLoWsdsw3ftiVVXuJC9V
EmSap+By5EEvhXFmFR6IJRoOSjy0L1/Oy9tMwWqlkvLbcvLpb7QMzlgIWDqF0MnA
hDm0hVn/Xm/OJUjA4kQJXLzTIhOeXJE7ikXzHKVZ/OhtXAp/XZJ0mNQVabZa9m5+
q+coCd/oSTFubUmEivVIokEd+C/lmgUFGkNQdK/ARmCU13zsg0fM3yZ0+AIbbShY
3LKuWvOimSnR8m9kLnWvIqjagy/DNDyr/OcwmD5G79nEiKQ8dr5z2Q/InCfBD/oQ
VWtCmLdJfEIyE8ZqEDlJlWJT3KNevYetfWfBWAz/f7fzLZ7pn3/BqlmlSWDrArbm
K9OS5+ppIiHqeJVLTz+3ihNU6g0A0CTSkNvQmzA1P+fg7i5c/xDmsxJ8ZpaGM1qq
H5cQ21BqPKVt9ZAvpPav9lodSeUGrWbjx0zMr6qJfwbtSujI1cUKlVRTPxCM55rF
Wid2hp3MgdsWOAOb1CrL14UxvwFpSLrECPKAvOwG4E8WJtu+UEQhqkgojQOwg7H0
7cOAaJ/+oD4w/hfOOJsuZnnKQyTs800D7MWCxW3tQR4ULhS5htMrp+QIIOsb+qwZ
HuXmeyIhJI6GopsXdf4XiSCpOucqY5rIXSyZJwLdRCW8I/2tPHG1DJ1m1TWRhgvA
aALZRaPQIQ8unuB73ppvMtsIKwaimzG/rpQznEFQ/Be+bsYH1OMHyjg+ByYPh8ka
wj2Yv5FGY0DCpzRIZs+uMHNmh2bGDmnqJUsffksbcjT49iT6r8He62D/2RAUxuNM
yM/oGNJVIRq4AZ+t1H4QZcwzA2BUt7PwVsMk4aZxaOreQJNBXLPcnFMVKBoGgnVz
H1Ssno1Zfw2P7IpOgpFUeyND5dAT9d8eOqC6D+51U9YODFfZ12edi8DAaXOjJiBF
uVAb9uzKpKk6I3DR5JIkov/GB4Du85/L54eIIdwnng7apCXiBsjW4e7msN0WKvRz
tEyYyrxsU9NJrujOx9dLNOPkoxHhZKTk1LusustDmaPNQx+6XZpepjekBsu3lOBU
WCy1I9EwhA1pIVzZEGzbx4zozrDRP8l3polE+StcUZdSAPVP6Owws9aCteGYP+TQ
KeAFhYhBpIpFleWLP0CVJa5M9NZhg1EKxbSGjTVke5Sw3nZjLhLP/dDgj+wL9c9A
cd/e5PImHV4kVcH665JkJAP6WaqBLcaI5UFSx0/+lQhotk5MxiU5YgmtlvhhPDGe
Uf9xxkQ2ex3UEmFBG/BV1LrXTLSu6IJ1jgjO5b/Pw1rl+6wVjdfezF/ujriJTpS/
/UmMa9o/WsGzyd5o1lDltCZYX8bFrKDvEtf9ewwAEcC2uSYH4timr57e1OFBWwB3
t5PHh+ox3q7YDdGMyhD93vamZkzvOzOaQNSPctNEK017IPJFuIJqkoNB3TvyVoqV
h2kr5ebSWGEA9EymuULTaRqzl7A+0EeWipoF3BXtcvt8TM0JvlbqNN8ivt+zrycl
H/DHortz2TRvoWXJyRfUVyEFu4n0olFcF7oX+1LMY3ZfUythwTo/+cbYWwK1psfB
VEImgx7uF7krfyEuIsEPzD2FGvPVS0nO7jqWE4X5Ifdqsl3Zuklb/tRzCBJsC/LU
KXqmy7XFbcpLoK4+RSrmS3VM1v3aTek5TdVr1fk4h3Wf6caB2sFKnR8D6Q892zpR
UqQf5/+DXX66J3XZJFiJK8bH+x8vX3oYDHMu2dZ6idpG02XWVLcHvKeD4jU/6n+v
X6VdboS8I6JRUpTW8T2m3qJZYUhdfXS0k2ooDXUrMMdCN7/buslGmFN0rH/f6il8
aSJgQmj/J92/9EaEHatP6RsHqPEPpcDVBsfP5CHRXnd2xNoDERHP4I12/CgK0nDH
SI6A95O02jntN4On0rxVLmLefBUgkg5rZLYJp4i6pBQkfPbWPKGk443eTCle1PtB
r4mHhK28QyoUo530uJQ9e4KZS6NvEYq2i9/cxPJY39CkqX95ivftQZ/MXcnt1oij
reDxpQ1MG9Pz4ZqwliAD+4THluxImDJZyZa+V2DOfm5Ejmb7yT7NFWLwq70dwNFW
viOgTk5vajFChEL/kG/9xEmvI8QtygpTXpKNzkVHI87cRnia4/oh2sPLhXZIqFO/
BbHkmlgz/Ekv9/sgKE68kVXiQWzF3IMDpq3H8xjpjyWUvi4RihOer9NEHrBxVK7Z
GOoDJAPx6WZkGxlZ0VnnYcvubFkcBjdhCgrKEU8wnbOJsS9ZxfwRW42QiqW3DvMh
/Mbu93jruCG/mF0unczYcvCmKKEI8q5SIG2O8bcUEV5lK0kjzEeKL+GMx1f24uyV
h3J1ZBp3ePlncqCOJfxwcP6txVhf6T2dRB8DUAFGGk05YiWNns5MaaHpXZAi5OnM
47qc1C9D3KRPJj66EK2m9TVzrLKgthw/zp941S8oQpLQiA/Slty3xdeufJciXkNU
gniUmMWUUcD1ziaVNgHcKSPHcZQe/wo475dzlkkOeKMjKW3p0efHxSdxU2Wh1g26
Z+qPIFo3mpZUiF6WqHFRU/OGCdnbBlhKTpbf4K9JsRw5Rj/sxKfbiB6WgIN22gqb
4QAYTK9pvWeifA/wKujAyzovMAYHorGyTslkjKGXc8hGT2gFy1Dh0zFFlmw2Wh7P
h3YUBjf6kEEKMOPXNtAn08XxzOCZD2iGrHOTFWjwwzlP40cbBOmyHf2jzTBDHYEB
EIEQUuQBYr9LyJIqk7lb6yDQ7qTheevnm0KdAgUoMTx+DW4Of9uI9yVRRYVQPyP5
iGqlNmqPJ1f/oPqeuHGKJ5Fv8zD96glu9Ke7+y2Dl/wk3NPZshDzZ3OrA+SW0TGA
Z2s//V3qERbzZbRm4QklEVIVNoUoFl5e8fNrZAk8Qas2cESlTolOQTTC9kLb5JQR
3+vrIQ4xR5RBl5z/2w5Rk7NHoGv7Wn16gdahhEbWfr3tHvrfGtqJD/0938R0NIVX
S2UfRrLZhglOsGrLDcanxLfQkiAeYPPOGwad/f02DzK62TvhNMdVShsioj9HoVQE
JdxvRD08oHiaPs3GmRSgD1jRDWuTS4lr6bQ/9+MWl81pwyg9UchQXgLR9s4w6/Y/
b/vro8pbVQ31SkNo2sct45/tD0qeYTGv4cm7urLEiHs2I39d2zAlnf4ZOTzBGlJd
Sa57HhP33QNVa13zB4/RzqKzA+BIFPgHdtfOcFP/Jw9wBDUh2NTRM4Isnpz8jCDq
f+jj+1c3ex4r3Fu4cuN97UXx+xprBbL1mgnH1UZDcly+0bv/j0CyvrM+vT9wUVuH
HQxMkqxG4aLOwbNO0MC3/WTQdrlzQ0d/TwsSJDkpeqjih5f/gTMEyT5tXfEjcKHa
LyepgluinmV7r54bf59IU4GyWJzI8SlGTz1H4uI6AF5OzkTlG38jDUP9hjGXU7HR
Me+06su9zzMj49fpUp1FrLzwYOtyhqd/KyzpEQWIlhjdXea2Rd5OyEesZBb8+Ryx
HY4hp6lpYlxeuHl/KPJh8ZcdDTRV5TAtQs8sKOKkc2qpVlrg38S+rZ2BShsu41le
gSz/s26oOp8lZ4p4fgcObf+dCxndXF7G/N0a9DCdnr8A1gSi1nD1oYdot/a+bpgL
cYHUCPWhlgIJvoHX5ZErtqacWjy6454sHduVkaEOIFBXjF2BkIKlypHeOpMKgLso
jcMSV2J52hno3alLyx5ubNg/8CiBX2SiCx1WSnLMQAmjrWh9yiDO5H3c2ERvYS8F
yb78HxeCGjvnm7ykx6fYYLckW+VQNFju3lJFf7RJGVTqS7PpLP6QyyHVkFl0tpPw
fVdkZ9FX4Hi2yhh2LpKRSJoaumBmfulN+TBnjSjB7XmmucZrmUxy5J0WAKrjtskY
0gAVcgXrsqdxHDIs9qwcFUTd+tHtFLMpI6KV4WejqPJPgs567oL0+Z4l0ai7ntZx
dydDBMrHgbMc0ud/DqowDMVqVf7Lr+jQbggMLylOj2XcXvYL9BTwFto4wW+ZMOBC
Tlc2uwpoks6LPOi5D0eHHPrx3LX2IJ5rGX3jx7sEJy0uH1mGqu/6BGvFaOgL6Wxb
TuLbx0lKja4M7mFIwN/9UmpaE+QfORO7j5Tjz1viYC3Z5jHSzizcEth/vbSF1WD8
Kh384lQhzfOyVzM30Qvnv1Vq8DOuZ51JlKtOv6vsb40TN1DYc7WlLNLKnwVUrBFW
cxEzerkZIpDpq/8H8kV6wBAYct0M6xdtbxgYQwWn13qYu5eINqpVgtcabAbe33mr
HkiFN161E000itdaYg/lbPFjo2NiaMCSQRisoAufrHtrndJYpmhxB5RWPVpLWbye
84AROIWssoc9zjb7mdyzpAalnkG2Tl9qxXLV6KPtyP/8TrFLfIZVCQBI2+0d8SAk
/pe702YANZSYyPmhcnZDFvCeHpOg8Iwd15h+oXHMIQJjWGs4UNjUTHNVKIzwndKR
vYbApkUZJDAAauUvMgC015hCI1e9KgF4ggB8ERZWfmzE/AkCoFtKaFs8GWE3tVA7
VzWe/rvfVjzcjjE/Upw3f5keQVHvWfs4jq7cVsJus1wovA9S3RoS2stdKe5YSaZk
LbzfMTpBBbBbEDLOvqLdXvsM59XPGp6GPbLjoppdMtWIttWwEqimEpLoKHW2ioFv
YCnU14KC8YAtdDlzHFP5/1xBwv7c5m45+OnAr0q5bP5tLQhELWZXsJGWA6OD26bU
cagm3+nQy6wXfbRQ+Hj2lj9y7rjXEAawwucLtsKXL7MO9vqP2IJViZDx5jh+jgLW
DOme4S/X1EUNJKDlPWg1mY1Wy4T3XERv6Sft4uI4GHUxZ7icozuyI8QU/iR2Oxvq
1qTNJb62OEQTwEB7crz2E2AJDvn2IBXodAHR30YGezY02F4Sb1E0wP9qlK1hteUf
XyFhnDj7+eEsA3Izc6s25Vnyf3fVogjxlwW+ndrgVCwFmx+rMhze/rag8kEimQ9u
qDbR9UrhRqJlv962V+qnIGjmMiqilWNWMj8MMN01j7rXjh7+kgR8biS9dUaD5pUY
czloM5UM6G5DYGqLHCM2S28bY7m2ShAGDA75LhAFbEJ984rTtqAv3R4WjC2BR/c4
w6qDF+B+uMHXDWr/9EUC0pLkp6MzLHEAKqC+TszwVaZ2MEJrKI/ypsInHO7NCF7T
6VtHV5JElW/vFw4+WJHWAQmVdXkvdtRFTNLpXHiGpj2BKT7EJGEb0LltVr45PtMx
FkwwMGQ9ADr+lIrFohHCiZjr67lo/klgy6eZunigqga3OZGAoEoAIjMJ2jHvlXOz
rYooSuOnL//qGWl0BFI6Lu9PjrOX/63ouxR1R9rpTr3CgiZWEIDsTwCcG21qTMjn
e0J4XJKlWUDDW+g7BHSWD5Weba9I0/Z7gOUr5g9fpTtl8Ec7+RkTu8UsWUxdJ/st
pveqkkg3Qog0inBj1FxzKBX28juwH3NoAaxXA1G2IR1qfRx2VilBQDWShGmKRTUi
h0YTOjTQe1iAOfJvnMzkdUjJl24b9ssO9tyDPylzdarg51NbxotMU0ShloognSGB
L9D5OSiAI01IKdP7j79j7+84z9/BeYZf/5UVP0mqMjaEwGYiY3TxKUjvo7m3byWG
8LjzRwsWEvhFVvzURLXATLcwNecG2Iz+4fzW7lMYg4CrXMJbGeDTiokzEvkWo03o
+sn9WTzWVUhdZeVoQe8QLWOLOkK4HLoH9WLl5fuJtmw8MFFoFdNPSZWv3r+Y3D9m
NLGGTfCcY+AIjhHRKgopGMJP2GrtsTdUPRXUR6yPWnsD8gn1X2N1SoZY3MHBCvoc
pnN+44TOZsAX127k4yBlzrhGRMp86FymnJ5CzMAzvxfz/q0wpBb/+v/jgcYnxXlW
5zZSKSjJTFrq+q6BAfpBeSN1oTG3Onds0v3A4Ud4d9Ysg0FWSG7ao4xDR6AJ9Y7B
tqr9r60ynEVizP3/oKbeSyy9advBl8F6BYmoWtriqvPJk9SaNqEzUVrljhOC9l99
VDQVIVa6vM1hl35VC86XUkYQLu3luVn9yiLFHcvBik/DJ4mhv6vMlNVmz5T85OvF
u58xpdTKM7bXnClCGEydWTuhzTqZ5iVsa5FdVZET6HR63ot0TuSniTvfC2hZ+lQf
4+wcVkC7be4W1vmKfzlB/HVVJFaT2aQhAMhJoKZfAFPdU47xpJz3DpSEsCS5dgp7
1n7Uvu3bxyrz0Ct7FuVUvb3U7vjZFEjAFpNZT9XuV0u0ci7Uhf+fdgV/r3DYX8Ch
Q0ePnn3IwP0ogFDJ/CBPCrh0XnoEd2fOBviMvg41xSVQVJgqUJMbvB4gk6365YdP
IHSQCnsE1DidI/li94EwRVzZFl/C2wp8a0pN62bMXurBSiWU7CQNNJMdat/UabPg
CTHkezYioPSHiXox8kfOs/k7oQG3uBCZEmPeMkufUM5gT6hY735mPNjkvrZ+xZG7
2jH8xuYU/dsOIgCXd7xBczeJPDnEnu5eizXBf1Z1dANgAXSikmYj9HT7gIiiUzCg
uoqrqXCIX5s2Igv83YWUHD50Mb/O+6Dh20UalBkJkPJrEOGpOhIidAAT+V/H368F
LCOHxBJf3B04fmlnCuzclfP3GO8U3wjos/1n+2I0yKbOun+7s98bENdOm/wVcVch
aW52wvCEKqWOBH0LcWjX/lcyRRQQTf9CvulxQiyhOJzE0HYWUz4nHZKUEqgB3nRG
9axcTI+9C93cwbQgObc47LuJ89YLU+LS96hHNpfBSsFsGBj9nwQ+rdTZSW+GHZBf
sJPX4WFORxq8x8q8jByYTPu3Lo89L0c62WXJ1yQbdNyVZyeRyRfHJ8vx2J9h50fA
XwcRj22KbjdVG2+tRRZTm9CJ5sYOYYlX2kaxw16YgfphDQHhyeSm+lqT9xKgUheJ
c6STPxTnUlN/nIMfHhz7rDI26Oi+h5hcw1tauOe2u0xkO+7NEZTyFyIoiJh9im0z
88Rz4fb9Jce+V2aJSzOcJTXSxDqpEmR+WN30L/XEE2oQc7CVigT8TbWKfcP4PE6m
UGIIFrfyW+5Sr27FfbGX30ozqJRjQ3PzNLDHZBVipoXJy7PwXau0sYe8bLIJSZi9
jhO+h/gSu37WzrDYURfzxmwP+qUs+tbjNhB53ld6/8hsJkjY/u5taWSNG2AIDCaI
bMrxHNZvqGkkG7A/vtEAgco2vA7cuY154aylqk1JLQqk6QklpBirm1yU4tnT+Z+/
jzHPJu1Ci5KydDodirLkTQYZwa88VxPbReqasLLmIVZimosxzORWBQW0kIFDfZKc
1/zvups8OPISnxd+bMoxdbEWHgRxndTvXRy9SbCgzrlrFZmRiPAgtSRUb5U75yed
FdDT04Pge0U7Otr4m5T39vDSLFs3BtP9HeIYPbr4qrGkuJKM3Lav5VV+sVTh7wSa
3RmzBJzVGHFNz9cqliPyHxYhhhxXOwHFCzurB07oLt7NLTEPlDrU2h6OL5ttNW/J
KGcgvQswaF2HBQ1MMvKRqMzA5e9OhIkGQXiGLC3+LUpOk7BUPZksOjeZFKTVncn9
cN4J3tHiJ8c8SS8bVdyLfw3YLH5ZEmSCz808583nqPerKuACt4eMxck7fi0GVsCV
taj7CZz3wRxDdD0RkxFpMEN00M2YifvFk34KfqvOAf4mm0Rm0Kr0kp0UMP9QtqzV
R06F2MQ7Tv2wjUbRs5bXOddUa9fhXmvWAxA8dkLu9tXgu5p0ZcLRX6BrYRRIhkqy
Fbm4ht0WZBCRjbq73qwGjIb+/XO/kQ3hB+9adiGle1LBc9xYWsEuNPc1Aw/chzR9
1/S3qeuYEvNZOYTCptghmCicAYxZDU8I0jIzXwqI3fBmuCR9F68xIipKO2Ee5qNX
6ZvJnqOfKDANKiL8N9fk4711y8vJZwBNPgHyfre/5zLL2d4R/8E5D13gWQOu9M6D
IprgN+6euptiwBdLilBXz8PpQplCcHEmTjRPXMt0wK9Za3mttaG48z7f38bOMcyl
0ACYBAxh71HDZFaG4FcQTEMK9FzUIOSMrWmj3wyPFI0GjPYB0yOsblftOJc5NRFi
Af+pWJsdWDgECTBau6gshaNlX2AP2HQcnbbLsdOMUEc+yKLel5VtEBzMSIMJei2S
Wa0pQGY81uSJPH22h6/Pmwt8ZlfkfYnCJT5rpmUexjBEdbVg5raK7MS3cgxlIujV
n49WkAaBe2i5shRua20lUD+hvDsVyVjEuzwR+J0tzZNiPzKFkhZt6gVKXijwgM5z
8e8ORIMHEir5lxm8kSUtJYXOQeF24YWyW50YqezbRPU4QYWw4H4p3wWbuWet3NyC
wNEaPDS2qEwwrO2L93SaXxEkMH4Lmsb12FyliTAs5Z0QPPDS5DcwasHrOLiTUv36
xii4nsRkuO6oaW9JlA7xv1WYzrHQ39RrufLxn7lpNaCz5aZC/UxiXvczF/JvCgFZ
nf1dSiwGh62O3552/qFgUbR2ogSSgxXg+bL4hlBXZuqjQKACVjzbs7DtvkIMkvGB
/unCMxtgUO2FP3EFkyknFniU/bizSFFu0+nbH6Yibr/6nqQ2eqUd+ChqjhFKYfTT
TVTR4EIoqRdbXQKzBqivlwkow8JQMK012sEfAJY9j1VmhHheb2f52wcxZbAxDf4P
pqko6CK7X7bJp/iX5Au2iyYhXVncJVzY8f9isYDOak8WYkIJ29Xeug3Zf6e4+JzA
W506ELllrX4v3u1QtajUhzqpvNNe9IwzutyNOmZx9VocoDE3DyaLPSTqCF9osbBo
W9Qlvqq5b50hffwKZM4sH2UN9v8xgvL0Y7JRoOx4ndF/YJ1ANzriLOuRF0xj3xSL
sl0KgRdsVOIvUz6lqjk5u99NtG7SPCQ9qTDBnmwbgLEfY7YohB9zmTCyj2HjYz0k
teuLMym7p7ajOmkE0KUO7nQxINkpx5ewjO02bpdQgWuFCPshtETh00Xdrgb+VZ2p
rj6cOiNGQYg3X+V/3yxsHO1Hp0LRW7ZeLnQqzkoeSwhhwpG29sUGC1ILhqieM9Nd
5TOAKa7bLgQZFrQAy1tnYzMlP4IHdb3ffQ25AHJRFXlr+uAOqIGyGiTWleUdITHT
DBtaBFxYs4UbjBpcUMmbtIMghWI07ug6xPLfls6JmyNRAzHHTN6AKDsPMrDycQjs
9LowoqgFs/hQoKbUCSy07HOYgTkDxiFyNmCE3FBm55bFd4bZD5r1vBSMMU23UaWC
XfVeHP4CmDNyxElUSYuTVj7BKjsXZWuBlsgHgoREOLCMDXPFI3/gbzsxItNrfU4d
xtSexKNPxeFytUtvEDOCsgIbDTZWUYYPVEk1gDIOJlFhy34Yw4OIz8Fckw+oXoar
TkUtj0I+ToC/6OWYvpPCNMAOuS342mz0lQTsh8Wdhh27a8mqPhVzi6bdk0qZ+seV
Ky0nvfsOhPovWloFn0nE2Slpp5FqLvkeNmo2A4QiWUg3+4+ebVzpz9iwUezmeuvS
1KThckgBtOmkSVo3IbvRkArTwdQNeIrYH1RjNZmO/1vTVXjppSE+kzsNvx/7/S6q
7Mlx7drVxewCO7RzX59qlqRjDBg55aPn1KBKsXILZ/6TFZoT8KdT45IGfJpOi80V
3JWeJsg+GltBc9T/oZR6JKkve1Aoq1rnUlpXM/oMU3PRIArik03aoBnUA7tMwpFL
JsxRFW7RoRXglbiTU/ljwFpC8mc+k5qpogiaARClaDEN6odWFZLPcBUqrPGYjliU
+4i7zEdTu3ywN4NDE949jzcvo4ghrwOt4tnmtAKW1Rwgpgjc7aIUeYxqBoYpc5NT
TamZm4+5RqRaxkdScXW6FmWIs8tSil2HMm8TXs8kUh5rxq708WKm/gS2jdPxn1Hw
pFir3mav99TuhniHrr8YIMRaOMiTyvj25IgdFUlFzGR0VgTRN5Q7k3CyEDate5l4
D6S3Qi2KHey0Niod1JK0HhlUmfaX4ErwO/r+NvAq/a8bNsGwgRo39luNP56j4ant
+u7esIDwZjueSFbrmnjerQZE9ASgk+2kwTPaO2lSnJ/8VyUxWTnIGav8Wr01xLIH
PQvmbWQptW6npMxQrISkY8EhKTC68FcA7oaYphPojxyIxZPlFC4Ag1KyofVgTPAu
5xFqQGeQVctykVjXm9Ttv6ilAhFvbEQl9Nc/XMKNOctmanZ0NAEYAeTCAQmTsOq2
NHkdYMjdS8t8Q9TMwUrqsCgBo3a4kxhTb/bAxlpDtPwDItGXoUItbPE1kLhII+4S
hEBfyO66v5Rs5JeEL9MWel6m1zLrHYveyJAyc299spWzBJedCBs3zA2RYpbataVp
0W2m3VZs1qhounWlM60bQZMSaRvviLfICpLsWuzPWOLN9A8uava7/SipviY4QHBx
QvAJNyD0WiOtv8gXduB+/poXjP4WdrgQqW/scVUrl4m0tjBKMG3qdEv04IzRDvSb
wsJS6c5B3btik079j7zsvDojb30YjevLYIZhDxkpvzV+pLIdHCxRp+67wUA0x4P7
nveaWpMTDIeqD3KMqBWCUYWSYG4eeqyc3obd/5CyDp82NNIBs6lhYd1ASxg0ual6
5CF9e2jiuF+AB8es7K6bdX4pviAruDbjz+gYUtqnJ3SOxu+oLzgcbFITV+M1fQiQ
ahTGHjr4p7cWrt/5ArXjRx0SagYW4R9LAarUMM57lvH0nd9EJwClfQs7pPBNFY+n
zEqC1CAkRd9o0XMeddCKxsSjfomxK+lgB6a9Dq6R5wTzb9WCL74Wt2B7LyzTTVab
atkiAByEyi9GFLl5NKsqEIx1C+/9qSx3rd4NrLVN+GgKdtnyMND+sQQG407RJbtc
Knh8wY29SRMHFZGEI3aVyFveYp27T0G3qES1iOkEdJeAoJ743OWLW7eeNkLhvZcq
fq+NtdPxkzZqVk+kpt4e8Jx9+uv9PfGTUq14jlk7AGX4IsMghPkrjLMIi4d1H8M1
vAFpZwA/JXokEVMVYdj7KrEu8fvLedGXUKn1+OJQ41yFAe5aB33BJGqZ/Rx58ab3
9mVeKxDQ9MTmGiX2sg+Df4fCytdEZ/5wWiqWGzHBNvAfi9jk4S7xObeG+JukjNYR
60dV2WAhO4jHjMtYIhkMgXQmssGSUpjoUmM/wHxSvE3pDywRNoGJDYjtswexhvTR
asSX96E01LrW6xbq4YRsLfYLMNCeYgAUfXxN0qD4etzpri171wMhT5Ht7XHwoln4
SeSnyiVnxbPjII5G7TGxZ2Yz0qU0Rwhyq5qSVjsBcbYDuDXjPuz/YLI6N1ZRgYNS
MDmWakD/wVUq/4STkIH96TFm72OXWhU7OBzKchnoBoCDpBMEecBc173Q06buvSlo
Qnh7uZ0Bpzu/RgmSL4E/pY0szybMWuxZBX4Tsm7c+ysYMW3YisTBIrZA/uoh4RlX
thjeC8UU4mycknC/fgi4/UW9mzMWaFGI6GzchuPR/XT/T5UXG4Uj91/j5Uma6WcD
VBv8DUCXTS5InytxuMupogJ+wlNRzuoGg5dkXk9zndwHElk0mc794qCeXzdWX7zQ
+B0EcXWDcqnrDQZHXpyvgWAQprFg0Ixzidg2ZbOzVPBFkYgpLmxpkR162GRlQkle
QZREUmHCaUjMBaqXGgJDrS5V//K9c8MWfktWK/sQ3tyB9JJn3yKKEoLBtAVnvU8z
p8FufYQxOSPFd7KjnETvJk/ATsRuIn2Gif9Wh4WaOoQQABmncVVLJ0CBr8LCQbyb
vJIe+PxjtLTeSxDw2wXvag4+Tz74W/oqsExNQe72jvrfQewm0AZVkjMb8Qo/4FU2
1qVrSZllXZorFBz2zunFFZVAarN7yA5StmIX0YeZEg0eyinbk9GhuU795/ATbwkG
D8gothgIka3U3bSPjXuAH4ImU2k6AxZqacV0TCB2tXM3U0pjABJdnr+9oCzziRa0
8E3Ieprt2m+MNZ+0JlYCs4EnUXrU3+AvIY2q5t77WbzVfPi0Wd9kCqMl7NtZiQUN
XD5cGIar8vhzBQI//qgh/vVBVLqvuUiOXvVTRhtGuokiHUJILk7wRdPz2jjUxTm1
+8wUtdG+6izvGpB8fnk6EET9q0PaqsHZ9yqjXDHSTFhkpfdrBTMkiTXc7k3GYPU3
nVQDfHuuo1S1nzAcNdjdh2+0i60pohDBNDxelkmrKH++w0PirOQtrt1cjUCjnBZw
1FIrt7nk5apXR+UcIiArRn6xPAQr0ds1HD/ROCaOMcUSOusonyK47Ndy6vmV8xgQ
FqRqIq1E1WtEg7e84N2LzqwJ9DV8MwT6TdmsTjnPvaFgYSTam1Sqd8IdBfPo0Zte
R4n/WPAzRfkSDi64L9CPpLFzTaOOFvsMUPKNC1QzTKtBMg4AFDR0yxxeybdKbo6+
xhEUxPGpbCDSxp2U9pdG4MYEgdEuKz6bea/Bw9yqVnpkF+UwCby1MJZsD0fhUTCO
uJfWjvNd3+FZSwB1rdvna93p0diNJaR8XoXQRQ5DFicyWdAadgcKwadmTw5VTyac
W2OABEoNSZ1JfNxlT2716CuuI9xztmnu9C4wYBTm2KTbOtYsKahLmWvaWEdmMp+o
jI3Q0Ym0bkbJOogUseqquG8YUV/bPO5YMK3dLhC1ymX42URWQ3yjEIkZ7HhTblal
+LbYfldgkOizFGwlVnVpm4bQ3Mz19Vug28tZUlT6bGEvDCipapjiAPNajcdvLFPq
Ytef/eCbNyGSI8ugpbhqm1t+Bnhn8SThOWdKMn3KD5Qdt9vT9nzOKgT+5phDGoEP
fgJ6pM39FooeyBie1nxjw58xfAlegI3JBqTknQmu1ki3azP2GqzAx6dnpDz7jV9Y
5NqXCYdOl2ckCQhvWzfxwyDzposR/nk2z0pXrp9GTSmusVeznNNVS7UxN63+Ewv7
Swlmq+BAhi8qWq8dwdCXyKMHeeoWx+dCFBx7CNYHf0T8icj6XnGDEEhNP/66hJJM
A2ooZTmhoB7K/XR0dbdrj0z39usquSIeqP8lrFJPQgh34H1Ajl7xzVy4YRAr9G/R
CY6waB3ww/4c78RJxfMrmHYOaQ1mG8IrRku/fuwruiApzWf9DOCCylClyX3NRMcY
L+Csugak8F5JfFGJ+NIOMqAETjN28D27egkJatgEL2XtJLSY4jh3NodEERYbtRei
tnvo1dFXeowrimOglcI/ungzAL+L3Z2LrAZV4McwuGQ4n6EYLxddAKAHgg1LSzg8
77aqwlwtOj2VeM1r+funtYpWpTq3wVR/9gFGdN9XY93nQzCyuu/tbicPpkqVnAI/
FBHnWnTDoypXmfAarbwu49qh6dU16btIJiDhC6tvVWyrLXycAckGWS4kkzKjU8HF
RxSYWx/bDwEV5Jhl5g3m1ilrxc+ZNL3bdXTsXXJO4T9gJJpsuRIBgNtPFKUQ/zCK
eym8uFdXw5NgI/jxdsHe6wYTNIX0SyT69nW4+wy9FvPQxp8ke4sS+iqYDs/l7azw
7bhuatUEjiVa+FHd+TxWBVBLbFPHGgS7JppkY4K9uhminPRZwiNRBgfSE+ezrRLx
nFIRnq6s8TbEedjDGngO1L1/g1fDYvmAbNzqC17nlVbDdwSCvPaGLKyH7ZQFqaRJ
hv+QZHeVdafpIV4FlARlViLQjGEWfFwmMkE6u5BhFdCT1gHoBXlRH9z5kililAU0
dB/i0jZEthj2zizlGq9NzHN/OyaTxVktGX8Mjax/38AMJV918hqLcjCXdIU4Cbzc
lPzem2JSkIOibzH+u7rPzC06iEfYCskWCTpaUiLFw/LSg6KnwHTDOAo4gj2dz+bt
uQXsk8UTFlKA8VbD9+uTv1Rk8ZrCKgCf+2P+sSsyVt+j9Hg59shs76PFMVZnDdBn
A8T4fJVDpLGlGo8FdH+a0t7I12Dr+iDPEKVEUWO8VkClNXY0vDFZ+zilKmtQqiVL
InTk1pBGWLQg/6YVYRHevlgLLaHf6Xt289lEzAlVRjl4DdekWIVWzcu9ax6Lh6MC
jLoapMiw+My8Zg3oInFSsO9m58zNj9kdAmuD4JhY86DYcnIRqKnOMG+avLOoR3V9
VrFb/fN+Jj+R5AU9ieMlT+a8M5QFDhLQjwfOny7Viof56whro+m9Z53454V8yPkS
rMejK0CUrsv+JP0W+ISTItwOfzurnVOAEKbzS5q5BAr+uSvrFKkhm8T7afAcmJTj
NwdxADmkidG1JPPZqy4z4rI/ZrEYk4qXfm/5CVb9mX4hF2g/q49L4P4Ku2lwVVR+
Zrg6jrXYm1SI6kAz/BCb677ahrOCwAJ+WxwnSyjEywxIo2tlwkCHjKP0ATuVqMeL
Efkqm/JhpkZEZtHgjyHpSCBQYkV3J1RjUQSIiXNlFYqq9KlPi8PbKE+opI3BqCyI
R8bQBWW6gaPmeCVS/PEigjVpfF71SqDj+1JjcIXB8KrayPfiroHduaYleQ8QG/Rn
4Tb+61O7dg/XKBQKMS4W6lUetsYOF4H9PsVMpI+dAvsue+7x9JTDVvLYPX2Bgehr
5tkm/JhIiMIQG/C1P8TN4aO05i9PgXjXFnxSfCXZKbNyRUJQ6Ppa9/VCh214MLEI
mW2oZ1BnhkJb8blgxRJlfWRUh7GFLNirQL3fWOH8H+iKD1ffmTgiud2FZ8pdCBKL
5MLptL3yRDSbD0TCuCQLTzDFAJ4MsFvnz11o3pmmM/jUOQU/BVriaDiTM0b9rbxD
pS7MCxburT9R+U4t+8zGj2P6sNbqRI1OAyLJwPjwfgp1eRcJ2q1tEdiBRRcXIFyO
txAbYaBsTcDx+/voBvzEY1gcX6JSH+ICYy0oZEwS+YPsdIsjW0dUqdr4tYAFeNdu
sbLC9WvSgbUUF66A3g2gDEnpXF7IgMeIPQsSGY4dC5QerrcgH3ASJI71a8nzmRf7
TEFqxUFh5xQacg3b9/MgQJ4kyqvdsHpdWBDFD1P/q9kNE0B5XQLmKJbBrrEDGcCC
sExbyPCdbZbEeoUMCSLG5T4qiESx0o/fqV3tVpES3qO8cMUyy9O66TGUgkHCRiOV
hI4C5G2ULiodcW8An3BhBgrB85FADDFTQBIcrrHuX3bYVGRLqsyxNFLn8w5WxQ/x
AlDRzN8n240Upyc17JJdouYlx2eVjyG8TSJEgYGnh4P3RdDHNW/9bzrIsSdqrrWa
tP2EIYKm3xClyQ78XHhvo5y3wA82lfsZrtKV7oVOaT+eVG+QyGckRt1yT0WYgPJA
nCMRQD6mxCfUcDq5tOmAXFH66Z4+W2r7jpf0mvf+Q6tzVi8Jm3vBv2rYK+74TgBD
QjHFfcIv7/adyJXSfqh2Z0CzAzJzeha/fNNulv8QkUBo4Db5EyV8JdekEtPJXPLg
8mJoFwV5Sn/5yQrqx1GGxbWnTkb9QUQ5ILkJ2F3Djc03vdwDT3qCBHJ74h8zGEgy
X2Rryfv5kJ/shfZ/sEI12VmxOxqCf/gSbi1MiglcWlaNWtbwf7v4lOZOQnED2Ue3
m+RSuyOvz3ZwN2VpF4rMhZ1AsSax6JUR9eqHGTdUpBjW/IXjFuIokJS/IYLgQC7Z
QumMsMEwFPU4nNAmCz3ADK4Q/GrfZg6Ahz5SkjyCsoxr30FLlPG8fvbPukT7WXFl
xKTCs05Fb4pz1UYzcvyWxsdWvDBaeloiu11DJcUWFYgZz/3d5XqPu85XXiuZ3kGz
674eilQOVG95VGAHJQhRQAEbjy9imVrDhQ8qqKVuEFJFC5NQRqvRNrB1udOjB0KU
PcL91wgP14y07h0c5q1oeH47GALuevhaC2uk0VYW7RDTOCIN9wzUofAb7dHbSKuc
c1geVMEMcPXHxwXnikDVAny94zBze9/6Q2FWhhHoyH8dV4GiHpiz+bOqyqZpqLtw
RquKaqPHAU4kO9hXfP76knqmWtD5NjZYWSR0whAN+sAvEQMDC/finUEKTMa6B7tw
PRcOJCSfI45mC45QxokS0MrwQs/PKeA5SIuhWBv0bzHnyXFf3iDB5wJUA4Fig2XJ
k4bajYL4WPG1K40HVZO6d6/dnw6qm4edlxCBa+8qOddUovqsxPH2yIiIh4KWL2Ix
Zc6wtfBYNbP6319H8viGZSTshLedkW3ms1jpjA83iwus6I0vk/Fx8VOZ/WWUFEeI
RdFpnuk4l5WErG8lXfoPD1u59pdHXpEg6C7o4KQg93Uposi0Cc7ATpbujjQh+RxE
PmMmIsyYELtmWFcaLWnY4U0kmWFyhrzA86yatMnsdi0IKKmzx483SQJ5c0ibpkMb
ldAJmiMYsnKG8TxYQOZRQxyYK4Fw/UNv9JKqK6aB1p1F+piJY8NGiJXuaBNezYfF
FIPyM8S6yQRDJgvoSAjIGdUMW7aHpdyGicgfjZ1LGHVs4XG1Z0s7/hVkCtiG/JxO
qg7DIaLdvAFUeryCqJYrWwiVl3gmVHqUCfaP0lV+kgh4ELSFPnHwqA2hb0nJm/W8
ZXjahME5T5PPXgje8xqbKinQ7i+x5KJewwlgrTYuMe+JwShQ/I9H6WOPyGw8ODw6
mU2/vOYgo4cZ0ORijdD8DHZ5+WXblOH1DEzsy3fKegakVmMPc0l7GgUwWZnK16I6
9vT650RHLE/d0PJnCOW6lBKMiCnQIYrOq8EBzmkexywUvq4+8E8/Kk/tTzmBb6kt
nsj7bfL9X7H6qFLfyrqW/kd/z+gAEGVLHUGn0GVFI6DTSAjJ21ONuXeqYd2CAtsU
b0XFxQY0blUvh2YiPcsDtG4drgfq07EqSR5S/aPjZGfXBC9o0xRbbd5Tx+/2lD63
pUAsODzpRcxCWXsWrav2UZH4Kym1q+ifPuU97ay/zGsB26+OHQrnrcBFnuaZPVYG
76WxyCSKqmmjguQxn5JoaOHw+sjdyR9IJpwlIdYTfHlYEPw3st4DPIO+Nsgc1LSz
qSsGpMTZ4ehdolwlvVYugcGr9VmCkqAcX2KuVcJCEwdvckVJpOgBfDkbVzdHzR4U
UxTik49DnxVLOwAbqsNCxh4DCnBrcI99PrSugTd0RFNtXv6vj9mV00TJjgWXiz06
AjFYjOLZXTOEVedM79CAoF9mM0jmiNYCHj5Cy+H1nLWKgbRNgbTRgmYA4+3Lc6Mb
T8KNNk4ofIw1ZUfqz5lt8LZtaY3CmgGb6zShgc9+WBLBavvzzysggZv8ZR+69kfm
v/QLTxRTfR73ONWyxUIRPZ60Gv9v/Ax41aefTZ6wwqPvz5COJ+MHTdapAKEumukY
wu1SL5q9KfS1DOmJ6OZIGeJXzQIp5taA0xzpiuBhv6cqlcG/zrx198Wu5i8vBYcK
7DFJFqaDIKikOllkB2zbH/8TV6RbijtCWKKOJwj3AIhFy5yqgFL697Z3iPmCLNoq
aOx+qF028rZdv/7tbFFzGP3nPa6jvO2GvLF4N+KsSsvN/cM3g6jEx7N+Upwr5Sxp
HUKnhL21dCgSz3KVURrDUDwODDqOjgaGm29YE9HFb9vLJI/TImbZWR+8mXsxiyxh
9gKasl+q9e52UqEwDy1y+kezq7uhZopM1DFGxz0ItrYtOGv+yqRF9c2uQHh435IO
rPQ7n2MmHcfCH/mBQHO2EBHt0fqnd10BqHtX46V/Vb3E0SnUn30ZWXGuzA+L5p7l
NI7G4fJEBdl7oSug/9Pgu7BBDtazJ6m0b9w5lwr9RXtw78EaDp5wguLZRs+p9+sS
5z1ho0Ip2mz2QRGdniZYEByeCCGC2yvCti1JncsnLDZSNhcisqaNM/g+evXwqCo2
Sy1yLgMfHzWhZroIeMQHNlqh4awb0IP0S645L6jQkV9FIfOJ72dM46aB0yj/aLtV
IKSPXnmxtri/kbUy3LUySCqlamBiC0kZz8G3wdFrSIWoniFOFU49mqhKtTil2bge
SbntO36dpLH38Wc65eWcyMJ+wmfhuBJhlSlTPWLIbh15mUkGDLzOoaw2YDISoY2w
nCdIPvIxC78MI+HFxmUmnqHKwOoxdWyBh4xeCGAOTIPM3fbUmeKqDi72a2+hEx3a
F/CQ54HQaAjIVBUEM318tcwan7DJxkOT5KF9mAuyKSip2OwUwtCuxdobR6Jy0e8H
3jSeERSqJO1GIlDLAwpIAAUM03dyauloL9B7RJSsXcGIj471hDywKmfxqwBp3kX6
iDoRl4PtmKWKrmvjhyxkKpGJ+z/pxVm8ejEEqQUlxbFIbmVQk/+LdLor1iM/uVpX
Tp7VSwU1+bdWsAh2ycCxtRG3DvXZa2aaR7E6Hjuo19dtdS10b5RaT4M7kj9gTsTd
G/pzCiwR30yAqRsNi1sF0JF/LcpZOycWlPvzv0BiDiD8KrwkwNgFiV/eCaO0x/O/
mrqcZKqp5D4uoeHMq3vMeOv/P0Fm9xufCKWsrByDdoPV8TlyHzVo71fTd8yZ6BB+
C4aBT8KLCuvY6nrxMEQ+DX/gMYH/g4izIlPOBi1nFRTcX33BdO88qh2lpc1Yu9yP
VsdijzDpip5gRFVQBPPeQnpvPFMcXp5bwdM3pWKWtLkGVHYEiOKk5zsJwl3dp0HJ
ch2wzaKjWXi/pVFMG0FGdXWHHmvH3ygW5avQiFJz1GyWELHR8yyjYI3VhcATNj6i
Mzdi3Pd/AEsemy5djWdUkjbqg86PQmkW516T83tcju1CvQkWnFN2VMGb+x9tKHb2
fEH2egZ3tNk8laO5KNGU3/gnh3F+GglvFh1+/Np8fuYlywsOoWRmoDIkH8ck/v22
7241YoWemd1EoYKQgPFFtH5aaNWtt9OAjimGGqeepUUOHb0ebCh+aukbe0hKSoZ6
eE4fhgNyIe+nloTTRJBOmLUHOVTt33jUKduMdf+sXw0CT8tPNtmfsYLdtKi/BP/a
xdV5qNY02ll4RUwgT0tDv3mGgziWn6J+GpKEE2xErKLv4HtTFRZClGsWSF3Ysicj
Sn3VGU8mKpHhyRARBCVyrx1+kNCXsCsNQl5A9XMWTs3Rc+8MH4wCUPliT7kChAOI
EPdi4EUUnqB92wFHLaSOivgTdHlh9P8jHrJLjds9lPRABiPqNvG0ObMyzCJqVHz7
3MBpZdasJ1DoJAgEX0AOvl/OBYbgixaBu1gXrtTnXGKuElgbbS+NJFiIWat7fLYU
y+49AB8CP0s9VrlJOxk60akhkZEFo584+Lzro1sga+EfKqTRJlqzHjJH6t86SNlL
OgbbYjHfhB/XfLkOkatZMx1s6NHdlGq8lFB7veiBgW5/We18+Jd6sv/f41YxX8Nm
kUzvnyQQjO9ny1t9wfJTUKxLp2WdaBHy4AzsmtE/nR38XFTQf5w5d7Vu7rIq3kPg
kFRfGy4/5WSw39kOBir+wN+FIsFG+4Dp6gstiZ3chKBGJ7snX7/DumMz0iU5Ew0L
QuqSRscm/KuNLmTrgZ7PtP4C+jporuBbq+V+IL4Eh/9rgo5COA/brJ2hMZC8FOcg
gUlwJRuWM8PbbtmuaA537nyEJXmTTwJ7UpXXPeFw9HhySH1XaozNpTQlU7+LSMcI
qRrbJPIdew0XMUb1EQd9pw6nW7Ay25oI9ugL47EfmcaZWWc2Nqk/yg5AhNWaHbzi
V9KvrbqugeovkwxGJFCENC2u0uuuF1enQvXty+uu0oZfQJ8foUSqZaZw1ubH7gy1
FC6lFjGpP6/nYYUgiV51k0TudCx5sZ3mWxuRU2sN+rUekQVLW7SOpPD+jFmZuIIx
kyD42q7E8LhIWntMKWjVpFyM1Dr549/M3FJKABpoBx07CmM/tQqKRwyQxeEMrv+/
/QQbbNaapfloYcpzVjDMBSHVp2EDaIA4C8eW+1O6aUtjAzz9GDYHMgoPqv9x7Ytn
h0QyOCdqrV+iiPVCQYmXv4WSgv3YSfXxXi6HrAXLBHOubTk3uFklDuT96qg1GU1v
HRJ7sNS8D7RXJQ8kaXLqmu9byX7kb9ZMFJG/WcenrxtNLZj3b4TYsqqM1ijGh2mR
UYbnZhuEcvwAecjNDgFv4VOwVqamjsw2AXXkU44yy739fSU7o+MyTRRvgEQVsTYX
ZrE4t3zyGzhfdaq+A1IqboiFjspTH8QN+H21PKJvlIcy7BB3sCP3z7Cjym2WemLK
X4ujR3S8iYd4yOqBvcExxomMwaef5Hh5Koy2o3/2CPO+ZH5g/86y0sB7ARPkw2ms
MTnE/unSo/i/hvcHr6IUjwCa9m+plCshKwHXmpF72OUHjTVgHpcTUaqo9KbFT2iP
gTBmjYHBiX6peIPgcplQ3kHeEItweeXRqgZHY6NIGFPbsmV9KHy82pJ8B//3YhZ4
3pezkB8sMXmyUdZMc9o0vqG56gwzHWDvbVGHNt0eTc+5yF4k2ssMiy55SNGQEdAk
FroXg2g1rJU1SMTURzkhV6ULh9Fp9lwNeI3NUplhvLK1evdsJ8EqtAclQBnd9Si0
R/J51RZQLDcl0Jmy8sbibYQZH0hWSeV2d2PFUJkgx6Z0VdZpqjpGMWp69Cb8wW0w
i0gkc2YJkgY3oHv/yqr7n/rEFMCGjSBXnHvn/Wz6c+6BzcNfYcnDOTBzO6ar0D+O
9gfI/DuWbAfIT5aN1gogaV6dIVbQUBQr5AUEYq2j5F8CKQWz9PL+sSwtwyt7cf30
BL/psrl0Bb2dEWrjBxcz9qEhYL8QbYldyrv8j3YuFkJbNzSdkZqsgHQRWvLbdf02
ksNevtoc+kefAnUr4Z34eYe7hyDMZEFQBOvomiub7boXCaWClzbPqYiBb835OlsW
S7TNB9texBj3WG5IQJIIBHu3K/YY7SMInXRXdgteKudDEKht4W8GfoyCjUHNzXHy
CrisHnEOot6AKZKU5OvqCHa97X2A8Rhtnf9M+KxXZ+9AYPJlCsnTX/XqzW5AdeAl
wBdPzCj6mPIKQoalyqjPvlWFf8ij9ZZ+ZlG1GfYi0klSIMJnPutPMBzvW8WumeBg
+NAzh1jATSjhIOwEpkOTZ4vewGZIrQJ98DSqRVZ7E06FgA76kUn0uevDj4xrCMM0
OXVOvq4n6hlqar+61f1QxlX4XqvuUQd7LjrX2VxojIxWCjDfvFGkdIZtncjydZzn
GvHkeVgKPG/H32Ss4BcS0BKU4dclZnFAdtWkS2cd9Nr88h6rlglWsXVVdsFYJ45x
+eFuJuyec5fLC1+njsIGSIki+2l62HomtdpggrD0jNzwCsRgX9iITB4cx41PFi/X
4FK2nWIRjGsqXrXk+/rMP7j/ebNTejSdiio6EVB81cSgugMxqWupXdtBp724QDqw
8ZKYttBOSY9kOeUSbuQSvwazo3vh0ZBJVb8i4ROy4my7Z634FVWDxDb7BroZC3Ht
5Jg4UVvDqkpB+zNePygs7xXgvLu/PTDMUATyAsFkMTH0sxlg8m6VU14rSOic9rwr
+FT/xGhfBtxQXdSw4jX48PSVBwmdTp2DBM88xzoVq8/NyaUGv5BV2YlfMY4/xTds
Bv+7R2XKOND9KElkEHo/AU4hvQSDIClVDc/iwwpi3RiE9iqgjipv5+fMJXbpVBwn
FGl1/vvwOgdGrYV/f8PLAzcF4tVqqwO+8g78NWwEEzRvVz53iHrp4kk+kGT1d92+
egjd070KlwY8dOADr8TkoKOG0XQaEX8a5/BOZ4ekC4EGYPE5PklfmjPJ/W2YFVET
WtCpttgW4LBnE6xvzO0m3kjfy7uma+Zl3EJ1ga8vrYdePnk5+46P7GjdfzQOvf92
J+Yappxe4/RpusZ6OftSx5PlzovtzNfm2RQi8sspXTXECX1Yptk2QEPdhmuTKgvt
LQv/7LIkUGhH9J6AAPV2cGGxhRHSKv7Pg6Yt4HSjG1Jg+EkOU0vEKr4w6OTFh+ma
r5chWgnDYPMRTSmjGnjJe51m58dfJDUdLHT6TgK1dNgnIulyrWZpNyDzKPr4CwYI
cxBel4GWV4HhpQ9NWwtI2xX5UCi81PYP6G8m7JJh2xfhLpPy50uD4a/wWPUOny80
NWN53RGVVnWF1i42EUx8/lUTymwlnreGRYExoScfaIIi6F6pz6ZLNp0Ak8TX+6Lv
Xw0PCeM9eYhbVZC7G3S3vgII01hOg+ze9PaM9fnwALyVN9Vhtp18tsDGktoNGjDw
5IW0iVFiJ8D4EGCZQkAapXmhrVYI59wmP65CYw8sqa89tTLjwh5arwY/WoWO35Lz
mFley5fMyrjkhexXtRmhpHjdPhxFr6hleAuESFXX93XyukBVC9fIdQBtUXR+c9YI
hJDv1VyB3ayVXNh5liBdWjAurAjyqFsztrIWJ+wCRbCA5ntpgGgc+p7bMKVmQ38C
DGN7sa3EEzWQulSKfs4H6uQqV0Oh7Pfwu+OOpPYIXpJMKlHqZWrtp9EejW9fxdqY
QBazXDPH6jCMgxBSup6c5/F+FUaLkziHIrG/PEv9257DzbN8HtO5/XihbDWTTIq7
F5rggdAqoWJ3opvp8bCSQvZSQUdBHIxzJnpYzFktM2CPuUxPVUXjLe51hT0YliTW
2VVFFOe3WX+hZDjEIQ47atdrwu0U8flVRvroMSmeu8n85IFepWny4s1QSUTAEKoS
AeSXFH0c4etMc8ifibIAcqRMzGfiSdO1FMuI4G+hI2/Z3iAxgwJvhhhQuOBbIQYY
pHjz8yNvMIrN/e5l5VEYs0Uq6G8QzJbaCs9F6t6lH327Av5wJlErHzuibqy7aETe
h6J5iQACrVOTuaA3XbNxG2rj3BC645TgGf8AMxP8rAYkfNGxlpTu6Rtwb5AISQf3
Ha1zRXL+jVa9biJsNTrDc4dgcGArn7gsWyoqkw1RPL9Q9Mnc3KM0iXYaxIYbdiuW
Mlofw1g8RtG3TCOS7MkrvbA38/n2ely+Xy5OhRtN+c8XtgmLGOR1iLPTKp443lvq
hHlZdcRGL5JVGAoLRq29pgOd/NEoX7fCuhcv7VHcKoiOWuqVQSCdfEjXxmTE8mK8
BPu/cm+armrHXc+0LeuNQB1dJPMiI/o2Aof2XOGmFioP/kXM9CiDXO4b4iTHKK0+
dtJRxue2OHz+TTriQD7SotLnZSNgP4khHmdps8uyMt1D4LucqQxzezz5EsYjjgpF
mLwkmcBqE2VS3iWHoLP0uUGz8GIZ6EH3Y90N7+Kx7bcvYOMnx2/dgx0TNZFSTe5/
JtU6pmRvVvtSWdcBrNMy8URpXZiRDtaKWVamaZHgUYNJW2260WtP53L1GdSkgBtW
6WQLau61VzAx7QUrXZMr8P5xF6zIkt1y9yC+PM/GkgG8YrJ2dElWhWY0UU/dR26d
Y4mLlwF29ViGcWEAlXnNtrIUFdiN+NUZVGclCINOoWpc1jY0Cbk0Ito4kFHA9CS7
jkkW4PenenKa+aYkeAOuXck6VUvS9w5JRE8uAWTULuAY7ye5s7MZNmJvAvCNpA5n
YZQkM49FMNhHjceC2+XYD6fo/lzRLmbhLC2ZxbiSxNrixcc3qXXyvFl6yXY+OraX
u+NXxq84CBBoN2nwjsKgZrPWUkaC/qkibMim/+1p54MSP9SeHQpHdVpYfMh43WcI
Tt7O7UEqlkmFSPb9/OBeEfDLI4MajdsDrBC1JFGvnoiE11m6GakYvPYd8DptyXsr
D93t9kNrtEQCw2bg0DI3ZeiDwEVUMknAhK9dCuy0DZ0ZtSzwRSMhN6S6gdg/Sbrt
PTZ3CE7fi8Y9ge/4nqnx0i0nTOslO324eH3nWoMa1LKEM+HOAGIslL8o68kYlE+j
Vr0ZRMT7hT2HzP2TuzzxrEKkk+UKqZztBy9QgKXYvk/B9w3XohsoAVwjYL9d0aRk
z+QmHkGo6OzQGUYnVPVc91+JlZA1cLGu7Dkd85zXaECLhQdZECK7yXuw2/Clm31H
VIsyqR//fEdP+XGryzUx+S2PHM7MLhmCF6q3FsQ6sH7gb49ZxR+nzeX4Pd8oaGXT
1C+jWYiynrjEnN+yDcCSp5/wlAvexwI16EuMMUZXBlg9WBJbp4iadkgT79590uh5
GjJRL+miDIehceRCpjTWHoMDCIU8cnUE9KmoG4mbAGzet9tALFFbpvZ3StnCJAbs
R7rAs/bLP4/FCuGB8jKbzpAP9pjNtRxDBkSW9TB6fo+BAUqnMvjUrwYPGUtDenpU
5FmCBhu3XCblZaQxn+WR7oJZ1oscK7sOOgdjQ6PZ2p8WYZDwqeHn7nQGV8juuDZL
NSb2AEut6G8uV2OOKKdZ3lLl1pQgxlZJv22baKlk+i94ujbKbPZTy44qpxpFSuLe
xXyrzrP2REZ/9b7DoAwMsC8J1oNTDAPI/k2Dv4OVzCc2uASQ3r5K4jErby04at7d
Yy3l5kdPDnsSMJn8u+4+pJ7V09gUNrRzv/b31ZNTcDHLT1eVLd1KTUdSWG/+ZvrX
VTe+FLrcaSkGNa8fWLo7IpPqf6sZgSvSYzMtE4NC7/RJjxKx50l7Uc0Y6nrdXorA
pfWtD4RwtRLVVfMdlRuw+8gtQuJZoFg9VrgwzB8asI20ja4AyvQpvr4c5SVpMLqL
G3ovnPd7GJxd4RyE8c0DffM5DeF72Yi/AODkQ4+a/y7zEQP/WtUhQ2/WTrMuoIW3
VA+hzzvosMpxwC+IovKOYJbTtrLtBFbtSdA86nyJJHzJ29s3mhlk2b7oRa+jpLds
erMtfm6u1IBqj/2xpdKaoO0D0rgV26MyGKJPegO4W8ldWr1lG2yJnp65cI0GVsxW
b74dh7OnFNzqNbjddhr3fOy5oLXu/MzIgCqWi/iOvTwvH7vjlnOsi7vaAWKP9mse
wI6xzhdVm/LS9jXvmOiWG3Qn9o2uAglBKocfCfyEK19K966hYaqNbaYcoi5DwyKp
b4SyUt2XZ6HubAB9OynGOZAfu91nhkT6lQ7nalK7XVMVPpTJ8Wv1cEN6roDDRu6f
KMC0xCanRll0+NPDDylcvuJrxbwM/+PDmuQhYrfMKd+vT5Pbn66NFwvzx79FrEgL
hszW+bnBu5JAbqx2VBb+sXaGwWoeAQqZKLDwbDvL/Ki2gfNLMZV8OktTB2e9dnge
LsOb1YEjGrNhEL8kfX+DeHZcKbG2qV1z8wmrXgzsnePlbdl6OVM5RWiZaa6Cir9t
bXbvb/iPNidXqQ1boFRHlIKQ1PN9RCPHQBK+qtuXq17cYeaIXGBYOg3F2hWMBymz
PDM41XZjB+IAwKkk+xY6+kte//9C+I0jjsFQM5egTMD/8T64yT1VY9ZN7c2UXYhs
jaAelfjEwK7iT589Qfe0nhopkjCyrBcQy6bkqNN1sRz3sFYQWwB3/yg7Su5whCLn
8amuDelMpdYhC44+PJiXeKWGMccKoPWiU+6AkN7bXzGdW2Azom3nQ2zSeJyqcRn7
jyZl9CI/SljfVdH4VOTGOZalB8lq2V4SzLGq8DG90WLiFNThj0a34TwL+8zCFY/4
LqsFAAGRao8YmMwAqN2/p0hHL7cAuEalqgHRWqs/16Ao7iFb+fmMea9EqWDPJ9TH
PgCDJg6UdBLQgiIF1hjSN0Cbnyyh1yZlSriEtCn7n8hx6KjrF2fbfWDbew+xahJa
jU6ae6M3gA+Ngvv3uYwdx8AcIggZEXGPBgp/yj3fGOqSt8gtt0QxXzIrGFhcRVnK
cFR4+y/Bg/UUJdx1W/ZzrvhU55xsJUyEJbJmjzDiI7/rWyPMF9FRxGncwE0pJYJG
swmtkoJFeRgTMiKypwMtRuJqIZSDd1iqLRD7QFiHtf7qHp2mi/qADppKQNuZ9X/h
TZeMNLoTBShJjZku2BDNYs+A/uaxrZxfeWYH8miCafnPDP5K5Q3awQKUtK6hMQn9
oXHWQeu85jVfJjZ4hL78IBEo5juo3uxtTOVRrCe+1hiVUif+C9Alky3UgCt7+dWq
+cwFoV9din5mYrHpO6ZJwctDkNQxwyFVWJ7dRAQx6QfkQxvxkofh2daMpiZ7JXEg
45NGywy1Vi7EMt8CuQ6g1MUtst61T8M37Be2o0a3wQa9nVDZ/fE2LNQUE8+44maV
1Au+Aci4NzJJnBl2xYUcgT4IeogLwLKaIgdWOad8gVCAepez5j6Q9d9pHpk3V6ck
oSkBc6wToA/pe1nRvs0cAffoWddydBB/RXEqUQXy1Iq7guRPpteYMdiuLUTBMLOT
46hEjjyHiVEyZikJDIG/DGovquxgTLZIcJfqmKB7mQ7/OzjSVuXBLxSv6auoW9DO
ZuLgkQv23ocqolDtgBizhCEZiq91J3notOjlM/82QaZYl/SmfxbRaBpVLbouYb+i
lwLcwuPDq+pqocanLMV3qyA9ZCIIYwK1p8h540aC30XtKE8OjC9gpN41vnOYRS9d
OPAuMUrLqh53y7QQ4lBmdB0Se+Pr55iPmFNYbLcS/825q+vg62ANnIPqBbE0eeFS
si9/X4GiO02Q6Wl98cJjszSa0w3HOqPfNcXAnLWNM0BYHbKRn5/zagHKp8i4wL7E
OJE67Ye7WbVCuZ6fQSn11Cpc6A2ErP0Jul9nk69tEhdgLd6TzUj0czlclTeqQrFo
4BjO20zowYtsKU3oRB2IZKVCahVSdAXC87tZGeeTJlXyKLP5ATwlWqCxI61ncksH
7/or/yS6xS2gI98eJD33xUskzumvwk6juQJGx/ckKntlGTRNTH2ChSEeXiuXpixs
u9DYDFXY4JpZEujNnNCNG8ZzljJD6NlnCxRF4Y1Mqfb9aMEsvxHlltea3g4loB6l
aY1F/D++gH08PkMnSVzDRSBdLHgN6CZsVtlNCh0fddO1DcGE8aauEKJ5wKg5tmLg
dmvHpmykIXCMqaQK50+G1atC6Qa3NKPs2AOvq9nLEi10b/Oih14utwlI/yUpoG7m
lhmK2/qI2/rv6Jh/BgIHVsPiCyEtedrX83frRT8iLEXdLi0cFhCXzIXV4wtUNG+E
9mGYpuhl/c8FbLrV2ryKm13Y6lhRKjW8AyGefLWFI1IqeUd1r079nUzp8bPj2NZO
5e7FoxyL7amC19Y7RHGrGM1UC0qx5NjU7kE73zzBrNxDLSGAE2bkQukU/E8px0Fl
e11PDrzS+9ewufMmXA0MplNGwSxzveWLaSXSiU3D7uXsmhQFleM+p84GguNGaqTv
LrWFBXqEiinfMSaNNfSV5j0aErMKbX+eQoZu3m2j2cWpLVpyWJiCYQGY0jBo9QA2
fFftAHA5NBlrMctznD+ZAkA1RPh4XbbbIOzkufEoECQOPIzCTZsBw58wND5GzUGG
o5ngal1qpZmDRjGfgh/+eBbGZWhAK5A0FYFLcojIEwZjZu4J82IA/cOC8q6E3amr
0heZQsOpYbOagXAt5e3EquOFs8RBRQVV1oQfC519K9j4t21ejG67USnt4GKF0MiL
g3gPwTSvz5vjDbGajskq6sREonmfSiDlgo+t2CAr4cmSGHhKIcDhfjLmsCZPoy0R
TNBzIx80xb1WXRhC3HWjpDMSlysA8IwIPiklEnkAFF0iGpzEIgIfKYGlj4+LzLGi
5BAn81eYpbuxAw6FEXYS+fVuem4bGZJ+nzLGShK2NNGuIKqTHmuBNhxSoowimROZ
2Y0GdLCzxNZ+VbKCGFG6HINfF9zhcCeHguuG0vrp0TSq/AeRvHB1otMCRNovvZL3
EAvnQt9cQGvdxruaHYFfiD/HP9yC26xK+3Incsnzx4PpzCj+dXXljKRsUWhvN+cr
ukBshO4ioTCxj5sI34j14aqMFlKi0+PAqSn5lTgHs2kCKBNZRxPji9UKSAegGRvF
LrgM4Fih+jgtPZuB8SE3wZof8YfBgoc9MjWXUPtHLZg5jMZOMRhBhA1Zy2+pup4u
x2cFw1UJHGZ8PUkPvmfr4eGWdmfaduaH92AqpeiKUhvAroRt+W5j3MxNv75MOQqu
fHS3xzS39SEUA7tB4mk3jJL6wnAckS+EH7oWlskBPIRDOCOA2WL84vOweiA1Ps8/
0V2SFunn7E27k5OHjYL+8chI7JcX89qQjhKh+lwvdKIqOkwkbkM1xkYKnUrYrtey
+cVEs3Gz5tDeskdgj9cEF5F0zVGkwKI/Jogt5hEC6HedSQdpJ9+FRNgxpjsFNl5m
Ud7HhpMQ50DT5vwd9/zm2v58ALMJd7g2rSIlxqZp+hfQVAkpo1n1kH7dARNgM1jw
Xoxu7/yuRmngfLeu/dp7HqSnrNA/9G76XSWETsVFidOXTMxQyPhvQOy1QfmbhjeY
izJ8tYLj10hNS5SXjAqiKuxsuzOEXJAK/Ubrhjs3bJwiXRerSJlqZAq1AM9NOMgW
CYQvpKCziV2XVr+K1wK/cl8gGC7hXnnFyCkQ+oDFWzBm1i5IfJWblXDbQR1C8O/g
d0qbzRFtV5uwHE7wkmTZW5mw/iEDHQk5ZNlTJS7E1rlo4hX+2yLEuO9aX/nxpCQ4
J2T52zngcxzpTC580tMZeflmDOToR4c7Ttw5SWcG8QJMyE3HFLxf6uZP+V9R0x2/
R27mXjoe4fnuWYBH1myaiSe80kztnY60nTUCTcRxM4qLIzluVJsymBx9TrhdWHGg
8M/LfRAGF0NWe5wr8QTY1SLaW45vtjjlfthWApwituvxJUw7nUiOFIH7D2ZMtDbh
LABhKwPLobZfdnCU+zLa5TXYwHFb+BruktSZu8lZkCcMreGz64w9zzCMODwNdCDU
TvISF+VMwLvfdPlmy60/m77yVwZtoIPaVQNkXQUMACWWikd5xh54msR5sCHYHVzV
QCS/RUBDF6A4jwFrlnc0U7FTlX7WjepUEPkc+08940pFXw80SzsiT2FPnxm3vgF2
3OSssmEY57/Olmd362qyT6GtlByST5aRAetCSz2GDHFhZ8XMAdNlJxSCiR8POs/M
eiRFbCICGDb0fE2T8Tvlu52zFKNPBwOgrv7LwzaAMLWUGechfczfV8sxrDRVqgL6
5Z7ZGud2hohRZFXvXymXfcXCU47Bv+OZspKs6klWqsuTwaUzEeTQdqeoKUJuj/eO
wgkh0jmrLDvfXI8HLDJpzUNZ0Ivgl0I42ayagy/Jo4nDkJWQ/mnyAQ8kLBwDVyla
xx0L87bCZml52OGvAcMvEJ+WI8vKWb8zGqeFDv/EuB+Sj28Kyk2R8OH3KdWVLLK+
K9yZX6csaJ1/g0ca8NZm2i0DmIKkM1fE+TqocJm2a2+tzBCSZqdO/h9IjiSL6J6Q
gVuE8MgSJZTmoIHDixm+8bUUHT+rZzLim2Ipq7kXLPkPsed7FGlUDOm+iHfbU0I7
6b3Ebi73XohfkAfdNfLfg16+38tNdGeJueRMvZ44n8W+b+bRL5ttFEKSKyiObrg4
mKklq+UVac9e+eySu9i7Q+tq4gBAnAZR7RG6hCr+MKJLZz06G6aqcdAFngdTMdNo
1afR2UQmi7BSgRpKmYEo1yr/yayFW+2MF4myw0fEIhlHebuyu1EnCAhxXgiZbuCG
CMgv5AdWnNwaw/1oTvq5YPr6GKP24bXCGoqDyEys9zEIG98ZTcpcbki16OXqJUDC
GGxKUfZ+dZOJnu0ZBvEajkxkodugQksS+0eAx2osKTvS0tFPWmDV1Nuc4i5sE9TL
ryTTRX+3w3zBU9fSIdGbcJMTipdI1saEPACGc1d28zB0XQmmpYKrJ+D6AHUIdG8z
VuGl7siN1oJwR9j7RYK2BA0Ig1EbfmOy2DpEXDZCukYNnPczrGYGzTgqQjExuROT
lu0XWkr9Y9v4PCHyU2JHT+ajJj+eXuGSKoX+EKA+mkyCJofUsMK3VAZNbNtGKaYn
gdDWJsCFWsKd7qVdn7Nr7Ta9blH2VJ1zEZ1i+T8k477VaqQ8NMIkEqQPkRKr+Edp
xu7uamQo8ba8+0zAkEr3GZ7mp4yR8JsBvCYriGfd/3Rn5d1n1A1/rOt7XdJvimb/
nTMqvBdoLTFH5D0XdWYPHlcZUTyifDQO/bvcsq5eGOBDXW1lElx9P9miRCCSiyiR
AOMBZhS7J2gW6dktra72hDVxZVnKgwc4WvFsquvMvH12aq8m8LVB1DnZQ8XLWsEd
6CGqylmBIp2teC2TZ+S/50jfheKfcOw1fwUzs/mG3ix1gNBHVnxZGF6ptWleajFN
u3bn4P4gZJeaNUixRXSibBR2rsFClKNCfi6X2eKSSkd+H9Qv2dkgtAEo29jpzFOL
O94IixRJMhU5UQmKrnZlcmQnxdkaWe4N6MC5o65DrORTsYq7MkYQtEZWFKBD/iv8
z5evFnNcForY6N0Wil9BMU0lJJfcqL4Am2BGS3HtACrLPsbZn9ncaVEmB5iDbM3V
SIzCxld/PrIlVBDzl8uIEu7KRAqszgmWxnG9FEhF1kT6W8QhHpVH0YH1vYExx5Cb
d+cEIcZ/ARxeqRNYUVpAWwltSJE4pCy7GxINDOTg5PzuWKBfmuWGIBvVbmFkRUxy
KnDpG9XDRlu+UMZVaIeoF1NsNsZi4ZxQZ0VUHSrjJRLZY/DFfFmkb1e+qeWoBUBV
dAaIeHfNWaMXkFfQPsCluhcrlTA7qN8Y0Y7KKthtM7sr2Nzpt9b8yonUd87vIzlB
xaHxxxO5Oka2KJNppcF85hn1ELtF0XVXIvExrPsM5CWigFpoqF2tQFo1llXIAs8e
kwLi+HQuX1hzwah/SyFI2x0pK/zsRAb8jhM+YcnzNhecxObx3Gg60ec3xp7+nAy+
1BCOvtIr0k4/nKiUr8LoNcLYmmDLWVMkKaVsgL0cPwRoQwrNVzbfX4AjXl+YfU/k
JMypSzBID5XPQSplMEZr16RPChmhtqEPufZtAsI1Tshfh58z+pyt2CQAKnpwah7m
+6GcKdN6SRuyMWgukcZwemxbac8xj+tECn1C/dZyt1nDRR8OyfogNadA0vdK66m7
xdQ/6ojfo0DohXsVL1LwzLmqTZ+SQoIYyn6MgSuB2TBkFVAoA85dIe8ZpJ5GaW4c
`pragma protect end_protected
