// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.0std
// ALTERA_TIMESTAMP:Wed Apr 26 13:33:40 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
LRGZ6yqB8KFU99h7oalE50lIdp0FT9JedMJp4duRTaK+A22MgT8Qa9VBkOkrCZSN
I/pzsCg/R5GP3pm4M+DBSg2hcIWnp2zxgt5oo9NZpoYGIEYuzSGrLeVsfW4hpsVH
0o31GMFj8kJ/XJTjVQnuu83AeToLLFsfhLnHL58fThY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9840)
P8pYfB/hURQfgJW/RSyS4uSW4MEBQmu5IipbVLX5OfgZ6k4TiXo6O9kLazglf+4V
L5mdI7Xsuqp/tNH0rhn/6tJGHxymY4AXuAPM7qhYzCqaBQ66TeqYLt0Sk2df9WJm
myVWsv7Bomro46sZ06ZamNfHnuCPX5sivJgVAv63lfCOSahtKra2Wig5BLO4NywU
FU8D+MXYVAADnQI+b7B7+0xKnHogBfDUHpL4jbEsXP7jehEDPhfKXYmIPWBJH0bi
rfdiw2ab2GqmF+1ZK5VDAJmkbeunGJvPzT1pdcrEJRE5zqZuviHYOe9d5HdoGjPV
pg8xQSgJjdhPbd1q0BWUaip1kEhEeCE6YRXnSA9egVm6CLwwIhtoVa9a1/47oDrc
Pbu5vuHA/eLUxTn6FAufl3uZJ3P2i5z/LCoMBIPulntXk6PfRTVssZ5VKKuzMxmL
XqnyW9wbR74A8NeKFmtVCtc2CNJqXTozYdpFRBd1GKmJdJ3aACBFII47/HJzhuNp
Kxlg1opvBxOVP1DjmJAsy5DMzqO4lJWPYVrQuOyi7rH450tfymECoq2JfPFpKnXe
cjjcfAo04yL0Yh5nsDLIC+krjtVuH0S40J7B3WUDfprXYVVgZIAXzJG+dz7ScXcy
YznQXOONLhyndO4BUXmXZg/IB8Ek2vtjdE4Ud6GZzsRLYYdaKujSHvjdLukbS3tn
P5rukjiOY5pH82urRAYfT1EnJLvNuAvYxezzZeSOkSNd+JJwSoshAKXasJc5JmPj
zZCu9E3LPOUkmqmqz+I1/ZwxFlUunDxf9Zh/SRmk/vJFpjHPtaZ8CyMvvIMdr9Un
uLg8k4Ungf83ybp5XF8B+qGOqs0KSvxfqn38wdPAtr5EtLWZJ5iMtWAtj2hrbYYh
SblqubbEnrz1a9xFkaRZK0wiORk5/4n59TjQyIoRcq+PZzv/a0Kw4QJJFkE4brVs
oAi+qLbVSrQVbpWv0djW60KX/I5daTI7Zk/WJAO0BgvnkQ77pu0bSzGyy4nT7OSX
qUF6lOdUOzyYB9T+/ZQitm9GHsYuA3Crffv5cJ8YJ/5YbHBGcmSQCFhDDMWTw8aZ
CdnQFCaeBCB356rCgfITtYXcuJN4dBO42Be986i9SPzhoy9wuxFggyZQawW/MUz3
DRZyJ8PvYgjMJyAKHMuKGG8PDKnddDqucet1pdW1bo2jnZDsd7CUHraxKm+dsWuO
rjLnwAFwzNSeKGJdrBbPcaqYDkDn0xd0xOXx6TGLWVOccmhhnYlKz+/FsZhdiBOM
6QWFsoZ2Ze4MuLp+87kDgozurS+TGehU4WWAOgEqHMXNdq0PI8v7NiZnTnX5ms+m
yr2vuYAKAVV4vUJ9C8VIXcJ7fmc2iPPpaxzy5j4HA6OeR+pwdMfc2mb3VGhnXT7K
wSuB00PBWFtE7duGqEeaN05h+dauKZAP5Yjsr9SaZj80JaGw6DAl2Gx/SyIckWGt
EuMTs6KkqJt7pUAVG/VLwzCHzwIdWiqhktfIC14hzOMN18N1e1Xg5T8nj3JZIBxV
FJvStzr1gfP8H1QOPNvWppx/ZysQh60+/7qby176l87jSybeMG7Hg6YOdjMjRR1q
XlR52r8Lcc5uzbu82GUA4/00KHj3ZFKfsoy5YNNSWA6LzzTSzOkN7AfKeyrpKM1v
sUf+5PWEV5robwAIV0MV7+BCM7pYCCLcD8suhzszthJsuvFGXd8xElutpUc5qcFz
FIKWazNWYjUxWYV2KXy1XP1ihkPWBzFi9KvNnyd7oH7idgrbUGdqV88J29LUEIUc
G1UxpdLM0+oMF8RplcZtXCHcQddMIa57TLKOSEx9t1/1E6hioG8NzgatJ3GB6icL
ggHWlehLlYd8jPy8l86QK0y/3M3pWBZ2a/yRsUJO4WQdbzi0zaF6GrlZRI05yA9T
BklA5LNJIbMzyfLtdWZ71i68i0bFnoGcfvHG1dTBPR3hnKHr/ct/PZg/Ze/ZDy0h
RfuwASyjb9rzXPn59F6AdBhgipY71OVnCFSFkbTelvoVE7qjBsuOq2Qmgy+Ewdz+
vXydSlqNy9lXMppTX8UkouImpI1YiJG7iXvBmaKYWFwh3sQLRyFvux/35sFXOBI8
YK1CtlzYw0krXxfiYOxzuQGkBPYLVXd3tIapDPtMKVmHuS9qLwUKf5nUeMoACz4s
wlpgEQut4vyvc4n7TG5z9H4k1QjJURusHpeXWD0y4admxtHZQqT0fU/0U2jTxk7N
/jCunq6sRhlNXAO2GepdEIWw4uUOF+gRZ1NMk9m8biaUtMGo4vCeV9gqxLXxNagg
n+clcQI0RRya0swUGhNUjzaoOODi0DVnJDsZgwhjKQkOvzhzOE0cO0Iab4s/XiBX
1H4RAd8kDYvuVlfs8GW+x+5zLkV+ZU8hGs2HF0IA+infNxF1yxPyeDSdMD8WVIpm
tD+kH7otMsKSPDHD1ttv/WL2I+V1mj3m6tJ74A/Zntt5jtp4o9CMw5ZqRKm27q32
Ld3zbFKMamZ8Lx0JMYwrRqv3aOwsza98atJAkqbpgwhj+6fLGua09JjejWWfbn9g
rqqK2yTuP7BvOZnu3lCWynGNekHIeZkeSl9UZ5t5zQN86QEOR+KUS0xlGxzHgnl4
+afqQfcfdrMgkq8QdG6jwArY662X2Itadp0eoYElfzK19vqR9700MXxmqEGTk2Xu
SVJYQHD+kq4+rWdCCTx2ZU0IEEghEHx1kxU0EKdl642+6u69IONTDMTWHtTbX+ke
TI55SVvDx+CcFP4wNESYxsiTa76kZAscHpMRxMb5QNRnbmGzLsPikHJRecT/u6e5
AWPzTtTUKYuyojwozCDYpVL6jNyQw6PYC7UigJVoWmsmTFweU4SSq1qNpq68LXtW
anbE3M7v1+GeESfPJ4LGLAQLOtp0WIZYsvDcHZx002pgSca12BpDcY6i3hejRXLv
Py5JOSnFUWu52W0KWCj/RQN5h+v6RLr5T/p+zwmzzMF3RlY/hFEV8P+kjvJuowIk
nxAZKWEMDzBn8mBDrMjbjLvFey7GmemJvrdbs7E/Fkp6drbJJdM9ic6ZekZv4YRK
0QXFwkMIjvViPrHFZxufsnJoVOdJuAZS0eNcuHwBzOoor2Lw56ozeo5rmvplOCbL
aNPzj9STItBUv2PKO8eNMRLQ/HHVJNmP+5pOPb6L806pM4J9fHLrepYrzo+vd5Z1
A5qH7e+67CY16rBhxUW0Mo9iIAECnmDRSyF09Q8A6RWm5SDpKc1v0Q3LFvTKzHlN
XK3mCTowayt5ZSBnV1nRWRaXmmfK29fy3y8e4C78nPTeSbaOcKTtb9y+AYZ44HuR
9GLgpqyQyGUJu1D9BAjpVLacnXVnLMIYp1Jyg8liXfZJdQhpwZGbsEO9J5m3Ncak
1+zMBlq4y2JJVIGOKK4ohpjB1yd7CsE+BUkSzqr5QsvRnjisG55sqcavADqdv84S
jcPYvc4PWaxOV9oao49pMLCOb8y9fvDL+25ZoApABPmU0d+6hNdFugQNRqb3tFe4
lQr+Qdcjx0HBmqzV/hfc7UZybq8imPHpHqlF8ShMatCaLMc6W6zMRltLS4kSXW/J
5DGYStuJpr+ViHObv/eAbGKEGqMcprHysFXsQYpj+EQ28ZkWG44qRFwTW4UWoQio
KdDgb4oEHtXGeGqWOEBA86mG+jtiyWAjRjTwsB5EBxiDB4GVw/120RL0opPXpDli
tkvnlK5pYyFK2YcqzfNpB73kO5kRiFCnNzzj/wUYb8JlUlvcwYXjTkfvGq/eQpYc
3qYhUdm0a5yCNjrtOZg5naZyjrN6fa8x8t42p73SN6ucaF+YotU3xpdAl2rMQvtg
VzGiVEstZFWlHDG4OuGjPSODn5LmXbYNWdsdlWjNw/KSGHik8GJkWvvryajc8tLM
TRTgjI0DG+yAqMVQWgIKbcPZnxIGH8dOH0cJ9NGPNAK0gCesU1TEe9VK7j6ka/rJ
eCPBCTYShXCNGAb+9CokxnHubQkYC14f/CrWqt7nf/RZdZ8w0VgASwWiAK5sk5q9
zxlyVi4864hMzAIbs0CN3C0o8M6NXh/LPbgHoNo3CB7LDuuUfM3jnKsOqeRTiMTn
JRDBJql27g16XvxdFah2gikDPdiZXffglwlMxw3mTrzhqY+EUMtIJpqHIZbrlL25
u4muxFTQfepIBr0BYln53NqknSAbRzwfoy+lZ8J3rtuxVeCGsno79O9XH50VjHkO
ox6Y3N47zAFa7Fj7rd6SbCpqQeLcr+UU0Zn8LKNWbIehn94Eaf6FGxgElRyISGu3
eP/qmYCVWFwQ11Ekzsw72lbJlvYEvqFeroE0YWil/rPX7vfF4lkPCg5z8gdeZHNQ
0+2XzeD+t6oDhD6Sz4NebUnv9PJuGyXVdESd3mAUfkOOFgOCT0JxltUg/7BdR2iS
F5f/rXvSZaFohFHFj2aXMze+8pQh5v57+YAqC0s4ebiocZ/eE7etpyKC9BHd/oL2
lqn7shK3aM5gPhwRAQT8UvJuZYyqQ6+9kZMOXmBPDnW1Z5PmKZc/4LWOME+fpjkJ
zBBymPXMRAk/xNbk40RZDwUPByq9Go4bvYJTDez45BKGCTplNVSYr56nesBy99ed
q08acI7ctn/rToaGiS2RpWfnvC/SK45ligAY7z52lglAeyJFOON4aYnjjrGrVZRq
vJkBzsP+cG4LV05UVAoCnGLykq11SZAoCS1Z85xAj5SzR2V8JQyfBjiGhRbD4LUe
MDNqSYwyuFh6o5YuO0ckciF3d09vuA3o3esrj8k4y0YIn3F3oi2AFCIiOa6Ce0aQ
uUw/Im6XVPF6GFbztmB3w0zRpRhyjE7gxeCNKfbl+P7U5Zylgks5asH4W19k5EXl
FUZhdlkQSbxMlLuaoTIfwn5CLxcaJw+7wvfoVDg0HBhi0tnt78hqoBBfEv419kXG
wsOQQTRiJuVo16gpDcJyBeys1OtLlOFDDxHxPT3h1nuvkwyagzOcinGHQrdjOVEZ
lSX4Ekvl1TpbjyN+jvP1fb54k/w/O3NMYSvdwWmOM+wU4tq1ODKyIlJmqpVyVr7O
5i0f/oVEe948qBya+b/MvdsdZNmjlmRQjgbBf/B0mx6/XEW2cC7X6CsRXpFfyuMf
WAuzlseuOGiG+0S8QYkM3AHse/SnkeCTmnZ/wcyc+LnpJp4uRssJ3/+nIRdQ9WTn
WoBvwr01N9Gs7YllKqUEVAQH0y1DmtsI06bk3BEnY400406nQPJ/eQP9mqMC6DHa
0t7NdiSd22M65aNDH6gY047qmYKGt0uNXhQ89dAbMPTc9L4dhQw3zrzlOYa99c+f
nkwgX3hlDiONkSyfo4uobFW/taDlkZN6jMQTEhQWc3fC5ljkbowYssrFyn3xm5XO
pu7zcUFZ6YqrzYvCmJXtQqagcUFnI2IakUEI9C/if8+FgdRGbdDwxphoDOv8Xqnl
Oj8tQyUeVPlN2FcOq/o7cwPOB3ygTwLztPYm1BPtddncLYS/3DEfu+PEA3UC37D1
i/Tap9PGKEO8j32ZIy6Yaf7DARzg78DocoH+ApbnmaOlviRWKvaRHPJJ5if5RNsc
0AtWdKg62/1f5NXgpxA8f1mbsj6l91J4MU+ltKG45IYu3Qtu0xdzngNmf7Dv5WsP
Swdys4x1XLwcpdQDO+X/57etsFxZmGxGlJYrj8M+90aWyt2pr3+1+hX3YdxMuCZ8
GOnsfJF/1Rg9udJfMR8UzjoiwLskiYTCR1qETjiQ9ZmIUcDWHz9z07gioLANFP1n
CKc6H+YXo9rEqUcD2lVVHJ9l9zMfQcqI1zO65H8WYs9oBWTbbYN0fco00qYpeE31
Lc2NCPMaEhX+DiQqyjLf2K6rYb/vTQM8qW4MviuOdfA/oJQ83rPFzdf3GAWP/PTX
KYcLlU0O4NXk9B/Rh9DmwxfsEf4KDM5BC2T58gR+iv2eC3vFQ0azrKh0l2TY79ZN
uVFZnEK8fAClvPCOYORlYwedlJdBrn90l/iXcF2+bcfaiOFBS4zb/mmQXpRbTKyG
9At/F/jZ/Ovh3XMmHPamh/efuiGY6MgiKcjIjiHqtGq4VYBn6VBL0IeHaxlV/Jj2
OndYs50IrPvgB2G850kSB8ZGZKY1kBLiBaNKBn3auyitE7A4Y5k19OC4sfjZvHEh
6pD+VinHF9jVOuA7uUXLYYWPtTbPtli+K17qMbGlTWRjjxOvScPMiJYz7GHwwwbv
55UXyrOJ0oFhMGw2ogpnR4OEcSzLJrupvWGsTIuCYu8e3St6qd2dzxlX+rOh7iQD
qDzn/A5AZFxpe79V1yolunGhZVMF4efyLaFRP3Ep40FSGXdO5j2l769XeCYUYWPa
jU8QxjkvbyRWncJOpfObsG9ZNuuYFDexfW2eIJkvXFe4hWFC9itOLSc66K0HfNSF
lD+iE4rsUP9Df6fBIt69Kt+K+WmfYiecUFgoC/aR6LauO4X3H3WP7eqXaUdPhCi/
b8ICThHCJkoumRnCZU34SwAV/SwembiGDeOJ9pn8VuA9LLC1zHRPknOt+xxAKV38
gE/QMVzbpJ2QI++/B3QRAvjmuSglEozhqWZSQ0rMeIXoamIzxLC84AtXcl0lfM7E
8W03i2HyXWkB5eGyDVVAcDO7VJw6mb3ET8UbjIdVQfUUuemxYF6Zm9q+KqvkHky1
QIauuWwUMmxI7iHPaoC1xN4PhYu98flzsh6FNyKJiIoSmTwF+kfk9FiqbeWx3AeM
8zTgbrH3CMz4KUzzouEchad+Q0bqz4i76qu/eoSFOh299qzENdIqfASi1kZx+2cS
4zxNiWIzpXkGqslYcFaAPLBPL1rCLimAQQTh8313HbqMyiZuubqnVO5sjN0ZCHR1
r26A41PPI6N4CgDSR5TM6qUeSmlDpIMqj8ceVFSzFa2KRTIlXiDd6P4a52u7lHtv
1SwgvGBvr4H327bzX3xmcv//fVRzrQDN+wTX4vIyAVeL34K4/XTozGGCGgiHHxXh
wA2T3UWTQLJp828OVKBLynHUck4ZZyVQvwYDHq4+flqxD+D6y5Yw9tcfYeeqfhOi
eXDDuJ7oqg1NNDpf4KMbSQtOmUbxW3AzXTWB2UVB7gwC6aPf608FlJQ/VhuF7u/H
x2ZRMZYnt1NrDl60CXDkZRH079FxH8rphyF5gZiZx68H23+VHTOYY8E1WqGyuVaz
OYtbE75ifx3/zerps57jAQeGdalVNH7v6Eg3hORjUcOLffHuB6kmr30I0djeaPrB
we4M77Em/F8K78uLTH3RZeMVGV9fDoSHEWv10TM6JjGqTiU1sw+2gtqnBG2bL6BY
Grj+FkGec7yqYpTwoyslmFU4XNsV5KVRGClfNncn579XrcDdAmIm824NzE6Hwqw6
NYapGQjhUCiIJY7NsNRlSBdzFv6LV4yjkvjtkaG/Zb6lwb329S5zb6LSw8FEHAwX
c+eQKls9qZjsAJEZ1IkLqyO8EneryTY28vrGp956/z7anovYxwSrLSg1in1YG18m
7wowVeI/5s4R2kmcOwyhWemUqGtAVlvxReFdW/Ii0jql0S8fsK737Rnbxt0FFPuz
oopx2penjq24K5bE7bIlHJJ4V9wc5yhBE+xymu9RptCfUsPveqtzkF8LdzsIklDo
mGtrs+yY4hw0fg0k4S7tu3Uh+AN/tr+WENsX5o8jlPjPw+uDUREIl7eigbVFJks8
0+SRmDBpHd8XlZfSpgWvaA/HMnPU8skxs55w8MwyBGB8ZAiPonn8neVWMJPdnRO1
h8N44/u0tijcFM6pxW+A4W3rjWp+mRM2YIqaj5FBoItOISKkYgDTSF/HflKYD7pZ
Ccm2qDp4EkcdcXupKSQ8xZ7pCofpCICBPGcwOO/gm47pGd1cRuUgKc+f5GsawgoO
bzUK97ZwG/XSY+C3NUlDn3qn3uEeiyrsIw/Es/6f7MRHma7F3GRMYJ+h6EQpfzVt
O5SrGlkS60p6o3uxevfTjaXDbIs/aAs8Ry5OVAu6L0E1Sy8i14efS9HKmDcixleT
UBg+CrET6WI/UinDa5405+89loE9OZwUIhLmw/vUlcVNU30DN69IgSlIUBwivp28
Qn2wfoIgBu3ATScqbzC9HRFeQTHCxFNp6wfSBpXfGOAWg7qcQVVEwLUoW5peGsvL
38hpHhFLCVMRvXJtzyBg6lmZwfaC4YOF2jPG62PXD1qrHphBa7b7p9oUl+1dKZJp
BzFVvyt894sPyFID4iY4lXuYt7cT/Vn8Au/ZnRPKi3SGB+FsxqKd0tG1ACXgnuOI
lfyQBGi9/Igo6ywxH8CDy6BIITxdYdVHa53J3tl9v36zkm2GB33E/imPNEPoETNz
nkKDF49RrWjirdpyFsYA80uTJfjQ5BTHrerId6QgnoNKt5BhPET+TNF66LrUAxe/
V56osnZ9zSC9I5HAdnkMgIRUWcJDKNd9uuM7O/6lIIvKFkyUNDygMk0w2zJV0PG+
3zl0ywPMIPvwb6uuIS91XjzjUxTNWXA6qPObCdRsZJEOszoO0sEWOAxeba1RpjnH
e+OhuDA+4yi2PERJqPvfXG/Q1/8XmknhCTcR0+xCJBgy/XZ1HIy8Udgtz7+9LeJ1
isGw7gLkRQRxbCkCXjwOoqG2sVMt5wQ/Wi9OCCBFVEnSaS/SX8I8Ta1/pf98MuA3
08OyBWvXr7hxBUGB0pirmG8lV3aanajl/BZPjrgCs7MjsIejU6n+07hIAtmH9kAj
aLj8CdgL+cvu7RLs8CBKergTtENRXpMUUbTKevB4vjtzUKiil/88bLM2sk6MCkaK
cwmJzBfeNBPtTRqA/Gu7kR7BnQie12pZeeI4Fe+9xxB2VmJH1Uoxw+e1n8OcZCyq
do13M5YWMJ2ve42rkv+DRzZSP/JPCRnduFY7f3sz7Ds7i4g3DWah6fS0RB7H1o3O
F48AQuWJTgWKhgVpTzz0nDZ0RJR/S7LrYmRcLpwCTWV/LwVs9x6HXIkf8aaXxWSB
WMxzbYQ+Jfmkm0uaFxL9dEYCbuIK2h0E1YHmO7xukgPoKzWAX46XBtcyUF7eoy6o
leZj0rbgH8j+PNZbegEsk7YDfFSEVFxaZTONJA2fQ/PLlzow0F5LFfLGefrpxrWP
Eq9dsY9n61dNuk1Ll9B6Nr3XdO5QnsrbirtzwNPgXkGSiMrXBEpH+FJ3MilPM8xV
t/GP2eK6h0mJrg8PXsdf+0uw5S3COI0h+RTf5fdfNra6biyi8+ZA7jVZMJhBJcAG
vzdrdXyJpwZhaHIwEyv4DgHC8uEWDpK89R6VYK2TiBf0qd3SV3XuYS+/zY936XrN
my+cBPKTHJkj0lmPqe+7Z7StqbOTJty73BI0qlEiAGYNLGXTVCoYGoIbwBh43BA5
WLTaZtd1EtvWbAp31zkSVEr/jmjHKMeccRggmQaBiDAEAkNJv0uDf17Kl0cUrTrp
1Ns9W2HZ0LLZuB0fACen0iRRrVccRMnWnUMjrsDUJaMb7oD/m7ceTJUOMk/zDptM
fxhrbeHOv6n3nHKWw6WEKHg/bJUPunurEDY1xLgz2zo/iWEflRCkCOpMnrtz39tC
P/1f/9OYiSk5Z5z0zxa0tzSrkh1gtfymk6qFPOCDJYTLx22EtgP+dy5dIcgDhxD+
G2u6aNUmcQhEENPa02Ai38biePShVzqBA1iYpulmw9w8HoX6iWYERFcNkLlG8jUM
uj0K+gtaXK7vqniZN+sY9oyeortrZ4jQCbuRTTR8xV1VzbPh7u3fYqKh5nazL0dp
wcJrUigsISDuixJO83hKmXrendyu73IF3NnW9Rg3QkveBVrhPJvoPFJSPDy4eGMb
+KiFpgrK8ffgHuZAFkuREyDC96HhgVOAPWFzshqFT8D+IccxaMSNsLW1UppBh0e4
ME1V57BDwMnl2UEEjljSE0hEuwUS8Quvco546/dRlfiuYJUd5JbUYQbj31Iy6VKV
XxtiKvq82eAU8OM4L6VWUnqI7doIRwnhAemwap1oUMsWOobh7DwrJmirdnuph5n6
54gNLmwHuxuV3BednifzeuRK2qZIToSDqbYPbBpa8ukjbSF2t7SZNfQwNmokLhAu
rEdgQOVyljAAeYL8HAmC/KpauNu+n2TfMyuWBvVVvvtYtqnLr6+y3AJ8FiglPoxp
irq8oX6zG9tmvFvfK5UxBx8o47F0P5EEsy2WkIwi3FHfD5mj6FHkL+lmfSiJk0wr
zovUi8vpCCFwpVHHwZW+Rhf8QhJx4hsI+wVC8vzqz1js1uHP4HHrtHqgT9fx2UxB
NsMAH6jDhhUqKhck965cLN+Ga+SeO5SnHLyjpObb5V3ZTnwwfvW0mx68hoQRg/tH
tTxvMiwRJ9sPh+Q/6P2aZM8yGapKFD5LfOQtk573VxwpMrDPEEj1u4RBgrcsmy0f
v82dtfPhGImRcy5UeYMkHRFqqcBkVjCZfRQVCnfjaksbLc64UMGEIaiMGIfQUOSJ
hQMAr2GaAFULxyv0Ki37+5li483sUm2OS614HWUZvPB8A//5HhaBQSY+ws2k3dRC
0A69yH9d1XdxBYIO8aJ1NgEUokspId+o5kH7k51DH4M2Z03I3KyPUybmTyqAF7zW
C69v/EsVxk5X/3Rk32UuEFcUZ1fBLFCAPtXGjvCw5SNahULtuzJnNms0kZQiLz7r
RT5XIUUOa2AW//++kGCXQivQazrHDMht5S7aE+FDQGsaqhv8S0gp1JjBJZYtixtC
PPmz0L6oYMdg9HMoMJ6f11rDIGF4KdOjF5WphQfN8IPYzE3tE90PKe27MQ2Gt9T+
VQJ9b+PuZEEvQ70e5yO9ucyS7c3TcFWPU/32XAItUOkNFZxF+GJ7BQdCkuBdNIit
ydE3K42TchyOTxuMIrzVQ3oG1biRgNE1zhbZOJ/VHq8vGtzMghPQvPTDQFkQRlhm
6vbOpLu33l5CyJHxKH1PR0uMji6TfW6D3DRLzIU80Vx93E0BvqA/HhzvxX6AivgM
YSA3RVYtAqAPJgGjDol0V+2qgKiYq2d91k+ph3iutBhU10yn313aRgMmUmdV4kQM
5nKJYws7/GwuYPsGaKFDJF7+edm8VMXLeg7hBqOurEe1uZkQv3fG0pjIwmwkC7wJ
i6EsA6UnhsJRfilFxXOdw7KQ3AAzbFNAl0o2JTpVrGZp/OxhYK+DUkJDXi3i85ij
mqdAZqKFbaxtw2OKkhPF6m/pUqCZAtP2pUe7ktwmpHpdAmPWUd3zqbEMZzFT6sQh
zjTAY5WcsaFPajJ485rqiqvALLzflsl6RkNujiFnfWZWMZ1N82eZ9tvQ7VKjP1io
vKPhQ8qGvgvTuNwEdSa/+Ht6CvIb3WDPCxrqnIIKVAK+t69fHn1w9LHVub21HKTA
JGhK5D6OnwR3kJ1QbNkgq6Jdk+uVKFMSOh5GCVfwF2O9NF0asT+g3dddK57IGhTg
ah/+7LuVe3988/oLl2NDZNS/Bx6pHbHIVtybIyFlqEO2bSMroD6iEYC5DdyPDXMM
DkIgdotrQHLCdnTK6zNiCKvynCNIhshQRU3AlafYprgyI6ghhsEzGBkLPD/TisfW
S8JCObSFEscB3Cn3od/5yZUw8+qxEQQGcqQiTKMVBAoeqCA3Sahm7JhFDAVLkQA2
zf4KbB7d7IcOGT6GUspjT6d3ja9MoQn7gwjcaAwQ4rE4jdUE/+bjff+k4dbZEky1
r/ZnC4mM3WjodCZKJOP0qGxmTRG9qllQFaS64L9ak5G6VM3xoz4Vrpa0wI8iX27a
ndXvWzuYp8nlRG1EuO5ySfzhWk/Ht8tF2i4VzpGMjKrGxtTjuZhJSlcQqjLVl2Km
v/RSl+4GoYDbsuJjz1j2pqwX4CTQ3Whv5K0TvjIaJZO7Y1KOwSx32EstNoq6+NVb
5dRVLWuHUTQMYJMu0lT5gsxCg9QYzyTMSm1TbS3z/3InP2ia/K+uc/H0d5ieeEh3
Qw3DtvqoLa+BLKHT8r/3supoyWAxMUC83nqcCp9rNel+7gBkFE+e0zoNoRMvLTSm
KEarPEqcTBW62grKKzpMtDBlsXd1FYD9ZkVIaqXW4ZzqvHflueY0pPnfPA7amfLT
tPrex0EzUn4WZlvc99rAirqTtJfY574MxdGTux/it3dk+ip6T2ov18NpXqIYCI1f
SaDS/MijVpc7MygjE48t9PJOd9xBXnizyqLV95s+U1bzuqzk3ST/6J153t5aDeB0
04lGYynSkTl44fW3zPnxlf/t04lxW1tniQlHspf/fp0CbMQ/x/ls+txa8PRdvZkq
swZwkxcxguocdmMcj66/QOENdxCPO1NzUqYXm484D4Px6UVSYnRB/Gychqi2eRI+
CxrbBLE9VwqQyr8iprrTCGLNO6K/3o8vHOTGDrdxDR7+nUTgC3WH284XoSBeDZVE
U7endaxhlbkFfTY0BKIlOdWuGK9KPZJFlC6PoWHJPrbKvuRWzHUipSAT+IhObOqA
q8fKbHBfeRYCsNHZIOkrYwgmiu2+lESrJPyYhj4aKOydCcdFs/2L6sQiqg4OYn7m
bHtwLW+DukKk+OajPsElDfA5x1dPXvEOGhp3z82g4KcxGlWU/3UhWZgdR1s8lrZV
Ktfp5Rr53bXwt82HXJ672mltEDCTrowzzz87raoG/QMf6isa0FZwkXxBza6wyAH4
Z2l2AAGgvNMR8m7XcwHSWWqGo0JaGS9rSsmWTj/dyOSjd+9XeJn1oEqQYwAq0G83
whT6pamfEqqvW6AqUHbFZUtq6FvRUQnjDL1l39SYT6vK9lvBTdsDIm23EASnw+U1
ien6s6ueInJwHZIo1G9r3IXM8lSVaNioq1xpIv2N7HYmC5Jhlr6L4HmE809rODka
leQH9HTbffhWPrHdwJEtd5R4Wk4BcuxqiyzcDUgLgKEfvGK042Zw6DBUvpRhQ8gd
93VjysG+tVkkWuLALeqhkZYqA3ODOnLYsi4WSdHTdmkMV6FJZU2V6FoOO+URVTwv
ThO/UoqUaHPnJ8ABMmX2YTQPcnD2cMTbDeWHn3shN20RA+a/jacqu0heCgngKOQr
BBnoHESzW1RHV+osq4qc2BJGCsjiyy+Jkjo4vWE2pUgYMqDI7E7IudZtLS1afc9G
2SJD+WTQzyMtOoQPF8WlwMpNYJ0khvAKPnk9OcOCHzyyIAEMd80ethIaPysEHgWc
`pragma protect end_protected
