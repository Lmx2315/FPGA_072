// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.0std
// ALTERA_TIMESTAMP:Wed Apr 26 13:33:43 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
W4MqI4b660brfywGUtf4iI+AK1ndmyrbC9hwbF+Jvnvg8XTWqxezGqBIFIIBAYg6
5JLGKfVUcr49+cg+BIyCAqk0A183sCnlya82fjMYkRf+ZLRkd+hUp7F2ZaaINBY8
M9yRCy08g8fSNUq5iOIEvj8IWQjoSA7latdOZvf2LWk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5408)
6aXpSiVePKcQhqgiJhiM9/dDR0Josk5tsgy5Zowx4YfbHmqECWe0cXyCOX9dPHMr
uu6KgCyT1djuacTQEcu+M4Z6iBru1kh/KXdNU24FBGb/pxxQcIdBub5QX5NVzG9V
iVrb528a/15eHUapoYFj6OJOv2RAzNXD4vOjGFRg5SIiExuC+6fwamm9OrAHBVOY
l7wa2CX5DSUXGLywAf5m9IuQQtS9wCYUcqwWh2mIGgaykBz+PnS4nNz/9c00wCEt
Ov9B7gyR02SZrKI0rfKsNBYv+j2CvbT5+ITTK03Ndir0IQK0W1facpjV22EJqlJg
CORw9pB2xExvjX2280Y9OF0XHQhpye2/V23nUMMHxa04bcXJzVGhgo0zw6RBi6fN
pucSTzhGWipzqthIl1+3WliYQtljjgkpr5uNsrcUT+g4H0nhpUcilsdrJ+R9PQr6
u3pP2HxFvh2Vuf3h/MUhSz0Zu4U1IkfeGk/4TGGcsDPHzAEI2DXaw5sjDje65wAd
xmeCY2wlvst8m+rq6JKBmKmswovnZW8WdYcewTxr0Z2qf0qgbBS+LVbdkbru/oUI
oa8wyFEygcEwb9M0NGDv3MJ+oZaQoAnBO8suIoq8DRf3fYxEy1IkUpQVgBkmcWEG
o/K0U7PglZIbztlXq+2UXMNkRSf5L7FXVuzec0xe2WjJBHuK2ViOfYFSqhQOptd6
GBUj2Ra5souH89ukUb+J2XpO/9OBXdAfhyWvcWkTsri+n5JOWcXQNrW5CsUeBm/E
8GbJxP7LvWLN1viTvmvfpaZtR2Zb/sM0E1Abt9TFHt4t3cI0QfOUeS6Npvn/vvd2
lzn7o13dgp1pYmn/PVa/5qvCtrqwe/QBHNtEsKosPtF/m1s4hFbUu+XNA49WdEjz
/2q0me67OZze+KLMLc4nP9oY2rlQ/eFgcU5ly3l/5Q9ueJWuz8K9i/UIu5wlp6bK
C9DRV4hWRnsUVqJzTavjIsmIVPN4wrlsZdwp+2/fPvvb6qEs1keUY8U1rO8BReae
5uxTKOOELq5q5gnSMBDZCuuflPKrJUv6HeJXrrs7ufTl98VznqpSDIlsFaKl+ZCs
JnbmLYiRB7JY+zv/6EuZEyXU7YfS5AhmNRf8tEkczY6zQKq9UwIsfk84J2NHaenP
Hw2Q9DoRsA9aQvyzsmn0BY9oieLzEvFSEdangrH8VZ3v5SfXiMIaVfR9obYlCEBS
v0B7jjWzPDSQmi7wNeaarpjqFTYQghPGAiJLCHwyEB+np5p73jNfnrsIuqRn2iDT
eYsDhYeOmnrxlT4u53HDXmcwKcUm9ij/5shpYnrfTAvfoK6wrQ7c5nHzJbwEUBdG
oERQ4za9MTkJrkbkM1KAyWj3ipW8Vx3ok2acWQ/eG4pBfHROTGUkKWM+eKqtjuGQ
qtAFAnnXUiidZBD7ye6ksNFROZ5wIonYsQKxRYywRQISEDbrGDmwCWaRY1/t0VeU
n3j4DzFhcyR0C7nTJCvU5WJv9dTPf/x0eRGanqE5boJMIHlt9S8yQoSF4/aquldH
1jZZwg3BH4oIZUN6/WQZ36Y0eDU4aAhIYEyRo4mUXrzYKCno5A3PR8my/J7QBmG0
xIFvIdhKHIWp/Hc2V9oJb/58IB/bXxq9KcmVd/toDE3A8rKzz3LF4K+K3KoXumG7
+vKWDhlrhsURJVy0IR03w3wSER13r8IdEpScSIYyZiZwR3u0YMK7dQN9wrockX2i
SKXgAWVYjwm6Axbr62MLQX7xqM9mi7fazFQAL7H1pTazZ7Mq9eSW+n92KVbYGxdr
kqxYldX+pyMVQg42fr3e2GFJMNBUHbiIY3+1DsCKsxT/wysWHu2mJw5AxeW6aeSo
XDzEEYzkoZFCoyfPoTAllfiCht4dUG+nGRHc7Z2ED7cOMqF+ibKt00sgJGPCfSIS
LjCL3CSJfLiiBV8kj+NxK2t/qAkN9bXfOXOYXPCCbZWzzpqZew+5PCoAzxts05KT
VBtzNoIT3JU8k9HASlOFJLpJ4tvA+TbYTSOsES8EjDbN3R37RNDhH3sjrCeTuUxr
fZHa9QA5RISKkuEnGlUU3oabusR/eLddnwuD/omr4zpj2IwXCivAbv4Ao/JYEXCE
ZqV44WDEZAf7ljnAJN8s0l+FYtAdY6GDvQOyCvzmq89OmuLo9PpPkNHQOKn5QJ3Y
6ETH29/9+hgQv4vM4omF3JjJvrszLtwuas/cgT2JtgfexmxCk+fiD+kRWJ3pVecH
+Yb5dE8aaTJ67imX+mM2Hxdc9VEXShu6dG6K/dBAvB9yO4uIyjCDw04dfsF78i7c
v9sW8esC2/4nSvjaOBiQmQoI+TB96X6bm2nvBDU1AajKtxosnQqV2mLNehEBN63I
gOM3b9lcDlHoxJ1NsYodG2hhRP/EYdDzpdUFGoZ+qXXseDFra2TMUCvpBoWrd3Hi
x0CMw3VRPpkWkxgZwimT1UkKJNc6Kov8WnzEUi8vdLxo7jdn02FR1T2mHNCLKxPs
Iz4AHNHt5KgrPDmMkRrFN0Zv+Ja9vr/9A2aAyMFuXrLjMcptk1HwPjDYB8rF/k5a
Fp5rUuZWzBnPgMhQ18F+A83ECCU5HZ0EeIOwh457q+3hjpn99OR8mokqviMOQEP8
PcB//omfaHwljVyP1B2Yc/N2Nk9A/pY8dPW0ljiFdSjYdlpEPgZqkDpRcckuE+jf
+Vx/fTBOSRzrBBaBDmyHgg5babLCyyqbchMMh2SE/KGleNsg3C4zxNCnrU+AFmzB
mKOm2catEXPvH+kxI1m4/uJdBUM7jCJAlW349LkHRJWXusRwYpH99J++FvZz9R/m
1crNaHjfeK72dqghUU5AhBaGFrWB2CQ3EwtcNIo10LWlz7BBdVa68BUB2brITup8
d+0ZbmZJ09a2wSKDGi3kt5Tda7MHzCWLoLqT6ypQZTtQx+XVGunx7knMcVJuw+tn
BLVAdIRHGga6Q/GxmhXF3iirWk6PSdn63SWdG0dDYCXwm7xlvhE9e4Yh+O1pGVJu
aY6vUCxPTdF7ctqCUDrTqKXkVVMS1sIfnF0QScxq32FGFl3th2yHj4wy0L7vsj0c
ITOe9eu8PbT6Y4xHbNBXoaGrxMYQ7L4dpb071wkkF+XjPDLnMI3msTrZy2Pl9/cn
99qi+PdJESAAqvXKQgmhaD9jKhlSqPESKh7NYPcQTDi1mbZNlP5CYXqAlwf1FaOR
wbPE/hMrdUHJuBW2uVRrZDSMNP1pwCxWjAmS+xITbD0KNfesZfvEOm4O615IIeSX
N8Uj1GP/lu/l0Rild3hm1dDMIBo5dvhwhd9ASdxuaaShcNzSSeYzHKoHLAd5yr7j
TM9mquKJMXEFLC5lyYZVbuLpxbI3CGHG6zjqU4JkU3oS4i/ZndkZBXjNY8QJ326k
Po48aoWKf6qWTGxD1/TSUEHKy7d37kW66Cy34Tkse+L8cYovaTanJXl6ZX/mnfud
hIC9FDIEjfDiJAYQAscvrxRKJcBgNSIKhx7+kSVQ6f4oxi3thWNqZajhTsHhYk9/
vUts+KncgQHvooZB5lPZscLyZ3F44e2frYJGjkKRjTqLkRyO7DwWcSyrC8mahVFJ
sgk6iyToNhloL+SBYidVxcaMZnTHc6h6uTv6vG/kfWgIEEQdUaeI6nXn6aYhpCja
e/K7FrrCJJayXvR276RKGTNkP098eMu4OuDNn250qfGrWPIGUlxrkNQ6AOQ7SIOd
WSkedoRPfT33IPWImzi5dfEREM6MBHDT3flJsVKcOwKY4sqaPHWXyovkWNKxXanE
6IjkKsM9IL31IRdn9YbRcjotpJmB20bwxmVxD+nKdfDzt6CPMbXwZuYJJoqctKOa
iE+q7oRYy2IHZlaS6jFyVgCGM5A0hjq0BgUHrVJbZScE3mBcVH9mBk+vV478h+9R
gNi5HCC5ff9Lv59E10Sl2gsy/f9Y9z0UPBDvncN2S1xQuv23i7UKnS7JuLI0XVuM
tzCb+PH0neqzSLSBqy0YtMk6VJVWG+AaOX/03g3Kck8zemHuPUkelqWrmsOd78xS
IuEPliASfoeeKDFKoZuyidhq3+adk8D+XGrIx6E4i5k0/Ra7EKB5Xk1FesA6r0PT
dahvqRcAyBLEkva605yhqsIMoLuC6zNY8gOclMNc4ahsigX/bPwfYeyLVRCaKNXe
fBfcKPYna46xckFVVBWdiLv7OVh25P7NLG0gnsv96eXJetcOJbrUTQwBDX5O5yqN
H9qZX8W5xRZZbPABzb57/hWmFnyVaQQqia3//TInZ3wlxq9l9tUl/XuEoDJFJCyV
+f8yBz5P3pLUjlay+Sf9UiiENpIw1RbMK/nkq7Aa0RyIi96V8H4qiUoQMA/2G8xp
KociZ8nZTqgp+LrvuccQiowfXfD9HpiBl8zwb83C+oylLrGCVV52Lq0+7zLXgB8S
wxGZwjRibw29EKxWN8A0vT392OSQprS/SdFLsIAfhTjO2DsMSNURdSWjmEuXjDM3
UE1ftkou+abiJ82mVkocudNbfzs++XsuNUpqnjrV8UW1ElmClkWR52c5Kw/HwAC5
syGze+9eD06TjBWVdhLB88CKC8/mQj+JCDRfbApGqQXPkP3lZ9RlFhXi6JACo6t4
o19wzcmjNWVOfkH4p377NO+Djaewsk8+pBrRhqVR7/l08sL8krlbbAZMfq6++Snz
1LF2oHC351GfEHGhVj2IpeuvoeAC5JaupiH+tl1TO/f85UvBFLrrMxpLICbTzUN8
kSCLXxa2gK8yDxCfhfXm7ef+6unpOyI3PkCdybB60ksAFwXSoxE11QZTPpDQ6wGV
7qCALxLowxHAhBviPVYkWRAlOvevdW2uFfVIholob5BISyzCnc8jmw7sO5kVx4Y2
Oc3DHP4cN6/vSiXehV4VMThFTZrun1LmpNrlv4FinKIHQw7TxSfJkviTtFKTT9FT
azG3Yszfs54aT3gL40SvLRQl1tpd+VdA+/J2T4TTlR3+R/T6SklmU422abGKUokh
le6Lp5SVPo39JKeeUEYeTv7ifz81AmuvmdsmszVQ+eykdqMCQNGcTwr7578yUa5n
Bs9VSnQSOX8ydyQzXc5OTj1SSt0oT6WfpBYNoGjZQLd0EEr8tWXTV3c0Xavw3Rfa
ZNNJOR12VjgWZ4ZrRioiT15SpN9QMSVMiiSmax14vONXNuENEHaRJvWIwCglowrt
ZWN98SIiFOHaqPkSs4/7q7Cte4AwaiOl3Ijk95Aa88VWphyhNnW0GDjfGYllLn0+
Qbaq0VCCiUVLcktB3lkq8bEQYmq2Hc9A34/lsx9tcqd50iYr0+eMBuxyuTWlI0ca
RyTp5v4T7Mj0V5Vqu1UW15X6jRQSI5cuGufcBKGHvB06kCCxp1cOuVUssFwNDWpN
EVkZBX2P44IAKDfldLrtRus+MNdeiec3+bxiVWjzfGTpA0ESA97uPhmzSEh8KHPd
Um379Wgcl1LEE6XntfhVASdQK+aTsrtDqLxXCSq+UpoWE9eFz69TyggnBvvKZcyh
g57UfNEzjfww+W2kRuSkoW8U+ZHbLmJQfymezOC7bpqFsN+C6ynnY95xTN+uaCue
J4OO4OacK5vISk8rnkl2wxkNvB5Ei2DntdG4Xu804MCw8izZ9Fzxcv3LvV8ZH5Tn
/4LOJrmPgOTLh243z4aJXqhWqAmo0+zVy4WRvY3QyWGHYWbHuJbkUIowAvi27suk
fyCxjn18MRoFOH3EfdB9+meJiQXi+lyJEHmE75lzP0kWPlP3AUg+TgiZpv7r8ots
dDR8v3mzUrE8vMywPFUcG+M0jG4zkQ7F5LRvCT6yBmTUAcNAOEsg7kvLaZtJDSeV
WCZDTZy3rjrsOYdFRCEqtDYFptC2ITxdBTSCsFhpXnp1Q1/NflpddLqMTxLyYr4f
Zr93p5r3WVedOHLKkCpzer7E07PR4fwsCMKNLzgwaMlI37N4KtV8OU0cZn+u4kob
j31gQcnlpBpTFX5sDebhYJL7AfDT+rzqbL1AbXr5zM0kiFRqLNS4p7YyLpcH30CE
CScuxooviD8gPDbvq84SP/n1FJEutJ905tbphjPvL2555HMjlw5q4Q0aNKvXUMHx
zuqulL1oar9NezjZseseuFMCahhUSTyGyocZCTN0czx338yDxcHERC1IXYl9LcOA
f/5eQau8YNl+L7te1A9mDNqokkmQAtEAGacnn4KsqYgG0kMDJNUok60Qtm6mjMtE
i6dM2DDWpxUlVULqM4KGdeeg3Em6O9ZhCpu4yk9vZ/7LxnJB/TLPuEnK4X0Clcrx
80XYBN1qFCAB2Wh5ZlgJP/XQjwuRhcS57lCwsZUE+ID20pCsDxCjt+J0LtY0vl/F
4haGzAvzwOZ4KA2+vTkwe6vv+FAxIbi7IdcbId7Zdsl+k6glewMbFZyIgBi1ZDsL
GLQVRTePVG4dOShP3udi/MTPXnd89AYDf9H9+8gOzyOqCLal4Eptn15ZsRDRBpmZ
mqPPhdYxPCXuyfKb1RHxIF7UI6m/f+FrS4lJUWcnpe2nEhUoQjqwG5uDrDitnY1I
Qyl5czNmw1gtuBW4VtpCc7EZMbpf5AK9y2EuWjGpWFMfBMuZplFpcDfXk+I8w4BH
dw2KYTYVi3N8Weq7gsJSPS7AepX4sCr1CZgRSsYIDDCPZh871tP7V7DAjO718aia
RCh7TqTM4HvpGQrnlzDRhzN3FA6u3L7wCf6ubvyyWNSBHRQ+eiatRuynjQsMIseD
LCnwZfhQKctZoE9z2AhwzQmdy8g56qR4WBv9TMcZ4AYTeMrT5lqM7m6tsUXWZ7j9
UlSisF1M5XLycwinSArylzLNeumlmLPirGICMi2dP3WnyBaQmd8vqgYQmPKDDLHt
+z420OlIwS0Dn5eIhc2bgNFd7q7iO+mB1+xzE0Bt+s2Go+i161IWg6l6cwNmbOb8
j6iyu1AKLebcbUO8Ahy5AXjtd3o49pU+Y2ieenNTHL2luiilxqDQQP4GUtyXRt5f
uvVz+sWAumc4NhEImjk4Q/Lp/ilHjjXqfHiOIw+BVfWxzCmQaFjiYy4JJI85YzqI
mxVUKe14iz6YxoizoAatIStq9jZ3Mz6dLdv3eeuYbT9vXR8XMmiivB1wBBLY3Adl
J0aX8ykgB5Mnq3iBx779k1Fo41R8v2WJHgfIQ5+n+ArdiEHbCGXp2jO1Pbglu5vp
0mtNIuLzr0Q2ogY2XICKB6jikggPgBH8pEN+eaACU9w=
`pragma protect end_protected
