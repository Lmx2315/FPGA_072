// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:36:49 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
AU79K/6W28EpxABacgLWdVFYz3B+G7rCc/pQ6JgV7hM9Xvbsu4xiF3R9+48S7qNd
CEskRZYk6k7wIn/zzPBPTTL95KwBfJf4mX2RULVvZ8ecTbSHsRTFwQBuyFCHAYil
C2Za8SGUNLqH7pcV0rBFklxH3jWmWcmw3jd8OrDuQNI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6528)
uBTNDm/bdJw2U4prrw/Cg90Z4j64YLKfXCb2jDe1Iks6CuJ04VOW8egIGXIabl+E
a4n75bNpWNPJPKIT94yLLsVgCvQYKJPh4ped/XP7aIncJP1mH11ZSa+0MFt34yDG
2I59EECk+nAgeGoG+JY/qjy17sxKTSF52DCCfoAPvGc6/SZ6DeVCCIo1scbbROL3
4kg0PklK7NIV1OnqAW1B5knHlRzBHvI27zbrGfEQbYqbz1BbAMeVpJvYnqNITqba
OZdoj+qVgED1mzKfkgTkhyCsc1yxrHZbBwNi3BPvieHh0jxxM1kz+uENTDXSl6iB
EtvJ7pNvqia99VGkwQcKJD6N/eQK2rT9lV6jcHBfVw2ByDd5DNAMWapjJSgoOobw
A7QDRgpxB1KOddY1qPEsEDnVgSzA1go3IdfW80U1qbT5ukOM+iFnkbTOQnY1+GnZ
hxdEFv8o0e8a92am7KfiOaYSiVp0+tO5z6kD89KUmmYoK8+0lfBT1EKgiF1h12/a
405zfbr6fZekVFes3iGTH3SCzcPIWU45NnRrhlY6Bsshrl/vJHkcc0eK+XeYN7UL
8aJ1Uk2M6GCNFDmew40VVKKa1CYAWWOJ1UJLQdbDhQfY2xujahI+wFW8WyHQFjcp
hJgumU9ktk0smCnw5eBHlMgnOuD1LcDSS4r/1NVdX7ZC23yRyjEtQFjL9tFDpKSF
fKxPBmTCXJpN5lPS/hVumQ69XTYAmB4W3mg8knVuyIat0kx304VQWayH8UCdkps5
62SMXnHaTzO5SbJ6re498by/mQ1O0qYsPoF5A3NQQELrbiJCBci6jeqXAFk+NcmR
W85jupzvUtqzGBmFP4QoWO1D2ixEOp72SXVCzFUplaTgkiNPpuM+paY0+hhRKMn4
4Uffb1QM2u6Q//Zm26guT/JZcFlfmvWbp/5T9EQXSFIUM4s5XxqQBcQ11z1rTDDI
x33ihkF/8DeArfsiH2apqF1TT9qmP9+97hhbAAKadwH7PIOrDHwqik+qWePWnYyZ
0kOsyHkAgJD5GhEgczlw8nJCYJ1QKXo5B0dWxfLZH6cbqOrOPysanZtljOi4rsMl
v6u7eNzcbEJHEfRMLNfaYp1XUv7uF6b9rPzpG7ObCy/xiROXCScvmNPcjFt0uP2V
SgEC4CApzjx5dSXzPfO1cuEMMrCdU3bVom+OQPgcXxNQ9OHK40Ih1YtL2mMACT6g
U+QDOfom4+s0cY3fUM7y21IYYrwFReqqB0a1sEK5wiBV/TyKJgMLjZRFN6rDTCvI
gzyY0852gENRnXTvNprAxvw5uXN404KfCBZzc7D9ECFr0c99c5hKgnU1xgGO9b/h
MDWPABrpL2KNNU/j5N7AUOIEWvhU9qAJ+A+sxXDd0zNBUzCWqYXg+ZkVQoAey298
ZIwU8aF1bAEpE+U2/LB9jOoqGYP7GJP9raLueQQaQ1JkT+yEBW924OUKpFXV74LS
IA2bR81LVJfuwizBmDhmWLLNaPn+wsjUWTRGr1ypaeR7DSEqouPbhNniYV/1rbVI
nN0eMcbK0qPjJkRhZCf1Yr4dziDVPV9qhOrjLXYyGAwswOpgOYjbgOI7pPDjcuZ6
Ovb+WAL2RIWiG645nEa5dL0qa+0ELy310eqcjpOsV0yVBLSqBqOMd6+X7+/dHkmx
3GD7Q/Y9lbI/qWuWq+TMRnMOwdW12Qo9BTDRyqJxF0dLqTQzYNGWDHUQrBJUESIj
bSGRGSUW47eNbSkiucOxGXafSZqMKv7uE+53SzRuR0v59Cr7A43Top6kXMS47gfE
2dMliI7jQSGGZY5JWzMWeRL78AG+0JikaWWertgQHxJCOJPNWGFhOvYhdTrOZ+LJ
EWgwjL1MxaDpwrHYOxLtkIK1d7PSyjMAQsBdHIQqSf7tqUva0PNv0byO8zaXTHCo
R+hlrZaeLBH/k8L1fvZPVGIFJf4i6kIp5kbXSUZxF7m/R33yBx8iiMeBpyGwhumQ
+LLiKwZw58zcuEp9EgbqDhH2UttS76LAwp+xi8kILQgBE25JnMEi3H4JtlkSIAXf
72nBkTcqipJE1Rm1My0yxdAEqBsZnoliDn69YKh9x8WIp/9Yxk2LLI1Yb4Uesbc7
GkQcuIFRpMwL3dYUdJih30P2SSYxE6pr98ku6MEqR8URPXOmkKYDiA1zXqshY2DY
1bRpQciR4ec6c+qnXX7N0GF/C+2fkEj+amXm0AsQu4WnBawXHT8nUD7GD+wqNHY5
uKAJy7YGZdjsOqUw/vUV5Wd0YJrYYjNdjAIplai4CvX1cy2itIF28cTFPAgaNCtU
AAzBt9KckwkyK3Z6bbnh4QY1MJg7LYR4anekn9sLdVxiZVHzr4EH1Ale4+BpQS25
F+pqZ481jeAd2batuxMTlNXkmNG5T9uK95nFulvU8RTA34mxPmsZDr5OS672D+V7
d7ioDKZ2AaYuCtHQSdzOoW/Qw23uKNrwRl8cC5bvOH3SlprqfczHhdZ81A43RExC
L9839UivJcCQ/5Mgk7R+ZpzQ6CfCVcs5P3lEGXJu7N2gC4v4loZLOK5JH1K2qVbx
3lyW4qgjuK6CLprpeH+BjXpsw/+7taHkYq8DzkDzOTcxj2K+Swnd9K9i2a1YbiYi
giiL+pxx66zpIVYWD0kQqHGvqLO3TJqBdWTmux2gXB23qKOLSfc1V9U5bIpsSmUf
yqnhfHx15v1Issrbx6+JUms8+ABrU5zHtmhPf5b0tFiPzdG7PnjY3rI+t2r7HWP1
0OIfbJeel4fLkuU6nW2wYoKxdHdqC4px2Qnz5Fv1TnnrRdWom9g2mVaos8iTZEKK
3eIIMw9wgkEQrWNg5xp0WZnM7rqjh2hSdYoU6tSZMhqr0M9ub1qXKdkKwNygLA4X
kBpgab2qv4sHGPvYoXW4xj6FVZTqSKb2qVlkeuvbp+x+jNVNStRJGIbQrMrZLk5n
CVeE8kwPp8j1am/Fqucl6iRaJXoqG1clCLMCuc4AGMqiWyiKCxvS7ysAni8y9RDf
mFB6w1OZzTj15n2rvUC34nCopMGttBetgYa9HVEM5ZUrfpCUmaVQWSVsKHFXbHP/
Oj5Dg2OeIXuLrH1VK0E0J4HdY2ptgRIacfE8hf1Gq0nK+EEUQIXY1QNyvXNS3YLT
AfjSxyVQ8zqq0LfMho7pHXJj3RjiwSdT7ixqAXARTG7E+icNeS5S7Z464QR9dB1l
a8O3vhipq8aznKnMSBmwbmaIEagpzPVPoKOTdGI/onke+PqCZOnD+umOkX8YwUE9
BNEcPx9U1Jt4nyrtFNXa1kvXfHTJj8r8CpptHeq/YwP0xcHLibb9V6WEvYkqu4mB
7DlGSxELkbhKnEbJLVDWLwCFZPVhTp9KbTH6ZFTNq19vqNa+S95/csH3VCbdGHV6
WZ4OkORIkQUArEYIJw57kh8pKqeCXeigWFxEmIBel6+jhS6E9xAQygJXf0q//+wd
1u0vT+cj+2ky+UyqAwwM4oLe/SM9F5zhEA4IzbmhLrbn0UGmARvLcuFGZFrQXru4
HrEkUYsKFjHWFtAfQfv8ixZBFvvwrkPcHRWeopIf/BR5JoSTKz5gKGWjujnfE2tB
qLsee1fNm5hfYtSBRXr29Ke9CQhJJ1HFSWFEkjBZ24WaahiAazptWzPSsLf/ez11
a4SxewGrv33B6i7YTUq6gG+PGhGcG/eXFHF7HO/PD0cmgWy+kH8XtObep0VSALv8
pFowzkv3ayRmzEIDzoxzZBw/aJBDXtQ9P0Fc/bZU6Z6Ex06tViz5fgemgvFBWjGC
A8enFxxyyOxH4qU9Dha5QcUYb3d7Fltp4Wl1B7671shnPjQvWH8kDqmDhb5e4YcK
HTDqYhNjDSq7wHPzd1VskzOV0LxE2gMTG2pNu8NwAT8X9Q3c3F8yFTj3t7FcuyvH
wJxleI3XwGs+sGJ1Xa0k6OnDPh4/Y8TiTwiWdfNJVL9c3beRX179BgGZ/tabncw1
UwP4gjHnEgWCntkga0kULAxjbkfV2T3FOsmIJ8crXDl3eX2W06o7PpOjR9xMggpf
6+LgNVq9/QTVR7jmUOB/r7iI1mwd5XE5FdEWOPn9hDADP4pbEJOMM4jbF95Zemug
WgyZfzOe+VPQ6eiN3c00Uewm34hCxN7EJcwBzERFAH4jZWmL9ewDeVlRdwoAzAig
p8HHvusjCHr/sN7xLx4i+7ZWSwNTFLRs5BERyj19C/tKgeVpBOx0hROR0IULXQPk
wgfAHap8jl7wT6Jc1V5THC9d8VJ16scvGdrDEW6elW/3pom2ueH8Htwfva2iQuJ0
LQroYGYqrXKDhawSTbuWGEKGdlmg3R1Bx3vxPMpWB5bfpOI7mClNKAqYe7Yv5mA8
0TWtrxhOB2rAElggF+TJaJU7Qc4tbPgM2M4aiNZSAvy/qLSQbMcQHLaJXDJJmItR
QD3dbgvTN7mXsF+Lk0Nf0M9lDaWsS4Ma85yo05PsgkrJLUSIJsIkTz+zzSZOGybN
isj4Z7N37ZzZssbrwmkOw7u/aWqXi5hmLOuhEjqTXn0n23OqFbHjO03DJ+yMNQFN
o6xF0tCGRWRySQHiyjApuGyKYFY1Z2uI0hP4IFKJHZ4pa/NOujaMNlG6m9tCOy0W
g3webgGMfAiENrTGCMTys4keKtNeGO0u7u85kayegw09mdzdHEawtqa7onDR9VzL
Csksq+g5KfB11kC7jPoCqW40gIHrFhwG/Jgl1gWigH1rFXeHBkLk7gsr2fPYRklL
CTM+304ie2idbPWYjdQcGDVvVkEZX4mBVlggxCBW60tcjzLWE/w78rVGWbs2DDVh
/bcswNTVy90Hyi8dEQq5nu9hQpXOVI3DDjPmHYQdrQWgYqO3khugV0sYrTbqz8Bq
RfjeDXApWYTbuz3LjzXbDLXJ1E4GnaP2pkBcEkI13Z5Oj2qhOvo/SrMdw9UbycYc
pOHy6h2II5XYORqt1TtuJjoKQKsE5t8s2OcaNAQ46cRpkm2NuQ7p9AWNsIC4z3M5
pUOXXPbOcylztkxpfmadHMuiMqAVKEp0s7WmIyDnDZOtrYBFhQZ6SNYXYO34qZJX
sEF++rV0f22+2z+rSa3Gq+7kHyHqfTaSC2aWwS7XhKbXgm5u1hCqyS8TsorHxtiu
AKVDQghTTpklPVX/g3DtNaekYIGR1XYDaBvcGPZaUrZS5meumXLzDCdOYmfJOIN1
+i1zYbWYXt9CgNvjUZo1ghGzZFihYiCJQOLoWM7KOgTPcKdzU8935ELvxVP+iXZ2
W0y1lbUBchkY+z72pmWAL7MDaWFZ8QHLUJ8I1tEF1M6/v21EPcGca8h6yj6OlUig
t6JGQApEJqQmIugwQFBF2cFVYDHdBsBJqwm1yyZpVCsVkB284r8zzlCAIq2yLn3d
kUnFvx3X57U2DTtDGl6sUg0rE8bax63hJMwfeD6CU0JLYI3fPV7FHFQQJcA51kff
pxnKCiSQEW1XRPrp6Ai45xC4TNZWq2sK7q+Kpirsm6f7GvfS2+casCO6H8jJlyG4
UjNE1o8PdDcEMiBoa7oZvtBexMEKWIdIT0CjXfILYSk6J5aYfXzfoHSBdC8b2MBj
cEKvqNbNE6r1pIRbJnknT+LnhN1dyxx0EbRb2bzWu7A6XNTmtK7h4Z4AdtMfGM61
U4pjVYuYq+wc8pp9nIeWvflqJcVT7B4k9Mfg0zGXFSglUoTlwgu6Iu4B+zNuOofr
DuWwjGzd6vvxPuQrkwzBxJQK9gJamWRSJbkyq5ibJhXrDNhT5CNtsw3wvGSuWiIz
qrH0ztvgnjD9QnVxPkOhb3KcOXyEZPpmCwmkhO2+UqvYiUDcaJ6EoDSxAsxouPVk
tQvTUYqQRGk0pkDWuoP8BBBN/mEJkXjUBTWa4EMx+jLTC14rmzV64yz8OJDKQmwi
emPCMlY9SDyydC87I6T7tjqPt+ndA2LRzz1PH4L0aMs/hRyV+pyOaw+WDhBkimdC
UqhvONStvMgZ/2/fztF6lBxfLBRp9D3xyQv+9bZ91vMCX98WJBu2ip7FbRPnILKv
1LGUCI8nQ/5B/udz0+VQpe06Y3n2pBu6/pBasr7OzuOTuZJiVgfeoibw8m/E7ZsM
CHw6tB4OMnFcYZQbdGyauw3bya3Z1xCXfLDKbpQiVmA9xQeGDAYwGnhAyP3L+9cC
Q3hOUxjzZh4bTIADILjZonVq1zyCFXXzt9OJdYjAOpCmhTq1MpbtpxprlETOvaHK
8nZrXqzeEsUunnm1sm09xkvYII8UYbi3WPSrR+gXJhv4pPYQpSLUPl0Yi+XvLCV6
npXJxh3v4M9Mj1PHjB9Dcx02pXE//85aiwrVfRA0rn5RQ4ITNRS9JVzwFMCdcweC
HsgP2u/OT0iIsyFiGyrUep/YnjDDyONWbDCOBWQyvgL1kgK2sTvC1ZunL7PwkJWN
95akRERxgka9cw+WYUXmkUEioVzwY0y6u9iVVop10Lx7OoMOveL0OHpH3TWQpys6
y6vyOs+S5fsI4wbPwP2lig8+nngyRWCFTHrRwx027OjjRn3aMoGinmrcUTMg8U1f
a2kcc5wjA4xn4xpeAwrL/7gQxeReTFIYJRS/e7llF+8vwN4zz3NI18q8pVTkByjS
zc/DiymYTIyDZGcsiRQQT8vyUDPBrvkViox8HNvjXiPZzuDhjvc47ghonasy4CJ3
aTm9FWBY3YI1QpBykTE/TLBLD1+bVsVdfF76absHNBf2nX5HDmSS4Cd/7Jv28xQ5
Jvmp8VuFGvsQcQW6kY7iVT77MpGztakYH7Q6zu6UrqD7zXVj/DcC4sSoouXsr2wa
t9eeGj9VUSXimEfDLVPuzrDe64s9pcUb45KjtAhxAvyh0Ip5K6ab8+jZW8lu7L9J
wEBmmAc/ytf1hlUk8R/0IivXryZVM8k32hdWGOsBd/10Uwv0Fiw0QW8/rFMnY1S9
YkyADXcnF2i5a9J/T0uC34uyhOnW/5osEmNUI3KrXF62bgc9NqzaZKegRyTKLPzd
RGAOQINpQ6FskVjjA9N0i4F9nbXr+bYgw9qmup9SYTQ8SW/a0+OVt3TKBlHXzacP
3iv1ZAMMuYmbhTRiV4Eu727tHKoKK6eWJos10lTf2PJQWgGW3HoZXTjuEaPKVyfH
cV1/EXX0Ti48xY5j2YJCd2eFrSQtR5aX/ZhHjg4FlcFg/epITFbAvgqpl8A/1sBZ
RJO9RwCpl9I+5OrIfix92M94v9cC2q3cW+MhK41UZtw/FFmKQ6FY/ybPFpicVsrP
njbbIvs8TlFEt2udeIqjhn8Y1TrorqBtIdY7rX5gTP7RJqxathU/wOCs3rmyzTj4
TEEchyGx5XiJ5Nu6tJ+H0m6iwbtjkQYL0wFxzumtzxddwxzzLAXtJbngVWkzLU+m
A3Eo5gfFcJvW/bvUQG1xp2xE9WyyQ9cIrouuzTNzB6z7J49BLUE4LIFZ+Md4Z4CJ
k2BRC5M426ehPgC/8JPxXxHlmWwJ8xvYCjnJ5NvZ/exgMVlyhBa0hnWceEyaUlNg
5GXQWrsti1HwfkzgoDqjYUVVctomLG+Vi/emTMpyxGFpn72zwHCsjhZvNdpAVOYw
423TY7hFMZiTvdST0o764x4ZA1VS59O4uym1xENChaP4t1Sd2IeJkM4pYWZMjM7R
u2NXjpE1oqi61NtrO2YQSylWJew2TxSHei5XNIl545CXqKOkobEMd6PVtH/an5T+
qVYLL734K5Kw0Is0CktuDI/pgvnOVDjonC6dAYcz3hjs8c0fc08/4jbPJrljw660
dPmcLuD68kTmxdIhdgUDrBMg08J/b/58KCscL0pQemPdTIqL379/P+4K0NNf71Jd
B+SqjbCaCOiuu6AVwSkBuMM9NLEUwPIaDyyBgJ0HY2OCu7FaPjjTX5JmYoGLJwgw
auy2SXT+IRlqntiTPv2yCrKLdZl64BmxJT68Ti1Jzb2FYUAk91+F4kF02NXznusS
rGu0VVA0eGFh3JNPW+7+lVHTD2BYaAyrYAH9v1B+N7bJd5Nuex9InWk8jCWbP+dr
taaWiShG4rDukpLrCEm6JUpAy+ZEWrzj69n5oK9xyNpq9sCzlM/GkCnDxlzY1B87
7fabwLWMhi/K8cruvg4G+eUslu0RxE0zxcpGid/BauUub8IAqzC8m5xpHCg7JVwy
LOhJSUu1UNmgotgP/3d/+MD0TjxuWvc+y85pjOnKqvN2p0CdYhP53fu93oOJ+x7L
/oZBSGrmJmhHuqJiA2EKcyWgAk4oOcUyEQOotaDrcjORJYrE1j8pCkW4DflGqsIF
+FTJNqHSX2YNE1QRSuAS1lFFu3rfr2Ufqxy1MiMQukhiwk6LxedkJ/lEPDAclcW2
zkggTQ65iR+70fPa4CHN5vdh4pOvUQ5csBJ0Jh5XYaXm2vBv4CpvKDdpduktN74o
9halbeYgADN4/4cweXIfmujHGw0kcisTCH8laKX4pYquGOar1zggXrdX2zciNZV6
Dw0qImp6IO7s75dY0ZDqfS4+2uoIHoirF9AxbQfZwDLEeIWM5y6kMaL4+9GtIHEu
469+QrDo8V4mDOPhK0HFVFOIfN7rHJ40iPxwBwmBNiVwOEPfKykyQZYDzQT7Vrh9
0JzpLYrYz0p4Ns0SzEJKqxldXZu5r2npVNzp2KZpQcVtnwI3xvEdZl88IocwP5PK
+5mu1eBrHe9EEe8yz2CDo4J77wfUy6eOEyDppRHq2NsBy5gYecFMxsAkk8jKaGaE
`pragma protect end_protected
