// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.0std
// ALTERA_TIMESTAMP:Wed Apr 26 13:33:39 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
bXXyo/O/SP+L6SAPK62xJg0ojXNfw4wVJkfBd/gAeeUFopTXGhneccXZcnjEySlE
e2oztOPPAletT6wYYP/5qVqaLDlvmwnUjuwzsATRDazC4PaEvmbd40f+5IB9tqwX
pgNYfXSBEUps0c8Ajv3J5ia4TBNSdafcfatjKZsKSas=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 19936)
U0wAyiWSoBxFznjYoUjElgu+if+qiG7wNn3DAcXkfTrOBZnNyqPdBGvDmmxqAX1C
3/bS/IblwpcZ6iqAnoDsJRj8mhA3kSzxF9oHbsptvxag9VnqgndNBw+3m4UWYQc+
yNVqMd3+GVf43bIrhjtS919FVkiLwsLjTsBtf2WqB5a88q9TpHgX+urEg7ubMFXe
agPRnln3nDaHs/6UpkgKZMDWSZpgyNOs1c48jGhxyVryUNUS6dogDiK0nfu5c1uc
a7diuMtpE1Ecqoy2o7K7UZI/2ttY4zs2rF5qwtrKXrKJC2i9/tCplLGpiuPip5BK
q9nx8oAXZEI8xd5n2SbjbN3dwGATxlSeIPUKzqWPVoZMUGqoGUJRPSjU6msthYy2
v67XezE/JM5YK/O5fFOSScUQdhCNiZnncUriioJWYlwaX8tyQcJlYX7giUR8Cxh+
ZYJmc3ZqrDaoDppdBCX3oVN0XM7oKFruNnqI00xqAB+niK7EEopbsYgyneM1S7Xl
dh5JgYLU0KPjFUoKa5pzIHiYmWEhs1S9og5K5+Rn5hA44pm6/hv4AhKnjn1yNieV
rPWHhUpmLqjte1KKEVwT5pOksUOo5DeQBBjm0jnL4E6lCQkhkJ7E9nlOHLENG0Uu
UdDd+OX6bxEbiowj5p2cMD8GNnttwXCasiAEumZWJRW5rA+1a1mjzukr7j/mrj5U
K4j5oKHxR9i+xdqlicsvcA6fbxresNxBi9ZNbqN1IDMT7N/qkE234p5onmJrookB
GJpfBYc6Vy0giJlLxjUdqsFbXU65OQ0PMlV4NKPe/KnztOOjjKeA2eBSCllResTT
XEoxgnk/IXdAtrLvDllmPW8LiNvYG05oVgT45MxTsSmdh3cY6ql5GbjoT+4sgKc8
8cG2ZnF+xCwvdFyehd8RxRu7KHLmq/nsW90mX9MLr4SWYgLKOmc01lRyMefr2aHj
kYBxstQITu0VEZvrosezK3xaguc0LZucLhwhoBxdHUFDF1pIX48IoAlHSbTSRGzw
OGK1P8pSN04FtYQpz/Y4dTwuws4TKtTNZbQN9VIX/1pTgQba2eqE9MNlFHg8h7LH
hwB/mRjPJajpn8TwPdlie7fFj//hplhAb7LLJb8Boh0IbYTye/rbGwqdoVJPVe/c
Tt4QyhGoWsA+CWLnSQhrnt/74uTEWdhYqlEsOpy4nAPROgc5btfLBWkCz1gn/o52
4b4NuHH3SkPmkhB4462HRDRFYAt6rx5hUXnpxXXeaOXvIC4/JQn7GbQrjzqPc24v
1/0jH3vsGeMY4xrh8ea/uDKxC+Y8nC/dfhdQGJsp3WyC3CCkfoO69G7Mv5r2vuy3
otPAHfIug3cyBA4LHG6/XiUCSQh+hNxKu2BgVFySuwSVwXXTLsgVXcADrc4I+3OS
RHZCf3UG60863k/ojyjdx5N8NYCrIxZ6zWoSUi6cWmiIP2hQjImsmxlgJvEMdGWp
O2B80zbwYEoxec+O4k1v2d9ALYNMZHcA8rMC+AXHdM6Hrb7YC92lMzQEjD1pz5z3
FAaxf85/fSi7o5kwsEUA0uv690N9YUsYFVcbFTqrhW2tITnOfMjbJkbFBc2TXUkk
cVBOSMCiW3PwhGaNH3Yc2u/FuCwir3P0Prfxsraq0UqdVk5gpbIIiAw6ppTk/uO4
A4R0lEopqocWy9O30esDsARiveJ69vPlHlGYf5+wuXlZjf2VuiNObpjm8XG17XJF
Dt70N3L2qI7Hig59fdFjl0gOc6cbdnap8VaUNE4H+QfxTgGHV7eUqBG2qeEDjta6
NKflfvohyuzMiJZ93TTKr846+yqnNb5Hvh/1Lmo4X+YAc3939FWATkYTejTZGKrd
ORwVTj3Kx5Xf/pzmUd2Nk0G2WUMx2fQV+l7Aj011lFUqR6sOak0OU5DDr8M0cVbt
0jBruLNJIlh/P4Tt+jUYRXL4+CLJohZIL0aaxggndug3auLAfT/ZhJjTDyv0EqZA
ZolDcfdzV0RKADIyI7rw4H+JZABPGC98cTNJ60Q1CXVgBpFI0KTwN0Gn2lBjpHv+
xyq6aklQWERAV6IDmiHGsmSql0/+mOkgssVFObCxp2LtzJj10kJgE9Zhb0xGeaJe
pxxVmQVLFw8VjUZShhUusU6s71/hHodF/ewgbtQAR3Q1Aa+LoJmIS5UWimgzNfr+
Ku1Vxq1nYFPB6m6flD3pS5l9UUYMWiQ4bUqr8e3B925cTM9IniRcpX2uVaYh35XH
tEbxFKjOvbKMObBYA13NHJ0XdYMaI7pDls5Ktv/P9HS0ieU+ROthLK+asJTFz6Ej
sJQTopYgS9HEO5LuY23nVdrL3RGTgXohw63bCU6Yg1nRC4vVA/fDqhIM0J0hWtIa
KNiud6W62ola1OFgfBzfmE0LOZOxRwgMKOVwXwVGKPTq3mdkwDAV9gaqRTNt8rXU
LWQXoZAGs7tZd5j2YzGtcvdsGp9Djo357M1Rnps2o3iFUaCZcgy0t1y+yc3hxTrQ
MfClk+/FhAoev1zH/pDMBTmXQSawOX2/VkZIPAytir7YK/X1+JWYyB4pDGxshL9y
4angwvkET6Co/HckcKrN4jaynbNq0ckPNuFjYN+cuNP6U6t3vZ4xjX8sbSLoxGc0
6qaqS+H0NW6RgH7ynT51HePxPaaCMgxWH0aBTL73QGciX0FmhAgGYl8TlMIeNMvC
AWpicnhJ90HgGFDzI8jRNG+C+xo/H1F3nEPH+Zum2ugVYkCNKWgwptT80tI3jqX5
C3ZNegr5JAlC2fWtBECg9sVi1j/YaVS6NabYDqezW5WamPQ3fhykIxSOcFngtpid
HnYovg3wPEGQir52TM3CbOJb/sjYNZYggDr7IpA/5sfDMliIXJK31mCkoVKtOVhX
b7byUCV1jtV/tmFc51N3meZU4Wv/PN73ioMAqi7lnEyi4jfo8/Ifoe6GqzajzuSO
cKO4jkUJJHSYzs0Ud0u7wZbnkG1WrqNozy0ecRvww1G01Lh48RNljONGoe1OF3Xv
MJ/D/L/f8c3dC9mIp4dvADTf+6S4JgaGV75scUIHsqvHzpiNOMZFJLjuZ4z6gc1q
WowkBnugvy8jWRdOMRbgZemNU+P2T+VxLY17tNW9hVGv+MKbBNHQCr/SDnkePwBM
8qjlQAk0Mk148x7ZK5jDMYU3HJFvtG5tvXrbei5623WtSVsqrokz8BYwhs8y1jfv
5YIq7WSj+Z+MlNrN8k8+XQaY6qVyJI+vMUxzIyliZdsbiC1CH/XMT7mWqYRd7OzS
ywTOP3Ma6UqeYarAF4e33P5AgHXSjEq3I8YrK4sm9PdjiIjd61rLFVH9s5FceRix
bJhNuzSu/BjPXdQMDxy6j+CNG3fZSnRsX8J1PztydP82F1vfyZE3wfMp9L8e8Fhx
brqTCdfKRt0wHeHYfIu9Aa9ZOFj2yCRwR5OrAoWhTYVvTL/VZtWtzYBf0cEEZ0Jd
BJqz0tJpsaIAI7JUcF+LbORbP2apSduXsl8B7+B/Z72Wr2MmqCBIeT+r/ZOs9j2K
UFGX6nJqPXmBKRPdfxC08IA3P/FUMPKGQ1NgbJ0c0KgvyOMTAKmHcl8kudZVA2JC
qmKyeXqKEOhgHvhQ8uY4VEjM6+AwlHD8FMdkAY65R8QAvvD4v0X8aMp5dt9rqlvm
j30L/U1ZGK7VsXzhJcjDwO/cRA8tBC8Lsq4mnQ0WxpvfZH43c3JOW60VNsAU0Ga6
FMy3Un9bOhH3Hc6M9AeiUXg5zJOUv71e16ERA3ObzXDvCpbRXENsWVdsQKIdswUo
03MBS45ViI1TQhh8NOqXd1Qe0X9bAeMbgA+iEzRKh+uL63Ej6EyTP8RD0tmnR7ea
6KN4Lji1Zf40l6eHGKAwXP0cRvXbs1cVsdug+ux+UDlThJC8YgGJHhESkAvJmuyu
8H+08C+Zy3ZToUhftc6exGCgr9KFdSDIMwHI/a6Rjbw0a7AIbR/F/M7DHX5o3fJv
kIeByFnY8BN3s0C2F790YePezotEYR525fsVJJtd+OBFpsXO3Y9hiS/ntGYx77dJ
PrQB6ez4LeiyY4S9iI8jAAhYKk900My37CkgVkXjtbtnNetCQCCAsCN4f8j1X2Dn
deQ+KI+1ypFbqPiEBuzs/mi4i5GezmkJnqYzBGp+oj3OFh7AIOBhbb6/ILZTmj8V
qZkFbguDRNEL705f8OxscaConmOTSdHMR7QdwlxAw8dkeDmAq2d5ThE/G8pjlmrH
nbcnoeISfZ2v9QWFm3i3RJZm++983D+a84W/XqY2Z4PQ424x0QRCK1ZwOE7hvHCD
P4dVJXLU43hgk9NOdfftYnqqlCwQUpgUI1zmSzM/RxDTqJbTfB+lNVIWilO3P2/k
7qUJzocO9OkVxuVq3MC89gum67oM1p+6nkEnN7uGK42Licm/mizI9VInJT7JwTug
kaPfPsBO6Od3x80fXmi28+eKBNyQjbO5OZigvElM9Yyn8FVLJykOCF8pEOb5Nqt4
jh5D6c421MXNwvvJlrdt8XJmZJ3viLieqEL5KP9MZkZsrBboSEXUQNwOJHebDPV8
7lhOR0uh5CmQq1lmyRyZlwzOGEpTqEQytGnFAWU3ycMAWXvJlMIJJPKT1fJGno/p
BIZpWr/KoBISIZCeH3Et4ptc+egaxyMTqw6vO1UxfkW0bydcH/ezKN12ND/7huw4
qk3BtYWnsZ1Pqie6BjsAdYgB8Soj5uHOZrhi83jQ+rrup4atln+vFZGBBxUQD/tk
ZrYcCXoldT3QIWne8D88YxfArPoPhjA+jMi8QmYRQoHa8MMIvOnYk+jTKe/DDkIh
/xHxyymesswxCkywIlWGaVAkUNJDaCxgJwBGk+ZW35HfJUrPCo4Mg6J7tc1oOdD4
njJ8JEnSAvbGRR7vSjted2QS9qp3V3KZAFwUHkboGXwZoPrgSR2YxL+BDxicqCWe
CTGn6CmRrRE7libUn+mqRXbi99LI6Voq608/J6qS2rduHnpJjM3cEupw6D7X6+Xb
PkNGPBrQbpuQCf6LiWFi0Y2q/qS4yFt/Ov8ugMPYl30YiN6mcRMTEGG8jzdUoeei
Xiew10egUwYLefDHxPlRW1tXgKAwwBwgVsts4YpE7YdLZN0ZwN9nUSggkTR2CB2V
yVgRB5Gjv6CPrNgFdvpE2d+YudNoNjZCwQNjLG4yuG0L0xrUA7HYd0RaKb2Zy8mS
VWzI/YrXN+/4udoR9/6fNw8242NDbMvUpDYfQrli/RwVWrDA0tIg9GTZKvNLPCDT
TsvFPizu/fWWbVBavINnmtF6Io8B9GCalmJbKpp83woCNKGj+tkCxq5cqzC/h+i4
j0mkgEKoPBtl9pl0XRwRBFDVoiKKKrF6R4UHfle38Se8KGUK6Vma2UAF7LoR2yvj
FK4KoOyjP0S9kkA3Fxqg+eUdS4w8RplVNPWW77ug9P3e+YKpp75IMZR/j62+VACP
KkhqlbcxVS0AFzHkkURQ0Sov7dy31f+8pM/NoR8OaWkN6gDEfTjW12yDnQlPz12Y
QB7Rcz56T6VGe6jeJRSGCaN657iUsnSOQQm6a6E3LK6YpC243OnYLUdqwTOxhC0s
IFOHR5QjQM526ZQoWrBubpF++Y1UDYYa3A+2waOqeW0Ivi1B6v4DxI10w87iFMl3
G5zQflts6Vv4LJbsxoq9fC8RROuUdiQz+YcYA7Fu+G4hlLZWEZ0K4zthHRNKJr7R
kR5op0IZN6E/i8Odw+guY1thnJRpLuKp91BPph6KESxIWW2mS8BYxMLplWg5Dksl
kt6TUl/OyA5OVu3jRP0XSxDt4FrnwRohNyoeeLze1EOpsGJI9ElTvdcxn+Qq8LxF
P04psrUD1GVBW8DYh6U6WA6keV/eWF9ejkae9lDROFt4M1mypwgxgGkvR0euh1ZJ
EPwPKN0GjyBVx8EdxrxxU08Mf0eFVUQ7nbgJMC4sQ9CrR6ze5sNWoQfpiR7KMEAS
xn/Br2DpQSDZri/GYJ9XMF2JSWn/ewsr90qP9fjeR/kXE9DWlemtjETDM/FVTZSu
4BSS8tMAyfy4Ur33GD9PgrH3sj8r8gyL9SbkEPawpplCGXEBQsHNatXH134CbykV
lbESdm/REo58iGPPsCU5SIp+xW5U/Y/Kd48m6U9W+0FxYMbe5OQFxhPReTLJDc8p
CicysVFR4gmYNAcs9paPHFwglON6eRVXfOohs/KfWiWk4v7CegfcxxN5vh//t3l5
7GtJTkpEM2TfZg2NxTi/rNyvIZTSsAhX4r9ZQoQfivBShJ5jc0CRtpNdA+Mqxj4a
FMRTFPe7uUk4o9i8JWi5DNpgZJKU+AmrEe4O5ejOH6VM4c+u83owUjiFbOGEJRwz
rUQe2bKU8ujk8sEh+wwuCCCX2qZnzro2t5ZjWW82BmyAmAtwpzHt9b9NE6GmF+7Z
FIZ08hwYdsYxSSRcto7SKVcdgunPIXqtMa+oFQG+NZ7nv6j6WtSrOg8bEbNMckbX
gWGIRLc+KvbxgCmi08Z4n9g+1T9sP7xSM9AXVr7hUs7hDPHFM9xF78toAr8UnPVx
4HeN8WbGKDmBKMEiXOMMeljP0gOMDa9H8eld2SAkQlXu9HXCS7Y+K+ATr2SFEU08
TJ4M4bZ72IrmXU6XTPdgJ08pKfxBeGNNA6ngS+JhfR/X3cOVGZ6W56eAFM9ll0uD
zIcn7o76pyBT7lle54kGFxpX8reet4ykw7lhhl7knE+SVZUyJ8q1JtGH5tDyZBXk
yNVFGkh73ft+zoPbyYmsHSQ18Zl6SX0B7UsWNgQtZjtJ2hXwNjzttRaYla1VyigK
ftZ5j8qLnssu7vAG+bkBJ9BHeR06ZvI6oAwM8++ukxcY1hXi0CmO8yMVidunT2UQ
TcfDDvjzABJZPxSSGkoagz2YS89uJJp2b9H0l3MaItprZKPqvVqoyN3kBdSH3Vms
K6fTLwGBOpkGFSIHkTD7BAbtuUQEBGoTDDqT58YJoPGwK5I8hW6tzZosxv7I15rR
8pnaHKAvZgdsNcZVi95kX3CHcFA+xJ3kKFk0hlV2TGgARA9xrPrejqTrdIDADrIj
VXQCM1aM0UiEdxW0jNTFEu8cMZxwTuvco5/X4pGAaGzQsJgJGfYO/YMvmdE3qiYS
SLYExwSdUHRXvNXIA53Tdcvshs+rTfPcBoE45CPvvas2IUDvmJcI8nowYl35uFP0
2yBYUfm/ZGsoMDQ+yp8qzSSOE7+vRoRIR3cYtioBkeFxcNTHX7RqjajX6GR663BD
S7ArTc0OsraCdDEYVTe2CVjM/46F3Adefmrc7Dh6aGSV83dcV93vCSpyjDsKByDd
faXlxPo5B3xZwlegduq8W+rqPN77/rnxj2iOanUohJgJCKEzwZo1FgF4D720jW/B
fhaVN4BjVkva6bbsX1f7rVXOMuUJbzVxfH85SpRDv1ozoU702hQDEE2IzUevZv56
0j7XHJVt+ZRKYnGlCDD8nhJdzhqUoo7PvFl+0XpKUDwWfBA2YgimACPwrE0HeYVr
WGsoU7A7XRiW8t0G5mTGFEUJptNQaAUmI7d1XX7LdQwt2K3fKzYHdVSt8efU/NfZ
+NE0weCYI74dbs5Bfn4P14LVFFTTbhT5Pxdt2NEH/TBnvYd1LzHJ/1uE3uoLzkjP
t1/WA+pwGmOdgzTMwxQfECMX19N5eflSkga0l9yfj5cbimb9dERiCfJj/Bjsb3f1
fbp3uuXutgjZk8MyMatac5xGP4m3zuSl3p5Hezty/btuYedfFXD5N0TZxlZV8zxf
0QXmt5rTKT78/1DFSIfaNncCX2t7Of2R9PLIvzbYbTICtyF/rDGl2+l/wXOcYgS4
wi0EjD9UOA1ySSPTk1NSHhMAXerB+iYsL+Y+pQduuxEoOPNOlKUiz4z+43HdZiom
l8oCgLh05Fpi+g7bKeYMRSoFIOpEw7G+wTLb6lyQSfhL4yO7F60sXIowMuQ4LfE7
kf2m7rjB6IpK+tjoZGSpnBVRFQbQiy47IWmMA4waX1ca+V0qvsZxg2nYmKl54jJ8
r3bzzgtnPFFB3fcoDbBTK24ewocX+j/TEZZFMiqBaBLaX1H8s4X8X2s/rpFYlu4O
tHSY8oe36ZRzsi8f/STf0IvnvcAJsxONgWXO2CUjMCLxTU58E5aoTPvU1f8rrgBt
KOGojUoXRQvfhMfDenan7dCBhZe0rL2x4LOuAgB2ePuS84t8T//0nPrHRXYmrhA9
YfDYarvdWPPUUCJPbqSEaXFeticvZa+QK8Z/iEDe5hRcDOorlesPBt/ykARNf/e3
2cqtqvFzmjLtKpm1mG1NPUEpNA3rkE78Hg4wnbd4YNTRQZfnX6Wonp2Nbrdji5lQ
oW10knqmEObFvjmkYM0/phlMI8vD3xSGQflZ1YYd1IfEOtRBFLAJru8cWjLPGo+i
+xd1wUhWpOlV4fvAZI7xr/GLmjrD4alRrvtP/F5NpI0PFy0z5QzAahsvo95ZFpVi
dUATobt6/f5WsTqG3Jrq/WH2JjX1QiTDV6S99Fh0iSbW0fxkGGhGKRQCMh/qdrny
ttR87lLSeQlr9qrGjgIUO8sXdCUF+1juhCrSg0dRNp+b3BLp4vn/NzvhpqNF2/H9
5qEdRBt1bYpRIIYut69OM6dp3Gl+/8KWHvOSRsC8dGBPSAj66ZOu6DGXbViV1oOM
8p5gF13bcY5HbN8l7i0YO/11fG/6ivoIWbIXbYFF8gM1dKileUF2nDHQjApSpQLh
a67Dwi0uhJCUgGn1pUay1/xuYowsT1iqzImhoCtHPtMJG+sqCd6Zr3VvbHr6MhX9
igJKxMibItG5mu6qvl9lIf/Zyjj+3hC4YGAqgnaotd7YWAQinz85jaZKK0RqmF/7
eOCGFA092YReSx1QTHYYc2zdgQNNw/kLGrCLk9YfffnU06P6xPOdtDMYoY7MrCS7
itMOcyICJ11VtyxJx0zY94rGy2uy2qC+Im4KYIDzIzCadIrLbCr31Pvx9E9AxjDZ
CQJnnQunBKSNsWL8o7CvIBU0nhb2lc7Mxrv1U4eG4GRSu1vHhgQdcCAjPUOqB0bc
E0jV3Fc+nm4Xe5Mu+jWTZekN+zrrz4bfF1xlFbXt6Iw5I/k1JMO4Aeu8mnhBB1Qi
IPE8PvMRJFqImj2pk5+W+y+7knwyd6n2Jxc6fS9wVrRbNoq2ZomtawFzrIBZM5kT
ymC0j9Z+AsbpjgBxIXjs0JSgyPIka9qjshAlwV3HUzF6V91vAIYQo2/D+Mhneh9Y
WhOO8T9+Z7tw1wgQr9IBWfI6UE04R66TGMgZG5SBaPlYruT3FW5QhEh/002gOnLu
m2jj3ELSGgEwQy6Y8h3bpOjVltPws183LKMS0KZQXA+zcF11DZ9oRktcIlV1Bq0W
sxPMXRvbDlnFfbpkaNnqUkZhNIw69NFIJWzImWe3jIXBc5YM2mtQ3HiWAVbNzzyx
/mZ9I5w0BoznaYXhwuEaWycL6gUhWvCCAqScuG7bMwQvEG9TwFwCSYb0y+ynabB1
Q19BYRN7qda5KEkERxguTk5xVtYLQRRizU1zszHN+RbTsYXmziOhelYhcqurculO
6lDxtaye9TUoouKDRehKmcDSYpDlFFneAHWNxWwmcccyuYFJ3tnA9f/RaN7ldBdi
FFbs/qoW0dcQsx8I04E5EWaaAJZLHukTf1qVX8PdPjF84PJEatdhjxnQpOJbXOcJ
hfOFM1za4v6W2inSQtMsI8G7blPbFetxEaFd6fJTpMwZFC8gEa+DuEbqAGvM6gGE
0b9jYm3vWmgjOwT+EHSc+cRlX31Fvjrb1/SicArPX2G9F9naTBR/T2NnKedzQJDG
YiSeMrwvkIpLnkKHMa1mIyAlCBvWP5FxO2Gam4cYfSNu9u3CxhtCCQp00fbEvhpK
pCWBGHEkNX8PtRWUq2VG3pZRSCne9RbE8RV0gY8ZcIobT2uihbgmFWPEDAXaYOHo
aKObjAoX2BRKrqlcpB1ETdnzEW9SQMd2lKp3gh7JJ7GXnkRHbdFCchxFiaydc4Lb
eDXx2VtLbaKSrte1hx2Ied0wxFHyBm51mhJKYPCBJwFnuZhNIHlXGQnRShBgl8HG
wB/YLhbBxUK/pDK+wiAOGS6fMSaUPf84UYS6nVntTUEirYfkVqkZQ/oLBuvGiNzl
9nzXuYQTLfpuDImfL4fr/8VHI2oUVI7bA0LJNcg7gZXP401EdkbGyzFXvJk0AvAI
XYOd/O2JZGCUJnAnlmgLk++xAgMMaPF+IAQvBjar8br6OX3I3hy035mBnAk9Qqej
xhQbrZ6Y/BSzUH71+9KFB9xq7nPyN/Apc2kGUcsHmNDglSlOKcR70YFUUDyw48AV
Xc1cRI9NnE0uEpSSTZmFo0CNlLtLoBx2Zp1RnRGZYNcNZw21v4CjFkZJNAOKDleL
NPzp3DBvRY1hVVChjPIjlifSdA7w1VnewHvY1jhsQU5As/GrO3GeqggKip1Xlrjl
FISYHRtnbUJ6rrSJ5AkTHO2rf8iG/WWoJ/n9mDp2mZ6kUXAkmm/hkFPbhghB2t39
HiqqrBJDeSOTnIQZM7U6Iv1m/wXkBUfbX+xAFSsqoK5aJEDSwoZXLXky372Hncym
s6WxdLNVCvDFRFoSjKjunir5UsU6eDLoWPhCGcDMNJvZa5amQpDtCP1ZDRwGHqtH
7Mx9JlJicwtU4K8GCAuWHK85P+CQGdI/usjUtudPPMlimZ5I9M09pm+vc47BccMq
54OmFbi01b9p6NtjlMFnuSaxLP3FXnJRD5At8WCrEdW1H72JG0uhQ+t7H+zuO0ac
vdvDc/QLzltTc3qi6eZfXaj9kCby2PmpXCLhHV+exZ+OfkIZVuXW9EPG0119MukB
kWGdkfutFTj/FbctV2QsWK8Nq9MAlpIV7uxUCatML+s0MIsvmIum1F8GEv5xNOIL
Gmt86k+qhzQ8Z6IbaUR6BMh4HDx1iUUdKIDYDQau6Ars8/WfTGf5+YL8goE8rSgY
A5cPUJljrdhk5w6mS/6RGbwH+U+V4EE23ix1pm3NATYy1RcCd6Z+PsbqN18sE/X0
NsgYE4eR1VTh5kq75Rq4xvdI93hhmKXw1HU37ag6ixfjmE805S/X83vyHCFDaQ2V
EsGvHPyrqP87/ruyT9VmbhGoeomFK3WiR1icK08Cy5Zi02XyNS+L+pZ7VLp9mAyh
1TzNILKOIcJ01MumWskIcSl+m1wlpVDF+9paj2Rgdlx9ROALJaoWbez0PkuqBC9I
cf8iI0Nc99anTTeG3i/UjfM7MGil9Zl/xl0iAlT/TaLayj2ibIU5OxVZTl5CKS9O
F4TcUZdKsKYYX/rcr2hlNIAbt4Fbi3JcyETbouzvQ+QnYgwla9l9Q52u32xavyha
085fx5yc26z5hJ0DPb/rBk7fU5coz6E0jCNCRxy80EKdDwmofml0WRF8573qum7l
ngDXmMaRkOsTi18ra6k8tessDGxAinJTf7MDJY1dlzJM7O6pgaiMcpHYH3mN0gTf
OViCGKEcV+/d3q9SSUefVutxcBhhyYBcKwuYtrnzu3XXbNc4Hxykf+2ug3FQFX+M
VVhIPlppwQxUEMONzCClPfVoaK8c2iH4WksKPZikNfKCNWPthGENi+WWgml2XHMP
NlnOvNl4UfRr3dkcJ0Ut4zdBclL3M+Cv2ST9Pg5bNbagdNU408+eYwaMBYCedX21
7zgoQ9IuEZ0njduQD9KrnYLRf7koV34I2LI8WsQp0JS4uX9WWww49g7UtrT4pLPl
a7cO8vnscrqzz9fZ/guc7EFaSI2gW47MrNPMs4jRZu0LmClkRAl1eGa5WWLvRE9N
/nF6MfeDoMDmsZoveryIv0owhQkrKfmAELFIMn0wNLgryRytrHOyGHdTeWbKaTrY
Ip6OnprSJIWBBkbxbGdJcpQbwibCsy+QDw+OXUOdbaOrVtSeD5Nfu6AKw21xfyhI
Fo1yp5EKUGCPFVHyYwkyTpIQ2QbgTtZmpEHBRMMyGDauq0GAjM0y8Dr2obdrim0Z
92tsx3fr0Ol5GbL3b591D0+dKXiZ3fjMpXiXjjVLaqCgh9YyyrS+RnQ+AqVWrxOQ
6C3hoxkiJhBwaDPmZWc4rL+vVEm7zmAAd1d8atNUlZe81FmuSzY99xzFti9RRkwA
4KhN44JaQNNcw11HpHZkAwOiBqHSTgfhm7Da/YK8iLlmK/DlAwWjGjJZRQHc3MmH
7auI0eFOyQnYA6QeQq040Qdk7BwyfxCS9Wc29iPK9kNrU800Ewy8awsrfGWo8c5x
SIy7cbX+t+7hHL84tbzDKffOBhzpI0VA4QLMDk6Oq0TqWVgWAJqxvI/vvxOwFVK1
PgPn7vuVNzBH7xHykYPYVf7N9aMW7K6ty9gzH8/OTgVrx/18Vk+9qz+9/En1Azew
F+HYtS/JnkXBOcNN/JqdOyMscl5z06r2MhlheoYcS4l9Mj9dzXd30303Qf7lrfKV
PNE3u65F4+gIRxzCbjNWcpbUCubZR35A/pSvrDEIAKi/6davEW8PN3yOtIg9bH1N
pqvdbFBr11+Syg94j/tagz+pp5RCtcKS/OxL8ox0YCuKlLwBP/GLopobW3Knzjo8
PXFypYE2p7I4ZpipAn/U2iR4wPoPKbAwd8h5Z7P7Ox0/nZwnN2W0KEVodmXlwk7b
xUiIb2SeIyRHrDoeE0yQrOWl+GYoLPiZoDQCpy83Zqkojuf757yctAm3aObjhBc9
cNy4fx6t0yv8Bt+FY/8QeZAGsKh0JXOXsz2SwCgIzw6WeHWWMixbQHu2vsuSBtRK
dMxOBbRRCPWccPQ0gyYcgk8B/EaMwyuZhIrfIxaDx9A22V+zq//ApAiaomYVatdp
Odbz+NDm48p9pGvQfpekO6LSZEB4BoYhC/QkvknaHo3F4F09zBiO4YzhnQUyYUvh
A93iBy7+2ggCYxwEg2Bcq5bixkKrWEsYYZOPBlzjiDkxhnvkagvI0STsZizYGojv
u/rR3BQDZOOG2NA6cyWYJdEe59E5UycVzIvHIJmqI+VXtQ4CPnViQAhhr68YLzoF
agkvetLO7VQl0XAcpVi5DT+5Qd4A0lHHGfoZPcCc/1NotzJHfLrpBgt0ka7pWkf2
nTt2cVCldJs8S4eF5KmZ/EIBNp0+4NRr4Q0aVHbMUWZuKwTfGuDO+Sr/m7pUFOKP
w+12VpspW28pl8Sp4V8ZOx3ircs5xesSf/hR5QyuriVg/iBa94N+spomKgiUyO4j
2Ez8rPYe1Cpy7+DyacYW6hXwX5V1RSoAmxLsDSKwZ8hFfr61//A64OuwPseWhczV
3TZHwKxRCnks3frD0oU1DkRnXuTbsMY7EM0iWZfyFQFkW8KHijFTK5t/2ESneMVg
jTCdhpWKQK7Z4xSAlTKSw8TlaCrxobNAC3kwWMhup1bhOOFMKPyw5+jPQeTez9aF
85yyTOAmcWe31fYmxX7HOcxk/xU+ShA4P0OL8gqZtjXkEm1ieCk2B0WCyC959qnw
waSjST1/EXCD+gmGzlXZtts400CHnSdEfBrsHxucsfFPjwM/qNWo742ZUIYtehA5
R4QdmWlIGpbAhRzIOZXralmGk4pY5+hXOk6hUnOGnypqI9WS+UZrCAHRNSCXYhL5
J+Rv6ynyqSF18xuDyJ6ty8i07Q+tB9xplAHgfALAw/Vc29xxlQm1EcrjVupQ1ahS
N6iWx+rK15kKLK9VPUz3ygWab5RG3sjUrZOwyU8nFdsMXWR3Re1VoXlvjqJYzEUz
sxtFmawRBH2OS5vsx6vR3OZQT3uXmx9q2ScuVld5VzIwa3GTJopoU/OR8IQWu6jD
LjCYoiykx34uUDC2BBajXQss9ZkMYlQZF6Gmoa1QujRBnLRfk8wD0WCNFevHOlwF
AyDd3DqqF4pxqyJ5kL66g1G+QJFbdTre7d/fNSLrdI/9/Jpt0sCQW/JP2dGOnl6i
KXkPNsGZP3UV780eJ3aVnVe5Ajvu2nzDL3EpIjcw5nFx73XSpweRtsHqkQ3vn4rx
T+6LQ0zQysyWYaeLormxuz5BBjGlb6HFj8Ob5C61lXpg1+zmYnsKBkL2iy0j+iv4
ofcfGkqVai9MupLYb01XGwykuGybEJFHV1xfdxQ9j+3p29RHxsEe9U8ERU38TEYZ
N/iM8ArOkFOxyi9mlvO+Tau963yQQr/yzHfWFEPTu2GslA0H0QwRaChkGafD1zRu
ppICclKfffPnqjEHYDk9YINUATsJ6PtoIPF/efxDh2W4ZRuF3B0pLWZn5U43zNm8
2il4+0zZt03ICXXzvRDmppqLkORhjiKRiHqNH4tyfDrYp7tQei6FcB+/Fr31TQRQ
4v/vJIuoeUTJo42ywGrX2P+uwe99ST4fS7kKNVEa1YP/ROftJ1ursoYmAbQl2KiE
37tioGfgUMjfLRa4crxawvyqrQzxvf3AUhWIpJAukcc68hh/cTHcjWFzUosRPlZw
c+cw4qRKhhLI7qcHP/Dc5JCwXqjyg9T7bUEr8ojqVfp2TRmukSBJDwKGi2GIQCjp
GfqZlcuFMSj2rxejRoJ8hSQilOnClOBTBSZro6D1NtY+E3OdcLbfB1RRYYPpWlyd
z96DUx6QMMwqES/KxGoiIAet3MDiUQcE+d58a+Ja7lGL1+dKDcXFx3SJS6sW+nOC
dYXU7DpWNRHZL7X9rSLD+lzhmW6l8Wrul0zsYbJZj6MWlv2QMVsQ1V7XO2lfxMuh
sabBZpfKyRQgXi3KlID7IzUe9O663Pea16T0OHvEQzFvIVtOyp8Od3NeZL66NCZK
edPyqsJJoua+bBRoBnRwVo5hDnjJkWH0+h7YbfmfUxSO5sZQ9YXlJ5qACDu3VFCU
WZa30eXmbg1RyB/9iM7gLcyObbxPoWlvYcjA4ZHlwQamUlYs26pSAmHXEauyFBmd
4TIKz6dFASGsFyZRTc7k806RGVvNtsCHYAT3dMlu/SUjM8oQaCqjxsos/sTZMZJB
0IH06UdtySynoYzh+LGKwJ79j8HQ/m9PkloueYGKLZEGTinKviXEtT/39JSMYHTt
G5Hkg86erkhKDzw8U8cQ21dpXWLrpJ3JHR47DhY5E7vVME8ov226MnB8rYKgAJFK
FohGVZ0bEdNRWZMyvxF/lKUK0VHIuZZZqevRYa58gNjp0KHLIKLsdqveKlMK09Hw
DUmvRfce6gY6Tz8Knp07TVEcqLi3YP+1J7leYb6WC1mcwTQ+0Xs22KaNP3PiEAUN
aDsZvOValD+fiyyPuWgUauKsU4/uBRpS88f5cc7ezc1RSu9QHRfxhEGROeVi44BC
XGrYrDj9Mmz45wbQVqxZns2wiNCL5izhWgljExg7cggJb6ul9bOOiGCrglfm5EcG
N6j5z92kVWaC27++SQyWSZb6GKvc5H6/3Q+7l4qMOECjpK59bqPgQ6mJ9c+7Luzr
nBwnbJ3m8OL7O+ifkwLIXzPZgbmg5UKT5taL4f6gUAk0jG0wGqZGICWm8XuEjagl
N9aYpFkl3+nQysJN1Stx2Rr8Nd5MIGPMhexrra4Q8cjZcHgO8yXDUCXu7NYvo0lF
TvNYABl8ntHF3KxhE6hrkU9mdyUOP/rtZG+Med/FTsHRYx3ut1APKomI41yze6FT
ea3LtUhpJIc7DslIJSgBP05eRP0rd5HknxS7VJxWr33s6Nvc/wRJHh39uoSZeXVv
G96k6YORiXvgzEfwqTD78sAsYkVNQOkRYhUaf5ivSEQJWMusIcoc4j4VxPoEWn7h
4fuh3H72MwljunoKeIFSa+umoz1VNWU1OEcBZ2kQ8DGYDQFwuZztTr+evydtjZbp
7NyD/h283JDDSQ+y9q4ang/VEAfTZRULWRzNhugXQNIFYc2vvXmQsVmCEQ89aDyd
/NMBQtgib+IJ/CVOCcQIjuAGyg9BTX8fiSGnD7WjhM0dh7PMHwUK7Qs4Qbr3TSBU
ui85LM3eJAlqbPbNUdDNp8yVPPgiEmP7vSCxYo18Xiu/XBN7kDBnHIK5hWqEP7de
Uqy4ZkQokH1s2X6xq4rLJQF+cbsvSF+szxFU+RLMIvuT09kO4n5DNbC8GGFXylA1
2kgC/l269wO5/RJQbvq078qtebGRHLUvg8KvTeDib4gJmlp0h+4gmHBbiQG9EUYj
NDeMjqIFrJDyBUoj7DmyqpI7Qheh+syn+Cpfq3hn8NmZOlAeK9/aocq619M3V1xj
zQLjZVPSWA4zuIi9qWvNIU2wO8m/0jzuzPxdEgQJwZGvr8VjJOdoJ/MjgBOrUNR5
7nmxzFupoI/9BBtk4S7zxTc5EEHjGI9U5xe4j3BhohkGyKHUxPS/dU7pe8lNmbRe
4JTmf4qnm2UTkqGflAMWSHx7jilbjF7YlptycSSTbTGS/vrMlv0VP6ppj69S7t24
7rX+ETTmvKonPSS7KmuIu4P1n11CnMJ+oAlucS6PX9klX7yIAIKChKnIJUSzRMDQ
ViFv7fL6J3BFMF3Pj+m9+KUOGkOIrEgPNnisZtR4zquEtlUtU3S/4ehemoznhKSF
7f8+fdy4DHEzBBYOghUMxolkNCbkBbzNVnzjh8YyN/MUr34m6Px2XPhMgrZQ05Jk
MtDXUg2YX8uikV+LBMonaOdNiV8azotfCmStsTeWscecc1u0f3V3edRPtRHQan2E
OEC+FSsJZd8jQ5QhZ1BxM+xft/kj8k3sZuRENcvYu9idLrhTOICp0ukqq2iDt4CZ
fkuF308ftqyKKxgaunZ9EZmxawpZ9yjPHlAZ9g2TBQn38gqR4wAByg5PJuLaGHCS
62Lw9tNeBALa3Y0KZOr8WunfNBico/ZOWdhqoSSwaymK1tgdf61e/vPMcLazQJ0n
ng9dq8r8fNq15kh/Napd7zLr38EqbCFECeje2RAw68shWXhgBwn/px0G3hLwRmX7
IbACDPr15AH/dmE3Vx1F0TwBwclKbPcMyfMX0bFyuihch0F7+Qs6quNOpHyi/Y3D
jsEJ66dJ+vBetL7S6oEH6pxpWn8rsRvvBggeNjWUFt2M64aSagFgKS5U0X+pHHSY
u0VI6/rpIRQnzHBkJAWipy2RSNHz6A4s4T1d+ElzCk2x8ZzoNv/fEeG6qkhz6slu
0Vnyl+0sdLCXyb9dyAHUa14tlLLcUzbtXwX3jIf3WEb2Iz134GrNwXnPHtfKtNbS
8s28HLe6SP9uKFxvbrWDMrbivae6FyWf0zod2utzmLTctNAjW3Rx2D5ITpMZ26Y1
1okMrHc5IgMVF0FIWDwEpLxFtDXCum3QklIrSGJzGIDCDWaC2w7oSn0DhDqpY90H
J3FErTYArdvXye0PHKRIEBgXNF1uIHjF/5/m+huXcbBafjl6XOBVOhXTQOvb5BPA
7tVZbdAZysSLVOQkG6jzuJ9N/0rYX19DYKfWegazUY54byQPW2I9VGakd9DbdoGk
DfORN6yfygOhicZSEm04Mpkg2cjgorw7DuxRrsV4P7Yd4AreUKy4JAyvz9bDkG3W
7A5qn5W8XjY/0CVGhdmM90brDUiC3Xu/+Luos/ar64TF9NtTRO01ai3c4FkP4FHR
VG0R1QL+yWLOvBepd0R0z2n2tb96TGbCqzEL7HjbAdbsv86sYOHEphrIsnmVWUU+
N5w9ceeerGD9aE95UKSLf/+nAcQv5epC5DsxQcXHoHWBBB6xC5Imo7yCBccszPi6
GRL2YvXZg0tj5/rzwmw3CHz4IVKFCgq1xf1Lwgu3GDW7vQ6dGwyKR+T5ej780Mwj
k21dA+1GNWpWUiMbOeYkuim0ok+w6cpd4czzsYrggpnLMdhvyuUIN+xdje3pxd4I
S0+/LpdxTwV0kDepM360nYjc91LRPShw5LWgya2fFGkgo1pc3JyU39vNa1Hb8lPo
5lIHawLjOPcc36j4INQKu3259yRmLvihskMEpsK96KSvKWgqijCDqLEH5VjDdqNP
vTwwANHiCh6ZAkbAAIAra0S1YQpGgiDRERac0lrLJL9hG7TnDtlXAd1FCox0TMtY
b3tGMdfRpFEBp1Xu2FiPCC6gSsmrYt9Ap6sOUU175C44n6OZFe/EaSxN91m1z+Gk
o10BYy6ShQEEDsXsZq4UekCw+WNo814aCOUPnvIrS3eyZAaCTABdFsGixuXPNrKD
nxrYhFbtLGUPEeSLPcLxyZuh6RIHovlYZ9o0oYnKGxnA3WuA9k6gtaeuKSR6ySRr
uxv9NPWE/hjFUylGTPlCmgLttmAs71Z8R3TL4LhJuEEayjhi3o1lHfVFTr1xBolc
U5RtOYP56OZ/NAU4kmQ/zihlAEYmY/DNB1JpgIrMv1J5AcMCRIKUIYQ7u5w9saFE
4rL61auB+MDAPFDGnoGnKHy2Biq5GT2RGagu9bzb9LjqMEZfuhJokahhU9b9GTe8
25q2ra25NpCGMN+MhCdZ4ytKYUYOfug757dsrKkfTMf9iGYF/gHP5Ig0p9WvQ+9T
8v3kswPydZa1/ISTeuQ0dhQJFeqVXuf3G5v9m8iG9bkYDiwtjZ5m4nWi72WVqkYO
A5EKYLW8uRrBIwHTEHe6ZJVAo+/JMqspf7UB21Odc+WWWWItxeuLPPzZNJYttgxO
6ZmWnKJh6Kwq6ECi022X06BdzVgPW5BAxmVeU9UWxLRNKe5vSxJpzGzYk42TmPGF
B7qicY6yNQWLk7LEBwXMmMGrTPrkjimGZFLK90TKF36u+sDJrIItrvyqew1TpUGx
jHYzEEqBrc2Cb70RO2vZONFone1u87YPInNhAL7ajlVo97zpiCGHfqlNo4XmCK6g
GCVYE1dsCHCoUuV4QnaUJ3HPrssHivf55G6iJpwFOgwD6doQpzpUfZICT9k1r5Il
oXSQCkzIbhtcpDhIECgTXhMABqbpYUh6pSahWDODENKU5Zt0wKGhqH6lPC2YIooo
Y5rEW1i8iyl1gSmUQ8A0STXupTrkfZc10ho8+HKmnTO9kFQI2l/aWz+MtzRZ6B6f
aQ8ecSGDqdZWinDS7Xb5j80N5jI+wGu302HhdiDMJ9SO4f8MWvk5ychc96iXhjeW
M+aSTrkb3BsB04YGd0tn3nGa+4HNllfiSLimjMb4EwkCy3n1/bUe2+Qc45MJCllI
efw/K6dVnZPuhsMSPz06xx2SmHkyFlpPI9EAyXLsJei1nVdBGtT9oaXeKv8Q3TT2
spCarjbkQUzdR2bSfptlC1wWrru4t3qS2A/WdSi4whqQyQTkWpBxGaey4J0EfONI
F3deWgg802YoIWoOJrpZYLr5fm27R0x4ISumzZdfDrU9HekCFN0wIaaT1XPsy1JR
kpsLFwTkTBB1iAmh0cS+kBbmWGXWMA4h21ieahNo9LC9yexUV0YPP5wAaeMWnlZl
SZf/1UnDu3CrXqh4b2lIDheL3lBqFirKx6LlXoPK1XV3dvbDtHsEuqY26OQWDURP
62xRTdP0Ehoe1g9uwCNRvS8YYn6e1oeBsI7CVAGDheiLBUqudobjLlWHp4+HxPAw
eI84XuxcoF/lNAQ3WAL3klu4KxCfAATjP79f6T3drOQodUuxZ0DRxaML1bVqg36t
exiV83HmyAdWy7PoItAXOicgS2eu052eZxVf48bpmyDRWvS+Z0WcEfqfaPf2KxrX
Fecg2Rmqe42xPubBoOMqpqze48ZtEeJwf6WQTFpjb5J1ccW0HoSkredaY4zAy4nX
k/YuR2xzkhrXaFhLRsJIV1HIeopwcheHDzGafAd9rICHDMAGQH5P4FKZXUKkMh+R
33bDtgkbLi3hsLgpPxn+6m2lTxcbD7Wsco2apPnXl0vIr4PwAbY+ffwsydb5D9Cr
tGfO3RK67ueLxPU5B7DuE+C8Hn7klyrz5q4a0K3ptKuPv9fBl8soc34f2JjpXOGP
2/rDYjpTakOqeTTMIu6g6eJPEoBESIQ8GdseT+FADt5hqvuHiwvlodLuzsoQo5sM
RDaF75uVyFo+4/TdthPSFeAgP7m7UFbuz2OAdkvwJArtLGW6MevwwM0Dj0u+meNK
o3XP9ov1k3yJiMd4h7SD40S/oBhViZR16x8fyStmeeR1NXUWJd4mwqD1YoHIxPYq
h86+DaKW9X8QPLkjhx0CSn0rqTfFPjfuROzk2xZS+u8Szs9qp+J1FfiYZMBzXe7U
BhRuVy2bfwWCyoqvnbn9eKVQa2HjkKVM8TQwFhv3WRYZqUcbw/Bs/W3v0nwtxZi4
NDtM1Lk2WJpK8lbdIoj/Tj0LlErMDzRm8qbgKyq2jAV3FtqkoqQGqi1xK356ttX0
+jPUIZyXLHDrcl/1UKZdsOXUgiN/I9cP00B9jKAyvZwMJc0ezS2ksZW/JsWWkOs8
CxFn5zfvPdorBSpT4N6S8My4HicUkh7EUZPGb5X/Qfm5zN8iTWjq/o+KLf/zku2M
uT4nTMGeOAMQXMviz02iY4dhVUhVo7Wd7i6oZSvZPLwFIaUgtuBNuAvItdpCB5mT
UItYV/69Lg40wN719L0aSunCBOBFEOnJsUOYMRlhwZpEvZ9QGIeaRP7J3bNu2cdi
QnEHNI3SArMmuNkIP7ef4DpjDeqepP6FCodmuGVZbu5WRidYLPVMZLF3gMNK6rst
BNX2Q69MP/BVEKpXdlqdVaWF42ZzTw9UmreNI7j5Dz05hKd0Ikmj5xcQ8VqJK7T/
9/JrITIkYVZGzRk7+LcTilgwpqHG7+YyXCG2CD/exSAuvXtsUexlrl/sxnEJ4tPy
e6pIR3RiO8MHi/13QRvfRJO1ewNZ2oI26Ge1ZB6pLX1und+TwAhIQvapPWHFYNPg
A65PbE/G56xYQ9zJTPotkRIq0lKbzrnFN1IG473LhltkTw9xs1z9vMKT4G8Z08v5
7EVl0iIFPNMYYKAoOOdCGMfshrHX+9A7TNIG7C04R3biSKi17LP8N51aAGQTChQE
2cGr2zIT+WqA6hKHtuGGO36kiKH1DvUpZGgJb/30/9r3bhB1NJyYimrJzCX/7N2e
rTXuOUCvsbTtE1iMW7nueYK/Fbskk60MY7WQOto/4Z/O0sWJKsBsKgfKSddu32w5
PpcG0y9kOUShg/Bm4jBRoiNtUuEA3svG9bye+yEhYjfU6LxDCg76/k2J2mpkzdEu
oXBFSTOFtvyqZi0KgUmKUd1/B9M+T9DRE0jdgpxZw+VFPp8vVURVZIk+A/ThxJ6w
ywp9GqzcAqPUQ+b9+oKItmJbnAXKx3N9QZibBOG7aAaHROacMDzhDGHdJYIE50ga
zCnJeoUZ5VFqKBg2WJukhTucteBjli+cHj5z9D2gn9zHA9e7oLL8+LKj2nCThytC
NVNDkB1pGzf1VI6rZGtretBlYv7g3y8Qym9nAMGUpfBCxeIWjhi7yuDnc4LpW/NA
8BfAjgV2QDFdRBRXapFonronUPKYYsRvWouQ7J12e6mIG/I0Cd3BSYDruO2yQNDG
lyMC5h90cajg/w2eJGKgzYmdnlZHJW4p4wZTVNUw91fHagbONaJWsFnafOVYgAB0
meODWdLbg5AkJL8v2bSWUmFcCnJbSQ3Qey0xCg+x58dsQsbp78cs2io65QUA9i6Q
IIpkT2eEw90m+M52q3K6vVnt3Vr5REpL7bLYo+H1iLGGoL7S4ofx92tn2UZpOO/X
yrJnY4q9e8IpgNpIQajJ5Fg0IZ3itMcxz/sJx2PtHGfQmAB215G1e5EwqmESKhFJ
AzIru5qx/Qat28R2l7QwLfHapVr3QKiCimbmGPASxddwsdf6wezRM1/6P/Pzfl+X
Ao0MCeRWXkWOA5RtSPgqEeffg3Z6uYb7ZkQ5ZYy63AmZMkupZMQjZ2Aju+iW6nha
SaTa0NICUFDlwLHdLvPx/8RzJevrBo2MEi+gXFKQCUoqp8CBTJ2V3jqrGuSXusLL
lQsE3HvMSHyi6+rfYK19sELz3WqkWMY7QUetGma1tL4hDxO5jPWJi2CPNpspEVSv
aRauO0njxc/Pui9HkBr15+wfhn9VGyDpb073NIqGsBEqRjSsSfds4jnMpPr1Zvi6
RBg7ZYVPP0RFJF5ixQV4/cQKSQMfmPsD2X4r9uXcr2ZZSqyl/l5wAdG8gp5oVl0f
NTt1griBX0x2KyAHnUOpONu7V/5l2GMfZA1AsGgdl5rlZTH47QlEQeIE0CD7us4H
NFco0ckqRWDfNF2ksxDSFU/8qcG0oNkxsXUu9tyTADfa7pbM57igXTjWAhsc5eKp
i+rWeX3W3RGEhBxq+hAKeH3sSv0XZMmPljzRaaRF8Y7pfAcF9RGEvCcpC/bC/y4P
CQmgkmYdRNFB/9RVZmGRoEPriYsBOleSwY4/F826krjELKflZPjQw0CidHssp8BR
cRXJ2vfh8BZpAIda92z7FIDTY6E2ddIGCJ5Ml8ewBALpfnPAZ+/fcUYmELPVFi/g
/2F5r4XQGmaA+fMnYufudcY1I9tO54ct8K9igvhC6AxrF09oCVCfbcgKeavSqhVM
TUbosXn9W+o82L4mEbMQqKB8VTbZW+KnIAza0NKjQGyMYpfhaXwmcZQ9yhuTb8/C
jbOJxdATgDe0TUwl29GFCvjzv3N8/izkygxJRIi7aQm3+q/DMUnuH36/hZ5M+BGV
F4Pfglzse7HDNd3OneGERYVzd3ima98eX+j0QiL57Vv15n1/N3lY9eVhUR5D2ZWU
W4n8j/C/uFYBjbCYJI332qVoDIiqeTB98qpnWnn1Q8D6LUjVMn8jKRGhpcxraXbY
ge6Z7E2R2GyRP+O7tJbQi9xFMVa859yQExj/o+8XTIeBUNn5L9lF8TiAa6QiTjuF
JaTOKWswcb9vEPeqLfSamZ8ZsS9x54Y1XBm8x6DkOpoOGoDWEMPm4tFNIC38cTTs
Q1sVKBfUOBjgoC35chyLHdwidg1i6vD21fTCenagm2HgdZjIe4T8jxE+ZZYTh/re
KzB2J+2EOqCa5VWPl1R4/Hrqzzw+vcVJdMbfetshqm0560N6wPB+rb7RXvfczGtd
o6Qc7B0JcIvWeEsOmAGn1HW4FKk67xn3reqpV5jVM3rQVJ00vcXPHBIiPKgjp00t
/L1cXqmIKOyeNu9mJo3w0kAGFcEVOZLnsAjZCrCtZ0NjJf3AxjG/IxVRhd63+qE9
J/jyS/NjOK1iSU3n/swMPAYqEVfwBkydpsKKzsCfRPlm2ZoLflcK8lewj7GgM9Fs
Fx7LfIH2Z5wZheoFSfYT+1kdb3eQBNcWVLdQxPIgQgjbHx8wzHkkFUil1BYVKAy+
js6xfTpadAlYugM4qYncpqaYsrzZmLyuQwBp4ULU9m2rkVkqftBTAKw17B+4Tr3r
h/fQYvwfepxeNdeoJrF1lQd4KML4Arg7KvGECALKFiPNTYZ+fwpy/9aZD0HX1wJQ
A5RSuoxm1O1rK/FP6/Ma19EPM7MQzFKkf1mdW/GsFW42AQCWh+3MYyfN283D/vDR
AuCid9CHvFwcc8MOXa7U6Wg6bId3iz7c44ysQsz7TJAKzXSjRHhs66pwLhfAOsQK
fBOScoH3UzvFuQpNnwH/w4dXC52btZM0/y/6E6k8bsQ2+HnEgM2XjgDtV+gLI5vz
Hus1AItMo2/dUVlKK+vuD4L4r01M+SHKBoIKP8Sgam/Hm5xNBDId5gdZ8RbzKLp4
94l+/7p187RrwMRL9RZZNkEG32Zu+F77ZW2VPCaUs4GbPZHYWBWElaA7DbvXT+wZ
29lQUGfu6A3/XE3xhgB3ejBw9/WmVREz5NWu4t/E25QUqYX/MMfy5m2L7em2Wt3m
bPLk0Rc/tRjMaInec8npB1IxQ1ur69Z03hOLeo7i8thEtiWtLluKAlCwoFxYqoOZ
AHJQP3PXEmDSwk7fEGkh++8ZApcnTql9ca7MdJO8YNamZ9VwvCz9c9IwQZo5FIPv
yN6DipVfJ0iyQ9r5ScvFXtsW+Ta+NQn8ZGOEjPbbFHpDe47ymVHY/KKImr2kilIf
cKhQ4MR4uMUG4ItXhMHrJxZzWxX9el7fhVeoiSTn56GDCMMThIEsKK1Rw+2SaMm+
jX7ROdp/NbPeC26CDCzSXMW0rPsUZcFdaLg4vjscuEGZ7mRKv1F1mIHtks/VKhjA
nCGOsNpM3PwpVxIA0dzMsYKSz4Ny4Y1ybdz0OyGySzVgMOwZMxl6HYbMH5pKrYMq
A1bB4+OpyGfqby6MFv7XDM5MiAif6pFj9Z3REnAoOuwoL4iBbz61nJyfKekdP6y8
tdWsxVBKMAZZWNTkmWgkqsE+jMEMPdXxklJzrXfa4pRLfYHfVDBpHIWv8oD0oDY4
PE/e7XdVxYyW7XpeqpSrJHlaQrXyLThu1LnBrvyqvkkI5OzmhWB9jgs8j5DjTqqd
d0VJV/NCfbgk49d8KrnJH3ZzdWuquw1MKAyLQAmc3E68Vtq9YdlQ9V6yHMp79Fd9
znRjLoenvIF3e+D7hCWJ1H8ZUBze4SxyC5gpA9CuufxDM5IBR5P3PvSlLIbQ8POW
tNgA19ep73R4Y2FOEPcdNEgf8XdIEMrrtD4gZxL099E7H7S82ligBgrPzR1/yAUz
Ll8kdtJYz5TyQlPEA8zSft4kyYY630qiXquVkPGUG+AqB9l7MlJx8/r5H5WRW0xL
eXOC1oOD+rOvaHVCe1+5qhUtTQJJS2IMvVbjMgjm8PC9zAxfYPhakJsedE0H2/ZY
cInYOChLpbAyfDxsiMQsUbirUXRyheC9BqtQ7JnzZ/XfJDsn9k1OnZxtTs56zHn2
ZMmBMLXoWGpausT9Pw6m3wiu/F9fjLCOxrnPvc0vAEo5aCUbIIRKJvipCSA0bYJG
v3a+xXRXHNK0Kx208s2jTDZ8jRcHtP+PKSXMhMOaS46zEflZzKneVgOFV+58G09w
RNJ7pfexUCcZLenk0jLItrHVltKarslwRU3eYAktCpoolOC2W7AmoM4Ooxz2QW/M
rmqVh3fK8dYx6i/g2hlgSCfuhiWoCa4cPz6dsUnMKSTp/Kl25JHtxXwxbZVtTiHr
h/5W7enTcTxVLMQlWLnlvIZ3x6dsW5kwjSZiFhGFR6JAhguu3Ki6mi/21FP1s7/+
gNPAE71XVQdgm4kzs9ta/UQdluMyUAExoCaODVxfsNVCXIzrV5vvxMdajG36H0Mx
2ih7EK8pnEjR+VIIGD5GsoJ7YlhElZye4a4yK2CwuSCcr1dctFHpJls2hzW+gw9w
Gm19K1Z2QI0/zMCuO4k2DDvOvEAseDzUGrrnwxvsxAid7VtCnuk5Ws8vP2epFf4c
Hj91dthMC+yjM17FfhUQ1mtdH+OJY3NsJbT4/Vq7KatuT9eA/4G99GYfWsB7D0sT
WNPGb9D61iyryaG1MvPzQ29fcl9iw2H5DIlsJ3f9+l95uRpyn3PEj9yH91t6qKBD
3ge6Xh8Qr3kPm966hfeX/rfL7JAOrls4TBZ0B4g2+HFDufV40Mn23I5Un8eVHDAf
VhDgEwGJlP7qesLRKShjMMKB0I1h6O37hEWb71lie9qWrdAS74f4ptyH51kjKn7K
VWFdFqUQ6Ogwi5/Z0Eze2OA0Ktgg/eQMGqYUS56hvBmliMnngoE2vsRoaa80nh4e
C55RYCb93h/NpsV0hxFpY/9dMWOjnReVbgjSQwYh/J3zUuKEevQ8FwgVmSoljwbk
wOMk70QixN7r/qSR7GOwJ8kM8kWXpGdRGcDpGzM8bYHOY48TruSPq/3kGQ3JZ98q
cxRvMpcbqnmdd3LA2G9afVkPoz3t3M2S7Ngsq48srOk6CHJyv+u/WziL5l3iJZ27
H6XUWckEaaibkrdB4MZzhgKeGuuhVcwptoGNPSBY2hAcV0d9KYIrSpYnUBJv0XvF
F2F6wULlK38vggtDBKJUJZBchlIvs5hd/ZSHDWeEFozdsfQQvOIzzJhhHucTTw5H
+2u+Hg8OIOa33ttN6/isMNGBkdbfz9+aWsieq3pKO8EtDUACTyDoEJaHfIsJbIYZ
PYSMj+loDGVC3tkR7awPdGX3pa6o4BwCqDfxDTKtwpjmVKBnfEbgeCzUC9T7L/Yt
kLGwrYQkt1Lo8DAdB4+ahAdTqJHeCNfIFJBoBLbGlKnhZxiLQsu7Od03YG/fs84z
Kdvdowe92QcTDWEgwz3WgLM73Ui/0ODxxZa4KDNEJjl71mZsdApqyM/6JNEG0PLG
qnZPzpLGjY8DqaAumV5Tlr1kuHD89IOrHfJZIfV+/vQnHOMUGVd9unsdG8fszqjQ
hdoy1LMNuc1/A+3WZth7mRz8/PM6an0PpI0ZaYM4IsOj/8/tir4LXSAi3JxytnHf
Z0eXoTfAxDkgPZI+Rnu+d9SObY4l7O1cKU6CD0qKsaShRiZ2yqz2IrgOicch/yl1
iPWAh4gKjxSPNGW1tQ5RBWRzjZhYsiflRVPgTh49q/QAdq+AlqF4IYc3MRQqkvvY
3Sn1uGit78DvOKu0mlCGEw5XxUxpkn2ziAxzCWHx+wQmJTiPv+rnDfuWsIQTDakP
wMFQ1WFUue2nlMsQddjovUqKASGyG+UBgpLCirOZUjEI5aTXk9RuE+5MCGp38lTB
dQ549PzSoHffObQZtJmcbrtnJz9TJdEgOuX+2WCr+u+XHMK5J+x5BCEsnxQLX4dP
8DEl37xOrk8P1opUuwA/hKxpkAqzO55BxTIhe93MzHQU8h5Zhq86cH+tglCHdUnX
w85cLjdN0crfeViO1voD5tgHfT1uhUVMO2Bs2M/TsHgwojFCrQeO9ceCEovGlKOY
YHxoKf5Ch/Ps/3cLea8PSA==
`pragma protect end_protected
