// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.0std
// ALTERA_TIMESTAMP:Wed Apr 26 13:33:43 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
dTqp/7lYtZisEQqv2KkxXIXx2CoTY3rM4muDS3J+zJL271252HmJkjaU9idxcPY9
Trju2oFu4aUOhNaZDrlbIygD+It32OyQr2MQJPJL8QkVrBtZVsDcyWGpBJYvVa7a
cAKySPjdoO5xJ8znC7SvI1YiSIB+DDHP2c292jjw3sw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2288)
ki8x6jniq8QP9nlbGSFmggh1zo0vInXxsdS5u/sorOZdqE14a9bKbZZA8xk6XbOE
c9C+ifjqa+VLkCnAXGL1XqSN+E2vft7BJ9tB9XFhGsX/HZt6yE66KwKrVWYMdlsB
+ZxDHLn3wDAfdMvs3XmrNRdc6NX6c2pG421m4qBnzZ+YY7kGm6r8hFVul1kA7JUU
LoHxOucs+iftFhD1x0SL8EkChZZIy1OZOIXGSyAQfu+15/p04cJ6k3M7Re2xTLrt
uWk2YYVFa3rYhxVlSBUOCy0qHLXWL7rEW5e6l3gDrYiwJMrI4Yg24QKFJUCySrAC
3cHbDsP/M5ibK2TnVOj6HJg2HyGAT0m3ZibAu6kXb5k6/Zn80Ylue0TQOufoAaCz
Bf/2VGlbn6t3NNOWL52s57jL7LKEoTpSZVwoyNspyJZJh/d9gPKCMA8sb5LASHxn
I9fkzOqo8zm7qDEW6Zn3BHQrs18WzpPM6gwOTZ9G8ybWCxE426ybyI/QvPCZEU9H
Ox9NSvAenWhgbHv7m3hfaiaAW4jbNtVgqkZT22xmQqEJ8pRx/OjaX73CpzHJ95N2
b+Y0w6wcVaJonK/v82JmOyhP/ODbvX7uoECzcRsRK077XziUh+8l9S8sLrafOihS
pkASq+NbQLsFxnYHPyA39Hn7Tc5fycEzr3VSM+jxbOqvYQJYqUuuKdMmqLe+eex+
8Wzvoyn5GmgHlxir8pgFP8zuLelIazZXo3VuUl+EQf+YxAesB02UFwtEepZRmVMe
eObK4ZOypmzIvN38+tt2uypsQGoBZBvk9SHoKJLt92f3DhsnFZ1mAxRRHcWGVyQ2
rgVdbcDUphRfdY8MjsUB4L3GPIizQUxmH6XoZxbk6Km9CaTY01dcj0K8w4AjJ1fV
bfI3w4LKXvukidZ/nEeukAM7zvgOmwO4sBoaTbtX4sctdDdFhMXOvFYqKOYbwJOC
jvJJfO9as1FGBGLcs7DNX0/iLAjEqhaJehQ2w61F/YQoooNmoWQNE9ufVvAa9302
NAPqORfM5wRX8ynshC9AurCfVjuG2/VlSmDBUJkWi+AvIAHd/wllhGIxqb1I6WST
XF5z29qWd/JCkB7AtluKvy66NKMoWnKJFvJHb01bVGJwsOVcLcgvFoOJhdLHQLnr
U7r/n+X86cwPrkwT3wDfkdf/LA7X9v8HDDvUew0m9Mhntc80rzl0wSceb8OUarhz
Ld9DkN71MADrIWeSbn+/vbE9mzbcn2CZZAmDwBpHLx7E39ITBbK9SpVBZ5hYaK1e
t3z4hetK5QPrn4/uL+6XTDMphZdoQtX3Q8uveu7Ko4nIKSgCQ42NSPH1phZHDtEH
6I4bzFR5phNhFhqbwuiSSYpLWMuBT1vSqvAH1CmsiL7RBKs4RFj/kbCYLERo/DeL
uEUosCQH5Xdd+DvTPz1vWxMoaSKjHVxypc31kT0K5gje4rjd3u9kfp2W0l2QW0Cu
30MzpU0ORH1iVqkdfwhrN10tTjji0ToQ3NiR+74EugYT6LaFzGaI7+38KgIfdutA
nY47LKDkTcNHYe/sg5zVYlpeExN3gGmTeN9t7xWFlKW2wCPjsR6lPkWbhaSm7VsG
KV3OkFvicWCr6Cw0d4W5Cqx4aAF9XVpcN5HUF2EdD6m4qeSIESqcv6LDXvmeXXhM
XYffLEfAgsGQZQWJdNzvspHI7YE+ju7vybsgMiduVukS4zaJ/9dbAuLLD8BFi8eO
oqGY1nzOs5FR8e/RFU6k4tpHevnLBvQ0m17iFbPt3uvqFNRGNUfCOagKM6DY2lMs
roOS2GbEDKKQl8/Mv10Yhpv9TCtctm3Gg8npVZTbf4pgjmTSBJ+VcO95nDc+BZhx
Ugn/OWta1i0crF1lro+CQgXT370deZFr/37r63acbXZZreXIeafumNqHZYyawydt
jhsM0Xi/xrNSykVgFl9xUuSrA/DLO+F1xfspKnfCnM4/yV47m4vKb4Taj1hWYLf+
Z2M4Eydz7LpD8YC61AqSpPgX8z6hnoA9tQURj5ZZei7lCBEIuIx07EFanpRBgkMK
acpNsdLL8Caradxyp+dCh5H/cFKu1AKuVZVUd6fg+n0N+etuPfOuLeZtk0r7P8pB
9WjZAZuYCeRKX0doMjSFCuzy9KdVHtb0Ji95q/kGT20zKYztHWSbQbsm6dZUFS0z
M1uJgRDeb82U6jWzhttjN/g6yFjbnyyaKVR/WNYYM0EViDnNSVHsMQll34zUYkCv
09M76ivzKdCRyny5CVadxe7BxfLymkJ11bpadRddCWF4isrj72KsZDDcPOMmJIiL
iC2mmgslDOc5o3/7s5q2+ILP/N+bj/vOpAJ9rKIt3SuY8JwX5CkqKfRUIYdpHBXT
C37z3AfeSda/J2X2NBbB/59RRqXErwIldwI/DwbwdSvGczYjbv2RsyZpUh7lRcOu
/+6bKamtL8JPdbkBytcMoGKvEmsIpkVGhp3GFXLHK2VLOyP6buuvSJmSohgTtFGO
041zNdoR78OppJZVEdyX+2lfOx6m+Qoq9YgccAFBBSPKg/o64wMqozFXOT3Fized
RxBBWW7QaxTfDlEv7IuT7EIwYzYab6ig0wg1D2NuvHvLzKsXbciKiPFTMbKvLrtO
kZ/zphwmlDyoRvQJah/neZ+jEYkxLMcOfxH+v5+cHUDFDcgMYBX/QTcUibtLYqsK
dwZRog6PdS4anGD9mDRtkwNrVgr6s21wtBpXeeN3/EiHIuCiPE1FQHTxBS0kSAaI
joh4DVhdk0QMDTyhfV0Qj4wCASNc/IuEiwiF27PBmxbeoEqc+A3StNG85A1IelKH
eOcH0cUbSRLcDx3oKmujUzWtNWJ7jsZNxeBqYRBuD0EF7pihBNkIrPQ03tMbh/AJ
CZ1rWuuIgmF28xKfluYfkgkQTZ2Rkclg/L3b+ynhYeqdRKEeAOprZW09Im+fNTU8
zVbrwJ+VNPYa+nLdgjHI+L5TwDhtqC/3TMm9boMmlRR+GGXCX/Smy9ioR7WM17Qb
B3m0sw5osccTkyp2YtQhPqO5k6scDMGjdeqVnWEH+b4=
`pragma protect end_protected
