-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
CeW1ZsRcM1lCwIPqtTdfRRgybOHtAWHr4OjC6uN32aO5LlwDwHC+rci3+/9ZcZHp6y/1qrv7N/8q
6BO4BqmnKnY3koPy6D6fJFZ99EIAvkt3UlySQdK0y8rwH7DRyGo0coiPPw4OvAgGFGP+NG2lr4lm
hCtQdIy+clR91Ef8NpeKP6Bi94BhDIABqnYaZND9JLlqP3qid47pzhvBfKkDFl140rRvstABjPdp
2WkBWMqWxgPFKXYJyu6nkKvDRkFZD8ds+6Z6Q1BWJ4Nb2qRyRIf5/kOLPokN8bPXANQ4+cbqo9Yu
V1cuMzAQgrDZVB/e0QqC73/gHj+8HUbc2un+0w==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 3792)
`protect data_block
H2nlDbM3gitmkRIyXXbC0YEqK8rz01aGUYO/XCJto27iw9HvBfmBbafExBCh3zvDKPZWw40kTx6p
LmRZmcGlyve/uMkGx4Vgxc6Edrps9d2xgzuApoT5lfTGxVENQnSKCrMzZ+QRslKV/0GvdXOJXNeP
9+FwAf5um6oJvnFR1IRszmhJNBz01NkjY4Uxfb3SpGfc/Xuh0Uhh5mTlfVk638XfewXnpCTGrnTk
hmLRH0r0ggLiUpwk+99A9xf0ZRhDoVBF2mF4xuiZAKnBPy6Pa97RG315gULWgF6BNXJx0QutqZUt
0bdYsv6QwwUex6U9lW/bIplAEwlqhb+scMa0Y6UTd/mgQz4gn0tn2DzAaS/ZVdu7YlSxwGrvhufT
kck5ExqT4BscIAtU5j6Gc0YB9btO7assyd4iNlYr47WGFS/d9MULODINoTOm7FdXpZswQwVro+Xz
Hr2IvPQcc0sO6nJqWT3Gwmf73Zr4qlbVAqfeIuBR5WdJlVf3WDHoG4jXpyPjmEXz0/FtkPT4cS9X
fAyX7yB6mfsGQqrKR1AclSRk+q1W4HZGlxQQFHiVOmZRbl0n/4I+U1yoLbZdSa2aeN9yxn/OKoQJ
0AF7GZsGL2iJcz+i1Be8eMufTmA8PrYbKZq4Nb1phzZLDgHTdbuccJ6FMojabGRg78g/O+6N+UCX
73jYddk+1sxlwT5gQO8ot6RIJUpcg8IgTUkBY/SnG0xnkADx6mpLI0sh9v+KXERFJd2Q0jd/m/0y
H9RVAg3+1xz/8stCC532b8tvGfDdHy4VuUBtEkPQXoKzVxcdyzddd/Qwty5Osr0MRhzEpJMeuI8K
nU8qskgJB/TK05P7wq/0Alv9L09OB6w5h58SfLXPB4NdJXQQ8FHmsYw3ccq+vwEh+AByT5RU9iCF
8k8h0g5W/bstpXQgE0YLyF4uDGZXh7+AtW/VptL3UcehqsBWQGMQV4yHyo8EcrxwsrvjJHD/TdUr
xbEfrPTfvus3xjPmjjPZOMdxyLX22BzS+56s/3AQxKDDCBsynnYlNClljZcixYTFvvu7nnzWchvi
VSTD9sZEAyMaancuNsXXCGvYgk7jp9U7DfI/eP+VW6pbP0FRncQ2agmZ4n932YAZCpVVVBMyR1Ht
sCD8rSR/TvC9V/eTk1Oo8s3foZ8/+pdnN2iKBVcujyrs7jAVvYW9YYcL8JqozJ/yU2+a4ocwjkJ0
CdvbIfc6mV4/YjBJfrzxMRrO4Ky3xlr48WU3up0HN6UGcfhiP/HRgz6aBnZLTAFWy5lHwxMZ2n1a
qKYtYgBulOUarqW8et6hseQFv7duaTTi+4YbYP5VYDHLXcTogs4g9VwN7iSVPQTYE6e6dEI6qJ05
tNczDRCECOvL87DKh9VcDDwSH06mFuV8wKk2LrZt8wZHLZyQ/4//XsDnbtR0tGV1EclCDA/8SByT
mXtB6LkraXWv0HDlcuRyHK4ro39LGDv9VcX8PBjBzP7QaI6tRXQHygeMRhRKPW05W4BPgHlON64g
2bLja8Yu2DyngTx6x5OHk3lDWmsZX+NAl6ZqgiYCmOxjpC8s7REzeDvEIY6wxvuSOWqj8THFOa2N
coXypaX699y37Qp3b9zY4BXy3CkH6okE35qpYOHswrQAX4PaaeCYgW8jAlN6S+4PIOv2+vSCSQAI
ayJO/5siZl37RaG8Ekzcz5o5Cwl/ZZxKna1AJ1CeUpqxCiOiyoRzZtEY5GUPipCsxF+cd0q+3rKe
RL94vPO4sPvEhBjeLbGu4bxGnk5outUoR+U6Z8JCVC2g0ds11o/gqxnnecO7FVl1Q6vHfxzr8PD9
GmhInpNnhlMAURBvR7nCRzHDkeoW3GEwiS/3RgP+yAkB5UUM9Zwbompm0PdE6iW9hsTaEA4FtaPs
kvwSxAa5/InrOe3yXxTDtg1dbyBVEFKrKMGHG2TalQ0MuUiDiobv/dGheCdivQ5ZaTFZSR1yHd/S
3/nNT9UF3GsE0LSTIKNgQFEdFbMZYNxDtir4aVydaH4MIIfkpwZb4FhGhrFXCHuDHnh1x8nh4NHU
MAMgtPGkKjEnVO8gqA4hbEgf/AeDA+uB05qwNDh7UVJ67NBhiiD9JAjJuu8SwC+iaoiftWCSHJ3g
fmMYXom5OwwgGWIyR8AlOU+IuoQq9op65a8mqx18SNdpD2EunTC4pdgjBh1FN6V2M6uum7iH1HHF
bqU4GujZlELoWagfYAJmYjFL1/nCbtQHlrr29G6JmOjN4O3+UETIdcZhME9SXv/q5+n1o1N9huzm
ao3uS8DIDwfV9p6ahxM4tc3CvHZOhhTd/wBI/fVTiojOTZZIO5/QUd5gReZyeKkGl0tj4kn35klX
HMWfziPfUdU2UedW6fs5JbiNc7CYRxqfdv34+5DwBT9JhPlLRoFFMoReo8DUGnwCYli44zv/wsGd
sK4lCjrkXFaKui+1q+qFpeYrjLf4yUB9A59yw76yZ7X4Wl4pKbsvuW4dL0dAGfEEZyhR+DNSOeZt
uR57jYYY6Hc5sM+qJ7HkM4Z2zwR+Rpd7O66otZrz4hbfJmLS9rky6GSyaD7pOCO95zqj2dKiOlQs
wf12diAB/xgqYf4BELnIqWtL95FHYpa1lncwF7Hwe92FSfPf6z9sqmjJhI8TpldvywthfS2QwxGi
T3Zm8Tk4ycnOMSpDSPL/xsfoyHwcFm1LfzwegQ0tzff0kIqfMouKzvoQePTTb8cFqdxP3W8fhZff
2W4q84NutzdevrOZfog/Kj7uwQXmZeUwI7HilDBvT0VhTePIwEN/NaLYFhMfTT82iuoXxa0up7Ir
nnokV6oU+Sq95LU3f2D34UfvZmW6iTzBZAkdyHFTWTLvNhkn+DG3EWjWTdbGxcjPNq0JHaLSgJTc
6RgK4Khh9I+8UazTtfTAmDaXkD2D4U22P8rKOJve7PBjw7tWLKa4r7yu/+8zlGrFGzG547AkaJWT
GTtlNzcxbgYymxr1zq9cK0JRzQhvQ36OAHr0sAVYVamv0OdDgxyA9TYq7RG/Hn8Vsi+0qsN9nOih
Qa+SNLXqBgezDo4cCbmOZcIdVu27dshac3ku9WC53CZIRgB2BXjDnH6ObJ9K7PbMuyOpF5zh2g9S
dPTqAEe4aj+pd9twd132V1dvH3m7lQo363Yg/oEnPI9RGkmdkzBInBDha9pdUy5IDP/DigCDM1ta
cgD5TDqaUFLxd8HYZ6Pee/sdH97qjKIkNnp2bHrim/sZu+Y65djEcVP+Tm0dACMmyf8o3zmxnAQk
McxTorwuRgVS1FEkq8GVGs54x9e6M+W/qiAtOAPAy7D0L5J1SkH3DFc2gqspvYuocxl1xAjM3YaN
OpRHWKjqiuSaloq8aoPmccSVJvQesl3Nt8fL7lZs4DikXlnQz8OpgZ6QK/64yDsQe6tVfsk+U+h+
dXU6Qx3KjbwqJyE7npCeBpMn0SttbgAJMXB+WmaLv6wbhzlg/KGiL5H0uNbz/BeOz12JIZr5V7dB
oAvoRdwzd9NueuDO48adNSfcw07Cl+1gN9WDKGrIsxDkZZLMsHukOahBcXNT9eiJ281/04RSao/b
+nPVunFmPy6+nPUOAILztbE/oIXLsGwC4V3vLvY+6bPO3i9IGIv6By8TlawNtXxGPMIJb+5qeXJG
I6sbp3wtLK5m4czl6mVoWW/iQwq5f3daGrds6m9J4pFdmHGePp/t4GYvMUaSfX3mejQ6wrb6OM86
LBwvLzRdWicSbauT4QNHCjhXjNjmyJbM1qiRmNwClIps4JzqAWJ3aYC41c52461HW6SfVIKeusz3
PBxQTVhTUfIj3iG+NEtMMbGw5r0TIxIzmRzwNhpoZuavgXta7IfIq2Zi3QNBjpOYEk9ec2mrMOOS
d2UG/tnBb1tZw2+U+ugUXuV7L9RrRQTPGcPbvhg7msGdpHqCYoVbXg3CqBlWqMMyA4AuS+mW71Pb
5vMXr+v5nbPaeZTVfMAaNG7csTKLXnJ7AMmFF+ScoR9++xKtt+JgNMNjm8rA2TrfeA/4hoWDsJtk
xONQnKwkiUopiQgKzgMxDxT64eIQ+/fmeitFiVVsQYjgQ9Vi37u53K+trhLBQ+bUrejLvYBDYhD2
6maw3fh2Q7M+mrLZ8DQe+QUz4AtEW0rTfAt8dKcH/owpgrYX+t663xxU4G03i1x3gsSk+neXPH4H
nbchT5540PUlWAS4CC6YMUMlgULAYkEJJlqu2MiyOZ3N+JXF2rAXwfeMmxZAOfxR9GZUAJ4sGE4U
s6nkWfgAjT6JzMiiFE5n/0Ocsr/epeUIZoDjDQJXE2enrFXdBpjG8+ksYlb/PPgWLxZP77MbvOIM
+a482ZxUziCACCyFgfL9yT+2AnBwYLMyywCUEfitv/vSzQOBbYWqo6CEoBYY6kYdHmTPyymAuHAr
4cGRf046HLrmn/Kiiz/4+DEhBvisCzPvvOaDJsdZ1VTuREayIPN0eNXfp3WLKOHo/dmnEJdkD9yt
SMqMzRtBhhX8vDuzB7ojSkSSKQAKUsdJIzakVnzk7YtY64OHwFcTiv9e2hYs28G0FNF04uUJhjaC
/EkpBjPsNHSOKGp/ibQoi+Y8bvkZNjBsp5Z2+UHMJIsys5msT/BVrIcIq/2iBuqlcBm6AehOYHrf
jK7iYkQvHaFCIH+p+uP8nOdBEJkLRW5rzH20Eso4lqGWkZ4nC/Ws94yZBfLuje9OY0xUe2qsnXLL
FWPirytUXjL9EU0W2V7/z1RbYJl+vsIOEtK902um0Ly7xBi43ot6SIWh3/qiad9uWUhMiQJH+S90
+z3yGCdAxzMlhtiVIoW56A9VhHdDHcj1j1ajguo+udR6txin8GcQZwGlNtnYOoSy7xnT9MMOTJOy
dd6cfrY4j+rjsH0fTrdRK9WsIayA24ceGkEQEBFs6FgisFRLiijjdITFbFTQd3UYdgzzL5WVK0bz
Mx7y4afTA/i35BN8bXjcpqQ2E/vwlcLBXx5pqcT24pkiFYjHs+o8FHPW5hH0MyFFvXBCOirmy0Fr
/Ud/ZFNbVfMibY0H0K63sf4uQwb8IBa0eUIFWDiF
`protect end_protected
